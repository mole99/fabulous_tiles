module RegFile (UserCLK,
    UserCLKo,
    E1BEG,
    E1END,
    E2BEG,
    E2BEGb,
    E2END,
    E2MID,
    E6BEG,
    E6END,
    EE4BEG,
    EE4END,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    NN4BEG,
    NN4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    SS4BEG,
    SS4END,
    W1BEG,
    W1END,
    W2BEG,
    W2BEGb,
    W2END,
    W2MID,
    W6BEG,
    W6END,
    WW4BEG,
    WW4END);
 input UserCLK;
 output UserCLKo;
 output [3:0] E1BEG;
 input [3:0] E1END;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 input [7:0] E2END;
 input [7:0] E2MID;
 output [11:0] E6BEG;
 input [11:0] E6END;
 output [15:0] EE4BEG;
 input [15:0] EE4END;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [15:0] NN4BEG;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 output [15:0] SS4BEG;
 input [15:0] SS4END;
 output [3:0] W1BEG;
 input [3:0] W1END;
 output [7:0] W2BEG;
 output [7:0] W2BEGb;
 input [7:0] W2END;
 input [7:0] W2MID;
 output [11:0] W6BEG;
 input [11:0] W6END;
 output [15:0] WW4BEG;
 input [15:0] WW4END;

 wire AD0;
 wire AD1;
 wire AD2;
 wire AD3;
 wire A_ADR0;
 wire BD0;
 wire BD1;
 wire BD2;
 wire BD3;
 wire B_ADR0;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net411;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net814;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire \Inst_RegFile_32x4.AD_comb[0] ;
 wire \Inst_RegFile_32x4.AD_comb[1] ;
 wire \Inst_RegFile_32x4.AD_comb[2] ;
 wire \Inst_RegFile_32x4.AD_comb[3] ;
 wire \Inst_RegFile_32x4.AD_reg[0] ;
 wire \Inst_RegFile_32x4.AD_reg[1] ;
 wire \Inst_RegFile_32x4.AD_reg[2] ;
 wire \Inst_RegFile_32x4.AD_reg[3] ;
 wire \Inst_RegFile_32x4.BD_comb[0] ;
 wire \Inst_RegFile_32x4.BD_comb[1] ;
 wire \Inst_RegFile_32x4.BD_comb[2] ;
 wire \Inst_RegFile_32x4.BD_comb[3] ;
 wire \Inst_RegFile_32x4.BD_reg[0] ;
 wire \Inst_RegFile_32x4.BD_reg[1] ;
 wire \Inst_RegFile_32x4.BD_reg[2] ;
 wire \Inst_RegFile_32x4.BD_reg[3] ;
 wire \Inst_RegFile_32x4.mem[0][0] ;
 wire \Inst_RegFile_32x4.mem[0][1] ;
 wire \Inst_RegFile_32x4.mem[0][2] ;
 wire \Inst_RegFile_32x4.mem[0][3] ;
 wire \Inst_RegFile_32x4.mem[10][0] ;
 wire \Inst_RegFile_32x4.mem[10][1] ;
 wire \Inst_RegFile_32x4.mem[10][2] ;
 wire \Inst_RegFile_32x4.mem[10][3] ;
 wire \Inst_RegFile_32x4.mem[11][0] ;
 wire \Inst_RegFile_32x4.mem[11][1] ;
 wire \Inst_RegFile_32x4.mem[11][2] ;
 wire \Inst_RegFile_32x4.mem[11][3] ;
 wire \Inst_RegFile_32x4.mem[12][0] ;
 wire \Inst_RegFile_32x4.mem[12][1] ;
 wire \Inst_RegFile_32x4.mem[12][2] ;
 wire \Inst_RegFile_32x4.mem[12][3] ;
 wire \Inst_RegFile_32x4.mem[13][0] ;
 wire \Inst_RegFile_32x4.mem[13][1] ;
 wire \Inst_RegFile_32x4.mem[13][2] ;
 wire \Inst_RegFile_32x4.mem[13][3] ;
 wire \Inst_RegFile_32x4.mem[14][0] ;
 wire \Inst_RegFile_32x4.mem[14][1] ;
 wire \Inst_RegFile_32x4.mem[14][2] ;
 wire \Inst_RegFile_32x4.mem[14][3] ;
 wire \Inst_RegFile_32x4.mem[15][0] ;
 wire \Inst_RegFile_32x4.mem[15][1] ;
 wire \Inst_RegFile_32x4.mem[15][2] ;
 wire \Inst_RegFile_32x4.mem[15][3] ;
 wire \Inst_RegFile_32x4.mem[16][0] ;
 wire \Inst_RegFile_32x4.mem[16][1] ;
 wire \Inst_RegFile_32x4.mem[16][2] ;
 wire \Inst_RegFile_32x4.mem[16][3] ;
 wire \Inst_RegFile_32x4.mem[17][0] ;
 wire \Inst_RegFile_32x4.mem[17][1] ;
 wire \Inst_RegFile_32x4.mem[17][2] ;
 wire \Inst_RegFile_32x4.mem[17][3] ;
 wire \Inst_RegFile_32x4.mem[18][0] ;
 wire \Inst_RegFile_32x4.mem[18][1] ;
 wire \Inst_RegFile_32x4.mem[18][2] ;
 wire \Inst_RegFile_32x4.mem[18][3] ;
 wire \Inst_RegFile_32x4.mem[19][0] ;
 wire \Inst_RegFile_32x4.mem[19][1] ;
 wire \Inst_RegFile_32x4.mem[19][2] ;
 wire \Inst_RegFile_32x4.mem[19][3] ;
 wire \Inst_RegFile_32x4.mem[1][0] ;
 wire \Inst_RegFile_32x4.mem[1][1] ;
 wire \Inst_RegFile_32x4.mem[1][2] ;
 wire \Inst_RegFile_32x4.mem[1][3] ;
 wire \Inst_RegFile_32x4.mem[20][0] ;
 wire \Inst_RegFile_32x4.mem[20][1] ;
 wire \Inst_RegFile_32x4.mem[20][2] ;
 wire \Inst_RegFile_32x4.mem[20][3] ;
 wire \Inst_RegFile_32x4.mem[21][0] ;
 wire \Inst_RegFile_32x4.mem[21][1] ;
 wire \Inst_RegFile_32x4.mem[21][2] ;
 wire \Inst_RegFile_32x4.mem[21][3] ;
 wire \Inst_RegFile_32x4.mem[22][0] ;
 wire \Inst_RegFile_32x4.mem[22][1] ;
 wire \Inst_RegFile_32x4.mem[22][2] ;
 wire \Inst_RegFile_32x4.mem[22][3] ;
 wire \Inst_RegFile_32x4.mem[23][0] ;
 wire \Inst_RegFile_32x4.mem[23][1] ;
 wire \Inst_RegFile_32x4.mem[23][2] ;
 wire \Inst_RegFile_32x4.mem[23][3] ;
 wire \Inst_RegFile_32x4.mem[24][0] ;
 wire \Inst_RegFile_32x4.mem[24][1] ;
 wire \Inst_RegFile_32x4.mem[24][2] ;
 wire \Inst_RegFile_32x4.mem[24][3] ;
 wire \Inst_RegFile_32x4.mem[25][0] ;
 wire \Inst_RegFile_32x4.mem[25][1] ;
 wire \Inst_RegFile_32x4.mem[25][2] ;
 wire \Inst_RegFile_32x4.mem[25][3] ;
 wire \Inst_RegFile_32x4.mem[26][0] ;
 wire \Inst_RegFile_32x4.mem[26][1] ;
 wire \Inst_RegFile_32x4.mem[26][2] ;
 wire \Inst_RegFile_32x4.mem[26][3] ;
 wire \Inst_RegFile_32x4.mem[27][0] ;
 wire \Inst_RegFile_32x4.mem[27][1] ;
 wire \Inst_RegFile_32x4.mem[27][2] ;
 wire \Inst_RegFile_32x4.mem[27][3] ;
 wire \Inst_RegFile_32x4.mem[28][0] ;
 wire \Inst_RegFile_32x4.mem[28][1] ;
 wire \Inst_RegFile_32x4.mem[28][2] ;
 wire \Inst_RegFile_32x4.mem[28][3] ;
 wire \Inst_RegFile_32x4.mem[29][0] ;
 wire \Inst_RegFile_32x4.mem[29][1] ;
 wire \Inst_RegFile_32x4.mem[29][2] ;
 wire \Inst_RegFile_32x4.mem[29][3] ;
 wire \Inst_RegFile_32x4.mem[2][0] ;
 wire \Inst_RegFile_32x4.mem[2][1] ;
 wire \Inst_RegFile_32x4.mem[2][2] ;
 wire \Inst_RegFile_32x4.mem[2][3] ;
 wire \Inst_RegFile_32x4.mem[30][0] ;
 wire \Inst_RegFile_32x4.mem[30][1] ;
 wire \Inst_RegFile_32x4.mem[30][2] ;
 wire \Inst_RegFile_32x4.mem[30][3] ;
 wire \Inst_RegFile_32x4.mem[31][0] ;
 wire \Inst_RegFile_32x4.mem[31][1] ;
 wire \Inst_RegFile_32x4.mem[31][2] ;
 wire \Inst_RegFile_32x4.mem[31][3] ;
 wire \Inst_RegFile_32x4.mem[3][0] ;
 wire \Inst_RegFile_32x4.mem[3][1] ;
 wire \Inst_RegFile_32x4.mem[3][2] ;
 wire \Inst_RegFile_32x4.mem[3][3] ;
 wire \Inst_RegFile_32x4.mem[4][0] ;
 wire \Inst_RegFile_32x4.mem[4][1] ;
 wire \Inst_RegFile_32x4.mem[4][2] ;
 wire \Inst_RegFile_32x4.mem[4][3] ;
 wire \Inst_RegFile_32x4.mem[5][0] ;
 wire \Inst_RegFile_32x4.mem[5][1] ;
 wire \Inst_RegFile_32x4.mem[5][2] ;
 wire \Inst_RegFile_32x4.mem[5][3] ;
 wire \Inst_RegFile_32x4.mem[6][0] ;
 wire \Inst_RegFile_32x4.mem[6][1] ;
 wire \Inst_RegFile_32x4.mem[6][2] ;
 wire \Inst_RegFile_32x4.mem[6][3] ;
 wire \Inst_RegFile_32x4.mem[7][0] ;
 wire \Inst_RegFile_32x4.mem[7][1] ;
 wire \Inst_RegFile_32x4.mem[7][2] ;
 wire \Inst_RegFile_32x4.mem[7][3] ;
 wire \Inst_RegFile_32x4.mem[8][0] ;
 wire \Inst_RegFile_32x4.mem[8][1] ;
 wire \Inst_RegFile_32x4.mem[8][2] ;
 wire \Inst_RegFile_32x4.mem[8][3] ;
 wire \Inst_RegFile_32x4.mem[9][0] ;
 wire \Inst_RegFile_32x4.mem[9][1] ;
 wire \Inst_RegFile_32x4.mem[9][2] ;
 wire \Inst_RegFile_32x4.mem[9][3] ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Inst_RegFile_switch_matrix.E1BEG0 ;
 wire \Inst_RegFile_switch_matrix.E1BEG1 ;
 wire \Inst_RegFile_switch_matrix.E1BEG2 ;
 wire \Inst_RegFile_switch_matrix.E1BEG3 ;
 wire \Inst_RegFile_switch_matrix.E2BEG0 ;
 wire \Inst_RegFile_switch_matrix.E2BEG1 ;
 wire \Inst_RegFile_switch_matrix.E2BEG2 ;
 wire \Inst_RegFile_switch_matrix.E2BEG3 ;
 wire \Inst_RegFile_switch_matrix.E2BEG4 ;
 wire \Inst_RegFile_switch_matrix.E2BEG5 ;
 wire \Inst_RegFile_switch_matrix.E2BEG6 ;
 wire \Inst_RegFile_switch_matrix.E2BEG7 ;
 wire \Inst_RegFile_switch_matrix.E6BEG0 ;
 wire \Inst_RegFile_switch_matrix.E6BEG1 ;
 wire \Inst_RegFile_switch_matrix.EE4BEG0 ;
 wire \Inst_RegFile_switch_matrix.EE4BEG1 ;
 wire \Inst_RegFile_switch_matrix.EE4BEG2 ;
 wire \Inst_RegFile_switch_matrix.EE4BEG3 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG0 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG1 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG2 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG3 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG4 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG5 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG6 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG7 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG0 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG1 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG2 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG3 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG4 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG5 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG6 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG7 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG0 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG1 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG2 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG3 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG4 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG5 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG6 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG7 ;
 wire \Inst_RegFile_switch_matrix.N1BEG0 ;
 wire \Inst_RegFile_switch_matrix.N1BEG1 ;
 wire \Inst_RegFile_switch_matrix.N1BEG2 ;
 wire \Inst_RegFile_switch_matrix.N1BEG3 ;
 wire \Inst_RegFile_switch_matrix.N4BEG0 ;
 wire \Inst_RegFile_switch_matrix.N4BEG1 ;
 wire \Inst_RegFile_switch_matrix.N4BEG2 ;
 wire \Inst_RegFile_switch_matrix.N4BEG3 ;
 wire \Inst_RegFile_switch_matrix.NN4BEG0 ;
 wire \Inst_RegFile_switch_matrix.NN4BEG1 ;
 wire \Inst_RegFile_switch_matrix.NN4BEG2 ;
 wire \Inst_RegFile_switch_matrix.NN4BEG3 ;
 wire \Inst_RegFile_switch_matrix.S1BEG0 ;
 wire \Inst_RegFile_switch_matrix.S1BEG1 ;
 wire \Inst_RegFile_switch_matrix.S1BEG2 ;
 wire \Inst_RegFile_switch_matrix.S1BEG3 ;
 wire \Inst_RegFile_switch_matrix.S4BEG0 ;
 wire \Inst_RegFile_switch_matrix.S4BEG1 ;
 wire \Inst_RegFile_switch_matrix.S4BEG2 ;
 wire \Inst_RegFile_switch_matrix.S4BEG3 ;
 wire \Inst_RegFile_switch_matrix.SS4BEG0 ;
 wire \Inst_RegFile_switch_matrix.SS4BEG1 ;
 wire \Inst_RegFile_switch_matrix.SS4BEG2 ;
 wire \Inst_RegFile_switch_matrix.SS4BEG3 ;
 wire \Inst_RegFile_switch_matrix.W1BEG0 ;
 wire \Inst_RegFile_switch_matrix.W1BEG1 ;
 wire \Inst_RegFile_switch_matrix.W1BEG2 ;
 wire \Inst_RegFile_switch_matrix.W1BEG3 ;
 wire \Inst_RegFile_switch_matrix.W6BEG0 ;
 wire \Inst_RegFile_switch_matrix.W6BEG1 ;
 wire \Inst_RegFile_switch_matrix.WW4BEG0 ;
 wire \Inst_RegFile_switch_matrix.WW4BEG1 ;
 wire \Inst_RegFile_switch_matrix.WW4BEG2 ;
 wire \Inst_RegFile_switch_matrix.WW4BEG3 ;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net811;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net815;
 wire net282;
 wire net817;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net593;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net816;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net813;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net812;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire UserCLK_regs;
 wire clknet_0_UserCLK;
 wire clknet_1_0__leaf_UserCLK;
 wire clknet_0_UserCLK_regs;
 wire clknet_4_0_0_UserCLK_regs;
 wire clknet_4_1_0_UserCLK_regs;
 wire clknet_4_2_0_UserCLK_regs;
 wire clknet_4_3_0_UserCLK_regs;
 wire clknet_4_4_0_UserCLK_regs;
 wire clknet_4_5_0_UserCLK_regs;
 wire clknet_4_6_0_UserCLK_regs;
 wire clknet_4_7_0_UserCLK_regs;
 wire clknet_4_8_0_UserCLK_regs;
 wire clknet_4_9_0_UserCLK_regs;
 wire clknet_4_10_0_UserCLK_regs;
 wire clknet_4_11_0_UserCLK_regs;
 wire clknet_4_12_0_UserCLK_regs;
 wire clknet_4_13_0_UserCLK_regs;
 wire clknet_4_14_0_UserCLK_regs;
 wire clknet_4_15_0_UserCLK_regs;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net408;
 wire net409;
 wire net410;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;

 sky130_fd_sc_hd__inv_1 _1041_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ),
    .Y(_0933_));
 sky130_fd_sc_hd__inv_1 _1042_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q ),
    .Y(_0934_));
 sky130_fd_sc_hd__inv_1 _1043_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ),
    .Y(_0935_));
 sky130_fd_sc_hd__inv_2 _1044_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ),
    .Y(_0936_));
 sky130_fd_sc_hd__inv_1 _1045_ (.A(\Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ),
    .Y(_0937_));
 sky130_fd_sc_hd__inv_1 _1046_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ),
    .Y(_0938_));
 sky130_fd_sc_hd__inv_2 _1047_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q ),
    .Y(_0939_));
 sky130_fd_sc_hd__inv_2 _1048_ (.A(\Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q ),
    .Y(_0940_));
 sky130_fd_sc_hd__inv_2 _1049_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ),
    .Y(_0941_));
 sky130_fd_sc_hd__inv_1 _1050_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ),
    .Y(_0942_));
 sky130_fd_sc_hd__inv_2 _1051_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ),
    .Y(_0943_));
 sky130_fd_sc_hd__inv_2 _1052_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q ),
    .Y(_0944_));
 sky130_fd_sc_hd__inv_2 _1053_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q ),
    .Y(_0945_));
 sky130_fd_sc_hd__inv_2 _1054_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q ),
    .Y(_0946_));
 sky130_fd_sc_hd__inv_1 _1055_ (.A(net103),
    .Y(_0947_));
 sky130_fd_sc_hd__inv_1 _1056_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ),
    .Y(_0948_));
 sky130_fd_sc_hd__inv_1 _1057_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q ),
    .Y(_0949_));
 sky130_fd_sc_hd__inv_2 _1058_ (.A(net131),
    .Y(_0950_));
 sky130_fd_sc_hd__inv_2 _1059_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ),
    .Y(_0951_));
 sky130_fd_sc_hd__inv_1 _1060_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q ),
    .Y(_0952_));
 sky130_fd_sc_hd__inv_1 _1061_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_0953_));
 sky130_fd_sc_hd__inv_2 _1062_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ),
    .Y(_0954_));
 sky130_fd_sc_hd__inv_1 _1063_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ),
    .Y(_0955_));
 sky130_fd_sc_hd__inv_1 _1064_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q ),
    .Y(_0956_));
 sky130_fd_sc_hd__inv_1 _1065_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ),
    .Y(_0957_));
 sky130_fd_sc_hd__inv_2 _1066_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q ),
    .Y(_0958_));
 sky130_fd_sc_hd__inv_1 _1067_ (.A(\Inst_RegFile_32x4.mem[22][0] ),
    .Y(_0959_));
 sky130_fd_sc_hd__inv_1 _1068_ (.A(\Inst_RegFile_32x4.mem[22][2] ),
    .Y(_0960_));
 sky130_fd_sc_hd__inv_2 _1069_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ),
    .Y(_0961_));
 sky130_fd_sc_hd__inv_1 _1070_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q ),
    .Y(_0962_));
 sky130_fd_sc_hd__inv_1 _1071_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ),
    .Y(_0963_));
 sky130_fd_sc_hd__inv_1 _1072_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q ),
    .Y(_0964_));
 sky130_fd_sc_hd__inv_2 _1073_ (.A(\Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q ),
    .Y(_0965_));
 sky130_fd_sc_hd__inv_2 _1074_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q ),
    .Y(_0966_));
 sky130_fd_sc_hd__inv_2 _1075_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q ),
    .Y(_0967_));
 sky130_fd_sc_hd__inv_2 _1076_ (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ),
    .Y(_0968_));
 sky130_fd_sc_hd__inv_2 _1077_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ),
    .Y(_0969_));
 sky130_fd_sc_hd__inv_1 _1078_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q ),
    .Y(_0970_));
 sky130_fd_sc_hd__inv_1 _1079_ (.A(net75),
    .Y(_0971_));
 sky130_fd_sc_hd__inv_1 _1080_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ),
    .Y(_0972_));
 sky130_fd_sc_hd__inv_2 _1081_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q ),
    .Y(_0973_));
 sky130_fd_sc_hd__inv_1 _1082_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ),
    .Y(_0974_));
 sky130_fd_sc_hd__inv_1 _1083_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q ),
    .Y(_0975_));
 sky130_fd_sc_hd__inv_1 _1084_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q ),
    .Y(_0976_));
 sky130_fd_sc_hd__inv_2 _1085_ (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ),
    .Y(_0977_));
 sky130_fd_sc_hd__inv_1 _1086_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ),
    .Y(_0978_));
 sky130_fd_sc_hd__inv_1 _1087_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q ),
    .Y(_0979_));
 sky130_fd_sc_hd__inv_1 _1088_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q ),
    .Y(_0980_));
 sky130_fd_sc_hd__inv_1 _1089_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ),
    .Y(_0981_));
 sky130_fd_sc_hd__inv_1 _1090_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q ),
    .Y(_0982_));
 sky130_fd_sc_hd__inv_2 _1091_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ),
    .Y(_0983_));
 sky130_fd_sc_hd__inv_2 _1092_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ),
    .Y(_0984_));
 sky130_fd_sc_hd__inv_1 _1093_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q ),
    .Y(_0985_));
 sky130_fd_sc_hd__inv_2 _1094_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ),
    .Y(_0986_));
 sky130_fd_sc_hd__inv_2 _1095_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q ),
    .Y(_0987_));
 sky130_fd_sc_hd__inv_1 _1096_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0988_));
 sky130_fd_sc_hd__inv_1 _1097_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q ),
    .Y(_0989_));
 sky130_fd_sc_hd__inv_1 _1098_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ),
    .Y(_0990_));
 sky130_fd_sc_hd__inv_1 _1099_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q ),
    .Y(_0991_));
 sky130_fd_sc_hd__inv_2 _1100_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ),
    .Y(_0992_));
 sky130_fd_sc_hd__inv_1 _1101_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q ),
    .Y(_0993_));
 sky130_fd_sc_hd__inv_1 _1102_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ),
    .Y(_0994_));
 sky130_fd_sc_hd__inv_1 _1103_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q ),
    .Y(_0995_));
 sky130_fd_sc_hd__inv_1 _1104_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ),
    .Y(_0996_));
 sky130_fd_sc_hd__inv_1 _1105_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q ),
    .Y(_0997_));
 sky130_fd_sc_hd__inv_1 _1106_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ),
    .Y(_0998_));
 sky130_fd_sc_hd__inv_1 _1107_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q ),
    .Y(_0999_));
 sky130_fd_sc_hd__inv_2 _1108_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q ),
    .Y(_1000_));
 sky130_fd_sc_hd__inv_1 _1109_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q ),
    .Y(_1001_));
 sky130_fd_sc_hd__inv_1 _1110_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ),
    .Y(_1002_));
 sky130_fd_sc_hd__inv_2 _1111_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ),
    .Y(_1003_));
 sky130_fd_sc_hd__inv_1 _1112_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q ),
    .Y(_1004_));
 sky130_fd_sc_hd__inv_2 _1113_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ),
    .Y(_1005_));
 sky130_fd_sc_hd__inv_1 _1114_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q ),
    .Y(_1006_));
 sky130_fd_sc_hd__inv_1 _1115_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ),
    .Y(_1007_));
 sky130_fd_sc_hd__inv_1 _1116_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q ),
    .Y(_1008_));
 sky130_fd_sc_hd__inv_1 _1117_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ),
    .Y(_1009_));
 sky130_fd_sc_hd__inv_1 _1118_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q ),
    .Y(_1010_));
 sky130_fd_sc_hd__inv_1 _1119_ (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q ),
    .Y(_1011_));
 sky130_fd_sc_hd__inv_1 _1120_ (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q ),
    .Y(_1012_));
 sky130_fd_sc_hd__inv_1 _1121_ (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q ),
    .Y(_1013_));
 sky130_fd_sc_hd__inv_1 _1122_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q ),
    .Y(_1014_));
 sky130_fd_sc_hd__inv_2 _1123_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .Y(_1015_));
 sky130_fd_sc_hd__inv_2 _1124_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ),
    .Y(_1016_));
 sky130_fd_sc_hd__inv_2 _1125_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q ),
    .Y(_1017_));
 sky130_fd_sc_hd__inv_2 _1126_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q ),
    .Y(_1018_));
 sky130_fd_sc_hd__inv_2 _1127_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ),
    .Y(_1019_));
 sky130_fd_sc_hd__mux4_2 _1128_ (.A0(net647),
    .A1(net679),
    .A2(net636),
    .A3(net641),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1020_));
 sky130_fd_sc_hd__or2_4 _1129_ (.A(_0966_),
    .B(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__mux4_1 _1130_ (.A0(net689),
    .A1(net672),
    .A2(net660),
    .A3(net653),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1022_));
 sky130_fd_sc_hd__o21a_1 _1131_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q ),
    .A2(_1022_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q ),
    .X(_1023_));
 sky130_fd_sc_hd__mux4_1 _1132_ (.A0(net25),
    .A1(net87),
    .A2(net89),
    .A3(net97),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1024_));
 sky130_fd_sc_hd__mux4_1 _1133_ (.A0(net61),
    .A1(net69),
    .A2(net780),
    .A3(net11),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1025_));
 sky130_fd_sc_hd__mux2_1 _1134_ (.A0(_1024_),
    .A1(_1025_),
    .S(_0966_),
    .X(_1026_));
 sky130_fd_sc_hd__a22o_1 _1135_ (.A1(_1021_),
    .A2(_1023_),
    .B1(_1026_),
    .B2(_0967_),
    .X(\Inst_RegFile_switch_matrix.E2BEG5 ));
 sky130_fd_sc_hd__a221o_1 _1136_ (.A1(_1021_),
    .A2(_1023_),
    .B1(_1026_),
    .B2(_0967_),
    .C1(_0965_),
    .X(_1027_));
 sky130_fd_sc_hd__o21a_1 _1137_ (.A1(net101),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q ),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q ),
    .X(_1028_));
 sky130_fd_sc_hd__o21ba_1 _1138_ (.A1(net73),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q ),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q ),
    .X(_1029_));
 sky130_fd_sc_hd__o21a_1 _1139_ (.A1(net15),
    .A2(_0965_),
    .B1(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__a21o_1 _1140_ (.A1(_1028_),
    .A2(_1027_),
    .B1(_1030_),
    .X(_1031_));
 sky130_fd_sc_hd__a211o_1 _1141_ (.A1(_1027_),
    .A2(_1028_),
    .B1(_1030_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_1032_));
 sky130_fd_sc_hd__mux4_2 _1142_ (.A0(net74),
    .A1(net16),
    .A2(net102),
    .A3(net130),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q ),
    .X(_1033_));
 sky130_fd_sc_hd__o21ba_1 _1143_ (.A1(_0968_),
    .A2(_1033_),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q ),
    .X(_1034_));
 sky130_fd_sc_hd__mux4_2 _1144_ (.A0(net687),
    .A1(net670),
    .A2(net657),
    .A3(net651),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_1035_));
 sky130_fd_sc_hd__or2_4 _1145_ (.A(_1035_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ),
    .X(_1036_));
 sky130_fd_sc_hd__mux4_2 _1146_ (.A0(net679),
    .A1(net636),
    .A2(net668),
    .A3(net640),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ),
    .X(_1037_));
 sky130_fd_sc_hd__o21a_1 _1147_ (.A1(_0957_),
    .A2(_1037_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_1038_));
 sky130_fd_sc_hd__mux4_1 _1148_ (.A0(net61),
    .A1(net67),
    .A2(net79),
    .A3(net9),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_1039_));
 sky130_fd_sc_hd__mux4_1 _1149_ (.A0(net21),
    .A1(net95),
    .A2(net114),
    .A3(net123),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_1040_));
 sky130_fd_sc_hd__mux2_1 _1150_ (.A0(_1039_),
    .A1(_1040_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ),
    .X(_0128_));
 sky130_fd_sc_hd__a22o_4 _1151_ (.A1(net414),
    .A2(_1038_),
    .B1(_0128_),
    .B2(_0958_),
    .X(\Inst_RegFile_switch_matrix.E2BEG3 ));
 sky130_fd_sc_hd__a221o_2 _1152_ (.A1(_1038_),
    .A2(_1036_),
    .B1(_0128_),
    .B2(_0958_),
    .C1(_0969_),
    .X(_0129_));
 sky130_fd_sc_hd__o21a_1 _1153_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ),
    .A2(net109),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _1154_ (.A0(net85),
    .A1(net7),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_0131_));
 sky130_fd_sc_hd__a221o_1 _1155_ (.A1(_0130_),
    .A2(_0129_),
    .B1(_0131_),
    .B2(_0970_),
    .C1(_0968_),
    .X(_0132_));
 sky130_fd_sc_hd__mux4_2 _1156_ (.A0(net66),
    .A1(net8),
    .A2(net94),
    .A3(net138),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q ),
    .X(_0133_));
 sky130_fd_sc_hd__or2_1 _1157_ (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ),
    .B(_0133_),
    .X(_0134_));
 sky130_fd_sc_hd__a32oi_4 _1158_ (.A1(_0132_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q ),
    .A3(_0134_),
    .B1(_1032_),
    .B2(_1034_),
    .Y(_0135_));
 sky130_fd_sc_hd__a32o_1 _1159_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q ),
    .A2(_0132_),
    .A3(_0134_),
    .B1(_1032_),
    .B2(_1034_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _1160_ (.A0(\Inst_RegFile_32x4.mem[26][0] ),
    .A1(\Inst_RegFile_32x4.mem[27][0] ),
    .S(net625),
    .X(_0137_));
 sky130_fd_sc_hd__mux4_1 _1161_ (.A0(net689),
    .A1(net672),
    .A2(net660),
    .A3(net654),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_0138_));
 sky130_fd_sc_hd__or2_1 _1162_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ),
    .B(_0138_),
    .X(_0139_));
 sky130_fd_sc_hd__mux4_1 _1163_ (.A0(net647),
    .A1(net680),
    .A2(net636),
    .A3(net641),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_0140_));
 sky130_fd_sc_hd__o21a_1 _1164_ (.A1(_0972_),
    .A2(_0140_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_0141_));
 sky130_fd_sc_hd__mux4_1 _1165_ (.A0(net61),
    .A1(net69),
    .A2(net780),
    .A3(net11),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_0142_));
 sky130_fd_sc_hd__mux4_1 _1166_ (.A0(net89),
    .A1(net97),
    .A2(net113),
    .A3(net115),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _1167_ (.A0(_0142_),
    .A1(_0143_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ),
    .X(_0144_));
 sky130_fd_sc_hd__a22oi_4 _1168_ (.A1(_0141_),
    .A2(_0139_),
    .B1(_0144_),
    .B2(_0973_),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_4 _1169_ (.A(_0145_),
    .Y(\Inst_RegFile_switch_matrix.JS2BEG5 ));
 sky130_fd_sc_hd__mux4_2 _1170_ (.A0(_0971_),
    .A1(_0950_),
    .A2(_0947_),
    .A3(_0145_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_0146_));
 sky130_fd_sc_hd__inv_2 _1171_ (.A(_0146_),
    .Y(_0147_));
 sky130_fd_sc_hd__mux4_2 _1172_ (.A0(net76),
    .A1(net18),
    .A2(net104),
    .A3(net132),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q ),
    .X(_0148_));
 sky130_fd_sc_hd__a21oi_1 _1173_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_0148_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q ),
    .Y(_0149_));
 sky130_fd_sc_hd__o21ai_1 _1174_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_0146_),
    .B1(_0149_),
    .Y(_0150_));
 sky130_fd_sc_hd__mux4_2 _1175_ (.A0(net687),
    .A1(net671),
    .A2(net658),
    .A3(net652),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0151_));
 sky130_fd_sc_hd__or2_4 _1176_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ),
    .B(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__mux4_1 _1177_ (.A0(net676),
    .A1(net635),
    .A2(net666),
    .A3(net409),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0153_));
 sky130_fd_sc_hd__o21a_1 _1178_ (.A1(_0974_),
    .A2(_0153_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q ),
    .X(_0154_));
 sky130_fd_sc_hd__mux4_1 _1179_ (.A0(net67),
    .A1(net9),
    .A2(net780),
    .A3(net26),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0155_));
 sky130_fd_sc_hd__mux4_1 _1180_ (.A0(net778),
    .A1(net95),
    .A2(net107),
    .A3(net123),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _1181_ (.A0(_0155_),
    .A1(_0156_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ),
    .X(_0157_));
 sky130_fd_sc_hd__a22o_4 _1182_ (.A1(_0154_),
    .A2(_0152_),
    .B1(_0157_),
    .B2(_0975_),
    .X(\Inst_RegFile_switch_matrix.JS2BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1183_ (.A0(net80),
    .A1(net123),
    .A2(net112),
    .A3(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q ),
    .X(_0158_));
 sky130_fd_sc_hd__mux4_1 _1184_ (.A0(net68),
    .A1(net10),
    .A2(net112),
    .A3(net124),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q ),
    .X(_0159_));
 sky130_fd_sc_hd__inv_1 _1185_ (.A(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__o21ai_1 _1186_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_0160_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q ),
    .Y(_0161_));
 sky130_fd_sc_hd__a21o_1 _1187_ (.A1(_0158_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ),
    .B1(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__and2_4 _1188_ (.A(_0150_),
    .B(_0162_),
    .X(_0163_));
 sky130_fd_sc_hd__nand2_1 _1189_ (.A(_0150_),
    .B(_0162_),
    .Y(_0164_));
 sky130_fd_sc_hd__mux2_1 _1190_ (.A0(\Inst_RegFile_32x4.mem[24][0] ),
    .A1(\Inst_RegFile_32x4.mem[25][0] ),
    .S(net624),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _1191_ (.A0(_0137_),
    .A1(_0165_),
    .S(net396),
    .X(_0166_));
 sky130_fd_sc_hd__nand2_1 _1192_ (.A(net648),
    .B(_0166_),
    .Y(_0167_));
 sky130_fd_sc_hd__mux4_1 _1193_ (.A0(net687),
    .A1(net669),
    .A2(net656),
    .A3(net651),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0168_));
 sky130_fd_sc_hd__or2_1 _1194_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ),
    .B(_0168_),
    .X(_0169_));
 sky130_fd_sc_hd__mux4_2 _1195_ (.A0(net676),
    .A1(net633),
    .A2(net664),
    .A3(net638),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ),
    .X(_0170_));
 sky130_fd_sc_hd__o21a_1 _1196_ (.A1(_0170_),
    .A2(_0978_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0171_));
 sky130_fd_sc_hd__mux4_1 _1197_ (.A0(net61),
    .A1(net67),
    .A2(net86),
    .A3(net9),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0172_));
 sky130_fd_sc_hd__mux4_1 _1198_ (.A0(net778),
    .A1(net95),
    .A2(net107),
    .A3(net123),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _1199_ (.A0(_0172_),
    .A1(_0173_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ),
    .X(_0174_));
 sky130_fd_sc_hd__a22o_4 _1200_ (.A1(_0171_),
    .A2(_0169_),
    .B1(_0174_),
    .B2(_0979_),
    .X(\Inst_RegFile_switch_matrix.JW2BEG3 ));
 sky130_fd_sc_hd__mux2_4 _1201_ (.A0(net138),
    .A1(\Inst_RegFile_switch_matrix.JW2BEG3 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q ),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _1202_ (.A0(net26),
    .A1(net107),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q ),
    .X(_0176_));
 sky130_fd_sc_hd__o21a_1 _1203_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q ),
    .A2(_0176_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ),
    .X(_0177_));
 sky130_fd_sc_hd__o21ai_4 _1204_ (.A1(_0980_),
    .A2(_0175_),
    .B1(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__mux4_2 _1205_ (.A0(net85),
    .A1(net6),
    .A2(net92),
    .A3(net120),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q ),
    .X(_0179_));
 sky130_fd_sc_hd__nand2_1 _1206_ (.A(_0977_),
    .B(_0179_),
    .Y(_0180_));
 sky130_fd_sc_hd__mux4_1 _1207_ (.A0(net139),
    .A1(net672),
    .A2(net659),
    .A3(net653),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_0181_));
 sky130_fd_sc_hd__mux4_2 _1208_ (.A0(net646),
    .A1(net679),
    .A2(net636),
    .A3(net640),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_4 _1209_ (.A0(_0181_),
    .A1(_0182_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ),
    .X(_0183_));
 sky130_fd_sc_hd__mux4_1 _1210_ (.A0(net61),
    .A1(net69),
    .A2(net3),
    .A3(net11),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_0184_));
 sky130_fd_sc_hd__and2b_1 _1211_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ),
    .B(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__mux4_1 _1212_ (.A0(net87),
    .A1(net97),
    .A2(net89),
    .A3(net689),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .X(_0186_));
 sky130_fd_sc_hd__a21o_1 _1213_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ),
    .A2(_0186_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q ),
    .X(_0187_));
 sky130_fd_sc_hd__o22a_4 _1214_ (.A1(_0183_),
    .A2(_0976_),
    .B1(_0185_),
    .B2(_0187_),
    .X(\Inst_RegFile_switch_matrix.JW2BEG5 ));
 sky130_fd_sc_hd__mux4_1 _1215_ (.A0(net13),
    .A1(net127),
    .A2(net99),
    .A3(\Inst_RegFile_switch_matrix.JW2BEG5 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q ),
    .X(_0188_));
 sky130_fd_sc_hd__mux4_1 _1216_ (.A0(net72),
    .A1(net14),
    .A2(net100),
    .A3(net128),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q ),
    .X(_0189_));
 sky130_fd_sc_hd__a21o_1 _1217_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ),
    .A2(_0189_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q ),
    .X(_0190_));
 sky130_fd_sc_hd__a21oi_1 _1218_ (.A1(_0977_),
    .A2(_0188_),
    .B1(_0190_),
    .Y(_0191_));
 sky130_fd_sc_hd__a31o_4 _1219_ (.A1(_0178_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q ),
    .A3(_0180_),
    .B1(_0191_),
    .X(_0192_));
 sky130_fd_sc_hd__clkinv_2 _1220_ (.A(_0192_),
    .Y(_0193_));
 sky130_fd_sc_hd__mux2_1 _1221_ (.A0(\Inst_RegFile_32x4.mem[28][0] ),
    .A1(\Inst_RegFile_32x4.mem[29][0] ),
    .S(net624),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _1222_ (.A0(\Inst_RegFile_32x4.mem[30][0] ),
    .A1(\Inst_RegFile_32x4.mem[31][0] ),
    .S(net624),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _1223_ (.A0(_0194_),
    .A1(_0195_),
    .S(net663),
    .X(_0196_));
 sky130_fd_sc_hd__a21oi_1 _1224_ (.A1(net408),
    .A2(_0196_),
    .B1(net395),
    .Y(_0197_));
 sky130_fd_sc_hd__mux2_1 _1225_ (.A0(\Inst_RegFile_32x4.mem[16][0] ),
    .A1(\Inst_RegFile_32x4.mem[17][0] ),
    .S(net631),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _1226_ (.A0(\Inst_RegFile_32x4.mem[18][0] ),
    .A1(\Inst_RegFile_32x4.mem[19][0] ),
    .S(net631),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _1227_ (.A0(_0198_),
    .A1(_0199_),
    .S(net662),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _1228_ (.A0(\Inst_RegFile_32x4.mem[22][0] ),
    .A1(\Inst_RegFile_32x4.mem[23][0] ),
    .S(net627),
    .X(_0201_));
 sky130_fd_sc_hd__or2_1 _1229_ (.A(net675),
    .B(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _1230_ (.A0(\Inst_RegFile_32x4.mem[20][0] ),
    .A1(\Inst_RegFile_32x4.mem[21][0] ),
    .S(net627),
    .X(_0203_));
 sky130_fd_sc_hd__o211a_1 _1231_ (.A1(net661),
    .A2(_0203_),
    .B1(_0202_),
    .C1(net650),
    .X(_0204_));
 sky130_fd_sc_hd__a211o_1 _1232_ (.A1(_0164_),
    .A2(_0200_),
    .B1(_0204_),
    .C1(_0193_),
    .X(_0205_));
 sky130_fd_sc_hd__mux4_1 _1233_ (.A0(net117),
    .A1(net672),
    .A2(net659),
    .A3(net653),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_0206_));
 sky130_fd_sc_hd__or2_1 _1234_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ),
    .B(_0206_),
    .X(_0207_));
 sky130_fd_sc_hd__mux4_1 _1235_ (.A0(net646),
    .A1(net679),
    .A2(net636),
    .A3(net640),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_0208_));
 sky130_fd_sc_hd__o21a_1 _1236_ (.A1(_0961_),
    .A2(_0208_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q ),
    .X(_0209_));
 sky130_fd_sc_hd__mux4_1 _1237_ (.A0(net11),
    .A1(net89),
    .A2(net97),
    .A3(net115),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_0210_));
 sky130_fd_sc_hd__mux4_1 _1238_ (.A0(net61),
    .A1(net85),
    .A2(net69),
    .A3(net780),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _1239_ (.A0(_0210_),
    .A1(_0211_),
    .S(_0961_),
    .X(_0212_));
 sky130_fd_sc_hd__a22o_4 _1240_ (.A1(_0209_),
    .A2(_0207_),
    .B1(_0212_),
    .B2(_0962_),
    .X(\Inst_RegFile_switch_matrix.JN2BEG5 ));
 sky130_fd_sc_hd__mux4_2 _1241_ (.A0(net63),
    .A1(net91),
    .A2(net24),
    .A3(net119),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q ),
    .X(_0213_));
 sky130_fd_sc_hd__mux4_1 _1242_ (.A0(_0213_),
    .A1(\Inst_RegFile_switch_matrix.JN2BEG5 ),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG5 ),
    .A3(\Inst_RegFile_switch_matrix.JW2BEG5 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q ),
    .X(_0214_));
 sky130_fd_sc_hd__mux4_1 _1243_ (.A0(net688),
    .A1(net672),
    .A2(net659),
    .A3(net653),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_0215_));
 sky130_fd_sc_hd__or2_1 _1244_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ),
    .B(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__mux4_1 _1245_ (.A0(net422),
    .A1(net680),
    .A2(net667),
    .A3(net641),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_0217_));
 sky130_fd_sc_hd__o21a_1 _1246_ (.A1(_0938_),
    .A2(_0217_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q ),
    .X(_0218_));
 sky130_fd_sc_hd__mux4_1 _1247_ (.A0(net62),
    .A1(net70),
    .A2(net779),
    .A3(net12),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_0219_));
 sky130_fd_sc_hd__mux4_1 _1248_ (.A0(net24),
    .A1(net88),
    .A2(net90),
    .A3(net98),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _1249_ (.A0(_0219_),
    .A1(_0220_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ),
    .X(_0221_));
 sky130_fd_sc_hd__a22o_1 _1250_ (.A1(_0216_),
    .A2(_0218_),
    .B1(_0221_),
    .B2(_0939_),
    .X(\Inst_RegFile_switch_matrix.E2BEG6 ));
 sky130_fd_sc_hd__a221o_1 _1251_ (.A1(_0216_),
    .A2(_0218_),
    .B1(_0221_),
    .B2(_0939_),
    .C1(_0937_),
    .X(_0222_));
 sky130_fd_sc_hd__o21a_1 _1252_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ),
    .A2(net129),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q ),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _1253_ (.A0(net73),
    .A1(net101),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ),
    .X(_0224_));
 sky130_fd_sc_hd__a22o_1 _1254_ (.A1(_0222_),
    .A2(_0223_),
    .B1(_0224_),
    .B2(_0940_),
    .X(_0225_));
 sky130_fd_sc_hd__mux4_1 _1255_ (.A0(net76),
    .A1(net18),
    .A2(net104),
    .A3(net132),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q ),
    .X(_0226_));
 sky130_fd_sc_hd__mux4_1 _1256_ (.A0(net64),
    .A1(net92),
    .A2(_0225_),
    .A3(_0226_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q ),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_2 _1257_ (.A0(_0227_),
    .A1(_0214_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ),
    .X(_0228_));
 sky130_fd_sc_hd__inv_2 _1258_ (.A(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__a21oi_1 _1259_ (.A1(_0167_),
    .A2(_0197_),
    .B1(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__mux2_1 _1260_ (.A0(\Inst_RegFile_32x4.mem[0][0] ),
    .A1(\Inst_RegFile_32x4.mem[1][0] ),
    .S(net627),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _1261_ (.A0(\Inst_RegFile_32x4.mem[2][0] ),
    .A1(\Inst_RegFile_32x4.mem[3][0] ),
    .S(net627),
    .X(_0232_));
 sky130_fd_sc_hd__or2_1 _1262_ (.A(net675),
    .B(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__o211a_1 _1263_ (.A1(net661),
    .A2(_0231_),
    .B1(_0233_),
    .C1(_0164_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _1264_ (.A0(\Inst_RegFile_32x4.mem[4][0] ),
    .A1(\Inst_RegFile_32x4.mem[5][0] ),
    .S(net630),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _1265_ (.A0(\Inst_RegFile_32x4.mem[6][0] ),
    .A1(\Inst_RegFile_32x4.mem[7][0] ),
    .S(net630),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _1266_ (.A0(_0235_),
    .A1(_0236_),
    .S(net662),
    .X(_0237_));
 sky130_fd_sc_hd__a211o_1 _1267_ (.A1(net650),
    .A2(_0237_),
    .B1(_0234_),
    .C1(_0193_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _1268_ (.A0(\Inst_RegFile_32x4.mem[10][0] ),
    .A1(\Inst_RegFile_32x4.mem[11][0] ),
    .S(net629),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _1269_ (.A0(\Inst_RegFile_32x4.mem[8][0] ),
    .A1(\Inst_RegFile_32x4.mem[9][0] ),
    .S(net629),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _1270_ (.A0(_0239_),
    .A1(_0240_),
    .S(net675),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_4 _1271_ (.A0(\Inst_RegFile_32x4.mem[12][0] ),
    .A1(\Inst_RegFile_32x4.mem[13][0] ),
    .S(net632),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _1272_ (.A0(\Inst_RegFile_32x4.mem[14][0] ),
    .A1(\Inst_RegFile_32x4.mem[15][0] ),
    .S(net626),
    .X(_0243_));
 sky130_fd_sc_hd__or2_1 _1273_ (.A(net396),
    .B(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__o21a_1 _1274_ (.A1(net663),
    .A2(_0242_),
    .B1(net649),
    .X(_0245_));
 sky130_fd_sc_hd__a221o_1 _1275_ (.A1(net648),
    .A2(_0241_),
    .B1(_0245_),
    .B2(_0244_),
    .C1(net395),
    .X(_0246_));
 sky130_fd_sc_hd__a32o_1 _1276_ (.A1(_0246_),
    .A2(_0238_),
    .A3(_0229_),
    .B1(_0230_),
    .B2(_0205_),
    .X(\Inst_RegFile_32x4.AD_comb[0] ));
 sky130_fd_sc_hd__mux2_4 _1277_ (.A0(\Inst_RegFile_32x4.AD_comb[0] ),
    .A1(\Inst_RegFile_32x4.AD_reg[0] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ),
    .X(AD0));
 sky130_fd_sc_hd__mux2_1 _1278_ (.A0(\Inst_RegFile_32x4.mem[10][1] ),
    .A1(\Inst_RegFile_32x4.mem[11][1] ),
    .S(net629),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _1279_ (.A0(\Inst_RegFile_32x4.mem[8][1] ),
    .A1(\Inst_RegFile_32x4.mem[9][1] ),
    .S(net629),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _1280_ (.A0(_0247_),
    .A1(_0248_),
    .S(net675),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _1281_ (.A0(\Inst_RegFile_32x4.mem[14][1] ),
    .A1(\Inst_RegFile_32x4.mem[15][1] ),
    .S(net626),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _1282_ (.A0(\Inst_RegFile_32x4.mem[12][1] ),
    .A1(\Inst_RegFile_32x4.mem[13][1] ),
    .S(net626),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _1283_ (.A0(_0250_),
    .A1(_0251_),
    .S(net396),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _1284_ (.A0(_0249_),
    .A1(_0252_),
    .S(net649),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _1285_ (.A0(\Inst_RegFile_32x4.mem[0][1] ),
    .A1(\Inst_RegFile_32x4.mem[1][1] ),
    .S(net627),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _1286_ (.A0(\Inst_RegFile_32x4.mem[2][1] ),
    .A1(\Inst_RegFile_32x4.mem[3][1] ),
    .S(net627),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _1287_ (.A0(_0254_),
    .A1(_0255_),
    .S(net661),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _1288_ (.A0(\Inst_RegFile_32x4.mem[4][1] ),
    .A1(\Inst_RegFile_32x4.mem[5][1] ),
    .S(net630),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _1289_ (.A0(\Inst_RegFile_32x4.mem[6][1] ),
    .A1(\Inst_RegFile_32x4.mem[7][1] ),
    .S(net628),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _1290_ (.A0(_0257_),
    .A1(_0258_),
    .S(net661),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _1291_ (.A0(_0256_),
    .A1(_0259_),
    .S(net650),
    .X(_0260_));
 sky130_fd_sc_hd__or2_1 _1292_ (.A(_0193_),
    .B(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__o21a_1 _1293_ (.A1(_0192_),
    .A2(_0253_),
    .B1(_0229_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _1294_ (.A0(\Inst_RegFile_32x4.mem[24][1] ),
    .A1(\Inst_RegFile_32x4.mem[25][1] ),
    .S(net624),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _1295_ (.A0(\Inst_RegFile_32x4.mem[26][1] ),
    .A1(\Inst_RegFile_32x4.mem[27][1] ),
    .S(net625),
    .X(_0264_));
 sky130_fd_sc_hd__or2_1 _1296_ (.A(net396),
    .B(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__o21a_1 _1297_ (.A1(net663),
    .A2(_0263_),
    .B1(net648),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _1298_ (.A0(\Inst_RegFile_32x4.mem[28][1] ),
    .A1(\Inst_RegFile_32x4.mem[29][1] ),
    .S(net624),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _1299_ (.A0(\Inst_RegFile_32x4.mem[30][1] ),
    .A1(\Inst_RegFile_32x4.mem[31][1] ),
    .S(net624),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _1300_ (.A0(_0267_),
    .A1(_0268_),
    .S(net663),
    .X(_0269_));
 sky130_fd_sc_hd__a221o_1 _1301_ (.A1(_0265_),
    .A2(_0266_),
    .B1(net408),
    .B2(_0269_),
    .C1(net395),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _1302_ (.A0(\Inst_RegFile_32x4.mem[16][1] ),
    .A1(\Inst_RegFile_32x4.mem[17][1] ),
    .S(net631),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _1303_ (.A0(\Inst_RegFile_32x4.mem[18][1] ),
    .A1(\Inst_RegFile_32x4.mem[19][1] ),
    .S(net631),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _1304_ (.A0(_0271_),
    .A1(_0272_),
    .S(net662),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _1305_ (.A0(\Inst_RegFile_32x4.mem[22][1] ),
    .A1(\Inst_RegFile_32x4.mem[23][1] ),
    .S(net628),
    .X(_0274_));
 sky130_fd_sc_hd__or2_1 _1306_ (.A(net675),
    .B(_0274_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _1307_ (.A0(\Inst_RegFile_32x4.mem[20][1] ),
    .A1(\Inst_RegFile_32x4.mem[21][1] ),
    .S(net628),
    .X(_0276_));
 sky130_fd_sc_hd__o211a_1 _1308_ (.A1(net661),
    .A2(_0276_),
    .B1(_0275_),
    .C1(net650),
    .X(_0277_));
 sky130_fd_sc_hd__a211o_1 _1309_ (.A1(_0164_),
    .A2(_0273_),
    .B1(_0277_),
    .C1(_0193_),
    .X(_0278_));
 sky130_fd_sc_hd__a32o_1 _1310_ (.A1(_0228_),
    .A2(_0278_),
    .A3(_0270_),
    .B1(_0261_),
    .B2(_0262_),
    .X(\Inst_RegFile_32x4.AD_comb[1] ));
 sky130_fd_sc_hd__mux2_4 _1311_ (.A0(\Inst_RegFile_32x4.AD_comb[1] ),
    .A1(\Inst_RegFile_32x4.AD_reg[1] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ),
    .X(AD1));
 sky130_fd_sc_hd__mux2_1 _1312_ (.A0(\Inst_RegFile_32x4.mem[10][2] ),
    .A1(\Inst_RegFile_32x4.mem[11][2] ),
    .S(net629),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _1313_ (.A0(\Inst_RegFile_32x4.mem[8][2] ),
    .A1(\Inst_RegFile_32x4.mem[9][2] ),
    .S(net629),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _1314_ (.A0(_0279_),
    .A1(_0280_),
    .S(net675),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _1315_ (.A0(\Inst_RegFile_32x4.mem[12][2] ),
    .A1(\Inst_RegFile_32x4.mem[13][2] ),
    .S(net626),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _1316_ (.A0(\Inst_RegFile_32x4.mem[14][2] ),
    .A1(\Inst_RegFile_32x4.mem[15][2] ),
    .S(net626),
    .X(_0283_));
 sky130_fd_sc_hd__or2_1 _1317_ (.A(net396),
    .B(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__o21a_1 _1318_ (.A1(net663),
    .A2(_0282_),
    .B1(net408),
    .X(_0285_));
 sky130_fd_sc_hd__a221o_1 _1319_ (.A1(net648),
    .A2(_0281_),
    .B1(_0284_),
    .B2(_0285_),
    .C1(_0192_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _1320_ (.A0(\Inst_RegFile_32x4.mem[0][2] ),
    .A1(\Inst_RegFile_32x4.mem[1][2] ),
    .S(net627),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _1321_ (.A0(\Inst_RegFile_32x4.mem[2][2] ),
    .A1(\Inst_RegFile_32x4.mem[3][2] ),
    .S(net627),
    .X(_0288_));
 sky130_fd_sc_hd__or2_1 _1322_ (.A(net675),
    .B(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__o211a_1 _1323_ (.A1(net661),
    .A2(_0287_),
    .B1(_0289_),
    .C1(net648),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _1324_ (.A0(\Inst_RegFile_32x4.mem[4][2] ),
    .A1(\Inst_RegFile_32x4.mem[5][2] ),
    .S(net630),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _1325_ (.A0(\Inst_RegFile_32x4.mem[6][2] ),
    .A1(\Inst_RegFile_32x4.mem[7][2] ),
    .S(net630),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _1326_ (.A0(_0291_),
    .A1(_0292_),
    .S(net661),
    .X(_0293_));
 sky130_fd_sc_hd__a211o_1 _1327_ (.A1(net408),
    .A2(_0293_),
    .B1(_0290_),
    .C1(_0193_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _1328_ (.A0(\Inst_RegFile_32x4.mem[26][2] ),
    .A1(\Inst_RegFile_32x4.mem[27][2] ),
    .S(net625),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _1329_ (.A0(\Inst_RegFile_32x4.mem[24][2] ),
    .A1(\Inst_RegFile_32x4.mem[25][2] ),
    .S(net625),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _1330_ (.A0(_0295_),
    .A1(_0296_),
    .S(net674),
    .X(_0297_));
 sky130_fd_sc_hd__nand2_1 _1331_ (.A(net648),
    .B(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__mux2_1 _1332_ (.A0(\Inst_RegFile_32x4.mem[28][2] ),
    .A1(\Inst_RegFile_32x4.mem[29][2] ),
    .S(net624),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _1333_ (.A0(\Inst_RegFile_32x4.mem[30][2] ),
    .A1(\Inst_RegFile_32x4.mem[31][2] ),
    .S(net624),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _1334_ (.A0(_0299_),
    .A1(_0300_),
    .S(net663),
    .X(_0301_));
 sky130_fd_sc_hd__a21oi_2 _1335_ (.A1(net408),
    .A2(_0301_),
    .B1(net395),
    .Y(_0302_));
 sky130_fd_sc_hd__mux2_1 _1336_ (.A0(\Inst_RegFile_32x4.mem[16][2] ),
    .A1(\Inst_RegFile_32x4.mem[17][2] ),
    .S(net630),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _1337_ (.A0(\Inst_RegFile_32x4.mem[18][2] ),
    .A1(\Inst_RegFile_32x4.mem[19][2] ),
    .S(net630),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _1338_ (.A0(_0303_),
    .A1(_0304_),
    .S(net662),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _1339_ (.A0(\Inst_RegFile_32x4.mem[22][2] ),
    .A1(\Inst_RegFile_32x4.mem[23][2] ),
    .S(net628),
    .X(_0306_));
 sky130_fd_sc_hd__or2_1 _1340_ (.A(net674),
    .B(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _1341_ (.A0(\Inst_RegFile_32x4.mem[20][2] ),
    .A1(\Inst_RegFile_32x4.mem[21][2] ),
    .S(net628),
    .X(_0308_));
 sky130_fd_sc_hd__o211a_1 _1342_ (.A1(net661),
    .A2(_0308_),
    .B1(_0307_),
    .C1(net650),
    .X(_0309_));
 sky130_fd_sc_hd__a211o_1 _1343_ (.A1(net648),
    .A2(_0305_),
    .B1(_0309_),
    .C1(_0193_),
    .X(_0310_));
 sky130_fd_sc_hd__a21oi_1 _1344_ (.A1(_0302_),
    .A2(_0298_),
    .B1(_0229_),
    .Y(_0311_));
 sky130_fd_sc_hd__a32o_1 _1345_ (.A1(_0229_),
    .A2(_0286_),
    .A3(_0294_),
    .B1(_0310_),
    .B2(_0311_),
    .X(\Inst_RegFile_32x4.AD_comb[2] ));
 sky130_fd_sc_hd__mux2_4 _1346_ (.A0(\Inst_RegFile_32x4.AD_comb[2] ),
    .A1(\Inst_RegFile_32x4.AD_reg[2] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ),
    .X(AD2));
 sky130_fd_sc_hd__mux2_1 _1347_ (.A0(\Inst_RegFile_32x4.mem[10][3] ),
    .A1(\Inst_RegFile_32x4.mem[11][3] ),
    .S(net626),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _1348_ (.A0(\Inst_RegFile_32x4.mem[8][3] ),
    .A1(\Inst_RegFile_32x4.mem[9][3] ),
    .S(net629),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _1349_ (.A0(_0312_),
    .A1(_0313_),
    .S(net674),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _1350_ (.A0(\Inst_RegFile_32x4.mem[12][3] ),
    .A1(\Inst_RegFile_32x4.mem[13][3] ),
    .S(net626),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _1351_ (.A0(\Inst_RegFile_32x4.mem[14][3] ),
    .A1(\Inst_RegFile_32x4.mem[15][3] ),
    .S(net626),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _1352_ (.A0(_0315_),
    .A1(_0316_),
    .S(net663),
    .X(_0317_));
 sky130_fd_sc_hd__a21o_1 _1353_ (.A1(net649),
    .A2(_0317_),
    .B1(_0192_),
    .X(_0318_));
 sky130_fd_sc_hd__a21oi_1 _1354_ (.A1(net648),
    .A2(_0314_),
    .B1(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__mux2_1 _1355_ (.A0(\Inst_RegFile_32x4.mem[0][3] ),
    .A1(\Inst_RegFile_32x4.mem[1][3] ),
    .S(net627),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _1356_ (.A0(\Inst_RegFile_32x4.mem[2][3] ),
    .A1(\Inst_RegFile_32x4.mem[3][3] ),
    .S(net627),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _1357_ (.A0(_0320_),
    .A1(_0321_),
    .S(net661),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _1358_ (.A0(\Inst_RegFile_32x4.mem[4][3] ),
    .A1(\Inst_RegFile_32x4.mem[5][3] ),
    .S(net630),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _1359_ (.A0(\Inst_RegFile_32x4.mem[6][3] ),
    .A1(\Inst_RegFile_32x4.mem[7][3] ),
    .S(net630),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _1360_ (.A0(_0323_),
    .A1(_0324_),
    .S(net661),
    .X(_0325_));
 sky130_fd_sc_hd__a21bo_1 _1361_ (.A1(net649),
    .A2(_0325_),
    .B1_N(_0192_),
    .X(_0326_));
 sky130_fd_sc_hd__a21oi_1 _1362_ (.A1(net648),
    .A2(_0322_),
    .B1(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__mux2_1 _1363_ (.A0(\Inst_RegFile_32x4.mem[26][3] ),
    .A1(\Inst_RegFile_32x4.mem[27][3] ),
    .S(net625),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _1364_ (.A0(\Inst_RegFile_32x4.mem[24][3] ),
    .A1(\Inst_RegFile_32x4.mem[25][3] ),
    .S(net625),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_4 _1365_ (.A0(_0328_),
    .A1(_0329_),
    .S(net674),
    .X(_0330_));
 sky130_fd_sc_hd__nand2_4 _1366_ (.A(net648),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__mux2_1 _1367_ (.A0(\Inst_RegFile_32x4.mem[28][3] ),
    .A1(\Inst_RegFile_32x4.mem[29][3] ),
    .S(net624),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _1368_ (.A0(\Inst_RegFile_32x4.mem[30][3] ),
    .A1(\Inst_RegFile_32x4.mem[31][3] ),
    .S(net624),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _1369_ (.A0(_0332_),
    .A1(_0333_),
    .S(net663),
    .X(_0334_));
 sky130_fd_sc_hd__nand2_1 _1370_ (.A(net649),
    .B(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__mux2_1 _1371_ (.A0(\Inst_RegFile_32x4.mem[18][3] ),
    .A1(\Inst_RegFile_32x4.mem[19][3] ),
    .S(net630),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _1372_ (.A0(\Inst_RegFile_32x4.mem[16][3] ),
    .A1(\Inst_RegFile_32x4.mem[17][3] ),
    .S(net631),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _1373_ (.A0(_0336_),
    .A1(_0337_),
    .S(net675),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _1374_ (.A0(\Inst_RegFile_32x4.mem[22][3] ),
    .A1(\Inst_RegFile_32x4.mem[23][3] ),
    .S(net628),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _1375_ (.A0(\Inst_RegFile_32x4.mem[20][3] ),
    .A1(\Inst_RegFile_32x4.mem[21][3] ),
    .S(net628),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _1376_ (.A0(_0339_),
    .A1(_0340_),
    .S(net674),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _1377_ (.A0(_0338_),
    .A1(_0341_),
    .S(net650),
    .X(_0342_));
 sky130_fd_sc_hd__nor2_1 _1378_ (.A(_0193_),
    .B(_0342_),
    .Y(_0343_));
 sky130_fd_sc_hd__a31o_1 _1379_ (.A1(_0331_),
    .A2(_0193_),
    .A3(_0335_),
    .B1(_0229_),
    .X(_0344_));
 sky130_fd_sc_hd__o32a_4 _1380_ (.A1(_0228_),
    .A2(_0319_),
    .A3(_0327_),
    .B1(_0344_),
    .B2(_0343_),
    .X(_0345_));
 sky130_fd_sc_hd__inv_1 _1381_ (.A(_0345_),
    .Y(\Inst_RegFile_32x4.AD_comb[3] ));
 sky130_fd_sc_hd__nand2_1 _1382_ (.A(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ),
    .B(\Inst_RegFile_32x4.AD_reg[3] ),
    .Y(_0346_));
 sky130_fd_sc_hd__o21ai_4 _1383_ (.A1(_0345_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ),
    .B1(_0346_),
    .Y(AD3));
 sky130_fd_sc_hd__a221o_1 _1384_ (.A1(_0222_),
    .A2(_0223_),
    .B1(_0224_),
    .B2(_0940_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ),
    .X(_0347_));
 sky130_fd_sc_hd__mux4_2 _1385_ (.A0(net74),
    .A1(net16),
    .A2(net102),
    .A3(net130),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q ),
    .X(_0348_));
 sky130_fd_sc_hd__o21ba_1 _1386_ (.A1(_0941_),
    .A2(_0348_),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q ),
    .X(_0349_));
 sky130_fd_sc_hd__mux4_1 _1387_ (.A0(net116),
    .A1(net673),
    .A2(net660),
    .A3(net654),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0350_));
 sky130_fd_sc_hd__or2_1 _1388_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ),
    .B(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__mux4_2 _1389_ (.A0(net421),
    .A1(net637),
    .A2(net667),
    .A3(net641),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0352_));
 sky130_fd_sc_hd__o21a_1 _1390_ (.A1(_0943_),
    .A2(_0352_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_0353_));
 sky130_fd_sc_hd__mux4_2 _1391_ (.A0(net26),
    .A1(net88),
    .A2(net90),
    .A3(net96),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0354_));
 sky130_fd_sc_hd__mux4_2 _1392_ (.A0(net60),
    .A1(net68),
    .A2(net2),
    .A3(net10),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_4 _1393_ (.A0(_0354_),
    .A1(_0355_),
    .S(_0943_),
    .X(_0356_));
 sky130_fd_sc_hd__a22o_1 _1394_ (.A1(_0351_),
    .A2(_0353_),
    .B1(_0356_),
    .B2(_0944_),
    .X(\Inst_RegFile_switch_matrix.E2BEG4 ));
 sky130_fd_sc_hd__a221o_1 _1395_ (.A1(_0351_),
    .A2(_0353_),
    .B1(_0356_),
    .B2(_0944_),
    .C1(_0942_),
    .X(_0357_));
 sky130_fd_sc_hd__o21a_1 _1396_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(net121),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _1397_ (.A0(net81),
    .A1(net113),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_0359_));
 sky130_fd_sc_hd__a221o_1 _1398_ (.A1(_0358_),
    .A2(_0357_),
    .B1(_0359_),
    .B2(_0945_),
    .C1(_0941_),
    .X(_0360_));
 sky130_fd_sc_hd__mux4_2 _1399_ (.A0(net66),
    .A1(net8),
    .A2(net111),
    .A3(net122),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q ),
    .X(_0361_));
 sky130_fd_sc_hd__or2_1 _1400_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ),
    .B(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__a32o_2 _1401_ (.A1(_0360_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q ),
    .A3(_0362_),
    .B1(_0347_),
    .B2(_0349_),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _1402_ (.A0(\Inst_RegFile_32x4.mem[0][0] ),
    .A1(\Inst_RegFile_32x4.mem[1][0] ),
    .S(net606),
    .X(_0364_));
 sky130_fd_sc_hd__mux4_1 _1403_ (.A0(net688),
    .A1(net672),
    .A2(net659),
    .A3(net653),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_0365_));
 sky130_fd_sc_hd__or2_1 _1404_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ),
    .B(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__mux4_2 _1405_ (.A0(net646),
    .A1(net679),
    .A2(net668),
    .A3(net640),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_0367_));
 sky130_fd_sc_hd__o21a_1 _1406_ (.A1(_0948_),
    .A2(_0367_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q ),
    .X(_0368_));
 sky130_fd_sc_hd__mux4_1 _1407_ (.A0(net62),
    .A1(net70),
    .A2(net4),
    .A3(net12),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_0369_));
 sky130_fd_sc_hd__mux4_1 _1408_ (.A0(net90),
    .A1(net98),
    .A2(net112),
    .A3(net116),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _1409_ (.A0(_0369_),
    .A1(_0370_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_0371_));
 sky130_fd_sc_hd__a22o_4 _1410_ (.A1(_0366_),
    .A2(_0368_),
    .B1(_0371_),
    .B2(_0949_),
    .X(\Inst_RegFile_switch_matrix.JS2BEG6 ));
 sky130_fd_sc_hd__mux4_2 _1411_ (.A0(net17),
    .A1(net103),
    .A2(net131),
    .A3(\Inst_RegFile_switch_matrix.JS2BEG6 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q ),
    .X(_0372_));
 sky130_fd_sc_hd__a21o_1 _1412_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q ),
    .A2(_0226_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ),
    .X(_0373_));
 sky130_fd_sc_hd__a21oi_1 _1413_ (.A1(_0946_),
    .A2(_0372_),
    .B1(_0373_),
    .Y(_0374_));
 sky130_fd_sc_hd__mux4_1 _1414_ (.A0(net118),
    .A1(net673),
    .A2(net660),
    .A3(net654),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0375_));
 sky130_fd_sc_hd__or2_1 _1415_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ),
    .B(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__mux4_2 _1416_ (.A0(net647),
    .A1(net637),
    .A2(net667),
    .A3(net641),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ),
    .X(_0377_));
 sky130_fd_sc_hd__o21a_1 _1417_ (.A1(_0377_),
    .A2(_0951_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q ),
    .X(_0378_));
 sky130_fd_sc_hd__mux4_1 _1418_ (.A0(net88),
    .A1(net96),
    .A2(net114),
    .A3(net116),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0379_));
 sky130_fd_sc_hd__mux4_1 _1419_ (.A0(net60),
    .A1(net68),
    .A2(net2),
    .A3(net10),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _1420_ (.A0(_0379_),
    .A1(_0380_),
    .S(_0951_),
    .X(_0381_));
 sky130_fd_sc_hd__a22o_4 _1421_ (.A1(_0378_),
    .A2(_0376_),
    .B1(_0381_),
    .B2(_0952_),
    .X(\Inst_RegFile_switch_matrix.JS2BEG4 ));
 sky130_fd_sc_hd__mux2_1 _1422_ (.A0(net140),
    .A1(\Inst_RegFile_switch_matrix.JS2BEG4 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q ),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _1423_ (.A0(net22),
    .A1(net108),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q ),
    .X(_0383_));
 sky130_fd_sc_hd__o21a_1 _1424_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0383_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q ),
    .X(_0384_));
 sky130_fd_sc_hd__o21ai_1 _1425_ (.A1(_0953_),
    .A2(_0382_),
    .B1(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__mux4_2 _1426_ (.A0(net84),
    .A1(net10),
    .A2(net96),
    .A3(net124),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q ),
    .X(_0386_));
 sky130_fd_sc_hd__nand2_1 _1427_ (.A(_0946_),
    .B(_0386_),
    .Y(_0387_));
 sky130_fd_sc_hd__a31oi_1 _1428_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ),
    .A2(_0385_),
    .A3(_0387_),
    .B1(_0374_),
    .Y(_0388_));
 sky130_fd_sc_hd__a31o_1 _1429_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ),
    .A2(_0385_),
    .A3(_0387_),
    .B1(_0374_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _1430_ (.A0(\Inst_RegFile_32x4.mem[2][0] ),
    .A1(\Inst_RegFile_32x4.mem[3][0] ),
    .S(net606),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _1431_ (.A0(_0364_),
    .A1(_0390_),
    .S(net682),
    .X(_0391_));
 sky130_fd_sc_hd__and2_1 _1432_ (.A(_0389_),
    .B(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__mux4_1 _1433_ (.A0(AD3),
    .A1(net634),
    .A2(net665),
    .A3(net638),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0393_));
 sky130_fd_sc_hd__or2_4 _1434_ (.A(_0955_),
    .B(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__mux4_1 _1435_ (.A0(net140),
    .A1(net670),
    .A2(net657),
    .A3(net655),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0395_));
 sky130_fd_sc_hd__o21a_1 _1436_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ),
    .A2(_0395_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0396_));
 sky130_fd_sc_hd__mux4_1 _1437_ (.A0(net60),
    .A1(net68),
    .A2(net2),
    .A3(net10),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0397_));
 sky130_fd_sc_hd__mux4_1 _1438_ (.A0(net88),
    .A1(net96),
    .A2(net90),
    .A3(net116),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _1439_ (.A0(_0397_),
    .A1(_0398_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ),
    .X(_0399_));
 sky130_fd_sc_hd__a22o_4 _1440_ (.A1(_0396_),
    .A2(_0394_),
    .B1(_0399_),
    .B2(_0956_),
    .X(\Inst_RegFile_switch_matrix.JW2BEG4 ));
 sky130_fd_sc_hd__mux4_2 _1441_ (.A0(net83),
    .A1(net778),
    .A2(net119),
    .A3(\Inst_RegFile_switch_matrix.JW2BEG4 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q ),
    .X(_0400_));
 sky130_fd_sc_hd__mux4_2 _1442_ (.A0(net64),
    .A1(net92),
    .A2(net26),
    .A3(net120),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q ),
    .X(_0401_));
 sky130_fd_sc_hd__mux4_1 _1443_ (.A0(net138),
    .A1(net670),
    .A2(net657),
    .A3(net651),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_0402_));
 sky130_fd_sc_hd__nand2b_1 _1444_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ),
    .B(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__mux4_2 _1445_ (.A0(net645),
    .A1(net678),
    .A2(net665),
    .A3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_0404_));
 sky130_fd_sc_hd__a21boi_2 _1446_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ),
    .A2(_0404_),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q ),
    .Y(_0405_));
 sky130_fd_sc_hd__mux4_1 _1447_ (.A0(net62),
    .A1(net70),
    .A2(net779),
    .A3(net12),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_0406_));
 sky130_fd_sc_hd__and2b_1 _1448_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ),
    .B(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__mux4_1 _1449_ (.A0(net88),
    .A1(net98),
    .A2(net90),
    .A3(net688),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_0408_));
 sky130_fd_sc_hd__a21o_1 _1450_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ),
    .A2(_0408_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q ),
    .X(_0409_));
 sky130_fd_sc_hd__o2bb2a_4 _1451_ (.A1_N(_0403_),
    .A2_N(_0405_),
    .B1(_0407_),
    .B2(_0409_),
    .X(\Inst_RegFile_switch_matrix.JW2BEG6 ));
 sky130_fd_sc_hd__mux4_2 _1452_ (.A0(net71),
    .A1(net13),
    .A2(net127),
    .A3(\Inst_RegFile_switch_matrix.JW2BEG6 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q ),
    .X(_0410_));
 sky130_fd_sc_hd__mux4_1 _1453_ (.A0(net72),
    .A1(net14),
    .A2(net100),
    .A3(net128),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q ),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_2 _1454_ (.A0(_0400_),
    .A1(_0401_),
    .S(_0954_),
    .X(_0412_));
 sky130_fd_sc_hd__o21ba_1 _1455_ (.A1(_0954_),
    .A2(_0411_),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q ),
    .X(_0413_));
 sky130_fd_sc_hd__o21a_1 _1456_ (.A1(_0410_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ),
    .B1(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__a21oi_2 _1457_ (.A1(_0412_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q ),
    .B1(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__inv_2 _1458_ (.A(net619),
    .Y(_0416_));
 sky130_fd_sc_hd__mux2_1 _1459_ (.A0(\Inst_RegFile_32x4.mem[6][0] ),
    .A1(\Inst_RegFile_32x4.mem[7][0] ),
    .S(net609),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _1460_ (.A0(\Inst_RegFile_32x4.mem[4][0] ),
    .A1(\Inst_RegFile_32x4.mem[5][0] ),
    .S(net609),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _1461_ (.A0(_0418_),
    .A1(_0417_),
    .S(net683),
    .X(_0419_));
 sky130_fd_sc_hd__a211o_1 _1462_ (.A1(net643),
    .A2(_0419_),
    .B1(_0416_),
    .C1(_0392_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _1463_ (.A0(\Inst_RegFile_32x4.mem[8][0] ),
    .A1(\Inst_RegFile_32x4.mem[9][0] ),
    .S(net608),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _1464_ (.A0(\Inst_RegFile_32x4.mem[10][0] ),
    .A1(\Inst_RegFile_32x4.mem[11][0] ),
    .S(net608),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _1465_ (.A0(_0421_),
    .A1(_0422_),
    .S(net413),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _1466_ (.A0(\Inst_RegFile_32x4.mem[12][0] ),
    .A1(\Inst_RegFile_32x4.mem[13][0] ),
    .S(net410),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _1467_ (.A0(\Inst_RegFile_32x4.mem[14][0] ),
    .A1(\Inst_RegFile_32x4.mem[15][0] ),
    .S(net410),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _1468_ (.A0(_0424_),
    .A1(_0425_),
    .S(net413),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _1469_ (.A0(_0423_),
    .A1(_0426_),
    .S(net642),
    .X(_0427_));
 sky130_fd_sc_hd__mux4_2 _1470_ (.A0(net398),
    .A1(net678),
    .A2(net665),
    .A3(net638),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0428_));
 sky130_fd_sc_hd__or2_4 _1471_ (.A(_0933_),
    .B(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__mux4_1 _1472_ (.A0(net688),
    .A1(net670),
    .A2(net657),
    .A3(net655),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0430_));
 sky130_fd_sc_hd__o21a_1 _1473_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ),
    .A2(_0430_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q ),
    .X(_0431_));
 sky130_fd_sc_hd__mux4_1 _1474_ (.A0(net62),
    .A1(net70),
    .A2(net84),
    .A3(net779),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0432_));
 sky130_fd_sc_hd__mux4_1 _1475_ (.A0(net12),
    .A1(net90),
    .A2(net98),
    .A3(net116),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _1476_ (.A0(_0432_),
    .A1(_0433_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ),
    .X(_0434_));
 sky130_fd_sc_hd__a22o_4 _1477_ (.A1(_0431_),
    .A2(_0429_),
    .B1(_0434_),
    .B2(_0934_),
    .X(\Inst_RegFile_switch_matrix.JN2BEG6 ));
 sky130_fd_sc_hd__mux4_2 _1478_ (.A0(_0179_),
    .A1(\Inst_RegFile_switch_matrix.JS2BEG6 ),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG6 ),
    .A3(\Inst_RegFile_switch_matrix.JW2BEG6 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ),
    .X(_0435_));
 sky130_fd_sc_hd__mux4_2 _1479_ (.A0(net15),
    .A1(net129),
    .A2(net101),
    .A3(\Inst_RegFile_switch_matrix.E2BEG3 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q ),
    .X(_0436_));
 sky130_fd_sc_hd__mux4_2 _1480_ (.A0(net76),
    .A1(net18),
    .A2(net104),
    .A3(net132),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q ),
    .X(_0437_));
 sky130_fd_sc_hd__mux4_2 _1481_ (.A0(net65),
    .A1(net93),
    .A2(_0436_),
    .A3(_0437_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q ),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_4 _1482_ (.A0(_0438_),
    .A1(_0435_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q ),
    .X(_0439_));
 sky130_fd_sc_hd__o21ba_1 _1483_ (.A1(net619),
    .A2(_0427_),
    .B1_N(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _1484_ (.A0(\Inst_RegFile_32x4.mem[16][0] ),
    .A1(\Inst_RegFile_32x4.mem[17][0] ),
    .S(net610),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _1485_ (.A0(\Inst_RegFile_32x4.mem[18][0] ),
    .A1(\Inst_RegFile_32x4.mem[19][0] ),
    .S(net610),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _1486_ (.A0(_0441_),
    .A1(_0442_),
    .S(net683),
    .X(_0443_));
 sky130_fd_sc_hd__nand2_1 _1487_ (.A(\Inst_RegFile_32x4.mem[23][0] ),
    .B(net606),
    .Y(_0444_));
 sky130_fd_sc_hd__o211ai_1 _1488_ (.A1(_0959_),
    .A2(net606),
    .B1(net682),
    .C1(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__mux2_1 _1489_ (.A0(\Inst_RegFile_32x4.mem[20][0] ),
    .A1(\Inst_RegFile_32x4.mem[21][0] ),
    .S(net606),
    .X(_0446_));
 sky130_fd_sc_hd__o211a_1 _1490_ (.A1(net682),
    .A2(_0446_),
    .B1(_0445_),
    .C1(net643),
    .X(_0447_));
 sky130_fd_sc_hd__a211o_1 _1491_ (.A1(_0389_),
    .A2(_0443_),
    .B1(_0447_),
    .C1(_0416_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _1492_ (.A0(\Inst_RegFile_32x4.mem[24][0] ),
    .A1(\Inst_RegFile_32x4.mem[25][0] ),
    .S(net603),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _1493_ (.A0(\Inst_RegFile_32x4.mem[26][0] ),
    .A1(\Inst_RegFile_32x4.mem[27][0] ),
    .S(net604),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _1494_ (.A0(_0449_),
    .A1(_0450_),
    .S(net412),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _1495_ (.A0(\Inst_RegFile_32x4.mem[30][0] ),
    .A1(\Inst_RegFile_32x4.mem[31][0] ),
    .S(net604),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _1496_ (.A0(\Inst_RegFile_32x4.mem[28][0] ),
    .A1(\Inst_RegFile_32x4.mem[29][0] ),
    .S(net603),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _1497_ (.A0(_0453_),
    .A1(_0452_),
    .S(net412),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _1498_ (.A0(_0451_),
    .A1(_0454_),
    .S(net642),
    .X(_0455_));
 sky130_fd_sc_hd__o21a_1 _1499_ (.A1(_0455_),
    .A2(_0415_),
    .B1(_0439_),
    .X(_0456_));
 sky130_fd_sc_hd__a22o_1 _1500_ (.A1(_0420_),
    .A2(_0440_),
    .B1(_0456_),
    .B2(_0448_),
    .X(\Inst_RegFile_32x4.BD_comb[0] ));
 sky130_fd_sc_hd__mux2_4 _1501_ (.A0(\Inst_RegFile_32x4.BD_comb[0] ),
    .A1(\Inst_RegFile_32x4.BD_reg[0] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .X(BD0));
 sky130_fd_sc_hd__mux2_1 _1502_ (.A0(\Inst_RegFile_32x4.mem[16][1] ),
    .A1(\Inst_RegFile_32x4.mem[17][1] ),
    .S(net610),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _1503_ (.A0(\Inst_RegFile_32x4.mem[18][1] ),
    .A1(\Inst_RegFile_32x4.mem[19][1] ),
    .S(net609),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _1504_ (.A0(_0457_),
    .A1(_0458_),
    .S(net683),
    .X(_0459_));
 sky130_fd_sc_hd__and2_1 _1505_ (.A(_0389_),
    .B(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _1506_ (.A0(\Inst_RegFile_32x4.mem[22][1] ),
    .A1(\Inst_RegFile_32x4.mem[23][1] ),
    .S(net606),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _1507_ (.A0(\Inst_RegFile_32x4.mem[20][1] ),
    .A1(\Inst_RegFile_32x4.mem[21][1] ),
    .S(net607),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _1508_ (.A0(_0462_),
    .A1(_0461_),
    .S(net682),
    .X(_0463_));
 sky130_fd_sc_hd__a211o_1 _1509_ (.A1(net643),
    .A2(_0463_),
    .B1(_0460_),
    .C1(_0416_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _1510_ (.A0(\Inst_RegFile_32x4.mem[24][1] ),
    .A1(\Inst_RegFile_32x4.mem[25][1] ),
    .S(net603),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _1511_ (.A0(\Inst_RegFile_32x4.mem[26][1] ),
    .A1(\Inst_RegFile_32x4.mem[27][1] ),
    .S(net604),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _1512_ (.A0(_0465_),
    .A1(_0466_),
    .S(net412),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _1513_ (.A0(\Inst_RegFile_32x4.mem[28][1] ),
    .A1(\Inst_RegFile_32x4.mem[29][1] ),
    .S(net603),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _1514_ (.A0(\Inst_RegFile_32x4.mem[30][1] ),
    .A1(\Inst_RegFile_32x4.mem[31][1] ),
    .S(net603),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _1515_ (.A0(_0468_),
    .A1(_0469_),
    .S(net412),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_4 _1516_ (.A0(_0467_),
    .A1(_0470_),
    .S(net642),
    .X(_0471_));
 sky130_fd_sc_hd__or2_1 _1517_ (.A(net619),
    .B(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _1518_ (.A0(\Inst_RegFile_32x4.mem[2][1] ),
    .A1(\Inst_RegFile_32x4.mem[3][1] ),
    .S(net606),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _1519_ (.A0(\Inst_RegFile_32x4.mem[0][1] ),
    .A1(\Inst_RegFile_32x4.mem[1][1] ),
    .S(net606),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _1520_ (.A0(_0474_),
    .A1(_0473_),
    .S(net682),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _1521_ (.A0(\Inst_RegFile_32x4.mem[6][1] ),
    .A1(\Inst_RegFile_32x4.mem[7][1] ),
    .S(net607),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _1522_ (.A0(\Inst_RegFile_32x4.mem[4][1] ),
    .A1(\Inst_RegFile_32x4.mem[5][1] ),
    .S(net609),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _1523_ (.A0(_0477_),
    .A1(_0476_),
    .S(net682),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _1524_ (.A0(_0475_),
    .A1(_0478_),
    .S(net643),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _1525_ (.A0(\Inst_RegFile_32x4.mem[8][1] ),
    .A1(\Inst_RegFile_32x4.mem[9][1] ),
    .S(net608),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _1526_ (.A0(\Inst_RegFile_32x4.mem[10][1] ),
    .A1(\Inst_RegFile_32x4.mem[11][1] ),
    .S(net608),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _1527_ (.A0(_0480_),
    .A1(_0481_),
    .S(net413),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _1528_ (.A0(\Inst_RegFile_32x4.mem[14][1] ),
    .A1(\Inst_RegFile_32x4.mem[15][1] ),
    .S(net410),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _1529_ (.A0(\Inst_RegFile_32x4.mem[12][1] ),
    .A1(\Inst_RegFile_32x4.mem[13][1] ),
    .S(net410),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _1530_ (.A0(_0484_),
    .A1(_0483_),
    .S(net412),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _1531_ (.A0(_0482_),
    .A1(_0485_),
    .S(net642),
    .X(_0486_));
 sky130_fd_sc_hd__or2_1 _1532_ (.A(net619),
    .B(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__o21ba_1 _1533_ (.A1(_0416_),
    .A2(_0479_),
    .B1_N(_0439_),
    .X(_0488_));
 sky130_fd_sc_hd__a32o_1 _1534_ (.A1(_0464_),
    .A2(_0439_),
    .A3(_0472_),
    .B1(_0487_),
    .B2(_0488_),
    .X(\Inst_RegFile_32x4.BD_comb[1] ));
 sky130_fd_sc_hd__mux2_4 _1535_ (.A0(\Inst_RegFile_32x4.BD_comb[1] ),
    .A1(\Inst_RegFile_32x4.BD_reg[1] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .X(BD1));
 sky130_fd_sc_hd__mux2_1 _1536_ (.A0(\Inst_RegFile_32x4.mem[16][3] ),
    .A1(\Inst_RegFile_32x4.mem[17][3] ),
    .S(net609),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _1537_ (.A0(\Inst_RegFile_32x4.mem[18][3] ),
    .A1(\Inst_RegFile_32x4.mem[19][3] ),
    .S(net609),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _1538_ (.A0(_0489_),
    .A1(_0490_),
    .S(net683),
    .X(_0491_));
 sky130_fd_sc_hd__and2_1 _1539_ (.A(_0389_),
    .B(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _1540_ (.A0(\Inst_RegFile_32x4.mem[22][3] ),
    .A1(\Inst_RegFile_32x4.mem[23][3] ),
    .S(net607),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _1541_ (.A0(\Inst_RegFile_32x4.mem[20][3] ),
    .A1(\Inst_RegFile_32x4.mem[21][3] ),
    .S(net607),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _1542_ (.A0(_0494_),
    .A1(_0493_),
    .S(net682),
    .X(_0495_));
 sky130_fd_sc_hd__a211o_1 _1543_ (.A1(net643),
    .A2(_0495_),
    .B1(_0492_),
    .C1(_0416_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _1544_ (.A0(\Inst_RegFile_32x4.mem[24][3] ),
    .A1(\Inst_RegFile_32x4.mem[25][3] ),
    .S(net604),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _1545_ (.A0(\Inst_RegFile_32x4.mem[26][3] ),
    .A1(\Inst_RegFile_32x4.mem[27][3] ),
    .S(net604),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _1546_ (.A0(_0497_),
    .A1(_0498_),
    .S(net681),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _1547_ (.A0(\Inst_RegFile_32x4.mem[28][3] ),
    .A1(\Inst_RegFile_32x4.mem[29][3] ),
    .S(net603),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _1548_ (.A0(\Inst_RegFile_32x4.mem[30][3] ),
    .A1(\Inst_RegFile_32x4.mem[31][3] ),
    .S(net603),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _1549_ (.A0(_0500_),
    .A1(_0501_),
    .S(net681),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _1550_ (.A0(_0499_),
    .A1(_0502_),
    .S(net642),
    .X(_0503_));
 sky130_fd_sc_hd__or2_1 _1551_ (.A(net619),
    .B(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _1552_ (.A0(\Inst_RegFile_32x4.mem[2][3] ),
    .A1(\Inst_RegFile_32x4.mem[3][3] ),
    .S(net607),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _1553_ (.A0(\Inst_RegFile_32x4.mem[0][3] ),
    .A1(\Inst_RegFile_32x4.mem[1][3] ),
    .S(net607),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _1554_ (.A0(_0506_),
    .A1(_0505_),
    .S(net682),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _1555_ (.A0(\Inst_RegFile_32x4.mem[6][3] ),
    .A1(\Inst_RegFile_32x4.mem[7][3] ),
    .S(net609),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _1556_ (.A0(\Inst_RegFile_32x4.mem[4][3] ),
    .A1(\Inst_RegFile_32x4.mem[5][3] ),
    .S(net609),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _1557_ (.A0(_0509_),
    .A1(_0508_),
    .S(net683),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _1558_ (.A0(_0507_),
    .A1(_0510_),
    .S(net642),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_4 _1559_ (.A0(\Inst_RegFile_32x4.mem[8][3] ),
    .A1(\Inst_RegFile_32x4.mem[9][3] ),
    .S(net608),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_2 _1560_ (.A0(\Inst_RegFile_32x4.mem[10][3] ),
    .A1(\Inst_RegFile_32x4.mem[11][3] ),
    .S(net410),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_4 _1561_ (.A0(_0512_),
    .A1(_0513_),
    .S(net681),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_2 _1562_ (.A0(\Inst_RegFile_32x4.mem[14][3] ),
    .A1(\Inst_RegFile_32x4.mem[15][3] ),
    .S(net605),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_2 _1563_ (.A0(\Inst_RegFile_32x4.mem[12][3] ),
    .A1(\Inst_RegFile_32x4.mem[13][3] ),
    .S(net605),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_4 _1564_ (.A0(_0516_),
    .A1(_0515_),
    .S(net684),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_4 _1565_ (.A0(_0514_),
    .A1(_0517_),
    .S(net642),
    .X(_0518_));
 sky130_fd_sc_hd__or2_4 _1566_ (.A(net619),
    .B(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__o21ba_1 _1567_ (.A1(_0416_),
    .A2(_0511_),
    .B1_N(_0439_),
    .X(_0520_));
 sky130_fd_sc_hd__a32o_1 _1568_ (.A1(_0439_),
    .A2(_0496_),
    .A3(_0504_),
    .B1(_0520_),
    .B2(_0519_),
    .X(\Inst_RegFile_32x4.BD_comb[3] ));
 sky130_fd_sc_hd__mux2_4 _1569_ (.A0(\Inst_RegFile_32x4.BD_comb[3] ),
    .A1(\Inst_RegFile_32x4.BD_reg[3] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .X(BD3));
 sky130_fd_sc_hd__mux2_1 _1570_ (.A0(\Inst_RegFile_32x4.mem[0][2] ),
    .A1(\Inst_RegFile_32x4.mem[1][2] ),
    .S(net606),
    .X(_0521_));
 sky130_fd_sc_hd__mux2_1 _1571_ (.A0(\Inst_RegFile_32x4.mem[2][2] ),
    .A1(\Inst_RegFile_32x4.mem[3][2] ),
    .S(net606),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _1572_ (.A0(_0521_),
    .A1(_0522_),
    .S(net682),
    .X(_0523_));
 sky130_fd_sc_hd__and2_1 _1573_ (.A(_0389_),
    .B(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _1574_ (.A0(\Inst_RegFile_32x4.mem[6][2] ),
    .A1(\Inst_RegFile_32x4.mem[7][2] ),
    .S(net609),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _1575_ (.A0(\Inst_RegFile_32x4.mem[4][2] ),
    .A1(\Inst_RegFile_32x4.mem[5][2] ),
    .S(net609),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_1 _1576_ (.A0(_0526_),
    .A1(_0525_),
    .S(net683),
    .X(_0527_));
 sky130_fd_sc_hd__a21bo_1 _1577_ (.A1(net642),
    .A2(_0527_),
    .B1_N(net619),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_1 _1578_ (.A0(\Inst_RegFile_32x4.mem[8][2] ),
    .A1(\Inst_RegFile_32x4.mem[9][2] ),
    .S(net608),
    .X(_0529_));
 sky130_fd_sc_hd__mux2_1 _1579_ (.A0(\Inst_RegFile_32x4.mem[10][2] ),
    .A1(\Inst_RegFile_32x4.mem[11][2] ),
    .S(net608),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_4 _1580_ (.A0(_0529_),
    .A1(_0530_),
    .S(net413),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _1581_ (.A0(\Inst_RegFile_32x4.mem[12][2] ),
    .A1(\Inst_RegFile_32x4.mem[13][2] ),
    .S(net605),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_1 _1582_ (.A0(\Inst_RegFile_32x4.mem[14][2] ),
    .A1(\Inst_RegFile_32x4.mem[15][2] ),
    .S(net605),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_1 _1583_ (.A0(_0532_),
    .A1(_0533_),
    .S(net684),
    .X(_0534_));
 sky130_fd_sc_hd__mux2_4 _1584_ (.A0(_0531_),
    .A1(_0534_),
    .S(net642),
    .X(_0535_));
 sky130_fd_sc_hd__o22a_1 _1585_ (.A1(_0524_),
    .A2(_0528_),
    .B1(net619),
    .B2(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__mux2_1 _1586_ (.A0(\Inst_RegFile_32x4.mem[16][2] ),
    .A1(\Inst_RegFile_32x4.mem[17][2] ),
    .S(net610),
    .X(_0537_));
 sky130_fd_sc_hd__mux2_1 _1587_ (.A0(\Inst_RegFile_32x4.mem[18][2] ),
    .A1(\Inst_RegFile_32x4.mem[19][2] ),
    .S(net610),
    .X(_0538_));
 sky130_fd_sc_hd__mux2_1 _1588_ (.A0(_0537_),
    .A1(_0538_),
    .S(net683),
    .X(_0539_));
 sky130_fd_sc_hd__nand2_1 _1589_ (.A(_0389_),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__nand2_1 _1590_ (.A(\Inst_RegFile_32x4.mem[23][2] ),
    .B(net607),
    .Y(_0541_));
 sky130_fd_sc_hd__o211a_1 _1591_ (.A1(_0960_),
    .A2(net607),
    .B1(net683),
    .C1(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_1 _1592_ (.A0(\Inst_RegFile_32x4.mem[20][2] ),
    .A1(\Inst_RegFile_32x4.mem[21][2] ),
    .S(net607),
    .X(_0543_));
 sky130_fd_sc_hd__nor2_1 _1593_ (.A(net682),
    .B(_0543_),
    .Y(_0544_));
 sky130_fd_sc_hd__o31a_1 _1594_ (.A1(_0389_),
    .A2(_0542_),
    .A3(_0544_),
    .B1(net619),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_1 _1595_ (.A0(\Inst_RegFile_32x4.mem[24][2] ),
    .A1(\Inst_RegFile_32x4.mem[25][2] ),
    .S(net603),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_1 _1596_ (.A0(\Inst_RegFile_32x4.mem[26][2] ),
    .A1(\Inst_RegFile_32x4.mem[27][2] ),
    .S(net604),
    .X(_0547_));
 sky130_fd_sc_hd__mux2_1 _1597_ (.A0(_0546_),
    .A1(_0547_),
    .S(net681),
    .X(_0548_));
 sky130_fd_sc_hd__mux2_1 _1598_ (.A0(\Inst_RegFile_32x4.mem[30][2] ),
    .A1(\Inst_RegFile_32x4.mem[31][2] ),
    .S(net603),
    .X(_0549_));
 sky130_fd_sc_hd__mux2_1 _1599_ (.A0(\Inst_RegFile_32x4.mem[28][2] ),
    .A1(\Inst_RegFile_32x4.mem[29][2] ),
    .S(net603),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_1 _1600_ (.A0(_0550_),
    .A1(_0549_),
    .S(net681),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_4 _1601_ (.A0(_0548_),
    .A1(_0551_),
    .S(net642),
    .X(_0552_));
 sky130_fd_sc_hd__o2bb2a_1 _1602_ (.A1_N(_0540_),
    .A2_N(_0545_),
    .B1(_0552_),
    .B2(net619),
    .X(_0553_));
 sky130_fd_sc_hd__mux2_4 _1603_ (.A0(_0536_),
    .A1(_0553_),
    .S(_0439_),
    .X(\Inst_RegFile_32x4.BD_comb[2] ));
 sky130_fd_sc_hd__mux2_4 _1604_ (.A0(\Inst_RegFile_32x4.BD_comb[2] ),
    .A1(\Inst_RegFile_32x4.BD_reg[2] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .X(BD2));
 sky130_fd_sc_hd__mux4_2 _1605_ (.A0(net688),
    .A1(net670),
    .A2(net657),
    .A3(net653),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0554_));
 sky130_fd_sc_hd__mux4_1 _1606_ (.A0(net644),
    .A1(net634),
    .A2(net668),
    .A3(net640),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ),
    .X(_0555_));
 sky130_fd_sc_hd__o21a_1 _1607_ (.A1(_0936_),
    .A2(_0555_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q ),
    .X(_0556_));
 sky130_fd_sc_hd__o21ai_4 _1608_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ),
    .A2(_0554_),
    .B1(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__mux4_1 _1609_ (.A0(net60),
    .A1(net68),
    .A2(net86),
    .A3(net2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0558_));
 sky130_fd_sc_hd__nor2_1 _1610_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ),
    .B(_0558_),
    .Y(_0559_));
 sky130_fd_sc_hd__mux4_1 _1611_ (.A0(net10),
    .A1(net88),
    .A2(net96),
    .A3(net116),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0560_));
 sky130_fd_sc_hd__nor2_1 _1612_ (.A(_0936_),
    .B(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__o31ai_4 _1613_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0559_),
    .A3(_0561_),
    .B1(_0557_),
    .Y(\Inst_RegFile_switch_matrix.JN2BEG4 ));
 sky130_fd_sc_hd__nor2_2 _1614_ (.A(\Inst_RegFile_switch_matrix.JN2BEG4 ),
    .B(_0935_),
    .Y(_0562_));
 sky130_fd_sc_hd__o21ai_1 _1615_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ),
    .A2(net110),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q ),
    .Y(_0563_));
 sky130_fd_sc_hd__mux2_1 _1616_ (.A0(net82),
    .A1(net23),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_0564_));
 sky130_fd_sc_hd__inv_1 _1617_ (.A(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__o221a_4 _1618_ (.A1(_0563_),
    .A2(_0562_),
    .B1(_0565_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q ),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ),
    .X(_0566_));
 sky130_fd_sc_hd__mux4_2 _1619_ (.A0(net70),
    .A1(net12),
    .A2(net98),
    .A3(net137),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q ),
    .X(_0567_));
 sky130_fd_sc_hd__o21ai_1 _1620_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ),
    .A2(_0567_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ),
    .Y(_0568_));
 sky130_fd_sc_hd__mux4_1 _1621_ (.A0(net77),
    .A1(net19),
    .A2(net105),
    .A3(\Inst_RegFile_switch_matrix.JN2BEG6 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q ),
    .X(_0569_));
 sky130_fd_sc_hd__nor2_1 _1622_ (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ),
    .B(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__mux4_1 _1623_ (.A0(net78),
    .A1(net20),
    .A2(net106),
    .A3(net134),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q ),
    .X(_0571_));
 sky130_fd_sc_hd__inv_2 _1624_ (.A(_0571_),
    .Y(_0572_));
 sky130_fd_sc_hd__a211o_1 _1625_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ),
    .A2(_0572_),
    .B1(_0570_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ),
    .X(_0573_));
 sky130_fd_sc_hd__o21ai_4 _1626_ (.A1(_0568_),
    .A2(_0566_),
    .B1(_0573_),
    .Y(B_ADR0));
 sky130_fd_sc_hd__mux4_1 _1627_ (.A0(net687),
    .A1(net669),
    .A2(net656),
    .A3(net651),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0574_));
 sky130_fd_sc_hd__mux4_2 _1628_ (.A0(net677),
    .A1(net633),
    .A2(net664),
    .A3(net638),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ),
    .X(_0575_));
 sky130_fd_sc_hd__or2_4 _1629_ (.A(_0575_),
    .B(_0963_),
    .X(_0576_));
 sky130_fd_sc_hd__o21a_1 _1630_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ),
    .A2(_0574_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q ),
    .X(_0577_));
 sky130_fd_sc_hd__mux4_1 _1631_ (.A0(net67),
    .A1(net79),
    .A2(net780),
    .A3(net9),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0578_));
 sky130_fd_sc_hd__mux4_1 _1632_ (.A0(net778),
    .A1(net95),
    .A2(net123),
    .A3(net140),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0579_));
 sky130_fd_sc_hd__mux2_1 _1633_ (.A0(_0578_),
    .A1(_0579_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ),
    .X(_0580_));
 sky130_fd_sc_hd__a22o_4 _1634_ (.A1(_0577_),
    .A2(_0576_),
    .B1(_0580_),
    .B2(_0964_),
    .X(\Inst_RegFile_switch_matrix.JN2BEG3 ));
 sky130_fd_sc_hd__mux4_1 _1635_ (.A0(net77),
    .A1(net19),
    .A2(net133),
    .A3(\Inst_RegFile_switch_matrix.JN2BEG5 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q ),
    .X(_0581_));
 sky130_fd_sc_hd__mux4_2 _1636_ (.A0(net78),
    .A1(net20),
    .A2(net106),
    .A3(net134),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q ),
    .X(_0582_));
 sky130_fd_sc_hd__mux4_2 _1637_ (.A0(net82),
    .A1(net8),
    .A2(net122),
    .A3(\Inst_RegFile_switch_matrix.JN2BEG3 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q ),
    .X(_0583_));
 sky130_fd_sc_hd__mux4_1 _1638_ (.A0(net70),
    .A1(net98),
    .A2(net25),
    .A3(net126),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q ),
    .X(_0584_));
 sky130_fd_sc_hd__mux4_2 _1639_ (.A0(_0581_),
    .A1(_0582_),
    .A2(_0584_),
    .A3(_0583_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q ),
    .X(A_ADR0));
 sky130_fd_sc_hd__mux4_1 _1640_ (.A0(net686),
    .A1(net669),
    .A2(net656),
    .A3(net644),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0585_));
 sky130_fd_sc_hd__or2_1 _1641_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ),
    .B(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__mux4_1 _1642_ (.A0(net677),
    .A1(net634),
    .A2(net665),
    .A3(net638),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .X(_0587_));
 sky130_fd_sc_hd__o21a_1 _1643_ (.A1(_0981_),
    .A2(_0587_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0588_));
 sky130_fd_sc_hd__mux4_1 _1644_ (.A0(net60),
    .A1(net66),
    .A2(net85),
    .A3(net8),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0589_));
 sky130_fd_sc_hd__mux4_1 _1645_ (.A0(net777),
    .A1(net94),
    .A2(net110),
    .A3(net122),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_1 _1646_ (.A0(_0589_),
    .A1(_0590_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ),
    .X(_0591_));
 sky130_fd_sc_hd__a22o_1 _1647_ (.A1(_0586_),
    .A2(_0588_),
    .B1(_0591_),
    .B2(_0982_),
    .X(\Inst_RegFile_switch_matrix.JW2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1648_ (.A0(net686),
    .A1(net669),
    .A2(net656),
    .A3(net644),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0592_));
 sky130_fd_sc_hd__nor2_1 _1649_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ),
    .B(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__mux4_1 _1650_ (.A0(net677),
    .A1(net633),
    .A2(net664),
    .A3(net638),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_0594_));
 sky130_fd_sc_hd__o21ai_1 _1651_ (.A1(_0983_),
    .A2(_0594_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q ),
    .Y(_0595_));
 sky130_fd_sc_hd__mux4_1 _1652_ (.A0(net66),
    .A1(net8),
    .A2(net2),
    .A3(net25),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_0596_));
 sky130_fd_sc_hd__nor2_1 _1653_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ),
    .B(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__mux4_1 _1654_ (.A0(net777),
    .A1(net94),
    .A2(net110),
    .A3(net122),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0598_));
 sky130_fd_sc_hd__nor2_1 _1655_ (.A(_0983_),
    .B(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__o32a_1 _1656_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q ),
    .A2(_0597_),
    .A3(_0599_),
    .B1(_0593_),
    .B2(_0595_),
    .X(_0600_));
 sky130_fd_sc_hd__inv_1 _1657_ (.A(_0600_),
    .Y(\Inst_RegFile_switch_matrix.JS2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1658_ (.A0(net136),
    .A1(net673),
    .A2(net659),
    .A3(net646),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0601_));
 sky130_fd_sc_hd__mux4_1 _1659_ (.A0(net679),
    .A1(net636),
    .A2(net667),
    .A3(net640),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .X(_0602_));
 sky130_fd_sc_hd__or2_1 _1660_ (.A(_0984_),
    .B(_0602_),
    .X(_0603_));
 sky130_fd_sc_hd__o21a_1 _1661_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ),
    .A2(_0601_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q ),
    .X(_0604_));
 sky130_fd_sc_hd__mux4_1 _1662_ (.A0(net777),
    .A1(net94),
    .A2(net113),
    .A3(net122),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0605_));
 sky130_fd_sc_hd__mux4_1 _1663_ (.A0(net60),
    .A1(net66),
    .A2(net82),
    .A3(net8),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_1 _1664_ (.A0(_0605_),
    .A1(_0606_),
    .S(_0984_),
    .X(_0607_));
 sky130_fd_sc_hd__a22o_1 _1665_ (.A1(_0603_),
    .A2(_0604_),
    .B1(_0607_),
    .B2(_0985_),
    .X(\Inst_RegFile_switch_matrix.E2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1666_ (.A0(net686),
    .A1(net672),
    .A2(net659),
    .A3(net646),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0608_));
 sky130_fd_sc_hd__or2_1 _1667_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ),
    .B(_0608_),
    .X(_0609_));
 sky130_fd_sc_hd__mux4_1 _1668_ (.A0(net680),
    .A1(net636),
    .A2(net668),
    .A3(net640),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ),
    .X(_0610_));
 sky130_fd_sc_hd__o211a_1 _1669_ (.A1(_0986_),
    .A2(_0610_),
    .B1(_0609_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q ),
    .X(_0611_));
 sky130_fd_sc_hd__mux4_1 _1670_ (.A0(net777),
    .A1(net94),
    .A2(net122),
    .A3(net139),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0612_));
 sky130_fd_sc_hd__mux4_1 _1671_ (.A0(net66),
    .A1(net2),
    .A2(net82),
    .A3(net8),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _1672_ (.A0(_0612_),
    .A1(_0613_),
    .S(_0986_),
    .X(_0614_));
 sky130_fd_sc_hd__a21o_1 _1673_ (.A1(_0987_),
    .A2(_0614_),
    .B1(_0611_),
    .X(\Inst_RegFile_switch_matrix.JN2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1674_ (.A0(net687),
    .A1(net671),
    .A2(net652),
    .A3(net645),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0615_));
 sky130_fd_sc_hd__or2_1 _1675_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ),
    .B(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__mux4_1 _1676_ (.A0(net676),
    .A1(net635),
    .A2(net666),
    .A3(net639),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0617_));
 sky130_fd_sc_hd__o21a_1 _1677_ (.A1(_0988_),
    .A2(_0617_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q ),
    .X(_0618_));
 sky130_fd_sc_hd__mux4_1 _1678_ (.A0(net59),
    .A1(net7),
    .A2(net65),
    .A3(net778),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0619_));
 sky130_fd_sc_hd__mux4_1 _1679_ (.A0(net93),
    .A1(net109),
    .A2(net112),
    .A3(net121),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_1 _1680_ (.A0(_0619_),
    .A1(_0620_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ),
    .X(_0621_));
 sky130_fd_sc_hd__a22o_1 _1681_ (.A1(_0616_),
    .A2(_0618_),
    .B1(_0621_),
    .B2(_0989_),
    .X(\Inst_RegFile_switch_matrix.JW2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1682_ (.A0(net687),
    .A1(net671),
    .A2(net423),
    .A3(net645),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0622_));
 sky130_fd_sc_hd__or2_1 _1683_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ),
    .B(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__mux4_1 _1684_ (.A0(net676),
    .A1(net635),
    .A2(net666),
    .A3(net639),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ),
    .X(_0624_));
 sky130_fd_sc_hd__o21a_1 _1685_ (.A1(_0990_),
    .A2(_0624_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q ),
    .X(_0625_));
 sky130_fd_sc_hd__mux4_1 _1686_ (.A0(net65),
    .A1(net7),
    .A2(net1),
    .A3(net778),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ),
    .X(_0626_));
 sky130_fd_sc_hd__mux4_1 _1687_ (.A0(net93),
    .A1(net109),
    .A2(net121),
    .A3(net138),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_1 _1688_ (.A0(_0626_),
    .A1(_0627_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_0628_));
 sky130_fd_sc_hd__a22o_1 _1689_ (.A1(_0623_),
    .A2(_0625_),
    .B1(_0628_),
    .B2(_0991_),
    .X(\Inst_RegFile_switch_matrix.JS2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1690_ (.A0(net680),
    .A1(net637),
    .A2(net667),
    .A3(net641),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ),
    .X(_0629_));
 sky130_fd_sc_hd__or2_1 _1691_ (.A(_0992_),
    .B(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__mux4_1 _1692_ (.A0(net687),
    .A1(net673),
    .A2(net654),
    .A3(net647),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0631_));
 sky130_fd_sc_hd__o21a_1 _1693_ (.A1(_0631_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q ),
    .X(_0632_));
 sky130_fd_sc_hd__mux4_1 _1694_ (.A0(net7),
    .A1(net93),
    .A2(net21),
    .A3(net121),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ),
    .X(_0633_));
 sky130_fd_sc_hd__mux4_1 _1695_ (.A0(net59),
    .A1(net65),
    .A2(net81),
    .A3(net84),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _1696_ (.A0(_0633_),
    .A1(_0634_),
    .S(_0992_),
    .X(_0635_));
 sky130_fd_sc_hd__a22o_4 _1697_ (.A1(_0632_),
    .A2(_0630_),
    .B1(_0635_),
    .B2(_0993_),
    .X(\Inst_RegFile_switch_matrix.E2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1698_ (.A0(net687),
    .A1(net669),
    .A2(net651),
    .A3(net644),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0636_));
 sky130_fd_sc_hd__or2_1 _1699_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ),
    .B(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__mux4_1 _1700_ (.A0(net677),
    .A1(net633),
    .A2(net664),
    .A3(net638),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ),
    .X(_0638_));
 sky130_fd_sc_hd__o21a_1 _1701_ (.A1(_0994_),
    .A2(_0638_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q ),
    .X(_0639_));
 sky130_fd_sc_hd__mux4_1 _1702_ (.A0(net65),
    .A1(net1),
    .A2(net81),
    .A3(net7),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ),
    .X(_0640_));
 sky130_fd_sc_hd__mux4_1 _1703_ (.A0(net24),
    .A1(net778),
    .A2(net93),
    .A3(net121),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0641_));
 sky130_fd_sc_hd__mux2_1 _1704_ (.A0(_0640_),
    .A1(_0641_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ),
    .X(_0642_));
 sky130_fd_sc_hd__a22o_1 _1705_ (.A1(_0637_),
    .A2(_0639_),
    .B1(_0642_),
    .B2(_0995_),
    .X(\Inst_RegFile_switch_matrix.JN2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1706_ (.A0(net137),
    .A1(net669),
    .A2(net656),
    .A3(net651),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_0643_));
 sky130_fd_sc_hd__or2_1 _1707_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ),
    .B(_0643_),
    .X(_0644_));
 sky130_fd_sc_hd__mux4_1 _1708_ (.A0(net644),
    .A1(net411),
    .A2(net664),
    .A3(net415),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_0645_));
 sky130_fd_sc_hd__o21a_1 _1709_ (.A1(_0996_),
    .A2(_0645_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q ),
    .X(_0646_));
 sky130_fd_sc_hd__mux4_1 _1710_ (.A0(net59),
    .A1(net1),
    .A2(net63),
    .A3(net5),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ),
    .X(_0647_));
 sky130_fd_sc_hd__mux4_1 _1711_ (.A0(net87),
    .A1(net91),
    .A2(net89),
    .A3(net115),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ),
    .X(_0648_));
 sky130_fd_sc_hd__mux2_1 _1712_ (.A0(_0647_),
    .A1(_0648_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ),
    .X(_0649_));
 sky130_fd_sc_hd__a22o_1 _1713_ (.A1(_0644_),
    .A2(_0646_),
    .B1(_0649_),
    .B2(_0997_),
    .X(\Inst_RegFile_switch_matrix.JW2BEG7 ));
 sky130_fd_sc_hd__mux4_1 _1714_ (.A0(net686),
    .A1(net652),
    .A2(net658),
    .A3(net645),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_0650_));
 sky130_fd_sc_hd__or2_1 _1715_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ),
    .B(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__mux4_1 _1716_ (.A0(net678),
    .A1(net635),
    .A2(net666),
    .A3(net639),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_0652_));
 sky130_fd_sc_hd__o21a_1 _1717_ (.A1(_0998_),
    .A2(_0652_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q ),
    .X(_0653_));
 sky130_fd_sc_hd__mux4_1 _1718_ (.A0(net62),
    .A1(net64),
    .A2(net6),
    .A3(net777),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0654_));
 sky130_fd_sc_hd__mux4_1 _1719_ (.A0(net92),
    .A1(net108),
    .A2(net111),
    .A3(net120),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_1 _1720_ (.A0(_0654_),
    .A1(_0655_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ),
    .X(_0656_));
 sky130_fd_sc_hd__a22o_1 _1721_ (.A1(_0651_),
    .A2(_0653_),
    .B1(_0656_),
    .B2(_0999_),
    .X(\Inst_RegFile_switch_matrix.JW2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1722_ (.A0(net644),
    .A1(net677),
    .A2(net664),
    .A3(net633),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0657_));
 sky130_fd_sc_hd__or2_1 _1723_ (.A(_1000_),
    .B(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__mux4_1 _1724_ (.A0(net689),
    .A1(net669),
    .A2(net656),
    .A3(net651),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0659_));
 sky130_fd_sc_hd__o21a_1 _1725_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q ),
    .A2(_0659_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q ),
    .X(_0660_));
 sky130_fd_sc_hd__mux4_1 _1726_ (.A0(net87),
    .A1(net91),
    .A2(net111),
    .A3(net115),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0661_));
 sky130_fd_sc_hd__mux4_1 _1727_ (.A0(net59),
    .A1(net1),
    .A2(net63),
    .A3(net5),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_1 _1728_ (.A0(_0661_),
    .A1(_0662_),
    .S(_1000_),
    .X(_0663_));
 sky130_fd_sc_hd__a22o_1 _1729_ (.A1(_0658_),
    .A2(_0660_),
    .B1(_0663_),
    .B2(_1001_),
    .X(\Inst_RegFile_switch_matrix.JS2BEG7 ));
 sky130_fd_sc_hd__mux4_1 _1730_ (.A0(net676),
    .A1(net635),
    .A2(net666),
    .A3(net639),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ),
    .X(_0664_));
 sky130_fd_sc_hd__mux4_1 _1731_ (.A0(net686),
    .A1(net652),
    .A2(net658),
    .A3(net645),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ),
    .X(_0665_));
 sky130_fd_sc_hd__or2_1 _1732_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ),
    .B(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__o211a_1 _1733_ (.A1(_1002_),
    .A2(_0664_),
    .B1(_0666_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q ),
    .X(_0667_));
 sky130_fd_sc_hd__mux4_1 _1734_ (.A0(net64),
    .A1(net6),
    .A2(net779),
    .A3(net777),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ),
    .X(_0668_));
 sky130_fd_sc_hd__mux4_1 _1735_ (.A0(net92),
    .A1(net120),
    .A2(net108),
    .A3(net137),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ),
    .X(_0669_));
 sky130_fd_sc_hd__mux2_1 _1736_ (.A0(_0668_),
    .A1(_0669_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ),
    .X(_0670_));
 sky130_fd_sc_hd__and2b_1 _1737_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q ),
    .B(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__or2_1 _1738_ (.A(_0667_),
    .B(_0671_),
    .X(\Inst_RegFile_switch_matrix.JS2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1739_ (.A0(net115),
    .A1(net669),
    .A2(net656),
    .A3(net651),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_0672_));
 sky130_fd_sc_hd__mux4_1 _1740_ (.A0(net644),
    .A1(net411),
    .A2(net665),
    .A3(net415),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_0673_));
 sky130_fd_sc_hd__or2_1 _1741_ (.A(_1003_),
    .B(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__o21a_1 _1742_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_0672_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q ),
    .X(_0675_));
 sky130_fd_sc_hd__mux4_1 _1743_ (.A0(net23),
    .A1(net89),
    .A2(net87),
    .A3(net91),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_0676_));
 sky130_fd_sc_hd__mux4_1 _1744_ (.A0(net59),
    .A1(net1),
    .A2(net63),
    .A3(net5),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_1 _1745_ (.A0(_0676_),
    .A1(_0677_),
    .S(_1003_),
    .X(_0678_));
 sky130_fd_sc_hd__a22o_1 _1746_ (.A1(_0674_),
    .A2(_0675_),
    .B1(_0678_),
    .B2(_1004_),
    .X(\Inst_RegFile_switch_matrix.E2BEG7 ));
 sky130_fd_sc_hd__mux4_1 _1747_ (.A0(net686),
    .A1(net423),
    .A2(net658),
    .A3(net645),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0679_));
 sky130_fd_sc_hd__or2_1 _1748_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ),
    .B(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__mux4_1 _1749_ (.A0(net676),
    .A1(net635),
    .A2(net666),
    .A3(net409),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0681_));
 sky130_fd_sc_hd__o21a_1 _1750_ (.A1(_1005_),
    .A2(_0681_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q ),
    .X(_0682_));
 sky130_fd_sc_hd__mux4_1 _1751_ (.A0(net6),
    .A1(net92),
    .A2(net777),
    .A3(net120),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0683_));
 sky130_fd_sc_hd__mux4_1 _1752_ (.A0(net62),
    .A1(net64),
    .A2(net80),
    .A3(net83),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_0684_));
 sky130_fd_sc_hd__mux2_1 _1753_ (.A0(_0683_),
    .A1(_0684_),
    .S(_1005_),
    .X(_0685_));
 sky130_fd_sc_hd__a22o_1 _1754_ (.A1(_0680_),
    .A2(_0682_),
    .B1(_0685_),
    .B2(_1006_),
    .X(\Inst_RegFile_switch_matrix.E2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1755_ (.A0(net644),
    .A1(net411),
    .A2(net664),
    .A3(net415),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ),
    .X(_0686_));
 sky130_fd_sc_hd__or2_1 _1756_ (.A(_1007_),
    .B(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__mux4_1 _1757_ (.A0(net689),
    .A1(net669),
    .A2(net656),
    .A3(net651),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ),
    .X(_0688_));
 sky130_fd_sc_hd__o21a_1 _1758_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ),
    .A2(_0688_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q ),
    .X(_0689_));
 sky130_fd_sc_hd__mux4_1 _1759_ (.A0(net59),
    .A1(net63),
    .A2(net83),
    .A3(net1),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ),
    .X(_0690_));
 sky130_fd_sc_hd__mux4_1 _1760_ (.A0(net5),
    .A1(net91),
    .A2(net87),
    .A3(net115),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_0691_));
 sky130_fd_sc_hd__mux2_1 _1761_ (.A0(_0690_),
    .A1(_0691_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ),
    .X(_0692_));
 sky130_fd_sc_hd__a22o_4 _1762_ (.A1(_0687_),
    .A2(_0689_),
    .B1(_0692_),
    .B2(_1008_),
    .X(\Inst_RegFile_switch_matrix.JN2BEG7 ));
 sky130_fd_sc_hd__mux4_1 _1763_ (.A0(net676),
    .A1(net635),
    .A2(net666),
    .A3(net409),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ),
    .X(_0693_));
 sky130_fd_sc_hd__or2_1 _1764_ (.A(_1009_),
    .B(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__mux4_1 _1765_ (.A0(net686),
    .A1(net423),
    .A2(net658),
    .A3(net645),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ),
    .X(_0695_));
 sky130_fd_sc_hd__o21a_1 _1766_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ),
    .A2(_0695_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_0696_));
 sky130_fd_sc_hd__mux4_1 _1767_ (.A0(net64),
    .A1(net80),
    .A2(net779),
    .A3(net6),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_0697_));
 sky130_fd_sc_hd__mux4_1 _1768_ (.A0(net23),
    .A1(net777),
    .A2(net92),
    .A3(net120),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_1 _1769_ (.A0(_0697_),
    .A1(_0698_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ),
    .X(_0699_));
 sky130_fd_sc_hd__a22o_1 _1770_ (.A1(_0694_),
    .A2(_0696_),
    .B1(_0699_),
    .B2(_1010_),
    .X(\Inst_RegFile_switch_matrix.JN2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1771_ (.A0(net85),
    .A1(net780),
    .A2(net113),
    .A3(net689),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .X(_0700_));
 sky130_fd_sc_hd__mux4_1 _1772_ (.A0(net670),
    .A1(net655),
    .A2(net657),
    .A3(net645),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_1 _1773_ (.A0(_0700_),
    .A1(_0701_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _1774_ (.A0(net75),
    .A1(net17),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q ),
    .X(_0703_));
 sky130_fd_sc_hd__nand2_1 _1775_ (.A(\Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q ),
    .B(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .Y(_0704_));
 sky130_fd_sc_hd__o21a_1 _1776_ (.A1(_0950_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q ),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q ),
    .X(_0705_));
 sky130_fd_sc_hd__a2bb2o_2 _1777_ (.A1_N(\Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q ),
    .A2_N(_0703_),
    .B1(_0704_),
    .B2(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__clkinv_2 _1778_ (.A(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__mux4_2 _1779_ (.A0(net75),
    .A1(net103),
    .A2(net17),
    .A3(\Inst_RegFile_switch_matrix.JS2BEG4 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q ),
    .X(_0708_));
 sky130_fd_sc_hd__mux4_2 _1780_ (.A0(_0707_),
    .A1(_0708_),
    .A2(_0147_),
    .A3(_0372_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .X(_0709_));
 sky130_fd_sc_hd__mux4_1 _1781_ (.A0(net678),
    .A1(net634),
    .A2(net665),
    .A3(net638),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_1 _1782_ (.A0(_0710_),
    .A1(_0709_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_0711_));
 sky130_fd_sc_hd__mux2_1 _1783_ (.A0(_0702_),
    .A1(_0711_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q ),
    .X(\Inst_RegFile_switch_matrix.W6BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1784_ (.A0(net84),
    .A1(net779),
    .A2(net112),
    .A3(net688),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .X(_0712_));
 sky130_fd_sc_hd__mux2_1 _1785_ (.A0(net651),
    .A1(net644),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_0713_));
 sky130_fd_sc_hd__mux2_1 _1786_ (.A0(net669),
    .A1(net656),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_0714_));
 sky130_fd_sc_hd__and2b_1 _1787_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .B(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__a21bo_1 _1788_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .A2(_0713_),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ),
    .X(_0716_));
 sky130_fd_sc_hd__o22a_1 _1789_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ),
    .A2(_0712_),
    .B1(_0715_),
    .B2(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__mux4_2 _1790_ (.A0(net74),
    .A1(net16),
    .A2(net102),
    .A3(net130),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q ),
    .X(_0718_));
 sky130_fd_sc_hd__mux4_2 _1791_ (.A0(net74),
    .A1(net16),
    .A2(net102),
    .A3(net130),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q ),
    .X(_0719_));
 sky130_fd_sc_hd__mux4_1 _1792_ (.A0(_0718_),
    .A1(_0719_),
    .A2(_1033_),
    .A3(net685),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .X(_0720_));
 sky130_fd_sc_hd__mux4_1 _1793_ (.A0(net411),
    .A1(net415),
    .A2(net664),
    .A3(net638),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _1794_ (.A0(_0721_),
    .A1(_0720_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ),
    .X(_0722_));
 sky130_fd_sc_hd__mux2_1 _1795_ (.A0(_0717_),
    .A1(_0722_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q ),
    .X(\Inst_RegFile_switch_matrix.W6BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1796_ (.A0(net67),
    .A1(net95),
    .A2(net23),
    .A3(net123),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q ),
    .X(_0723_));
 sky130_fd_sc_hd__mux4_2 _1797_ (.A0(net411),
    .A1(_0147_),
    .A2(_0372_),
    .A3(_0723_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q ),
    .X(_0724_));
 sky130_fd_sc_hd__mux4_1 _1798_ (.A0(net60),
    .A1(net88),
    .A2(net116),
    .A3(net670),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q ),
    .X(_0725_));
 sky130_fd_sc_hd__mux2_4 _1799_ (.A0(_0725_),
    .A1(_0724_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q ),
    .X(\Inst_RegFile_switch_matrix.WW4BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1800_ (.A0(net67),
    .A1(net9),
    .A2(net113),
    .A3(net123),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q ),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_1 _1801_ (.A0(net685),
    .A1(_0726_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ),
    .X(_0727_));
 sky130_fd_sc_hd__mux2_1 _1802_ (.A0(net638),
    .A1(_1033_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ),
    .X(_0728_));
 sky130_fd_sc_hd__mux2_1 _1803_ (.A0(_0728_),
    .A1(_0727_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ),
    .X(_0729_));
 sky130_fd_sc_hd__mux4_1 _1804_ (.A0(net59),
    .A1(net87),
    .A2(net115),
    .A3(net644),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _1805_ (.A0(_0730_),
    .A1(_0729_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q ),
    .X(\Inst_RegFile_switch_matrix.WW4BEG2 ));
 sky130_fd_sc_hd__mux4_2 _1806_ (.A0(net635),
    .A1(_0707_),
    .A2(_0708_),
    .A3(_0159_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q ),
    .X(_0731_));
 sky130_fd_sc_hd__mux4_1 _1807_ (.A0(net62),
    .A1(net90),
    .A2(net688),
    .A3(net423),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q ),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_4 _1808_ (.A0(_0732_),
    .A1(_0731_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q ),
    .X(\Inst_RegFile_switch_matrix.WW4BEG1 ));
 sky130_fd_sc_hd__mux2_1 _1809_ (.A0(_0719_),
    .A1(_0386_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _1810_ (.A0(net664),
    .A1(_0718_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _1811_ (.A0(_0734_),
    .A1(_0733_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q ),
    .X(_0735_));
 sky130_fd_sc_hd__mux4_1 _1812_ (.A0(net61),
    .A1(net89),
    .A2(net689),
    .A3(net656),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q ),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_1 _1813_ (.A0(_0736_),
    .A1(_0735_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q ),
    .X(\Inst_RegFile_switch_matrix.WW4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1814_ (.A0(net60),
    .A1(net2),
    .A2(net116),
    .A3(net673),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ),
    .X(_0737_));
 sky130_fd_sc_hd__or2_1 _1815_ (.A(\Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ),
    .B(net680),
    .X(_0738_));
 sky130_fd_sc_hd__a21oi_1 _1816_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ),
    .A2(_0146_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ),
    .Y(_0739_));
 sky130_fd_sc_hd__mux4_2 _1817_ (.A0(net63),
    .A1(net91),
    .A2(net5),
    .A3(net140),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q ),
    .X(_0740_));
 sky130_fd_sc_hd__mux2_1 _1818_ (.A0(_0372_),
    .A1(_0740_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ),
    .X(_0741_));
 sky130_fd_sc_hd__a22o_1 _1819_ (.A1(_0738_),
    .A2(_0739_),
    .B1(_0741_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ),
    .X(_0742_));
 sky130_fd_sc_hd__mux2_1 _1820_ (.A0(_0737_),
    .A1(_0742_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q ),
    .X(\Inst_RegFile_switch_matrix.SS4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _1821_ (.A0(net641),
    .A1(_1033_),
    .A2(net685),
    .A3(_0213_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ),
    .X(_0743_));
 sky130_fd_sc_hd__mux4_2 _1822_ (.A0(net59),
    .A1(net1),
    .A2(net115),
    .A3(net421),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ),
    .X(_0744_));
 sky130_fd_sc_hd__mux2_4 _1823_ (.A0(_0744_),
    .A1(_0743_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q ),
    .X(\Inst_RegFile_switch_matrix.SS4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1824_ (.A0(net62),
    .A1(net779),
    .A2(net688),
    .A3(net654),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ),
    .X(_0745_));
 sky130_fd_sc_hd__mux4_2 _1825_ (.A0(net637),
    .A1(_0707_),
    .A2(_0708_),
    .A3(_0179_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ),
    .X(_0746_));
 sky130_fd_sc_hd__mux2_4 _1826_ (.A0(_0745_),
    .A1(_0746_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q ),
    .X(\Inst_RegFile_switch_matrix.SS4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1827_ (.A0(net667),
    .A1(_0718_),
    .A2(_0719_),
    .A3(_0401_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ),
    .X(_0747_));
 sky130_fd_sc_hd__mux4_1 _1828_ (.A0(net61),
    .A1(net780),
    .A2(net689),
    .A3(net660),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ),
    .X(_0748_));
 sky130_fd_sc_hd__mux2_1 _1829_ (.A0(_0748_),
    .A1(_0747_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q ),
    .X(\Inst_RegFile_switch_matrix.SS4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1830_ (.A0(net86),
    .A1(net114),
    .A2(net780),
    .A3(net689),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .X(_0749_));
 sky130_fd_sc_hd__or2_1 _1831_ (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ),
    .B(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__mux4_1 _1832_ (.A0(net672),
    .A1(net653),
    .A2(net659),
    .A3(net422),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .X(_0751_));
 sky130_fd_sc_hd__inv_2 _1833_ (.A(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__a21oi_1 _1834_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ),
    .A2(_0752_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q ),
    .Y(_0753_));
 sky130_fd_sc_hd__mux4_2 _1835_ (.A0(_0707_),
    .A1(_0708_),
    .A2(_0147_),
    .A3(_0372_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .X(_0754_));
 sky130_fd_sc_hd__mux4_1 _1836_ (.A0(net679),
    .A1(net636),
    .A2(net667),
    .A3(net640),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .X(_0755_));
 sky130_fd_sc_hd__mux2_4 _1837_ (.A0(_0755_),
    .A1(_0754_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_0756_));
 sky130_fd_sc_hd__a22o_1 _1838_ (.A1(_0750_),
    .A2(_0753_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q ),
    .B2(_0756_),
    .X(\Inst_RegFile_switch_matrix.E6BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1839_ (.A0(net83),
    .A1(net111),
    .A2(net779),
    .A3(net688),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_0757_));
 sky130_fd_sc_hd__mux2_1 _1840_ (.A0(net653),
    .A1(net422),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_0758_));
 sky130_fd_sc_hd__mux2_1 _1841_ (.A0(net672),
    .A1(net659),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_0759_));
 sky130_fd_sc_hd__and2b_1 _1842_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .B(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__a21bo_1 _1843_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .A2(_0758_),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ),
    .X(_0761_));
 sky130_fd_sc_hd__o22a_1 _1844_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ),
    .A2(_0757_),
    .B1(_0760_),
    .B2(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__mux4_1 _1845_ (.A0(_0718_),
    .A1(_0719_),
    .A2(_1033_),
    .A3(net685),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .X(_0763_));
 sky130_fd_sc_hd__mux4_1 _1846_ (.A0(net679),
    .A1(net636),
    .A2(net667),
    .A3(net640),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_0764_));
 sky130_fd_sc_hd__mux2_1 _1847_ (.A0(_0764_),
    .A1(_0763_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ),
    .X(_0765_));
 sky130_fd_sc_hd__mux2_1 _1848_ (.A0(_0762_),
    .A1(_0765_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q ),
    .X(\Inst_RegFile_switch_matrix.E6BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1849_ (.A0(net60),
    .A1(net2),
    .A2(net88),
    .A3(net673),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ),
    .X(_0766_));
 sky130_fd_sc_hd__mux4_1 _1850_ (.A0(net69),
    .A1(net11),
    .A2(net114),
    .A3(net125),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q ),
    .X(_0767_));
 sky130_fd_sc_hd__mux2_1 _1851_ (.A0(_0372_),
    .A1(_0767_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ),
    .X(_0768_));
 sky130_fd_sc_hd__nor2_1 _1852_ (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ),
    .B(net679),
    .Y(_0769_));
 sky130_fd_sc_hd__a211oi_1 _1853_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ),
    .A2(_0146_),
    .B1(_0769_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ),
    .Y(_0770_));
 sky130_fd_sc_hd__a21bo_1 _1854_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ),
    .A2(_0768_),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q ),
    .X(_0771_));
 sky130_fd_sc_hd__o22a_1 _1855_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q ),
    .A2(_0766_),
    .B1(_0770_),
    .B2(_0771_),
    .X(\Inst_RegFile_switch_matrix.EE4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _1856_ (.A0(net86),
    .A1(net11),
    .A2(net97),
    .A3(net125),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q ),
    .X(_0772_));
 sky130_fd_sc_hd__mux4_1 _1857_ (.A0(net640),
    .A1(_1033_),
    .A2(net685),
    .A3(_0772_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ),
    .X(_0773_));
 sky130_fd_sc_hd__nand2b_1 _1858_ (.A_N(net1),
    .B(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ),
    .Y(_0774_));
 sky130_fd_sc_hd__o21ba_1 _1859_ (.A1(net59),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ),
    .X(_0775_));
 sky130_fd_sc_hd__mux2_1 _1860_ (.A0(net87),
    .A1(net422),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ),
    .X(_0776_));
 sky130_fd_sc_hd__a221o_1 _1861_ (.A1(_0774_),
    .A2(_0775_),
    .B1(_0776_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q ),
    .X(_0777_));
 sky130_fd_sc_hd__o21a_1 _1862_ (.A1(_1011_),
    .A2(_0773_),
    .B1(_0777_),
    .X(\Inst_RegFile_switch_matrix.EE4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1863_ (.A0(net62),
    .A1(net779),
    .A2(net90),
    .A3(net654),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ),
    .X(_0778_));
 sky130_fd_sc_hd__mux2_4 _1864_ (.A0(_0708_),
    .A1(_0584_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ),
    .X(_0779_));
 sky130_fd_sc_hd__or2_1 _1865_ (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ),
    .B(net637),
    .X(_0780_));
 sky130_fd_sc_hd__a21oi_1 _1866_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ),
    .A2(_0706_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ),
    .Y(_0781_));
 sky130_fd_sc_hd__a221o_1 _1867_ (.A1(_0779_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ),
    .B1(_0780_),
    .B2(_0781_),
    .C1(_1012_),
    .X(_0782_));
 sky130_fd_sc_hd__o21a_1 _1868_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q ),
    .A2(_0778_),
    .B1(_0782_),
    .X(\Inst_RegFile_switch_matrix.EE4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1869_ (.A0(net667),
    .A1(_0718_),
    .A2(_0719_),
    .A3(_0567_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ),
    .X(_0783_));
 sky130_fd_sc_hd__nand2b_1 _1870_ (.A_N(net780),
    .B(\Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ),
    .Y(_0784_));
 sky130_fd_sc_hd__o21ba_1 _1871_ (.A1(net61),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ),
    .X(_0785_));
 sky130_fd_sc_hd__mux2_1 _1872_ (.A0(net89),
    .A1(net659),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ),
    .X(_0786_));
 sky130_fd_sc_hd__a221o_1 _1873_ (.A1(_0784_),
    .A2(_0785_),
    .B1(_0786_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q ),
    .X(_0787_));
 sky130_fd_sc_hd__o21a_1 _1874_ (.A1(_1013_),
    .A2(_0783_),
    .B1(_0787_),
    .X(\Inst_RegFile_switch_matrix.EE4BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1875_ (.A0(net83),
    .A1(net93),
    .A2(net7),
    .A3(net121),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q ),
    .X(_0788_));
 sky130_fd_sc_hd__mux4_2 _1876_ (.A0(net679),
    .A1(_0147_),
    .A2(_0372_),
    .A3(_0788_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q ),
    .X(_0789_));
 sky130_fd_sc_hd__mux4_1 _1877_ (.A0(net60),
    .A1(net2),
    .A2(net116),
    .A3(net672),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q ),
    .X(_0790_));
 sky130_fd_sc_hd__mux2_4 _1878_ (.A0(_0790_),
    .A1(_0789_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q ),
    .X(\Inst_RegFile_switch_matrix.NN4BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1879_ (.A0(net65),
    .A1(net93),
    .A2(net7),
    .A3(net139),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q ),
    .X(_0791_));
 sky130_fd_sc_hd__mux4_1 _1880_ (.A0(net641),
    .A1(_1033_),
    .A2(net685),
    .A3(_0791_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ),
    .X(_0792_));
 sky130_fd_sc_hd__mux4_1 _1881_ (.A0(net59),
    .A1(net1),
    .A2(net115),
    .A3(net422),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ),
    .X(_0793_));
 sky130_fd_sc_hd__mux2_1 _1882_ (.A0(_0793_),
    .A1(_0792_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q ),
    .X(\Inst_RegFile_switch_matrix.NN4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1883_ (.A0(net62),
    .A1(net779),
    .A2(net688),
    .A3(net653),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ),
    .X(_0794_));
 sky130_fd_sc_hd__nor2_1 _1884_ (.A(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ),
    .B(net636),
    .Y(_0795_));
 sky130_fd_sc_hd__a211o_1 _1885_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ),
    .A2(_0706_),
    .B1(_0795_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ),
    .X(_0796_));
 sky130_fd_sc_hd__mux2_4 _1886_ (.A0(_0708_),
    .A1(_0133_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ),
    .X(_0797_));
 sky130_fd_sc_hd__a21bo_1 _1887_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ),
    .A2(_0797_),
    .B1_N(_0796_),
    .X(_0798_));
 sky130_fd_sc_hd__mux2_4 _1888_ (.A0(_0794_),
    .A1(_0798_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q ),
    .X(\Inst_RegFile_switch_matrix.NN4BEG1 ));
 sky130_fd_sc_hd__mux2_1 _1889_ (.A0(_0719_),
    .A1(_0361_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ),
    .X(_0799_));
 sky130_fd_sc_hd__mux2_1 _1890_ (.A0(net667),
    .A1(_0718_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ),
    .X(_0800_));
 sky130_fd_sc_hd__mux2_1 _1891_ (.A0(_0800_),
    .A1(_0799_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ),
    .X(_0801_));
 sky130_fd_sc_hd__mux4_1 _1892_ (.A0(net61),
    .A1(net780),
    .A2(net689),
    .A3(net659),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ),
    .X(_0802_));
 sky130_fd_sc_hd__mux2_1 _1893_ (.A0(_0802_),
    .A1(_0801_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q ),
    .X(\Inst_RegFile_switch_matrix.NN4BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1894_ (.A0(net86),
    .A1(net110),
    .A2(net137),
    .A3(\Inst_RegFile_switch_matrix.JN2BEG1 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q ),
    .X(_0803_));
 sky130_fd_sc_hd__mux4_1 _1895_ (.A0(net671),
    .A1(_0437_),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG2 ),
    .A3(_0803_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q ),
    .X(\Inst_RegFile_switch_matrix.W1BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1896_ (.A0(net409),
    .A1(net685),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG1 ),
    .A3(net394),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q ),
    .X(\Inst_RegFile_switch_matrix.W1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1897_ (.A0(net635),
    .A1(_0582_),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG0 ),
    .A3(_0158_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q ),
    .X(\Inst_RegFile_switch_matrix.W1BEG1 ));
 sky130_fd_sc_hd__mux4_2 _1898_ (.A0(net72),
    .A1(net14),
    .A2(net100),
    .A3(net128),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q ),
    .X(_0804_));
 sky130_fd_sc_hd__mux4_2 _1899_ (.A0(net81),
    .A1(net126),
    .A2(net7),
    .A3(\Inst_RegFile_switch_matrix.E2BEG2 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q ),
    .X(_0805_));
 sky130_fd_sc_hd__mux4_1 _1900_ (.A0(net666),
    .A1(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .A2(_0804_),
    .A3(_0805_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q ),
    .X(\Inst_RegFile_switch_matrix.W1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1901_ (.A0(net92),
    .A1(net687),
    .A2(net107),
    .A3(net421),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q ),
    .X(\Inst_RegFile_switch_matrix.S4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _1902_ (.A0(net91),
    .A1(net686),
    .A2(net110),
    .A3(net653),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q ),
    .X(\Inst_RegFile_switch_matrix.S4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1903_ (.A0(net778),
    .A1(net94),
    .A2(net109),
    .A3(net660),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q ),
    .X(\Inst_RegFile_switch_matrix.S4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1904_ (.A0(net22),
    .A1(net108),
    .A2(net93),
    .A3(net673),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q ),
    .X(\Inst_RegFile_switch_matrix.S4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1905_ (.A0(net641),
    .A1(_0437_),
    .A2(\Inst_RegFile_switch_matrix.E2BEG2 ),
    .A3(_0803_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q ),
    .X(\Inst_RegFile_switch_matrix.S1BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1906_ (.A0(net635),
    .A1(net685),
    .A2(\Inst_RegFile_switch_matrix.E2BEG1 ),
    .A3(net397),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q ),
    .X(\Inst_RegFile_switch_matrix.S1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1907_ (.A0(net666),
    .A1(_0582_),
    .A2(\Inst_RegFile_switch_matrix.E2BEG0 ),
    .A3(_0158_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q ),
    .X(\Inst_RegFile_switch_matrix.S1BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1908_ (.A0(net680),
    .A1(\Inst_RegFile_switch_matrix.E2BEG3 ),
    .A2(_0804_),
    .A3(_0805_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q ),
    .X(\Inst_RegFile_switch_matrix.S1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1909_ (.A0(net637),
    .A1(_0437_),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG2 ),
    .A3(_0803_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q ),
    .X(\Inst_RegFile_switch_matrix.E1BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1910_ (.A0(net666),
    .A1(net685),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG1 ),
    .A3(net394),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q ),
    .X(\Inst_RegFile_switch_matrix.E1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1911_ (.A0(net676),
    .A1(_0582_),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG0 ),
    .A3(_0158_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q ),
    .X(\Inst_RegFile_switch_matrix.E1BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1912_ (.A0(net421),
    .A1(\Inst_RegFile_switch_matrix.JN2BEG3 ),
    .A2(_0804_),
    .A3(_0805_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q ),
    .X(\Inst_RegFile_switch_matrix.E1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1913_ (.A0(net64),
    .A1(net79),
    .A2(net687),
    .A3(net409),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q ),
    .X(\Inst_RegFile_switch_matrix.N4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _1914_ (.A0(net63),
    .A1(net686),
    .A2(net82),
    .A3(net415),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q ),
    .X(\Inst_RegFile_switch_matrix.N4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1915_ (.A0(net66),
    .A1(net81),
    .A2(net778),
    .A3(net665),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q ),
    .X(\Inst_RegFile_switch_matrix.N4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1916_ (.A0(net65),
    .A1(net80),
    .A2(net777),
    .A3(net676),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q ),
    .X(\Inst_RegFile_switch_matrix.N4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1917_ (.A0(net664),
    .A1(_0437_),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG2 ),
    .A3(_0803_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q ),
    .X(\Inst_RegFile_switch_matrix.N1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _1918_ (.A0(net676),
    .A1(net685),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG1 ),
    .A3(net394),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q ),
    .X(\Inst_RegFile_switch_matrix.N1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1919_ (.A0(net645),
    .A1(_0582_),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG0 ),
    .A3(_0158_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q ),
    .X(\Inst_RegFile_switch_matrix.N1BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1920_ (.A0(net423),
    .A1(\Inst_RegFile_switch_matrix.JW2BEG3 ),
    .A2(_0804_),
    .A3(_0805_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q ),
    .X(\Inst_RegFile_switch_matrix.N1BEG0 ));
 sky130_fd_sc_hd__mux2_1 _1921_ (.A0(\Inst_RegFile_switch_matrix.JS2BEG7 ),
    .A1(\Inst_RegFile_switch_matrix.JW2BEG7 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ),
    .X(_0806_));
 sky130_fd_sc_hd__mux2_1 _1922_ (.A0(_0740_),
    .A1(\Inst_RegFile_switch_matrix.JN2BEG7 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ),
    .X(_0807_));
 sky130_fd_sc_hd__mux2_1 _1923_ (.A0(_0807_),
    .A1(_0806_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q ),
    .X(_0808_));
 sky130_fd_sc_hd__mux4_2 _1924_ (.A0(net63),
    .A1(net91),
    .A2(_1031_),
    .A3(_0148_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q ),
    .X(_0809_));
 sky130_fd_sc_hd__mux2_4 _1925_ (.A0(_0809_),
    .A1(_0808_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q ),
    .X(_0810_));
 sky130_fd_sc_hd__mux4_1 _1926_ (.A0(net71),
    .A1(net127),
    .A2(net99),
    .A3(\Inst_RegFile_switch_matrix.JW2BEG4 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q ),
    .X(_0811_));
 sky130_fd_sc_hd__and2b_1 _1927_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q ),
    .B(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__a21o_1 _1928_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(_0804_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ),
    .X(_0813_));
 sky130_fd_sc_hd__nor2_1 _1929_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q ),
    .B(_0213_),
    .Y(_0814_));
 sky130_fd_sc_hd__o21a_1 _1930_ (.A1(net135),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q ),
    .X(_0815_));
 sky130_fd_sc_hd__o21ai_1 _1931_ (.A1(_1019_),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG2 ),
    .B1(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__o21ba_1 _1932_ (.A1(net79),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q ),
    .X(_0817_));
 sky130_fd_sc_hd__o21ai_1 _1933_ (.A1(net111),
    .A2(_1019_),
    .B1(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__a31o_1 _1934_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(_0816_),
    .A3(_0818_),
    .B1(_0814_),
    .X(_0819_));
 sky130_fd_sc_hd__o2bb2a_1 _1935_ (.A1_N(\Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ),
    .A2_N(_0819_),
    .B1(_0813_),
    .B2(_0812_),
    .X(_0820_));
 sky130_fd_sc_hd__a2bb2o_1 _1936_ (.A1_N(_0812_),
    .A2_N(_0813_),
    .B1(_0819_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ),
    .X(_0821_));
 sky130_fd_sc_hd__nand2_1 _1937_ (.A(_0810_),
    .B(_0820_),
    .Y(_0822_));
 sky130_fd_sc_hd__mux4_1 _1938_ (.A0(net76),
    .A1(net18),
    .A2(net104),
    .A3(net132),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q ),
    .X(_0823_));
 sky130_fd_sc_hd__a21o_1 _1939_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q ),
    .A2(_0823_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ),
    .X(_0824_));
 sky130_fd_sc_hd__a21oi_2 _1940_ (.A1(_1018_),
    .A2(_0708_),
    .B1(_0824_),
    .Y(_0825_));
 sky130_fd_sc_hd__mux4_2 _1941_ (.A0(net84),
    .A1(net24),
    .A2(net108),
    .A3(\Inst_RegFile_switch_matrix.JS2BEG2 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q ),
    .X(_0826_));
 sky130_fd_sc_hd__or2_1 _1942_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q ),
    .B(_0726_),
    .X(_0827_));
 sky130_fd_sc_hd__o21ai_2 _1943_ (.A1(_1018_),
    .A2(_0826_),
    .B1(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__a21oi_4 _1944_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ),
    .A2(_0828_),
    .B1(_0825_),
    .Y(_0829_));
 sky130_fd_sc_hd__a21o_2 _1945_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ),
    .A2(_0828_),
    .B1(_0825_),
    .X(_0830_));
 sky130_fd_sc_hd__nor2_2 _1946_ (.A(_0822_),
    .B(_0829_),
    .Y(_0831_));
 sky130_fd_sc_hd__o21ba_1 _1947_ (.A1(_0667_),
    .A2(_0671_),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_0832_));
 sky130_fd_sc_hd__a21bo_1 _1948_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG0 ),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ),
    .X(_0833_));
 sky130_fd_sc_hd__mux2_1 _1949_ (.A0(_0401_),
    .A1(\Inst_RegFile_switch_matrix.JN2BEG0 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_0834_));
 sky130_fd_sc_hd__o22a_1 _1950_ (.A1(_0832_),
    .A2(_0833_),
    .B1(_0834_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ),
    .X(_0835_));
 sky130_fd_sc_hd__mux4_2 _1951_ (.A0(net73),
    .A1(net129),
    .A2(net15),
    .A3(\Inst_RegFile_switch_matrix.E2BEG4 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q ),
    .X(_0836_));
 sky130_fd_sc_hd__mux4_2 _1952_ (.A0(net66),
    .A1(net94),
    .A2(_0836_),
    .A3(_0823_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ),
    .X(_0837_));
 sky130_fd_sc_hd__mux2_4 _1953_ (.A0(_0837_),
    .A1(_0835_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q ),
    .X(_0838_));
 sky130_fd_sc_hd__a211oi_1 _1954_ (.A1(_0987_),
    .A2(_0614_),
    .B1(_0611_),
    .C1(_1016_),
    .Y(_0839_));
 sky130_fd_sc_hd__o21ai_1 _1955_ (.A1(net139),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q ),
    .Y(_0840_));
 sky130_fd_sc_hd__mux2_1 _1956_ (.A0(net8),
    .A1(net114),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ),
    .X(_0841_));
 sky130_fd_sc_hd__inv_1 _1957_ (.A(_0841_),
    .Y(_0842_));
 sky130_fd_sc_hd__o221a_1 _1958_ (.A1(_0839_),
    .A2(_0840_),
    .B1(_0842_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q ),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .X(_0843_));
 sky130_fd_sc_hd__o21ai_1 _1959_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(_0772_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ),
    .Y(_0844_));
 sky130_fd_sc_hd__o311a_1 _1960_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0559_),
    .A3(_0561_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q ),
    .C1(_0557_),
    .X(_0845_));
 sky130_fd_sc_hd__o21ai_1 _1961_ (.A1(net133),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q ),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q ),
    .Y(_0846_));
 sky130_fd_sc_hd__mux2_1 _1962_ (.A0(net19),
    .A1(net105),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q ),
    .X(_0847_));
 sky130_fd_sc_hd__inv_1 _1963_ (.A(_0847_),
    .Y(_0848_));
 sky130_fd_sc_hd__o221a_1 _1964_ (.A1(_0845_),
    .A2(_0846_),
    .B1(_0848_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q ),
    .C1(_1015_),
    .X(_0849_));
 sky130_fd_sc_hd__mux4_1 _1965_ (.A0(net78),
    .A1(net20),
    .A2(net106),
    .A3(net134),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q ),
    .X(_0850_));
 sky130_fd_sc_hd__nor2_1 _1966_ (.A(_1015_),
    .B(_0850_),
    .Y(_0851_));
 sky130_fd_sc_hd__o32a_1 _1967_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ),
    .A2(_0849_),
    .A3(_0851_),
    .B1(_0843_),
    .B2(_0844_),
    .X(_0852_));
 sky130_fd_sc_hd__nand2_8 _1968_ (.A(_0838_),
    .B(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__mux2_1 _1969_ (.A0(_0719_),
    .A1(_0836_),
    .S(_1017_),
    .X(_0854_));
 sky130_fd_sc_hd__a21bo_1 _1970_ (.A1(_1017_),
    .A2(_0791_),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ),
    .X(_0855_));
 sky130_fd_sc_hd__a21o_1 _1971_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(_0805_),
    .B1(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__o21ai_4 _1972_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ),
    .A2(_0854_),
    .B1(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__o21a_2 _1973_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ),
    .A2(_0854_),
    .B1(_0856_),
    .X(_0858_));
 sky130_fd_sc_hd__nor2_8 _1974_ (.A(_0853_),
    .B(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__nand2_4 _1975_ (.A(_0859_),
    .B(_0831_),
    .Y(_0860_));
 sky130_fd_sc_hd__mux2_1 _1976_ (.A0(net133),
    .A1(\Inst_RegFile_switch_matrix.JN2BEG3 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q ),
    .X(_0861_));
 sky130_fd_sc_hd__inv_1 _1977_ (.A(_0861_),
    .Y(_0862_));
 sky130_fd_sc_hd__mux2_1 _1978_ (.A0(net77),
    .A1(net105),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q ),
    .X(_0863_));
 sky130_fd_sc_hd__nor2_1 _1979_ (.A(\Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q ),
    .B(_0863_),
    .Y(_0864_));
 sky130_fd_sc_hd__a211o_1 _1980_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q ),
    .A2(_0862_),
    .B1(_0864_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ),
    .X(_0865_));
 sky130_fd_sc_hd__mux4_1 _1981_ (.A0(net78),
    .A1(net20),
    .A2(net106),
    .A3(net134),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q ),
    .X(_0866_));
 sky130_fd_sc_hd__a21oi_1 _1982_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ),
    .A2(_0866_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q ),
    .Y(_0867_));
 sky130_fd_sc_hd__mux2_1 _1983_ (.A0(_0767_),
    .A1(_0803_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ),
    .X(_0868_));
 sky130_fd_sc_hd__o2bb2a_2 _1984_ (.A1_N(_0865_),
    .A2_N(_0867_),
    .B1(_0868_),
    .B2(_1014_),
    .X(_0869_));
 sky130_fd_sc_hd__mux2_1 _1985_ (.A0(net599),
    .A1(net814),
    .S(_0860_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _1986_ (.A0(net420),
    .A1(_0718_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ),
    .X(_0870_));
 sky130_fd_sc_hd__mux4_1 _1987_ (.A0(net25),
    .A1(net126),
    .A2(net109),
    .A3(\Inst_RegFile_switch_matrix.E2BEG1 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q ),
    .X(_0871_));
 sky130_fd_sc_hd__mux2_1 _1988_ (.A0(_0788_),
    .A1(_0871_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ),
    .X(_0872_));
 sky130_fd_sc_hd__mux2_1 _1989_ (.A0(_0870_),
    .A1(_0872_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q ),
    .X(_0873_));
 sky130_fd_sc_hd__mux2_1 _1990_ (.A0(net615),
    .A1(net833),
    .S(_0860_),
    .X(_0001_));
 sky130_fd_sc_hd__mux4_1 _1991_ (.A0(net80),
    .A1(net686),
    .A2(net777),
    .A3(\Inst_RegFile_switch_matrix.JS2BEG1 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q ),
    .X(_0874_));
 sky130_fd_sc_hd__mux4_1 _1992_ (.A0(_0707_),
    .A1(_0723_),
    .A2(_0437_),
    .A3(_0874_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q ),
    .X(_0875_));
 sky130_fd_sc_hd__mux2_4 _1993_ (.A0(net620),
    .A1(net909),
    .S(_0860_),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_1 _1994_ (.A0(net107),
    .A1(\Inst_RegFile_switch_matrix.JW2BEG1 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ),
    .X(_0876_));
 sky130_fd_sc_hd__mux2_1 _1995_ (.A0(net79),
    .A1(net778),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ),
    .X(_0877_));
 sky130_fd_sc_hd__inv_1 _1996_ (.A(_0877_),
    .Y(_0878_));
 sky130_fd_sc_hd__o21ai_1 _1997_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q ),
    .A2(_0878_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ),
    .Y(_0879_));
 sky130_fd_sc_hd__a21o_1 _1998_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q ),
    .A2(_0876_),
    .B1(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__or2_1 _1999_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ),
    .B(_0740_),
    .X(_0881_));
 sky130_fd_sc_hd__mux4_1 _2000_ (.A0(net71),
    .A1(net13),
    .A2(net99),
    .A3(\Inst_RegFile_switch_matrix.JW2BEG3 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q ),
    .X(_0882_));
 sky130_fd_sc_hd__mux4_1 _2001_ (.A0(net72),
    .A1(net14),
    .A2(net100),
    .A3(net128),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q ),
    .X(_0883_));
 sky130_fd_sc_hd__inv_1 _2002_ (.A(_0883_),
    .Y(_0884_));
 sky130_fd_sc_hd__a21oi_1 _2003_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ),
    .A2(_0884_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q ),
    .Y(_0885_));
 sky130_fd_sc_hd__o21a_1 _2004_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ),
    .A2(_0882_),
    .B1(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__a31o_1 _2005_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q ),
    .A2(_0880_),
    .A3(_0881_),
    .B1(_0886_),
    .X(_0887_));
 sky130_fd_sc_hd__mux2_1 _2006_ (.A0(net611),
    .A1(net866),
    .S(_0860_),
    .X(_0003_));
 sky130_fd_sc_hd__nand2b_4 _2007_ (.A_N(_0852_),
    .B(_0838_),
    .Y(_0888_));
 sky130_fd_sc_hd__nor2_8 _2008_ (.A(_0858_),
    .B(_0888_),
    .Y(_0889_));
 sky130_fd_sc_hd__nand2_8 _2009_ (.A(_0831_),
    .B(_0889_),
    .Y(_0890_));
 sky130_fd_sc_hd__mux2_1 _2010_ (.A0(net599),
    .A1(net829),
    .S(_0890_),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_4 _2011_ (.A0(net615),
    .A1(net931),
    .S(_0890_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_4 _2012_ (.A0(net620),
    .A1(net932),
    .S(_0890_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_4 _2013_ (.A0(net611),
    .A1(net938),
    .S(_0890_),
    .X(_0007_));
 sky130_fd_sc_hd__nor2_8 _2014_ (.A(_0853_),
    .B(_0857_),
    .Y(_0891_));
 sky130_fd_sc_hd__nand2_4 _2015_ (.A(_0831_),
    .B(_0891_),
    .Y(_0892_));
 sky130_fd_sc_hd__mux2_1 _2016_ (.A0(net599),
    .A1(net826),
    .S(_0892_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_4 _2017_ (.A0(net615),
    .A1(net907),
    .S(_0892_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _2018_ (.A0(net620),
    .A1(net813),
    .S(_0892_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _2019_ (.A0(net611),
    .A1(net815),
    .S(_0892_),
    .X(_0011_));
 sky130_fd_sc_hd__nor2_8 _2020_ (.A(_0857_),
    .B(_0888_),
    .Y(_0893_));
 sky130_fd_sc_hd__nand2_2 _2021_ (.A(_0831_),
    .B(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__mux2_1 _2022_ (.A0(net599),
    .A1(net868),
    .S(_0894_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _2023_ (.A0(net615),
    .A1(net877),
    .S(_0894_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _2024_ (.A0(net620),
    .A1(net834),
    .S(_0894_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _2025_ (.A0(net611),
    .A1(net883),
    .S(_0894_),
    .X(_0015_));
 sky130_fd_sc_hd__nor2_2 _2026_ (.A(_0822_),
    .B(_0830_),
    .Y(_0895_));
 sky130_fd_sc_hd__nand2_8 _2027_ (.A(net593),
    .B(_0895_),
    .Y(_0896_));
 sky130_fd_sc_hd__mux2_4 _2028_ (.A0(net599),
    .A1(net902),
    .S(_0896_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_4 _2029_ (.A0(net615),
    .A1(net917),
    .S(_0896_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_4 _2030_ (.A0(net620),
    .A1(net905),
    .S(_0896_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_4 _2031_ (.A0(net611),
    .A1(net900),
    .S(_0896_),
    .X(_0019_));
 sky130_fd_sc_hd__or2_4 _2032_ (.A(_0810_),
    .B(_0820_),
    .X(_0897_));
 sky130_fd_sc_hd__nor2_8 _2033_ (.A(_0829_),
    .B(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__nand2_4 _2034_ (.A(_0891_),
    .B(_0898_),
    .Y(_0899_));
 sky130_fd_sc_hd__mux2_1 _2035_ (.A0(net600),
    .A1(net841),
    .S(_0899_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_2 _2036_ (.A0(net617),
    .A1(net923),
    .S(_0899_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_2 _2037_ (.A0(net621),
    .A1(net901),
    .S(_0899_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_2 _2038_ (.A0(net612),
    .A1(net885),
    .S(_0899_),
    .X(_0023_));
 sky130_fd_sc_hd__nand2_4 _2039_ (.A(_0891_),
    .B(_0895_),
    .Y(_0900_));
 sky130_fd_sc_hd__mux2_1 _2040_ (.A0(net599),
    .A1(net843),
    .S(_0900_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _2041_ (.A0(net615),
    .A1(net832),
    .S(_0900_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _2042_ (.A0(net620),
    .A1(net850),
    .S(_0900_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _2043_ (.A0(net611),
    .A1(net821),
    .S(_0900_),
    .X(_0027_));
 sky130_fd_sc_hd__or2_4 _2044_ (.A(_0821_),
    .B(_0810_),
    .X(_0901_));
 sky130_fd_sc_hd__nor2_8 _2045_ (.A(_0901_),
    .B(_0829_),
    .Y(_0902_));
 sky130_fd_sc_hd__nand2_4 _2046_ (.A(_0889_),
    .B(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__mux2_1 _2047_ (.A0(net600),
    .A1(net879),
    .S(_0903_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _2048_ (.A0(net616),
    .A1(net853),
    .S(_0903_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _2049_ (.A0(net621),
    .A1(net864),
    .S(_0903_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _2050_ (.A0(net614),
    .A1(net872),
    .S(_0903_),
    .X(_0031_));
 sky130_fd_sc_hd__nor2_8 _2051_ (.A(_0830_),
    .B(_0901_),
    .Y(_0904_));
 sky130_fd_sc_hd__nand2_4 _2052_ (.A(_0889_),
    .B(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hd__mux2_1 _2053_ (.A0(net602),
    .A1(net847),
    .S(_0905_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _2054_ (.A0(net618),
    .A1(net846),
    .S(_0905_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _2055_ (.A0(net623),
    .A1(net836),
    .S(_0905_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _2056_ (.A0(net611),
    .A1(net867),
    .S(_0905_),
    .X(_0035_));
 sky130_fd_sc_hd__nand2_1 _2057_ (.A(_0810_),
    .B(_0821_),
    .Y(_0906_));
 sky130_fd_sc_hd__nor2_2 _2058_ (.A(_0829_),
    .B(_0906_),
    .Y(_0907_));
 sky130_fd_sc_hd__nand2_4 _2059_ (.A(_0889_),
    .B(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__mux2_1 _2060_ (.A0(net601),
    .A1(net844),
    .S(_0908_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _2061_ (.A0(net617),
    .A1(net840),
    .S(_0908_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _2062_ (.A0(net623),
    .A1(net889),
    .S(_0908_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _2063_ (.A0(net613),
    .A1(net887),
    .S(_0908_),
    .X(_0039_));
 sky130_fd_sc_hd__nor2_2 _2064_ (.A(_0830_),
    .B(_0906_),
    .Y(_0909_));
 sky130_fd_sc_hd__nand2_4 _2065_ (.A(_0891_),
    .B(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__mux2_1 _2066_ (.A0(net601),
    .A1(net862),
    .S(_0910_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_4 _2067_ (.A0(net617),
    .A1(net919),
    .S(_0910_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_4 _2068_ (.A0(net622),
    .A1(net935),
    .S(_0910_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_4 _2069_ (.A0(net612),
    .A1(net927),
    .S(_0910_),
    .X(_0043_));
 sky130_fd_sc_hd__nand2_2 _2070_ (.A(_0893_),
    .B(_0909_),
    .Y(_0911_));
 sky130_fd_sc_hd__mux2_1 _2071_ (.A0(net601),
    .A1(net869),
    .S(_0911_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _2072_ (.A0(net617),
    .A1(net937),
    .S(_0911_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _2073_ (.A0(net622),
    .A1(net863),
    .S(_0911_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _2074_ (.A0(net612),
    .A1(net892),
    .S(_0911_),
    .X(_0047_));
 sky130_fd_sc_hd__nand2_4 _2075_ (.A(_0891_),
    .B(_0904_),
    .Y(_0912_));
 sky130_fd_sc_hd__mux2_2 _2076_ (.A0(net599),
    .A1(net891),
    .S(_0912_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_2 _2077_ (.A0(net615),
    .A1(net904),
    .S(_0912_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_2 _2078_ (.A0(net620),
    .A1(net884),
    .S(_0912_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_2 _2079_ (.A0(_0887_),
    .A1(net895),
    .S(_0912_),
    .X(_0051_));
 sky130_fd_sc_hd__nand2_4 _2080_ (.A(_0893_),
    .B(_0904_),
    .Y(_0913_));
 sky130_fd_sc_hd__mux2_1 _2081_ (.A0(net599),
    .A1(net831),
    .S(_0913_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _2082_ (.A0(net615),
    .A1(net857),
    .S(_0913_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _2083_ (.A0(net620),
    .A1(net859),
    .S(_0913_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _2084_ (.A0(_0887_),
    .A1(net817),
    .S(_0913_),
    .X(_0055_));
 sky130_fd_sc_hd__nand2_8 _2085_ (.A(_0859_),
    .B(_0907_),
    .Y(_0914_));
 sky130_fd_sc_hd__mux2_4 _2086_ (.A0(net602),
    .A1(net903),
    .S(_0914_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_4 _2087_ (.A0(net618),
    .A1(net911),
    .S(_0914_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_4 _2088_ (.A0(net622),
    .A1(net906),
    .S(_0914_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_4 _2089_ (.A0(net613),
    .A1(net934),
    .S(_0914_),
    .X(_0059_));
 sky130_fd_sc_hd__nand2_8 _2090_ (.A(_0907_),
    .B(_0891_),
    .Y(_0915_));
 sky130_fd_sc_hd__mux2_1 _2091_ (.A0(net601),
    .A1(net816),
    .S(_0915_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_4 _2092_ (.A0(net617),
    .A1(net929),
    .S(_0915_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_4 _2093_ (.A0(net622),
    .A1(net894),
    .S(_0915_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_4 _2094_ (.A0(net613),
    .A1(net910),
    .S(_0915_),
    .X(_0063_));
 sky130_fd_sc_hd__nand2_4 _2095_ (.A(_0898_),
    .B(_0889_),
    .Y(_0916_));
 sky130_fd_sc_hd__mux2_1 _2096_ (.A0(net600),
    .A1(net830),
    .S(_0916_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _2097_ (.A0(net617),
    .A1(net873),
    .S(_0916_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_2 _2098_ (.A0(net621),
    .A1(net908),
    .S(_0916_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _2099_ (.A0(net612),
    .A1(net871),
    .S(_0916_),
    .X(_0067_));
 sky130_fd_sc_hd__nand2_4 _2100_ (.A(_0859_),
    .B(_0909_),
    .Y(_0917_));
 sky130_fd_sc_hd__mux2_1 _2101_ (.A0(net600),
    .A1(net835),
    .S(_0917_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _2102_ (.A0(net616),
    .A1(net827),
    .S(_0917_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_4 _2103_ (.A0(net621),
    .A1(net897),
    .S(_0917_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _2104_ (.A0(net612),
    .A1(net849),
    .S(_0917_),
    .X(_0071_));
 sky130_fd_sc_hd__nand2_4 _2105_ (.A(_0889_),
    .B(_0909_),
    .Y(_0918_));
 sky130_fd_sc_hd__mux2_1 _2106_ (.A0(net600),
    .A1(net855),
    .S(_0918_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _2107_ (.A0(net616),
    .A1(net882),
    .S(_0918_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_4 _2108_ (.A0(net621),
    .A1(net926),
    .S(_0918_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _2109_ (.A0(net612),
    .A1(net865),
    .S(_0918_),
    .X(_0075_));
 sky130_fd_sc_hd__nand2_2 _2110_ (.A(_0893_),
    .B(_0907_),
    .Y(_0919_));
 sky130_fd_sc_hd__mux2_1 _2111_ (.A0(net601),
    .A1(net861),
    .S(_0919_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _2112_ (.A0(net617),
    .A1(net886),
    .S(_0919_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _2113_ (.A0(net622),
    .A1(net842),
    .S(_0919_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _2114_ (.A0(net613),
    .A1(net845),
    .S(_0919_),
    .X(_0079_));
 sky130_fd_sc_hd__nand2_4 _2115_ (.A(_0889_),
    .B(_0895_),
    .Y(_0920_));
 sky130_fd_sc_hd__mux2_1 _2116_ (.A0(net599),
    .A1(net838),
    .S(_0920_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _2117_ (.A0(net615),
    .A1(net860),
    .S(_0920_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _2118_ (.A0(net620),
    .A1(net878),
    .S(_0920_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _2119_ (.A0(net611),
    .A1(net876),
    .S(_0920_),
    .X(_0083_));
 sky130_fd_sc_hd__nand2_4 _2120_ (.A(_0893_),
    .B(_0895_),
    .Y(_0921_));
 sky130_fd_sc_hd__mux2_1 _2121_ (.A0(net599),
    .A1(net852),
    .S(_0921_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_4 _2122_ (.A0(net615),
    .A1(net928),
    .S(_0921_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _2123_ (.A0(net620),
    .A1(net858),
    .S(_0921_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_2 _2124_ (.A0(net611),
    .A1(net912),
    .S(_0921_),
    .X(_0087_));
 sky130_fd_sc_hd__nand2_4 _2125_ (.A(_0893_),
    .B(_0898_),
    .Y(_0922_));
 sky130_fd_sc_hd__mux2_1 _2126_ (.A0(net600),
    .A1(net848),
    .S(_0922_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_2 _2127_ (.A0(net616),
    .A1(net924),
    .S(_0922_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_2 _2128_ (.A0(net621),
    .A1(net913),
    .S(_0922_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_2 _2129_ (.A0(net612),
    .A1(net921),
    .S(_0922_),
    .X(_0091_));
 sky130_fd_sc_hd__nor2_8 _2130_ (.A(_0830_),
    .B(_0897_),
    .Y(_0923_));
 sky130_fd_sc_hd__nand2_2 _2131_ (.A(_0859_),
    .B(_0923_),
    .Y(_0924_));
 sky130_fd_sc_hd__mux2_1 _2132_ (.A0(net601),
    .A1(net819),
    .S(_0924_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _2133_ (.A0(net617),
    .A1(net828),
    .S(_0924_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _2134_ (.A0(net622),
    .A1(net825),
    .S(_0924_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _2135_ (.A0(net613),
    .A1(net820),
    .S(_0924_),
    .X(_0095_));
 sky130_fd_sc_hd__nand2_2 _2136_ (.A(_0889_),
    .B(_0923_),
    .Y(_0925_));
 sky130_fd_sc_hd__mux2_1 _2137_ (.A0(net601),
    .A1(net837),
    .S(_0925_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _2138_ (.A0(net617),
    .A1(net875),
    .S(_0925_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _2139_ (.A0(net622),
    .A1(net856),
    .S(_0925_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _2140_ (.A0(net613),
    .A1(net881),
    .S(_0925_),
    .X(_0099_));
 sky130_fd_sc_hd__nand2_4 _2141_ (.A(_0891_),
    .B(_0923_),
    .Y(_0926_));
 sky130_fd_sc_hd__mux2_1 _2142_ (.A0(net601),
    .A1(net822),
    .S(_0926_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _2143_ (.A0(net616),
    .A1(net818),
    .S(_0926_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _2144_ (.A0(net622),
    .A1(net824),
    .S(_0926_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _2145_ (.A0(net612),
    .A1(net854),
    .S(_0926_),
    .X(_0103_));
 sky130_fd_sc_hd__nand2_4 _2146_ (.A(_0893_),
    .B(_0923_),
    .Y(_0927_));
 sky130_fd_sc_hd__mux2_2 _2147_ (.A0(net601),
    .A1(net933),
    .S(_0927_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_2 _2148_ (.A0(net616),
    .A1(net925),
    .S(_0927_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_2 _2149_ (.A0(net622),
    .A1(net915),
    .S(_0927_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_2 _2150_ (.A0(net612),
    .A1(net936),
    .S(_0927_),
    .X(_0107_));
 sky130_fd_sc_hd__nand2_4 _2151_ (.A(_0859_),
    .B(_0902_),
    .Y(_0928_));
 sky130_fd_sc_hd__mux2_1 _2152_ (.A0(net600),
    .A1(net811),
    .S(_0928_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_2 _2153_ (.A0(net616),
    .A1(net896),
    .S(_0928_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_2 _2154_ (.A0(net621),
    .A1(net914),
    .S(_0928_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_2 _2155_ (.A0(net614),
    .A1(net920),
    .S(_0928_),
    .X(_0111_));
 sky130_fd_sc_hd__nand2_4 _2156_ (.A(_0859_),
    .B(_0898_),
    .Y(_0929_));
 sky130_fd_sc_hd__mux2_1 _2157_ (.A0(net600),
    .A1(net812),
    .S(_0929_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_4 _2158_ (.A0(net616),
    .A1(net898),
    .S(_0929_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_2 _2159_ (.A0(net621),
    .A1(net916),
    .S(_0929_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_2 _2160_ (.A0(net612),
    .A1(net890),
    .S(_0929_),
    .X(_0115_));
 sky130_fd_sc_hd__nand2_4 _2161_ (.A(_0891_),
    .B(_0902_),
    .Y(_0930_));
 sky130_fd_sc_hd__mux2_1 _2162_ (.A0(net600),
    .A1(net880),
    .S(_0930_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_2 _2163_ (.A0(net616),
    .A1(net899),
    .S(_0930_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_2 _2164_ (.A0(net621),
    .A1(net918),
    .S(_0930_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_2 _2165_ (.A0(net614),
    .A1(net922),
    .S(_0930_),
    .X(_0119_));
 sky130_fd_sc_hd__nand2_4 _2166_ (.A(_0893_),
    .B(_0902_),
    .Y(_0931_));
 sky130_fd_sc_hd__mux2_1 _2167_ (.A0(net600),
    .A1(net893),
    .S(_0931_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _2168_ (.A0(net616),
    .A1(net870),
    .S(_0931_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _2169_ (.A0(net621),
    .A1(net874),
    .S(_0931_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _2170_ (.A0(net614),
    .A1(net839),
    .S(_0931_),
    .X(_0123_));
 sky130_fd_sc_hd__nand2_4 _2171_ (.A(_0859_),
    .B(_0904_),
    .Y(_0932_));
 sky130_fd_sc_hd__mux2_2 _2172_ (.A0(net602),
    .A1(net930),
    .S(_0932_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _2173_ (.A0(net618),
    .A1(net851),
    .S(_0932_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _2174_ (.A0(net623),
    .A1(net823),
    .S(_0932_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _2175_ (.A0(net611),
    .A1(net888),
    .S(_0932_),
    .X(_0127_));
 sky130_fd_sc_hd__dfxtp_1 _2176_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0000_),
    .Q(\Inst_RegFile_32x4.mem[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2177_ (.CLK(clknet_4_1_0_UserCLK_regs),
    .D(_0001_),
    .Q(\Inst_RegFile_32x4.mem[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2178_ (.CLK(clknet_4_5_0_UserCLK_regs),
    .D(_0002_),
    .Q(\Inst_RegFile_32x4.mem[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2179_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0003_),
    .Q(\Inst_RegFile_32x4.mem[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2180_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0004_),
    .Q(\Inst_RegFile_32x4.mem[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2181_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0005_),
    .Q(\Inst_RegFile_32x4.mem[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2182_ (.CLK(clknet_4_5_0_UserCLK_regs),
    .D(_0006_),
    .Q(\Inst_RegFile_32x4.mem[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2183_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0007_),
    .Q(\Inst_RegFile_32x4.mem[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2184_ (.CLK(clknet_4_1_0_UserCLK_regs),
    .D(_0008_),
    .Q(\Inst_RegFile_32x4.mem[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2185_ (.CLK(clknet_4_1_0_UserCLK_regs),
    .D(_0009_),
    .Q(\Inst_RegFile_32x4.mem[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2186_ (.CLK(clknet_4_4_0_UserCLK_regs),
    .D(_0010_),
    .Q(\Inst_RegFile_32x4.mem[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2187_ (.CLK(clknet_4_4_0_UserCLK_regs),
    .D(_0011_),
    .Q(\Inst_RegFile_32x4.mem[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2188_ (.CLK(clknet_4_1_0_UserCLK_regs),
    .D(_0012_),
    .Q(\Inst_RegFile_32x4.mem[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2189_ (.CLK(clknet_4_1_0_UserCLK_regs),
    .D(_0013_),
    .Q(\Inst_RegFile_32x4.mem[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2190_ (.CLK(clknet_4_4_0_UserCLK_regs),
    .D(_0014_),
    .Q(\Inst_RegFile_32x4.mem[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2191_ (.CLK(clknet_4_4_0_UserCLK_regs),
    .D(_0015_),
    .Q(\Inst_RegFile_32x4.mem[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2192_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0016_),
    .Q(\Inst_RegFile_32x4.mem[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2193_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0017_),
    .Q(\Inst_RegFile_32x4.mem[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2194_ (.CLK(clknet_4_5_0_UserCLK_regs),
    .D(_0018_),
    .Q(\Inst_RegFile_32x4.mem[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2195_ (.CLK(clknet_4_5_0_UserCLK_regs),
    .D(_0019_),
    .Q(\Inst_RegFile_32x4.mem[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2196_ (.CLK(clknet_4_8_0_UserCLK_regs),
    .D(_0020_),
    .Q(\Inst_RegFile_32x4.mem[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2197_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0021_),
    .Q(\Inst_RegFile_32x4.mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2198_ (.CLK(clknet_4_8_0_UserCLK_regs),
    .D(_0022_),
    .Q(\Inst_RegFile_32x4.mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2199_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0023_),
    .Q(\Inst_RegFile_32x4.mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2200_ (.CLK(clknet_4_1_0_UserCLK_regs),
    .D(_0024_),
    .Q(\Inst_RegFile_32x4.mem[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2201_ (.CLK(clknet_4_1_0_UserCLK_regs),
    .D(_0025_),
    .Q(\Inst_RegFile_32x4.mem[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2202_ (.CLK(clknet_4_5_0_UserCLK_regs),
    .D(_0026_),
    .Q(\Inst_RegFile_32x4.mem[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2203_ (.CLK(clknet_4_4_0_UserCLK_regs),
    .D(_0027_),
    .Q(\Inst_RegFile_32x4.mem[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2204_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(_0028_),
    .Q(\Inst_RegFile_32x4.mem[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2205_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(_0029_),
    .Q(\Inst_RegFile_32x4.mem[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2206_ (.CLK(clknet_4_9_0_UserCLK_regs),
    .D(_0030_),
    .Q(\Inst_RegFile_32x4.mem[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2207_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(_0031_),
    .Q(\Inst_RegFile_32x4.mem[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2208_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0032_),
    .Q(\Inst_RegFile_32x4.mem[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2209_ (.CLK(clknet_4_3_0_UserCLK_regs),
    .D(_0033_),
    .Q(\Inst_RegFile_32x4.mem[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2210_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0034_),
    .Q(\Inst_RegFile_32x4.mem[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2211_ (.CLK(clknet_4_3_0_UserCLK_regs),
    .D(_0035_),
    .Q(\Inst_RegFile_32x4.mem[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2212_ (.CLK(clknet_4_12_0_UserCLK_regs),
    .D(_0036_),
    .Q(\Inst_RegFile_32x4.mem[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2213_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0037_),
    .Q(\Inst_RegFile_32x4.mem[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2214_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0038_),
    .Q(\Inst_RegFile_32x4.mem[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2215_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0039_),
    .Q(\Inst_RegFile_32x4.mem[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2216_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0040_),
    .Q(\Inst_RegFile_32x4.mem[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2217_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0041_),
    .Q(\Inst_RegFile_32x4.mem[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2218_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0042_),
    .Q(\Inst_RegFile_32x4.mem[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2219_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0043_),
    .Q(\Inst_RegFile_32x4.mem[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2220_ (.CLK(clknet_4_9_0_UserCLK_regs),
    .D(_0044_),
    .Q(\Inst_RegFile_32x4.mem[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2221_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0045_),
    .Q(\Inst_RegFile_32x4.mem[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2222_ (.CLK(clknet_4_9_0_UserCLK_regs),
    .D(_0046_),
    .Q(\Inst_RegFile_32x4.mem[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2223_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0047_),
    .Q(\Inst_RegFile_32x4.mem[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2224_ (.CLK(clknet_4_6_0_UserCLK_regs),
    .D(_0048_),
    .Q(\Inst_RegFile_32x4.mem[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2225_ (.CLK(clknet_4_6_0_UserCLK_regs),
    .D(_0049_),
    .Q(\Inst_RegFile_32x4.mem[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2226_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0050_),
    .Q(\Inst_RegFile_32x4.mem[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2227_ (.CLK(clknet_4_6_0_UserCLK_regs),
    .D(_0051_),
    .Q(\Inst_RegFile_32x4.mem[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2228_ (.CLK(clknet_4_6_0_UserCLK_regs),
    .D(_0052_),
    .Q(\Inst_RegFile_32x4.mem[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2229_ (.CLK(clknet_4_6_0_UserCLK_regs),
    .D(_0053_),
    .Q(\Inst_RegFile_32x4.mem[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2230_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0054_),
    .Q(\Inst_RegFile_32x4.mem[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2231_ (.CLK(clknet_4_6_0_UserCLK_regs),
    .D(_0055_),
    .Q(\Inst_RegFile_32x4.mem[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2232_ (.CLK(clknet_4_12_0_UserCLK_regs),
    .D(_0056_),
    .Q(\Inst_RegFile_32x4.mem[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2233_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0057_),
    .Q(\Inst_RegFile_32x4.mem[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2234_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0058_),
    .Q(\Inst_RegFile_32x4.mem[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2235_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0059_),
    .Q(\Inst_RegFile_32x4.mem[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2236_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0060_),
    .Q(\Inst_RegFile_32x4.mem[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2237_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0061_),
    .Q(\Inst_RegFile_32x4.mem[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2238_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0062_),
    .Q(\Inst_RegFile_32x4.mem[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2239_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0063_),
    .Q(\Inst_RegFile_32x4.mem[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2240_ (.CLK(clknet_4_8_0_UserCLK_regs),
    .D(_0064_),
    .Q(\Inst_RegFile_32x4.mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2241_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0065_),
    .Q(\Inst_RegFile_32x4.mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2242_ (.CLK(clknet_4_8_0_UserCLK_regs),
    .D(_0066_),
    .Q(\Inst_RegFile_32x4.mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2243_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0067_),
    .Q(\Inst_RegFile_32x4.mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2244_ (.CLK(clknet_4_9_0_UserCLK_regs),
    .D(_0068_),
    .Q(\Inst_RegFile_32x4.mem[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2245_ (.CLK(clknet_4_9_0_UserCLK_regs),
    .D(_0069_),
    .Q(\Inst_RegFile_32x4.mem[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2246_ (.CLK(clknet_4_9_0_UserCLK_regs),
    .D(_0070_),
    .Q(\Inst_RegFile_32x4.mem[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2247_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0071_),
    .Q(\Inst_RegFile_32x4.mem[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2248_ (.CLK(clknet_4_9_0_UserCLK_regs),
    .D(_0072_),
    .Q(\Inst_RegFile_32x4.mem[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2249_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0073_),
    .Q(\Inst_RegFile_32x4.mem[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2250_ (.CLK(clknet_4_9_0_UserCLK_regs),
    .D(_0074_),
    .Q(\Inst_RegFile_32x4.mem[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2251_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0075_),
    .Q(\Inst_RegFile_32x4.mem[21][3] ));
 sky130_fd_sc_hd__dlxtp_1 _2252_ (.D(net751),
    .GATE(net56),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2253_ (.D(net748),
    .GATE(net56),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2254_ (.D(net747),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2255_ (.D(net746),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2256_ (.D(net745),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2257_ (.D(net744),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2258_ (.D(net743),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2259_ (.D(net742),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2260_ (.D(net775),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2261_ (.D(net774),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2262_ (.D(net773),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2263_ (.D(net772),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2264_ (.D(net770),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2265_ (.D(net769),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2266_ (.D(net767),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2267_ (.D(net766),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2268_ (.D(net765),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2269_ (.D(net764),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2270_ (.D(net762),
    .GATE(net729),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2271_ (.D(net761),
    .GATE(net729),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2272_ (.D(net760),
    .GATE(net729),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2273_ (.D(net759),
    .GATE(net729),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2274_ (.D(net758),
    .GATE(net729),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2275_ (.D(net757),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2276_ (.D(net756),
    .GATE(net729),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2277_ (.D(net44),
    .GATE(net729),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2278_ (.D(net754),
    .GATE(net729),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2279_ (.D(net45),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2280_ (.D(net47),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2281_ (.D(net48),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2282_ (.D(net27),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2283_ (.D(net763),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2284_ (.D(net751),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2285_ (.D(net748),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2286_ (.D(net747),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2287_ (.D(net746),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2288_ (.D(net52),
    .GATE(net732),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2289_ (.D(net53),
    .GATE(net732),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2290_ (.D(net743),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2291_ (.D(net55),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2292_ (.D(net28),
    .GATE(net730),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2293_ (.D(net29),
    .GATE(net732),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2294_ (.D(net30),
    .GATE(net732),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2295_ (.D(net31),
    .GATE(net732),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2296_ (.D(net771),
    .GATE(net730),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2297_ (.D(net769),
    .GATE(net730),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2298_ (.D(net767),
    .GATE(net730),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2299_ (.D(net766),
    .GATE(net730),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2300_ (.D(net34),
    .GATE(net730),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2301_ (.D(net764),
    .GATE(net730),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2302_ (.D(net37),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2303_ (.D(net38),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2304_ (.D(net760),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2305_ (.D(net759),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2306_ (.D(net41),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2307_ (.D(net42),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2308_ (.D(net43),
    .GATE(net730),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2309_ (.D(net44),
    .GATE(net730),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2310_ (.D(net753),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2311_ (.D(net752),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2312_ (.D(net750),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2313_ (.D(net749),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2314_ (.D(net776),
    .GATE(net737),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2315_ (.D(net763),
    .GATE(net737),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2316_ (.D(net751),
    .GATE(net734),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2317_ (.D(net748),
    .GATE(net734),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2318_ (.D(net50),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2319_ (.D(net746),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2320_ (.D(net52),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2321_ (.D(net53),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2322_ (.D(net54),
    .GATE(net737),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2323_ (.D(net55),
    .GATE(net737),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2324_ (.D(net775),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2325_ (.D(net29),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2326_ (.D(net30),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2327_ (.D(net31),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2328_ (.D(net771),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2329_ (.D(net769),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2330_ (.D(net32),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2331_ (.D(net766),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2332_ (.D(net765),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2333_ (.D(net764),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2334_ (.D(net762),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2335_ (.D(net38),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2336_ (.D(net39),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2337_ (.D(net759),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2338_ (.D(net758),
    .GATE(net734),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2339_ (.D(net757),
    .GATE(net734),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2340_ (.D(net756),
    .GATE(net734),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2341_ (.D(net755),
    .GATE(net734),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2342_ (.D(net753),
    .GATE(net734),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2343_ (.D(net752),
    .GATE(net734),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2344_ (.D(net750),
    .GATE(net734),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2345_ (.D(net749),
    .GATE(net734),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2346_ (.D(net776),
    .GATE(net691),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2347_ (.D(net763),
    .GATE(net691),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2348_ (.D(net751),
    .GATE(net691),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2349_ (.D(net748),
    .GATE(net690),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2350_ (.D(net747),
    .GATE(net690),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2351_ (.D(net746),
    .GATE(net690),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2352_ (.D(net745),
    .GATE(net691),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2353_ (.D(net744),
    .GATE(net691),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2354_ (.D(net743),
    .GATE(net691),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2355_ (.D(net742),
    .GATE(net690),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2356_ (.D(net775),
    .GATE(net690),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2357_ (.D(net774),
    .GATE(net690),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2358_ (.D(net773),
    .GATE(net691),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2359_ (.D(net772),
    .GATE(net691),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2360_ (.D(net771),
    .GATE(net691),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2361_ (.D(net768),
    .GATE(net691),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2362_ (.D(net767),
    .GATE(net690),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2363_ (.D(net766),
    .GATE(net690),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2364_ (.D(net765),
    .GATE(net690),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2365_ (.D(net764),
    .GATE(net692),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2366_ (.D(net37),
    .GATE(net693),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2367_ (.D(net38),
    .GATE(net693),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2368_ (.D(net760),
    .GATE(net693),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2369_ (.D(net759),
    .GATE(net693),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2370_ (.D(net758),
    .GATE(net692),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2371_ (.D(net757),
    .GATE(net692),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2372_ (.D(net756),
    .GATE(net692),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2373_ (.D(net755),
    .GATE(net692),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2374_ (.D(net754),
    .GATE(net693),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2375_ (.D(net752),
    .GATE(net693),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2376_ (.D(net750),
    .GATE(net693),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2377_ (.D(net749),
    .GATE(net690),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2378_ (.D(net776),
    .GATE(net58),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2379_ (.D(net36),
    .GATE(net697),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2380_ (.D(net46),
    .GATE(net697),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2381_ (.D(net748),
    .GATE(net697),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2382_ (.D(net50),
    .GATE(net697),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2383_ (.D(net746),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2384_ (.D(net745),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2385_ (.D(net53),
    .GATE(net696),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2386_ (.D(net54),
    .GATE(net696),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2387_ (.D(net742),
    .GATE(net696),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2388_ (.D(net775),
    .GATE(net696),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2389_ (.D(net774),
    .GATE(net696),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2390_ (.D(net30),
    .GATE(net696),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2391_ (.D(net31),
    .GATE(net696),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2392_ (.D(net770),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2393_ (.D(net768),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2394_ (.D(net767),
    .GATE(net695),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2395_ (.D(net766),
    .GATE(net695),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2396_ (.D(net34),
    .GATE(net696),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2397_ (.D(net35),
    .GATE(net696),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2398_ (.D(net762),
    .GATE(net697),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2399_ (.D(net761),
    .GATE(net697),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2400_ (.D(net760),
    .GATE(net695),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2401_ (.D(net759),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2402_ (.D(net758),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2403_ (.D(net757),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2404_ (.D(net756),
    .GATE(net695),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2405_ (.D(net755),
    .GATE(net695),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2406_ (.D(net753),
    .GATE(net695),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2407_ (.D(net45),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2408_ (.D(net750),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2409_ (.D(net749),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2410_ (.D(net27),
    .GATE(net701),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2411_ (.D(net763),
    .GATE(net701),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2412_ (.D(net46),
    .GATE(net700),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2413_ (.D(net49),
    .GATE(net700),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2414_ (.D(net50),
    .GATE(net699),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2415_ (.D(net51),
    .GATE(net699),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2416_ (.D(net745),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2417_ (.D(net744),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2418_ (.D(net743),
    .GATE(net699),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2419_ (.D(net742),
    .GATE(net700),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2420_ (.D(net28),
    .GATE(net700),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2421_ (.D(net29),
    .GATE(net700),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2422_ (.D(net773),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2423_ (.D(net772),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2424_ (.D(net770),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2425_ (.D(net768),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2426_ (.D(net767),
    .GATE(net700),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2427_ (.D(net33),
    .GATE(net700),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2428_ (.D(net34),
    .GATE(net700),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2429_ (.D(net35),
    .GATE(net701),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2430_ (.D(net762),
    .GATE(net701),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2431_ (.D(net761),
    .GATE(net701),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2432_ (.D(net760),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2433_ (.D(net759),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2434_ (.D(net758),
    .GATE(net699),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2435_ (.D(net757),
    .GATE(net699),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2436_ (.D(net756),
    .GATE(net701),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2437_ (.D(net755),
    .GATE(net701),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2438_ (.D(net753),
    .GATE(net700),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2439_ (.D(net45),
    .GATE(net700),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2440_ (.D(net750),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2441_ (.D(net749),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2442_ (.D(net776),
    .GATE(net705),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2443_ (.D(net763),
    .GATE(net705),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2444_ (.D(net751),
    .GATE(net704),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2445_ (.D(net748),
    .GATE(net704),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2446_ (.D(net50),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2447_ (.D(net51),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2448_ (.D(net745),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2449_ (.D(net744),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2450_ (.D(net743),
    .GATE(net705),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2451_ (.D(net742),
    .GATE(net705),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2452_ (.D(net775),
    .GATE(net704),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2453_ (.D(net774),
    .GATE(net704),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2454_ (.D(net773),
    .GATE(net705),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2455_ (.D(net772),
    .GATE(net705),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2456_ (.D(net770),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2457_ (.D(net768),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2458_ (.D(net767),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2459_ (.D(net766),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2460_ (.D(net765),
    .GATE(net704),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2461_ (.D(net764),
    .GATE(net704),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2462_ (.D(net762),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2463_ (.D(net761),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2464_ (.D(net760),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2465_ (.D(net759),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2466_ (.D(net758),
    .GATE(net704),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2467_ (.D(net757),
    .GATE(net704),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2468_ (.D(net756),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2469_ (.D(net755),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2470_ (.D(net753),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2471_ (.D(net45),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2472_ (.D(net750),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2473_ (.D(net749),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2474_ (.D(net27),
    .GATE(net709),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2475_ (.D(net36),
    .GATE(net709),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2476_ (.D(net46),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2477_ (.D(net49),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2478_ (.D(net747),
    .GATE(net707),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2479_ (.D(net746),
    .GATE(net707),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2480_ (.D(net745),
    .GATE(net706),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2481_ (.D(net744),
    .GATE(net706),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2482_ (.D(net54),
    .GATE(net709),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2483_ (.D(net55),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2484_ (.D(net775),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2485_ (.D(net774),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2486_ (.D(net773),
    .GATE(net707),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2487_ (.D(net772),
    .GATE(net707),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2488_ (.D(net770),
    .GATE(net706),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2489_ (.D(net768),
    .GATE(net706),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2490_ (.D(net32),
    .GATE(net709),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2491_ (.D(net33),
    .GATE(net709),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2492_ (.D(net765),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2493_ (.D(net764),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2494_ (.D(net762),
    .GATE(net706),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2495_ (.D(net761),
    .GATE(net706),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2496_ (.D(net760),
    .GATE(net706),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2497_ (.D(net759),
    .GATE(net706),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2498_ (.D(net41),
    .GATE(net709),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2499_ (.D(net42),
    .GATE(net709),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2500_ (.D(net43),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2501_ (.D(net755),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2502_ (.D(net753),
    .GATE(net707),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2503_ (.D(net752),
    .GATE(net707),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2504_ (.D(net750),
    .GATE(net706),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2505_ (.D(net749),
    .GATE(net706),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2506_ (.D(net776),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2507_ (.D(net763),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2508_ (.D(net751),
    .GATE(net711),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2509_ (.D(net748),
    .GATE(net711),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2510_ (.D(net747),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2511_ (.D(net746),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2512_ (.D(net745),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2513_ (.D(net744),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2514_ (.D(net743),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2515_ (.D(net742),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2516_ (.D(net775),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2517_ (.D(net774),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2518_ (.D(net773),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2519_ (.D(net772),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2520_ (.D(net770),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2521_ (.D(net768),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2522_ (.D(net767),
    .GATE(net712),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2523_ (.D(net766),
    .GATE(net712),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2524_ (.D(net765),
    .GATE(net712),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2525_ (.D(net764),
    .GATE(net712),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2526_ (.D(net762),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2527_ (.D(net761),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2528_ (.D(net39),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2529_ (.D(net40),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2530_ (.D(net758),
    .GATE(net712),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2531_ (.D(net757),
    .GATE(net712),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2532_ (.D(net756),
    .GATE(net712),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2533_ (.D(net755),
    .GATE(net712),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2534_ (.D(net753),
    .GATE(net711),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2535_ (.D(net752),
    .GATE(net711),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2536_ (.D(net47),
    .GATE(net711),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2537_ (.D(net48),
    .GATE(net711),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2538_ (.D(net776),
    .GATE(net714),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2539_ (.D(net763),
    .GATE(net714),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2540_ (.D(net751),
    .GATE(net714),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2541_ (.D(net748),
    .GATE(net714),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2542_ (.D(net747),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2543_ (.D(net51),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2544_ (.D(net52),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2545_ (.D(net53),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2546_ (.D(net743),
    .GATE(net717),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2547_ (.D(net742),
    .GATE(net717),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2548_ (.D(net28),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2549_ (.D(net29),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2550_ (.D(net773),
    .GATE(net717),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2551_ (.D(net772),
    .GATE(net717),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2552_ (.D(net770),
    .GATE(net714),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2553_ (.D(net768),
    .GATE(net714),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2554_ (.D(net32),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2555_ (.D(net33),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2556_ (.D(net765),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2557_ (.D(net35),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2558_ (.D(net762),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2559_ (.D(net761),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2560_ (.D(net760),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2561_ (.D(net759),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2562_ (.D(net41),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2563_ (.D(net42),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2564_ (.D(net43),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2565_ (.D(net44),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2566_ (.D(net753),
    .GATE(net714),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2567_ (.D(net752),
    .GATE(net714),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2568_ (.D(net750),
    .GATE(net714),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2569_ (.D(net749),
    .GATE(net714),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2570_ (.D(net776),
    .GATE(net718),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2571_ (.D(net763),
    .GATE(net718),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2572_ (.D(net751),
    .GATE(net718),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2573_ (.D(net748),
    .GATE(net718),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2574_ (.D(net747),
    .GATE(net718),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2575_ (.D(net746),
    .GATE(net718),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2576_ (.D(net745),
    .GATE(net718),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2577_ (.D(net744),
    .GATE(net718),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2578_ (.D(net743),
    .GATE(net720),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2579_ (.D(net742),
    .GATE(net720),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2580_ (.D(net775),
    .GATE(net720),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2581_ (.D(net774),
    .GATE(net720),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2582_ (.D(net773),
    .GATE(net719),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2583_ (.D(net772),
    .GATE(net719),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2584_ (.D(net770),
    .GATE(net718),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2585_ (.D(net768),
    .GATE(net718),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2586_ (.D(net767),
    .GATE(net719),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2587_ (.D(net766),
    .GATE(net719),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2588_ (.D(net765),
    .GATE(net57),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2589_ (.D(net764),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2590_ (.D(net37),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2591_ (.D(net38),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2592_ (.D(net760),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2593_ (.D(net40),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2594_ (.D(net758),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2595_ (.D(net757),
    .GATE(net720),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2596_ (.D(net756),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2597_ (.D(net755),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2598_ (.D(net754),
    .GATE(net720),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2599_ (.D(net752),
    .GATE(net720),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2600_ (.D(net47),
    .GATE(net720),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2601_ (.D(net48),
    .GATE(net720),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2602_ (.D(net776),
    .GATE(net722),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2603_ (.D(net763),
    .GATE(net722),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2604_ (.D(net751),
    .GATE(net725),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2605_ (.D(net748),
    .GATE(net725),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2606_ (.D(net747),
    .GATE(net722),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2607_ (.D(net746),
    .GATE(net722),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2608_ (.D(net745),
    .GATE(net722),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2609_ (.D(net744),
    .GATE(net722),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2610_ (.D(net743),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2611_ (.D(net742),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2612_ (.D(net775),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2613_ (.D(net774),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2614_ (.D(net773),
    .GATE(net722),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2615_ (.D(net772),
    .GATE(net722),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2616_ (.D(net770),
    .GATE(net722),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2617_ (.D(net768),
    .GATE(net722),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2618_ (.D(net767),
    .GATE(net724),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2619_ (.D(net766),
    .GATE(net724),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2620_ (.D(net765),
    .GATE(net724),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2621_ (.D(net764),
    .GATE(net724),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2622_ (.D(net762),
    .GATE(net726),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2623_ (.D(net761),
    .GATE(net726),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2624_ (.D(net39),
    .GATE(net726),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2625_ (.D(net40),
    .GATE(net726),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2626_ (.D(net758),
    .GATE(net724),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2627_ (.D(net757),
    .GATE(net724),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2628_ (.D(net756),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2629_ (.D(net755),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2630_ (.D(net753),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2631_ (.D(net752),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2632_ (.D(net47),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2633_ (.D(net48),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2634_ (.D(net776),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2635_ (.D(net763),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2636_ (.D(net46),
    .GATE(net740),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2637_ (.D(net49),
    .GATE(net740),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2638_ (.D(net747),
    .GATE(net738),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2639_ (.D(net746),
    .GATE(net738),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2640_ (.D(net745),
    .GATE(net738),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2641_ (.D(net744),
    .GATE(net738),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2642_ (.D(net54),
    .GATE(net741),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2643_ (.D(net55),
    .GATE(net740),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2644_ (.D(net775),
    .GATE(net740),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2645_ (.D(net774),
    .GATE(net740),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2646_ (.D(net773),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2647_ (.D(net772),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2648_ (.D(net770),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2649_ (.D(net768),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2650_ (.D(net32),
    .GATE(net740),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2651_ (.D(net33),
    .GATE(net740),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2652_ (.D(net34),
    .GATE(net741),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2653_ (.D(net35),
    .GATE(net741),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2654_ (.D(net762),
    .GATE(net738),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2655_ (.D(net761),
    .GATE(net738),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2656_ (.D(net760),
    .GATE(net738),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2657_ (.D(net759),
    .GATE(net738),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2658_ (.D(net758),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2659_ (.D(net757),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2660_ (.D(net756),
    .GATE(net741),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2661_ (.D(net44),
    .GATE(net741),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2662_ (.D(net753),
    .GATE(net740),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2663_ (.D(net752),
    .GATE(net740),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2664_ (.D(net750),
    .GATE(net738),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2665_ (.D(net749),
    .GATE(net738),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q ));
 sky130_fd_sc_hd__dfxtp_1 _2666_ (.CLK(clknet_4_12_0_UserCLK_regs),
    .D(\Inst_RegFile_32x4.BD_comb[0] ),
    .Q(\Inst_RegFile_32x4.BD_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2667_ (.CLK(clknet_4_12_0_UserCLK_regs),
    .D(\Inst_RegFile_32x4.BD_comb[1] ),
    .Q(\Inst_RegFile_32x4.BD_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2668_ (.CLK(clknet_4_12_0_UserCLK_regs),
    .D(\Inst_RegFile_32x4.BD_comb[2] ),
    .Q(\Inst_RegFile_32x4.BD_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2669_ (.CLK(clknet_4_12_0_UserCLK_regs),
    .D(\Inst_RegFile_32x4.BD_comb[3] ),
    .Q(\Inst_RegFile_32x4.BD_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2670_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(\Inst_RegFile_32x4.AD_comb[0] ),
    .Q(\Inst_RegFile_32x4.AD_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2671_ (.CLK(clknet_4_12_0_UserCLK_regs),
    .D(\Inst_RegFile_32x4.AD_comb[1] ),
    .Q(\Inst_RegFile_32x4.AD_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2672_ (.CLK(clknet_4_12_0_UserCLK_regs),
    .D(\Inst_RegFile_32x4.AD_comb[2] ),
    .Q(\Inst_RegFile_32x4.AD_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2673_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(\Inst_RegFile_32x4.AD_comb[3] ),
    .Q(\Inst_RegFile_32x4.AD_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2674_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0076_),
    .Q(\Inst_RegFile_32x4.mem[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2675_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0077_),
    .Q(\Inst_RegFile_32x4.mem[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2676_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0078_),
    .Q(\Inst_RegFile_32x4.mem[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2677_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0079_),
    .Q(\Inst_RegFile_32x4.mem[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2678_ (.CLK(clknet_4_3_0_UserCLK_regs),
    .D(_0080_),
    .Q(\Inst_RegFile_32x4.mem[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2679_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0081_),
    .Q(\Inst_RegFile_32x4.mem[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2680_ (.CLK(clknet_4_5_0_UserCLK_regs),
    .D(_0082_),
    .Q(\Inst_RegFile_32x4.mem[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2681_ (.CLK(clknet_4_5_0_UserCLK_regs),
    .D(_0083_),
    .Q(\Inst_RegFile_32x4.mem[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2682_ (.CLK(clknet_4_1_0_UserCLK_regs),
    .D(_0084_),
    .Q(\Inst_RegFile_32x4.mem[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2683_ (.CLK(clknet_4_1_0_UserCLK_regs),
    .D(_0085_),
    .Q(\Inst_RegFile_32x4.mem[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2684_ (.CLK(clknet_4_5_0_UserCLK_regs),
    .D(_0086_),
    .Q(\Inst_RegFile_32x4.mem[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2685_ (.CLK(clknet_4_4_0_UserCLK_regs),
    .D(_0087_),
    .Q(\Inst_RegFile_32x4.mem[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2686_ (.CLK(clknet_4_8_0_UserCLK_regs),
    .D(_0088_),
    .Q(\Inst_RegFile_32x4.mem[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2687_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0089_),
    .Q(\Inst_RegFile_32x4.mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2688_ (.CLK(clknet_4_8_0_UserCLK_regs),
    .D(_0090_),
    .Q(\Inst_RegFile_32x4.mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2689_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0091_),
    .Q(\Inst_RegFile_32x4.mem[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2690_ (.CLK(clknet_4_14_0_UserCLK_regs),
    .D(_0092_),
    .Q(\Inst_RegFile_32x4.mem[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2691_ (.CLK(clknet_4_14_0_UserCLK_regs),
    .D(_0093_),
    .Q(\Inst_RegFile_32x4.mem[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2692_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0094_),
    .Q(\Inst_RegFile_32x4.mem[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2693_ (.CLK(clknet_4_14_0_UserCLK_regs),
    .D(_0095_),
    .Q(\Inst_RegFile_32x4.mem[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2694_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0096_),
    .Q(\Inst_RegFile_32x4.mem[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2695_ (.CLK(clknet_4_14_0_UserCLK_regs),
    .D(_0097_),
    .Q(\Inst_RegFile_32x4.mem[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2696_ (.CLK(clknet_4_14_0_UserCLK_regs),
    .D(_0098_),
    .Q(\Inst_RegFile_32x4.mem[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2697_ (.CLK(clknet_4_14_0_UserCLK_regs),
    .D(_0099_),
    .Q(\Inst_RegFile_32x4.mem[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2698_ (.CLK(clknet_4_14_0_UserCLK_regs),
    .D(_0100_),
    .Q(\Inst_RegFile_32x4.mem[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2699_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0101_),
    .Q(\Inst_RegFile_32x4.mem[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2700_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0102_),
    .Q(\Inst_RegFile_32x4.mem[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2701_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0103_),
    .Q(\Inst_RegFile_32x4.mem[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2702_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0104_),
    .Q(\Inst_RegFile_32x4.mem[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2703_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0105_),
    .Q(\Inst_RegFile_32x4.mem[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2704_ (.CLK(clknet_4_14_0_UserCLK_regs),
    .D(_0106_),
    .Q(\Inst_RegFile_32x4.mem[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2705_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0107_),
    .Q(\Inst_RegFile_32x4.mem[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2706_ (.CLK(clknet_4_8_0_UserCLK_regs),
    .D(_0108_),
    .Q(\Inst_RegFile_32x4.mem[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2707_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(_0109_),
    .Q(\Inst_RegFile_32x4.mem[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2708_ (.CLK(clknet_4_8_0_UserCLK_regs),
    .D(_0110_),
    .Q(\Inst_RegFile_32x4.mem[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2709_ (.CLK(clknet_4_3_0_UserCLK_regs),
    .D(_0111_),
    .Q(\Inst_RegFile_32x4.mem[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2710_ (.CLK(clknet_4_8_0_UserCLK_regs),
    .D(_0112_),
    .Q(\Inst_RegFile_32x4.mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2711_ (.CLK(clknet_4_8_0_UserCLK_regs),
    .D(_0113_),
    .Q(\Inst_RegFile_32x4.mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2712_ (.CLK(clknet_4_8_0_UserCLK_regs),
    .D(_0114_),
    .Q(\Inst_RegFile_32x4.mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2713_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0115_),
    .Q(\Inst_RegFile_32x4.mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2714_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(_0116_),
    .Q(\Inst_RegFile_32x4.mem[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2715_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(_0117_),
    .Q(\Inst_RegFile_32x4.mem[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2716_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(_0118_),
    .Q(\Inst_RegFile_32x4.mem[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2717_ (.CLK(clknet_4_3_0_UserCLK_regs),
    .D(_0119_),
    .Q(\Inst_RegFile_32x4.mem[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2718_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(_0120_),
    .Q(\Inst_RegFile_32x4.mem[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2719_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(_0121_),
    .Q(\Inst_RegFile_32x4.mem[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2720_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(_0122_),
    .Q(\Inst_RegFile_32x4.mem[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2721_ (.CLK(clknet_4_3_0_UserCLK_regs),
    .D(_0123_),
    .Q(\Inst_RegFile_32x4.mem[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2722_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0124_),
    .Q(\Inst_RegFile_32x4.mem[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2723_ (.CLK(clknet_4_3_0_UserCLK_regs),
    .D(_0125_),
    .Q(\Inst_RegFile_32x4.mem[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2724_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0126_),
    .Q(\Inst_RegFile_32x4.mem[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2725_ (.CLK(clknet_4_3_0_UserCLK_regs),
    .D(_0127_),
    .Q(\Inst_RegFile_32x4.mem[12][3] ));
 sky130_fd_sc_hd__clkbuf_2 _2726_ (.A(\Inst_RegFile_switch_matrix.E1BEG0 ),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 _2727_ (.A(\Inst_RegFile_switch_matrix.E1BEG1 ),
    .X(net142));
 sky130_fd_sc_hd__buf_6 _2728_ (.A(\Inst_RegFile_switch_matrix.E1BEG2 ),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 _2729_ (.A(\Inst_RegFile_switch_matrix.E1BEG3 ),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 _2730_ (.A(\Inst_RegFile_switch_matrix.E2BEG0 ),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 _2731_ (.A(\Inst_RegFile_switch_matrix.E2BEG1 ),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 _2732_ (.A(\Inst_RegFile_switch_matrix.E2BEG2 ),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 _2733_ (.A(\Inst_RegFile_switch_matrix.E2BEG3 ),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 _2734_ (.A(\Inst_RegFile_switch_matrix.E2BEG4 ),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 _2735_ (.A(\Inst_RegFile_switch_matrix.E2BEG5 ),
    .X(net150));
 sky130_fd_sc_hd__buf_1 _2736_ (.A(\Inst_RegFile_switch_matrix.E2BEG6 ),
    .X(net151));
 sky130_fd_sc_hd__buf_4 _2737_ (.A(\Inst_RegFile_switch_matrix.E2BEG7 ),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_2 _2738_ (.A(net13),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 _2739_ (.A(net14),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 _2740_ (.A(net15),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 _2741_ (.A(net16),
    .X(net156));
 sky130_fd_sc_hd__buf_1 _2742_ (.A(net17),
    .X(net157));
 sky130_fd_sc_hd__buf_1 _2743_ (.A(net18),
    .X(net158));
 sky130_fd_sc_hd__buf_1 _2744_ (.A(net19),
    .X(net159));
 sky130_fd_sc_hd__buf_1 _2745_ (.A(net20),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 _2746_ (.A(E6END[2]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 _2747_ (.A(E6END[3]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 _2748_ (.A(E6END[4]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 _2749_ (.A(E6END[5]),
    .X(net166));
 sky130_fd_sc_hd__buf_1 _2750_ (.A(E6END[6]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 _2751_ (.A(E6END[7]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 _2752_ (.A(E6END[8]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 _2753_ (.A(E6END[9]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 _2754_ (.A(E6END[10]),
    .X(net171));
 sky130_fd_sc_hd__buf_1 _2755_ (.A(E6END[11]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 _2756_ (.A(\Inst_RegFile_switch_matrix.E6BEG0 ),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 clone18 (.A(net678),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_1 _2758_ (.A(EE4END[4]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 _2759_ (.A(EE4END[5]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 _2760_ (.A(EE4END[6]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 _2761_ (.A(EE4END[7]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 _2762_ (.A(EE4END[8]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 _2763_ (.A(EE4END[9]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 _2764_ (.A(EE4END[10]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 _2765_ (.A(EE4END[11]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 _2766_ (.A(EE4END[12]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 _2767_ (.A(EE4END[13]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 _2768_ (.A(EE4END[14]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 _2769_ (.A(EE4END[15]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 _2770_ (.A(\Inst_RegFile_switch_matrix.EE4BEG0 ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\Inst_RegFile_32x4.mem[24][0] ),
    .X(net814));
 sky130_fd_sc_hd__clkbuf_1 _2772_ (.A(\Inst_RegFile_switch_matrix.EE4BEG2 ),
    .X(net178));
 sky130_fd_sc_hd__buf_1 _2773_ (.A(\Inst_RegFile_switch_matrix.EE4BEG3 ),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 _2774_ (.A(net776),
    .X(net189));
 sky130_fd_sc_hd__buf_1 _2775_ (.A(net36),
    .X(net200));
 sky130_fd_sc_hd__buf_4 _2776_ (.A(net751),
    .X(net211));
 sky130_fd_sc_hd__buf_1 _2777_ (.A(net49),
    .X(net214));
 sky130_fd_sc_hd__buf_2 _2778_ (.A(net747),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 _2779_ (.A(net51),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 _2780_ (.A(net52),
    .X(net217));
 sky130_fd_sc_hd__buf_4 _2781_ (.A(net744),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 _2782_ (.A(net743),
    .X(net219));
 sky130_fd_sc_hd__buf_1 _2783_ (.A(net742),
    .X(net220));
 sky130_fd_sc_hd__buf_1 _2784_ (.A(net28),
    .X(net190));
 sky130_fd_sc_hd__buf_2 _2785_ (.A(net774),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 _2786_ (.A(net30),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 _2787_ (.A(net31),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 _2788_ (.A(net771),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 _2789_ (.A(net769),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 _2790_ (.A(net767),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_2 _2791_ (.A(net766),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 _2792_ (.A(net765),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 _2793_ (.A(net764),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_1 _2794_ (.A(net37),
    .X(net201));
 sky130_fd_sc_hd__buf_1 _2795_ (.A(net761),
    .X(net202));
 sky130_fd_sc_hd__buf_1 _2796_ (.A(net39),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 _2797_ (.A(net40),
    .X(net204));
 sky130_fd_sc_hd__buf_1 _2798_ (.A(net41),
    .X(net205));
 sky130_fd_sc_hd__buf_1 _2799_ (.A(net42),
    .X(net206));
 sky130_fd_sc_hd__buf_1 _2800_ (.A(net43),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 _2801_ (.A(net755),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 _2802_ (.A(net754),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_2 _2803_ (.A(net752),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 _2804_ (.A(net750),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 _2805_ (.A(net749),
    .X(net213));
 sky130_fd_sc_hd__buf_1 _2806_ (.A(net740),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_1 _2807_ (.A(net726),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 _2808_ (.A(net721),
    .X(net233));
 sky130_fd_sc_hd__buf_1 _2809_ (.A(net715),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 _2810_ (.A(net713),
    .X(net235));
 sky130_fd_sc_hd__buf_1 _2811_ (.A(net708),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 _2812_ (.A(net705),
    .X(net237));
 sky130_fd_sc_hd__buf_1 _2813_ (.A(net701),
    .X(net238));
 sky130_fd_sc_hd__buf_1 _2814_ (.A(net696),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 _2815_ (.A(net693),
    .X(net240));
 sky130_fd_sc_hd__buf_1 _2816_ (.A(net737),
    .X(net222));
 sky130_fd_sc_hd__buf_1 _2817_ (.A(net730),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_2 _2818_ (.A(net56),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_1 _2819_ (.A(FrameStrobe[13]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 _2820_ (.A(FrameStrobe[14]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 _2821_ (.A(FrameStrobe[15]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 _2822_ (.A(FrameStrobe[16]),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_1 _2823_ (.A(FrameStrobe[17]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 _2824_ (.A(FrameStrobe[18]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_1 _2825_ (.A(FrameStrobe[19]),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 _2826_ (.A(\Inst_RegFile_switch_matrix.N1BEG0 ),
    .X(net241));
 sky130_fd_sc_hd__buf_4 _2827_ (.A(\Inst_RegFile_switch_matrix.N1BEG1 ),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_2 _2828_ (.A(\Inst_RegFile_switch_matrix.N1BEG2 ),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_2 _2829_ (.A(\Inst_RegFile_switch_matrix.N1BEG3 ),
    .X(net244));
 sky130_fd_sc_hd__buf_4 _2830_ (.A(\Inst_RegFile_switch_matrix.JN2BEG0 ),
    .X(net245));
 sky130_fd_sc_hd__buf_1 _2831_ (.A(\Inst_RegFile_switch_matrix.JN2BEG1 ),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 _2832_ (.A(\Inst_RegFile_switch_matrix.JN2BEG2 ),
    .X(net247));
 sky130_fd_sc_hd__buf_1 _2833_ (.A(\Inst_RegFile_switch_matrix.JN2BEG3 ),
    .X(net248));
 sky130_fd_sc_hd__buf_1 _2834_ (.A(\Inst_RegFile_switch_matrix.JN2BEG4 ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\Inst_RegFile_32x4.mem[8][0] ),
    .X(net811));
 sky130_fd_sc_hd__buf_4 _2836_ (.A(\Inst_RegFile_switch_matrix.JN2BEG6 ),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 _2837_ (.A(\Inst_RegFile_switch_matrix.JN2BEG7 ),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_2 _2838_ (.A(net71),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_2 _2839_ (.A(net72),
    .X(net254));
 sky130_fd_sc_hd__buf_4 _2840_ (.A(net73),
    .X(net255));
 sky130_fd_sc_hd__buf_1 _2841_ (.A(net74),
    .X(net256));
 sky130_fd_sc_hd__buf_2 _2842_ (.A(net75),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_2 _2843_ (.A(net76),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_2 _2844_ (.A(net77),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_2 _2845_ (.A(net78),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_2 _2846_ (.A(N4END[4]),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_2 _2847_ (.A(N4END[5]),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_2 _2848_ (.A(N4END[6]),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_2 _2849_ (.A(N4END[7]),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_2 _2850_ (.A(N4END[8]),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_2 _2851_ (.A(N4END[9]),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_2 _2852_ (.A(N4END[10]),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_2 _2853_ (.A(N4END[11]),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_2 _2854_ (.A(N4END[12]),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_2 _2855_ (.A(N4END[13]),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_2 _2856_ (.A(N4END[14]),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_2 _2857_ (.A(N4END[15]),
    .X(net263));
 sky130_fd_sc_hd__buf_1 _2858_ (.A(\Inst_RegFile_switch_matrix.N4BEG0 ),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_1 _2859_ (.A(\Inst_RegFile_switch_matrix.N4BEG1 ),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 _2860_ (.A(\Inst_RegFile_switch_matrix.N4BEG2 ),
    .X(net266));
 sky130_fd_sc_hd__buf_1 _2861_ (.A(\Inst_RegFile_switch_matrix.N4BEG3 ),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_2 _2862_ (.A(NN4END[4]),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_2 _2863_ (.A(NN4END[5]),
    .X(net284));
 sky130_fd_sc_hd__buf_2 _2864_ (.A(NN4END[6]),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_2 _2865_ (.A(NN4END[7]),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_2 _2866_ (.A(NN4END[8]),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_2 _2867_ (.A(NN4END[9]),
    .X(net288));
 sky130_fd_sc_hd__buf_2 _2868_ (.A(NN4END[10]),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_2 _2869_ (.A(NN4END[11]),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_2 _2870_ (.A(NN4END[12]),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_2 _2871_ (.A(NN4END[13]),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_2 _2872_ (.A(NN4END[14]),
    .X(net278));
 sky130_fd_sc_hd__buf_2 _2873_ (.A(NN4END[15]),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_2 _2874_ (.A(\Inst_RegFile_switch_matrix.NN4BEG0 ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\Inst_RegFile_32x4.mem[26][3] ),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_2 _2876_ (.A(\Inst_RegFile_switch_matrix.NN4BEG2 ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\Inst_RegFile_32x4.mem[15][3] ),
    .X(net817));
 sky130_fd_sc_hd__buf_1 _2878_ (.A(\Inst_RegFile_switch_matrix.S1BEG0 ),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_2 _2879_ (.A(\Inst_RegFile_switch_matrix.S1BEG1 ),
    .X(net294));
 sky130_fd_sc_hd__buf_6 _2880_ (.A(\Inst_RegFile_switch_matrix.S1BEG2 ),
    .X(net295));
 sky130_fd_sc_hd__buf_4 _2881_ (.A(\Inst_RegFile_switch_matrix.S1BEG3 ),
    .X(net296));
 sky130_fd_sc_hd__buf_1 _2882_ (.A(\Inst_RegFile_switch_matrix.JS2BEG0 ),
    .X(net297));
 sky130_fd_sc_hd__buf_4 _2883_ (.A(\Inst_RegFile_switch_matrix.JS2BEG1 ),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_2 _2884_ (.A(\Inst_RegFile_switch_matrix.JS2BEG2 ),
    .X(net299));
 sky130_fd_sc_hd__buf_1 _2885_ (.A(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .X(net300));
 sky130_fd_sc_hd__buf_6 _2886_ (.A(\Inst_RegFile_switch_matrix.JS2BEG4 ),
    .X(net301));
 sky130_fd_sc_hd__buf_6 rebuffer200 (.A(_0859_),
    .X(net593));
 sky130_fd_sc_hd__buf_1 _2888_ (.A(\Inst_RegFile_switch_matrix.JS2BEG6 ),
    .X(net303));
 sky130_fd_sc_hd__buf_4 _2889_ (.A(\Inst_RegFile_switch_matrix.JS2BEG7 ),
    .X(net304));
 sky130_fd_sc_hd__buf_1 _2890_ (.A(net99),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_2 _2891_ (.A(net100),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_2 _2892_ (.A(net101),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_2 _2893_ (.A(net102),
    .X(net308));
 sky130_fd_sc_hd__buf_1 _2894_ (.A(net103),
    .X(net309));
 sky130_fd_sc_hd__buf_1 _2895_ (.A(net104),
    .X(net310));
 sky130_fd_sc_hd__buf_1 _2896_ (.A(net105),
    .X(net311));
 sky130_fd_sc_hd__buf_1 _2897_ (.A(net106),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_2 _2898_ (.A(S4END[4]),
    .X(net313));
 sky130_fd_sc_hd__buf_4 _2899_ (.A(S4END[5]),
    .X(net320));
 sky130_fd_sc_hd__buf_4 _2900_ (.A(S4END[6]),
    .X(net321));
 sky130_fd_sc_hd__buf_4 _2901_ (.A(S4END[7]),
    .X(net322));
 sky130_fd_sc_hd__buf_2 _2902_ (.A(S4END[8]),
    .X(net323));
 sky130_fd_sc_hd__buf_4 _2903_ (.A(S4END[9]),
    .X(net324));
 sky130_fd_sc_hd__buf_2 _2904_ (.A(S4END[10]),
    .X(net325));
 sky130_fd_sc_hd__buf_2 _2905_ (.A(S4END[11]),
    .X(net326));
 sky130_fd_sc_hd__buf_2 _2906_ (.A(S4END[12]),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_2 _2907_ (.A(S4END[13]),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_2 _2908_ (.A(S4END[14]),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_2 _2909_ (.A(S4END[15]),
    .X(net315));
 sky130_fd_sc_hd__buf_1 _2910_ (.A(\Inst_RegFile_switch_matrix.S4BEG0 ),
    .X(net316));
 sky130_fd_sc_hd__buf_1 _2911_ (.A(\Inst_RegFile_switch_matrix.S4BEG1 ),
    .X(net317));
 sky130_fd_sc_hd__buf_2 _2912_ (.A(\Inst_RegFile_switch_matrix.S4BEG2 ),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_2 _2913_ (.A(\Inst_RegFile_switch_matrix.S4BEG3 ),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_2 _2914_ (.A(SS4END[4]),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_2 _2915_ (.A(SS4END[5]),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_2 _2916_ (.A(SS4END[6]),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_2 _2917_ (.A(SS4END[7]),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_2 _2918_ (.A(SS4END[8]),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_2 _2919_ (.A(SS4END[9]),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_2 _2920_ (.A(SS4END[10]),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_2 _2921_ (.A(SS4END[11]),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 _2922_ (.A(SS4END[12]),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_2 _2923_ (.A(SS4END[13]),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_2 _2924_ (.A(SS4END[14]),
    .X(net330));
 sky130_fd_sc_hd__buf_1 _2925_ (.A(SS4END[15]),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_2 _2926_ (.A(\Inst_RegFile_switch_matrix.SS4BEG0 ),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\Inst_RegFile_32x4.mem[18][0] ),
    .X(net816));
 sky130_fd_sc_hd__buf_6 _2928_ (.A(\Inst_RegFile_switch_matrix.SS4BEG2 ),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_2 _2929_ (.A(\Inst_RegFile_switch_matrix.SS4BEG3 ),
    .X(net335));
 sky130_fd_sc_hd__buf_2 _2930_ (.A(clknet_1_0__leaf_UserCLK),
    .X(net345));
 sky130_fd_sc_hd__buf_2 _2931_ (.A(\Inst_RegFile_switch_matrix.W1BEG0 ),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_2 _2932_ (.A(\Inst_RegFile_switch_matrix.W1BEG1 ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\Inst_RegFile_32x4.mem[26][2] ),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_2 _2934_ (.A(\Inst_RegFile_switch_matrix.W1BEG3 ),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_2 _2935_ (.A(\Inst_RegFile_switch_matrix.JW2BEG0 ),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_2 _2936_ (.A(\Inst_RegFile_switch_matrix.JW2BEG1 ),
    .X(net351));
 sky130_fd_sc_hd__buf_4 _2937_ (.A(\Inst_RegFile_switch_matrix.JW2BEG2 ),
    .X(net352));
 sky130_fd_sc_hd__buf_1 _2938_ (.A(\Inst_RegFile_switch_matrix.JW2BEG3 ),
    .X(net353));
 sky130_fd_sc_hd__buf_1 _2939_ (.A(\Inst_RegFile_switch_matrix.JW2BEG4 ),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\Inst_RegFile_32x4.mem[0][0] ),
    .X(net812));
 sky130_fd_sc_hd__buf_2 _2941_ (.A(\Inst_RegFile_switch_matrix.JW2BEG6 ),
    .X(net356));
 sky130_fd_sc_hd__buf_1 _2942_ (.A(\Inst_RegFile_switch_matrix.JW2BEG7 ),
    .X(net357));
 sky130_fd_sc_hd__buf_1 _2943_ (.A(net127),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_1 _2944_ (.A(net128),
    .X(net359));
 sky130_fd_sc_hd__buf_4 _2945_ (.A(net129),
    .X(net360));
 sky130_fd_sc_hd__buf_1 _2946_ (.A(net130),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_2 _2947_ (.A(net131),
    .X(net362));
 sky130_fd_sc_hd__buf_1 _2948_ (.A(net132),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_2 _2949_ (.A(net133),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_2 _2950_ (.A(net134),
    .X(net365));
 sky130_fd_sc_hd__buf_1 _2951_ (.A(W6END[2]),
    .X(net366));
 sky130_fd_sc_hd__buf_1 _2952_ (.A(W6END[3]),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_1 _2953_ (.A(W6END[4]),
    .X(net370));
 sky130_fd_sc_hd__buf_1 _2954_ (.A(W6END[5]),
    .X(net371));
 sky130_fd_sc_hd__buf_1 _2955_ (.A(W6END[6]),
    .X(net372));
 sky130_fd_sc_hd__buf_1 _2956_ (.A(W6END[7]),
    .X(net373));
 sky130_fd_sc_hd__buf_1 _2957_ (.A(W6END[8]),
    .X(net374));
 sky130_fd_sc_hd__buf_4 _2958_ (.A(W6END[9]),
    .X(net375));
 sky130_fd_sc_hd__buf_4 _2959_ (.A(W6END[10]),
    .X(net376));
 sky130_fd_sc_hd__buf_4 _2960_ (.A(W6END[11]),
    .X(net377));
 sky130_fd_sc_hd__buf_1 _2961_ (.A(\Inst_RegFile_switch_matrix.W6BEG0 ),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_2 _2962_ (.A(\Inst_RegFile_switch_matrix.W6BEG1 ),
    .X(net368));
 sky130_fd_sc_hd__buf_1 _2963_ (.A(WW4END[4]),
    .X(net378));
 sky130_fd_sc_hd__buf_1 _2964_ (.A(WW4END[5]),
    .X(net385));
 sky130_fd_sc_hd__buf_1 _2965_ (.A(WW4END[6]),
    .X(net386));
 sky130_fd_sc_hd__buf_1 _2966_ (.A(WW4END[7]),
    .X(net387));
 sky130_fd_sc_hd__buf_1 _2967_ (.A(WW4END[8]),
    .X(net388));
 sky130_fd_sc_hd__buf_1 _2968_ (.A(WW4END[9]),
    .X(net389));
 sky130_fd_sc_hd__buf_1 _2969_ (.A(WW4END[10]),
    .X(net390));
 sky130_fd_sc_hd__buf_1 _2970_ (.A(WW4END[11]),
    .X(net391));
 sky130_fd_sc_hd__buf_1 _2971_ (.A(WW4END[12]),
    .X(net392));
 sky130_fd_sc_hd__buf_1 _2972_ (.A(WW4END[13]),
    .X(net393));
 sky130_fd_sc_hd__buf_1 _2973_ (.A(WW4END[14]),
    .X(net379));
 sky130_fd_sc_hd__buf_1 _2974_ (.A(WW4END[15]),
    .X(net380));
 sky130_fd_sc_hd__buf_1 _2975_ (.A(\Inst_RegFile_switch_matrix.WW4BEG0 ),
    .X(net381));
 sky130_fd_sc_hd__buf_6 _2976_ (.A(\Inst_RegFile_switch_matrix.WW4BEG1 ),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_2 _2977_ (.A(\Inst_RegFile_switch_matrix.WW4BEG2 ),
    .X(net383));
 sky130_fd_sc_hd__buf_8 _2978_ (.A(\Inst_RegFile_switch_matrix.WW4BEG3 ),
    .X(net384));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_831 ();
 sky130_fd_sc_hd__clkbuf_2 fanout599 (.A(net602),
    .X(net599));
 sky130_fd_sc_hd__buf_4 fanout600 (.A(net601),
    .X(net600));
 sky130_fd_sc_hd__buf_2 fanout601 (.A(net602),
    .X(net601));
 sky130_fd_sc_hd__buf_4 fanout602 (.A(_0869_),
    .X(net602));
 sky130_fd_sc_hd__buf_6 fanout603 (.A(net604),
    .X(net603));
 sky130_fd_sc_hd__buf_4 fanout604 (.A(net605),
    .X(net604));
 sky130_fd_sc_hd__buf_8 fanout605 (.A(B_ADR0),
    .X(net605));
 sky130_fd_sc_hd__clkbuf_4 fanout606 (.A(net607),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_4 fanout607 (.A(net608),
    .X(net607));
 sky130_fd_sc_hd__buf_6 fanout608 (.A(B_ADR0),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_4 fanout609 (.A(B_ADR0),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_2 fanout610 (.A(B_ADR0),
    .X(net610));
 sky130_fd_sc_hd__clkbuf_2 fanout611 (.A(_0887_),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_2 fanout612 (.A(net614),
    .X(net612));
 sky130_fd_sc_hd__buf_1 fanout613 (.A(net614),
    .X(net613));
 sky130_fd_sc_hd__buf_2 fanout614 (.A(_0887_),
    .X(net614));
 sky130_fd_sc_hd__clkbuf_2 fanout615 (.A(net618),
    .X(net615));
 sky130_fd_sc_hd__buf_4 fanout616 (.A(net617),
    .X(net616));
 sky130_fd_sc_hd__buf_4 fanout617 (.A(net618),
    .X(net617));
 sky130_fd_sc_hd__buf_4 fanout618 (.A(_0873_),
    .X(net618));
 sky130_fd_sc_hd__buf_2 fanout619 (.A(_0415_),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_2 fanout620 (.A(net623),
    .X(net620));
 sky130_fd_sc_hd__clkbuf_2 fanout621 (.A(net622),
    .X(net621));
 sky130_fd_sc_hd__clkbuf_2 fanout622 (.A(net623),
    .X(net622));
 sky130_fd_sc_hd__clkbuf_2 fanout623 (.A(_0875_),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_4 fanout624 (.A(net626),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_2 fanout625 (.A(net626),
    .X(net625));
 sky130_fd_sc_hd__buf_4 fanout626 (.A(net632),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_4 fanout627 (.A(net628),
    .X(net627));
 sky130_fd_sc_hd__clkbuf_4 fanout628 (.A(net629),
    .X(net628));
 sky130_fd_sc_hd__buf_2 fanout629 (.A(net632),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_4 fanout630 (.A(net632),
    .X(net630));
 sky130_fd_sc_hd__clkbuf_2 fanout631 (.A(net632),
    .X(net631));
 sky130_fd_sc_hd__buf_6 fanout632 (.A(A_ADR0),
    .X(net632));
 sky130_fd_sc_hd__buf_8 fanout633 (.A(net634),
    .X(net633));
 sky130_fd_sc_hd__buf_8 fanout634 (.A(BD2),
    .X(net634));
 sky130_fd_sc_hd__buf_2 fanout635 (.A(BD2),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_4 fanout636 (.A(net637),
    .X(net636));
 sky130_fd_sc_hd__clkbuf_2 fanout637 (.A(BD2),
    .X(net637));
 sky130_fd_sc_hd__buf_8 fanout638 (.A(net639),
    .X(net638));
 sky130_fd_sc_hd__buf_8 fanout639 (.A(BD3),
    .X(net639));
 sky130_fd_sc_hd__clkbuf_4 fanout640 (.A(net641),
    .X(net640));
 sky130_fd_sc_hd__buf_4 fanout641 (.A(BD3),
    .X(net641));
 sky130_fd_sc_hd__buf_4 fanout642 (.A(_0388_),
    .X(net642));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout643 (.A(_0388_),
    .X(net643));
 sky130_fd_sc_hd__buf_4 fanout644 (.A(net645),
    .X(net644));
 sky130_fd_sc_hd__buf_6 fanout645 (.A(AD3),
    .X(net645));
 sky130_fd_sc_hd__buf_8 fanout646 (.A(net647),
    .X(net646));
 sky130_fd_sc_hd__buf_6 fanout647 (.A(AD3),
    .X(net647));
 sky130_fd_sc_hd__buf_2 fanout648 (.A(_0164_),
    .X(net648));
 sky130_fd_sc_hd__buf_6 fanout649 (.A(_0163_),
    .X(net649));
 sky130_fd_sc_hd__clkbuf_2 fanout650 (.A(_0163_),
    .X(net650));
 sky130_fd_sc_hd__buf_2 fanout651 (.A(net652),
    .X(net651));
 sky130_fd_sc_hd__buf_8 fanout652 (.A(net655),
    .X(net652));
 sky130_fd_sc_hd__buf_6 fanout653 (.A(net654),
    .X(net653));
 sky130_fd_sc_hd__buf_2 fanout654 (.A(net655),
    .X(net654));
 sky130_fd_sc_hd__buf_8 fanout655 (.A(AD2),
    .X(net655));
 sky130_fd_sc_hd__buf_2 fanout656 (.A(net658),
    .X(net656));
 sky130_fd_sc_hd__buf_6 fanout657 (.A(net658),
    .X(net657));
 sky130_fd_sc_hd__buf_8 fanout658 (.A(AD1),
    .X(net658));
 sky130_fd_sc_hd__buf_2 fanout659 (.A(net660),
    .X(net659));
 sky130_fd_sc_hd__buf_2 fanout660 (.A(AD1),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_4 fanout661 (.A(net662),
    .X(net661));
 sky130_fd_sc_hd__clkbuf_2 fanout662 (.A(net663),
    .X(net662));
 sky130_fd_sc_hd__buf_4 fanout663 (.A(_0136_),
    .X(net663));
 sky130_fd_sc_hd__buf_6 fanout664 (.A(net668),
    .X(net664));
 sky130_fd_sc_hd__clkbuf_2 fanout665 (.A(net668),
    .X(net665));
 sky130_fd_sc_hd__buf_2 fanout666 (.A(net668),
    .X(net666));
 sky130_fd_sc_hd__buf_8 fanout667 (.A(net668),
    .X(net667));
 sky130_fd_sc_hd__buf_8 fanout668 (.A(BD1),
    .X(net668));
 sky130_fd_sc_hd__buf_2 fanout669 (.A(net671),
    .X(net669));
 sky130_fd_sc_hd__buf_8 fanout670 (.A(net671),
    .X(net670));
 sky130_fd_sc_hd__buf_8 fanout671 (.A(AD0),
    .X(net671));
 sky130_fd_sc_hd__buf_2 fanout672 (.A(net673),
    .X(net672));
 sky130_fd_sc_hd__buf_2 fanout673 (.A(AD0),
    .X(net673));
 sky130_fd_sc_hd__buf_6 fanout674 (.A(_0135_),
    .X(net674));
 sky130_fd_sc_hd__buf_6 fanout675 (.A(_0135_),
    .X(net675));
 sky130_fd_sc_hd__buf_2 fanout676 (.A(net678),
    .X(net676));
 sky130_fd_sc_hd__buf_8 fanout677 (.A(net678),
    .X(net677));
 sky130_fd_sc_hd__buf_8 fanout678 (.A(BD0),
    .X(net678));
 sky130_fd_sc_hd__buf_6 fanout679 (.A(net680),
    .X(net679));
 sky130_fd_sc_hd__buf_6 fanout680 (.A(BD0),
    .X(net680));
 sky130_fd_sc_hd__buf_8 fanout681 (.A(net684),
    .X(net681));
 sky130_fd_sc_hd__clkbuf_4 fanout682 (.A(net683),
    .X(net682));
 sky130_fd_sc_hd__clkbuf_4 fanout683 (.A(net684),
    .X(net683));
 sky130_fd_sc_hd__buf_8 fanout684 (.A(_0363_),
    .X(net684));
 sky130_fd_sc_hd__clkbuf_4 fanout685 (.A(_0348_),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_4 fanout686 (.A(net136),
    .X(net686));
 sky130_fd_sc_hd__clkbuf_4 fanout687 (.A(net135),
    .X(net687));
 sky130_fd_sc_hd__clkbuf_4 fanout688 (.A(net118),
    .X(net688));
 sky130_fd_sc_hd__clkbuf_4 fanout689 (.A(net117),
    .X(net689));
 sky130_fd_sc_hd__clkbuf_2 fanout690 (.A(net692),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_2 fanout691 (.A(net692),
    .X(net691));
 sky130_fd_sc_hd__buf_2 fanout692 (.A(net693),
    .X(net692));
 sky130_fd_sc_hd__buf_2 fanout693 (.A(FrameStrobe[9]),
    .X(net693));
 sky130_fd_sc_hd__clkbuf_2 fanout694 (.A(net695),
    .X(net694));
 sky130_fd_sc_hd__clkbuf_2 fanout695 (.A(net58),
    .X(net695));
 sky130_fd_sc_hd__buf_2 fanout696 (.A(net697),
    .X(net696));
 sky130_fd_sc_hd__clkbuf_2 fanout697 (.A(net58),
    .X(net697));
 sky130_fd_sc_hd__buf_2 fanout698 (.A(net699),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_2 fanout699 (.A(FrameStrobe[7]),
    .X(net699));
 sky130_fd_sc_hd__buf_2 fanout700 (.A(FrameStrobe[7]),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_2 fanout701 (.A(FrameStrobe[7]),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_2 fanout702 (.A(net704),
    .X(net702));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout703 (.A(net704),
    .X(net703));
 sky130_fd_sc_hd__buf_2 fanout704 (.A(net705),
    .X(net704));
 sky130_fd_sc_hd__clkbuf_2 fanout705 (.A(FrameStrobe[6]),
    .X(net705));
 sky130_fd_sc_hd__buf_2 fanout706 (.A(FrameStrobe[5]),
    .X(net706));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout707 (.A(FrameStrobe[5]),
    .X(net707));
 sky130_fd_sc_hd__buf_2 fanout708 (.A(FrameStrobe[5]),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_2 fanout709 (.A(FrameStrobe[5]),
    .X(net709));
 sky130_fd_sc_hd__clkbuf_2 fanout710 (.A(net711),
    .X(net710));
 sky130_fd_sc_hd__clkbuf_2 fanout711 (.A(net712),
    .X(net711));
 sky130_fd_sc_hd__buf_2 fanout712 (.A(net713),
    .X(net712));
 sky130_fd_sc_hd__clkbuf_2 fanout713 (.A(FrameStrobe[4]),
    .X(net713));
 sky130_fd_sc_hd__buf_2 fanout714 (.A(net717),
    .X(net714));
 sky130_fd_sc_hd__clkbuf_2 fanout715 (.A(net716),
    .X(net715));
 sky130_fd_sc_hd__buf_2 fanout716 (.A(net717),
    .X(net716));
 sky130_fd_sc_hd__clkbuf_2 fanout717 (.A(FrameStrobe[3]),
    .X(net717));
 sky130_fd_sc_hd__clkbuf_2 fanout718 (.A(net719),
    .X(net718));
 sky130_fd_sc_hd__clkbuf_2 fanout719 (.A(net720),
    .X(net719));
 sky130_fd_sc_hd__buf_2 fanout720 (.A(net721),
    .X(net720));
 sky130_fd_sc_hd__clkbuf_2 fanout721 (.A(net57),
    .X(net721));
 sky130_fd_sc_hd__buf_2 fanout722 (.A(net725),
    .X(net722));
 sky130_fd_sc_hd__buf_2 fanout723 (.A(net725),
    .X(net723));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout724 (.A(net725),
    .X(net724));
 sky130_fd_sc_hd__clkbuf_2 fanout725 (.A(net726),
    .X(net725));
 sky130_fd_sc_hd__clkbuf_2 fanout726 (.A(FrameStrobe[1]),
    .X(net726));
 sky130_fd_sc_hd__buf_2 fanout727 (.A(net729),
    .X(net727));
 sky130_fd_sc_hd__clkbuf_2 fanout728 (.A(net729),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_4 fanout729 (.A(net56),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_2 fanout730 (.A(net731),
    .X(net730));
 sky130_fd_sc_hd__buf_2 fanout731 (.A(net732),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_2 fanout732 (.A(FrameStrobe[11]),
    .X(net732));
 sky130_fd_sc_hd__buf_2 fanout733 (.A(FrameStrobe[11]),
    .X(net733));
 sky130_fd_sc_hd__buf_2 fanout734 (.A(net737),
    .X(net734));
 sky130_fd_sc_hd__buf_2 fanout735 (.A(net736),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_2 fanout736 (.A(net737),
    .X(net736));
 sky130_fd_sc_hd__clkbuf_2 fanout737 (.A(FrameStrobe[10]),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_2 fanout738 (.A(net739),
    .X(net738));
 sky130_fd_sc_hd__clkbuf_2 fanout739 (.A(FrameStrobe[0]),
    .X(net739));
 sky130_fd_sc_hd__buf_2 fanout740 (.A(FrameStrobe[0]),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_2 fanout741 (.A(FrameStrobe[0]),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_4 fanout742 (.A(net55),
    .X(net742));
 sky130_fd_sc_hd__buf_4 fanout743 (.A(net54),
    .X(net743));
 sky130_fd_sc_hd__buf_4 fanout744 (.A(net53),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_4 fanout745 (.A(net52),
    .X(net745));
 sky130_fd_sc_hd__clkbuf_4 fanout746 (.A(net51),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_4 fanout747 (.A(net50),
    .X(net747));
 sky130_fd_sc_hd__buf_4 fanout748 (.A(net49),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_4 fanout749 (.A(net48),
    .X(net749));
 sky130_fd_sc_hd__clkbuf_4 fanout750 (.A(net47),
    .X(net750));
 sky130_fd_sc_hd__buf_4 fanout751 (.A(net46),
    .X(net751));
 sky130_fd_sc_hd__clkbuf_4 fanout752 (.A(net45),
    .X(net752));
 sky130_fd_sc_hd__buf_4 fanout753 (.A(net754),
    .X(net753));
 sky130_fd_sc_hd__buf_2 fanout754 (.A(FrameData[28]),
    .X(net754));
 sky130_fd_sc_hd__buf_4 fanout755 (.A(net44),
    .X(net755));
 sky130_fd_sc_hd__buf_4 fanout756 (.A(net43),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_4 fanout757 (.A(net42),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_4 fanout758 (.A(net41),
    .X(net758));
 sky130_fd_sc_hd__buf_4 fanout759 (.A(net40),
    .X(net759));
 sky130_fd_sc_hd__buf_4 fanout760 (.A(net39),
    .X(net760));
 sky130_fd_sc_hd__buf_4 fanout761 (.A(net38),
    .X(net761));
 sky130_fd_sc_hd__buf_4 fanout762 (.A(net37),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_4 fanout763 (.A(net36),
    .X(net763));
 sky130_fd_sc_hd__buf_4 fanout764 (.A(net35),
    .X(net764));
 sky130_fd_sc_hd__buf_4 fanout765 (.A(net34),
    .X(net765));
 sky130_fd_sc_hd__buf_4 fanout766 (.A(net33),
    .X(net766));
 sky130_fd_sc_hd__buf_4 fanout767 (.A(net32),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_4 fanout768 (.A(net769),
    .X(net768));
 sky130_fd_sc_hd__buf_2 fanout769 (.A(FrameData[15]),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_4 fanout770 (.A(net771),
    .X(net770));
 sky130_fd_sc_hd__buf_2 fanout771 (.A(FrameData[14]),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_4 fanout772 (.A(net31),
    .X(net772));
 sky130_fd_sc_hd__clkbuf_4 fanout773 (.A(net30),
    .X(net773));
 sky130_fd_sc_hd__buf_4 fanout774 (.A(net29),
    .X(net774));
 sky130_fd_sc_hd__buf_4 fanout775 (.A(net28),
    .X(net775));
 sky130_fd_sc_hd__buf_4 fanout776 (.A(net27),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_4 fanout777 (.A(net22),
    .X(net777));
 sky130_fd_sc_hd__buf_2 fanout778 (.A(net21),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_4 fanout779 (.A(net4),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_4 fanout780 (.A(net3),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(E1END[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_6 input2 (.A(E1END[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(E1END[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(E1END[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(E2END[0]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(E2END[1]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(E2END[2]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(E2END[3]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(E2END[4]),
    .X(net9));
 sky130_fd_sc_hd__buf_6 input10 (.A(E2END[5]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(E2END[6]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(E2END[7]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(E2MID[0]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(E2MID[1]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(E2MID[2]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(E2MID[3]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(E2MID[4]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(E2MID[5]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(E2MID[6]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(E2MID[7]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(E6END[0]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(E6END[1]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(EE4END[0]),
    .X(net23));
 sky130_fd_sc_hd__buf_2 input24 (.A(EE4END[1]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input25 (.A(EE4END[2]),
    .X(net25));
 sky130_fd_sc_hd__buf_6 input26 (.A(EE4END[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_2 input27 (.A(FrameData[0]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(FrameData[10]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(FrameData[11]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input30 (.A(FrameData[12]),
    .X(net30));
 sky130_fd_sc_hd__buf_2 input31 (.A(FrameData[13]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input32 (.A(FrameData[16]),
    .X(net32));
 sky130_fd_sc_hd__buf_2 input33 (.A(FrameData[17]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(FrameData[18]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(FrameData[19]),
    .X(net35));
 sky130_fd_sc_hd__buf_2 input36 (.A(FrameData[1]),
    .X(net36));
 sky130_fd_sc_hd__buf_2 input37 (.A(FrameData[20]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 input38 (.A(FrameData[21]),
    .X(net38));
 sky130_fd_sc_hd__buf_2 input39 (.A(FrameData[22]),
    .X(net39));
 sky130_fd_sc_hd__buf_2 input40 (.A(FrameData[23]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(FrameData[24]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(FrameData[25]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(FrameData[26]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 input44 (.A(FrameData[27]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 input45 (.A(FrameData[29]),
    .X(net45));
 sky130_fd_sc_hd__buf_2 input46 (.A(FrameData[2]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(FrameData[30]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(FrameData[31]),
    .X(net48));
 sky130_fd_sc_hd__buf_2 input49 (.A(FrameData[3]),
    .X(net49));
 sky130_fd_sc_hd__buf_2 input50 (.A(FrameData[4]),
    .X(net50));
 sky130_fd_sc_hd__buf_2 input51 (.A(FrameData[5]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(FrameData[6]),
    .X(net52));
 sky130_fd_sc_hd__buf_2 input53 (.A(FrameData[7]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 input54 (.A(FrameData[8]),
    .X(net54));
 sky130_fd_sc_hd__buf_2 input55 (.A(FrameData[9]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(FrameStrobe[12]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(FrameStrobe[2]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(FrameStrobe[8]),
    .X(net58));
 sky130_fd_sc_hd__buf_4 input59 (.A(N1END[0]),
    .X(net59));
 sky130_fd_sc_hd__buf_12 input60 (.A(N1END[1]),
    .X(net60));
 sky130_fd_sc_hd__buf_4 input61 (.A(N1END[2]),
    .X(net61));
 sky130_fd_sc_hd__buf_4 input62 (.A(N1END[3]),
    .X(net62));
 sky130_fd_sc_hd__buf_2 input63 (.A(N2END[0]),
    .X(net63));
 sky130_fd_sc_hd__buf_2 input64 (.A(N2END[1]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 input65 (.A(N2END[2]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 input66 (.A(N2END[3]),
    .X(net66));
 sky130_fd_sc_hd__buf_2 input67 (.A(N2END[4]),
    .X(net67));
 sky130_fd_sc_hd__buf_6 input68 (.A(N2END[5]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_4 input69 (.A(N2END[6]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 input70 (.A(N2END[7]),
    .X(net70));
 sky130_fd_sc_hd__dlymetal6s2s_1 input71 (.A(N2MID[0]),
    .X(net71));
 sky130_fd_sc_hd__dlymetal6s2s_1 input72 (.A(N2MID[1]),
    .X(net72));
 sky130_fd_sc_hd__buf_2 input73 (.A(N2MID[2]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(N2MID[3]),
    .X(net74));
 sky130_fd_sc_hd__buf_2 input75 (.A(N2MID[4]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 input76 (.A(N2MID[5]),
    .X(net76));
 sky130_fd_sc_hd__buf_2 input77 (.A(N2MID[6]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(N2MID[7]),
    .X(net78));
 sky130_fd_sc_hd__buf_2 input79 (.A(N4END[0]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(N4END[1]),
    .X(net80));
 sky130_fd_sc_hd__buf_2 input81 (.A(N4END[2]),
    .X(net81));
 sky130_fd_sc_hd__buf_2 input82 (.A(N4END[3]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 input83 (.A(NN4END[0]),
    .X(net83));
 sky130_fd_sc_hd__buf_2 input84 (.A(NN4END[1]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 input85 (.A(NN4END[2]),
    .X(net85));
 sky130_fd_sc_hd__buf_2 input86 (.A(NN4END[3]),
    .X(net86));
 sky130_fd_sc_hd__buf_2 input87 (.A(S1END[0]),
    .X(net87));
 sky130_fd_sc_hd__buf_6 input88 (.A(S1END[1]),
    .X(net88));
 sky130_fd_sc_hd__buf_2 input89 (.A(S1END[2]),
    .X(net89));
 sky130_fd_sc_hd__buf_6 input90 (.A(S1END[3]),
    .X(net90));
 sky130_fd_sc_hd__buf_2 input91 (.A(S2END[0]),
    .X(net91));
 sky130_fd_sc_hd__buf_2 input92 (.A(S2END[1]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_4 input93 (.A(S2END[2]),
    .X(net93));
 sky130_fd_sc_hd__buf_2 input94 (.A(S2END[3]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(S2END[4]),
    .X(net95));
 sky130_fd_sc_hd__buf_6 input96 (.A(S2END[5]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(S2END[6]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 input98 (.A(S2END[7]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(S2MID[0]),
    .X(net99));
 sky130_fd_sc_hd__buf_2 input100 (.A(S2MID[1]),
    .X(net100));
 sky130_fd_sc_hd__buf_2 input101 (.A(S2MID[2]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 input102 (.A(S2MID[3]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 input103 (.A(S2MID[4]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 input104 (.A(S2MID[5]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 input105 (.A(S2MID[6]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 input106 (.A(S2MID[7]),
    .X(net106));
 sky130_fd_sc_hd__buf_2 input107 (.A(S4END[0]),
    .X(net107));
 sky130_fd_sc_hd__buf_2 input108 (.A(S4END[1]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 input109 (.A(S4END[2]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input110 (.A(S4END[3]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_4 input111 (.A(SS4END[0]),
    .X(net111));
 sky130_fd_sc_hd__buf_2 input112 (.A(SS4END[1]),
    .X(net112));
 sky130_fd_sc_hd__buf_2 input113 (.A(SS4END[2]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 input114 (.A(SS4END[3]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 input115 (.A(W1END[0]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 input116 (.A(W1END[1]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 input117 (.A(W1END[2]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 input118 (.A(W1END[3]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 input119 (.A(W2END[0]),
    .X(net119));
 sky130_fd_sc_hd__buf_2 input120 (.A(W2END[1]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_4 input121 (.A(W2END[2]),
    .X(net121));
 sky130_fd_sc_hd__buf_2 input122 (.A(W2END[3]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_4 input123 (.A(W2END[4]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input124 (.A(W2END[5]),
    .X(net124));
 sky130_fd_sc_hd__buf_1 input125 (.A(W2END[6]),
    .X(net125));
 sky130_fd_sc_hd__dlymetal6s2s_1 input126 (.A(W2END[7]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 input127 (.A(W2MID[0]),
    .X(net127));
 sky130_fd_sc_hd__buf_2 input128 (.A(W2MID[1]),
    .X(net128));
 sky130_fd_sc_hd__dlymetal6s2s_1 input129 (.A(W2MID[2]),
    .X(net129));
 sky130_fd_sc_hd__buf_2 input130 (.A(W2MID[3]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(W2MID[4]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 input132 (.A(W2MID[5]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 input133 (.A(W2MID[6]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 input134 (.A(W2MID[7]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 input135 (.A(W6END[0]),
    .X(net135));
 sky130_fd_sc_hd__dlymetal6s2s_1 input136 (.A(W6END[1]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_4 input137 (.A(WW4END[0]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_4 input138 (.A(WW4END[1]),
    .X(net138));
 sky130_fd_sc_hd__buf_2 input139 (.A(WW4END[2]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_4 input140 (.A(WW4END[3]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_4 output141 (.A(net141),
    .X(E1BEG[0]));
 sky130_fd_sc_hd__buf_4 output142 (.A(net142),
    .X(E1BEG[1]));
 sky130_fd_sc_hd__buf_4 output143 (.A(net143),
    .X(E1BEG[2]));
 sky130_fd_sc_hd__buf_4 output144 (.A(net144),
    .X(E1BEG[3]));
 sky130_fd_sc_hd__buf_4 output145 (.A(net145),
    .X(E2BEG[0]));
 sky130_fd_sc_hd__buf_6 output146 (.A(net146),
    .X(E2BEG[1]));
 sky130_fd_sc_hd__buf_6 output147 (.A(net147),
    .X(E2BEG[2]));
 sky130_fd_sc_hd__buf_6 output148 (.A(net148),
    .X(E2BEG[3]));
 sky130_fd_sc_hd__buf_6 output149 (.A(net149),
    .X(E2BEG[4]));
 sky130_fd_sc_hd__buf_6 output150 (.A(net150),
    .X(E2BEG[5]));
 sky130_fd_sc_hd__buf_4 output151 (.A(net151),
    .X(E2BEG[6]));
 sky130_fd_sc_hd__buf_4 output152 (.A(net152),
    .X(E2BEG[7]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(E2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(E2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(E2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(E2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(E2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(E2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(E2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(E2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output161 (.A(net161),
    .X(E6BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output162 (.A(net162),
    .X(E6BEG[10]));
 sky130_fd_sc_hd__buf_6 output163 (.A(\Inst_RegFile_switch_matrix.E6BEG1 ),
    .X(E6BEG[11]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net164),
    .X(E6BEG[1]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(E6BEG[2]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(E6BEG[3]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(E6BEG[4]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(E6BEG[5]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(E6BEG[6]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(E6BEG[7]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net171),
    .X(E6BEG[8]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(E6BEG[9]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net173),
    .X(EE4BEG[0]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net174),
    .X(EE4BEG[10]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net175),
    .X(EE4BEG[11]));
 sky130_fd_sc_hd__buf_2 output176 (.A(net176),
    .X(EE4BEG[12]));
 sky130_fd_sc_hd__buf_6 output177 (.A(\Inst_RegFile_switch_matrix.EE4BEG1 ),
    .X(EE4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output178 (.A(net178),
    .X(EE4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output179 (.A(net179),
    .X(EE4BEG[15]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net180),
    .X(EE4BEG[1]));
 sky130_fd_sc_hd__buf_2 output181 (.A(net181),
    .X(EE4BEG[2]));
 sky130_fd_sc_hd__buf_2 output182 (.A(net182),
    .X(EE4BEG[3]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net183),
    .X(EE4BEG[4]));
 sky130_fd_sc_hd__buf_2 output184 (.A(net184),
    .X(EE4BEG[5]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net185),
    .X(EE4BEG[6]));
 sky130_fd_sc_hd__buf_2 output186 (.A(net186),
    .X(EE4BEG[7]));
 sky130_fd_sc_hd__buf_2 output187 (.A(net187),
    .X(EE4BEG[8]));
 sky130_fd_sc_hd__buf_2 output188 (.A(net188),
    .X(EE4BEG[9]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net189),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output190 (.A(net190),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output191 (.A(net191),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output192 (.A(net192),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output193 (.A(net193),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output194 (.A(net194),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output195 (.A(net195),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output199 (.A(net199),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output201 (.A(net201),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output203 (.A(net203),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output204 (.A(net204),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output205 (.A(net205),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net206),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output207 (.A(net207),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net208),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output209 (.A(net209),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output210 (.A(net210),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output211 (.A(net211),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output212 (.A(net212),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output213 (.A(net213),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output214 (.A(net214),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output215 (.A(net215),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output216 (.A(net216),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output217 (.A(net217),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output218 (.A(net218),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output219 (.A(net219),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output220 (.A(net220),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output221 (.A(net221),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output222 (.A(net222),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output223 (.A(net223),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output224 (.A(net224),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output225 (.A(net225),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output226 (.A(net226),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output227 (.A(net227),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output228 (.A(net228),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output229 (.A(net229),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output230 (.A(net230),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output231 (.A(net231),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output232 (.A(net232),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output233 (.A(net233),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output234 (.A(net234),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output235 (.A(net235),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output236 (.A(net236),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output237 (.A(net237),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output238 (.A(net238),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output239 (.A(net239),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output240 (.A(net240),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__clkbuf_4 output241 (.A(net241),
    .X(N1BEG[0]));
 sky130_fd_sc_hd__buf_4 output242 (.A(net242),
    .X(N1BEG[1]));
 sky130_fd_sc_hd__buf_4 output243 (.A(net243),
    .X(N1BEG[2]));
 sky130_fd_sc_hd__buf_4 output244 (.A(net244),
    .X(N1BEG[3]));
 sky130_fd_sc_hd__buf_4 output245 (.A(net245),
    .X(N2BEG[0]));
 sky130_fd_sc_hd__buf_4 output246 (.A(net246),
    .X(N2BEG[1]));
 sky130_fd_sc_hd__buf_6 output247 (.A(net247),
    .X(N2BEG[2]));
 sky130_fd_sc_hd__buf_2 output248 (.A(net248),
    .X(N2BEG[3]));
 sky130_fd_sc_hd__buf_2 output249 (.A(net249),
    .X(N2BEG[4]));
 sky130_fd_sc_hd__buf_8 output250 (.A(\Inst_RegFile_switch_matrix.JN2BEG5 ),
    .X(N2BEG[5]));
 sky130_fd_sc_hd__buf_6 output251 (.A(net251),
    .X(N2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output252 (.A(net252),
    .X(N2BEG[7]));
 sky130_fd_sc_hd__buf_2 output253 (.A(net253),
    .X(N2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output254 (.A(net254),
    .X(N2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output255 (.A(net255),
    .X(N2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output256 (.A(net256),
    .X(N2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output257 (.A(net257),
    .X(N2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output258 (.A(net258),
    .X(N2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output259 (.A(net259),
    .X(N2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output260 (.A(net260),
    .X(N2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output261 (.A(net261),
    .X(N4BEG[0]));
 sky130_fd_sc_hd__buf_2 output262 (.A(net262),
    .X(N4BEG[10]));
 sky130_fd_sc_hd__buf_2 output263 (.A(net263),
    .X(N4BEG[11]));
 sky130_fd_sc_hd__buf_2 output264 (.A(net264),
    .X(N4BEG[12]));
 sky130_fd_sc_hd__buf_2 output265 (.A(net265),
    .X(N4BEG[13]));
 sky130_fd_sc_hd__buf_2 output266 (.A(net266),
    .X(N4BEG[14]));
 sky130_fd_sc_hd__buf_2 output267 (.A(net267),
    .X(N4BEG[15]));
 sky130_fd_sc_hd__buf_2 output268 (.A(net268),
    .X(N4BEG[1]));
 sky130_fd_sc_hd__buf_2 output269 (.A(net269),
    .X(N4BEG[2]));
 sky130_fd_sc_hd__buf_2 output270 (.A(net270),
    .X(N4BEG[3]));
 sky130_fd_sc_hd__buf_2 output271 (.A(net271),
    .X(N4BEG[4]));
 sky130_fd_sc_hd__buf_2 output272 (.A(net272),
    .X(N4BEG[5]));
 sky130_fd_sc_hd__buf_2 output273 (.A(net273),
    .X(N4BEG[6]));
 sky130_fd_sc_hd__buf_2 output274 (.A(net274),
    .X(N4BEG[7]));
 sky130_fd_sc_hd__buf_2 output275 (.A(net275),
    .X(N4BEG[8]));
 sky130_fd_sc_hd__buf_2 output276 (.A(net276),
    .X(N4BEG[9]));
 sky130_fd_sc_hd__buf_2 output277 (.A(net277),
    .X(NN4BEG[0]));
 sky130_fd_sc_hd__buf_2 output278 (.A(net278),
    .X(NN4BEG[10]));
 sky130_fd_sc_hd__buf_2 output279 (.A(net279),
    .X(NN4BEG[11]));
 sky130_fd_sc_hd__buf_2 output280 (.A(net280),
    .X(NN4BEG[12]));
 sky130_fd_sc_hd__buf_8 output281 (.A(\Inst_RegFile_switch_matrix.NN4BEG1 ),
    .X(NN4BEG[13]));
 sky130_fd_sc_hd__buf_4 output282 (.A(net282),
    .X(NN4BEG[14]));
 sky130_fd_sc_hd__buf_8 output283 (.A(\Inst_RegFile_switch_matrix.NN4BEG3 ),
    .X(NN4BEG[15]));
 sky130_fd_sc_hd__buf_2 output284 (.A(net284),
    .X(NN4BEG[1]));
 sky130_fd_sc_hd__buf_2 output285 (.A(net285),
    .X(NN4BEG[2]));
 sky130_fd_sc_hd__buf_2 output286 (.A(net286),
    .X(NN4BEG[3]));
 sky130_fd_sc_hd__buf_2 output287 (.A(net287),
    .X(NN4BEG[4]));
 sky130_fd_sc_hd__buf_2 output288 (.A(net288),
    .X(NN4BEG[5]));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .X(NN4BEG[6]));
 sky130_fd_sc_hd__buf_2 output290 (.A(net290),
    .X(NN4BEG[7]));
 sky130_fd_sc_hd__buf_2 output291 (.A(net291),
    .X(NN4BEG[8]));
 sky130_fd_sc_hd__buf_2 output292 (.A(net292),
    .X(NN4BEG[9]));
 sky130_fd_sc_hd__buf_4 output293 (.A(net293),
    .X(S1BEG[0]));
 sky130_fd_sc_hd__buf_4 output294 (.A(net294),
    .X(S1BEG[1]));
 sky130_fd_sc_hd__buf_4 output295 (.A(net295),
    .X(S1BEG[2]));
 sky130_fd_sc_hd__buf_4 output296 (.A(net296),
    .X(S1BEG[3]));
 sky130_fd_sc_hd__buf_4 output297 (.A(net297),
    .X(S2BEG[0]));
 sky130_fd_sc_hd__buf_4 output298 (.A(net298),
    .X(S2BEG[1]));
 sky130_fd_sc_hd__buf_6 output299 (.A(net299),
    .X(S2BEG[2]));
 sky130_fd_sc_hd__buf_2 output300 (.A(net300),
    .X(S2BEG[3]));
 sky130_fd_sc_hd__buf_8 output301 (.A(net301),
    .X(S2BEG[4]));
 sky130_fd_sc_hd__buf_6 output302 (.A(\Inst_RegFile_switch_matrix.JS2BEG5 ),
    .X(S2BEG[5]));
 sky130_fd_sc_hd__buf_6 output303 (.A(net303),
    .X(S2BEG[6]));
 sky130_fd_sc_hd__buf_4 output304 (.A(net304),
    .X(S2BEG[7]));
 sky130_fd_sc_hd__buf_2 output305 (.A(net305),
    .X(S2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output306 (.A(net306),
    .X(S2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output307 (.A(net307),
    .X(S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output308 (.A(net308),
    .X(S2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output309 (.A(net309),
    .X(S2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output310 (.A(net310),
    .X(S2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output311 (.A(net311),
    .X(S2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output312 (.A(net312),
    .X(S2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output313 (.A(net313),
    .X(S4BEG[0]));
 sky130_fd_sc_hd__buf_2 output314 (.A(net314),
    .X(S4BEG[10]));
 sky130_fd_sc_hd__buf_2 output315 (.A(net315),
    .X(S4BEG[11]));
 sky130_fd_sc_hd__buf_2 output316 (.A(net316),
    .X(S4BEG[12]));
 sky130_fd_sc_hd__buf_2 output317 (.A(net317),
    .X(S4BEG[13]));
 sky130_fd_sc_hd__buf_6 output318 (.A(net318),
    .X(S4BEG[14]));
 sky130_fd_sc_hd__buf_4 output319 (.A(net319),
    .X(S4BEG[15]));
 sky130_fd_sc_hd__buf_2 output320 (.A(net320),
    .X(S4BEG[1]));
 sky130_fd_sc_hd__buf_2 output321 (.A(net321),
    .X(S4BEG[2]));
 sky130_fd_sc_hd__buf_2 output322 (.A(net322),
    .X(S4BEG[3]));
 sky130_fd_sc_hd__buf_2 output323 (.A(net323),
    .X(S4BEG[4]));
 sky130_fd_sc_hd__buf_2 output324 (.A(net324),
    .X(S4BEG[5]));
 sky130_fd_sc_hd__buf_2 output325 (.A(net325),
    .X(S4BEG[6]));
 sky130_fd_sc_hd__buf_2 output326 (.A(net326),
    .X(S4BEG[7]));
 sky130_fd_sc_hd__buf_2 output327 (.A(net327),
    .X(S4BEG[8]));
 sky130_fd_sc_hd__buf_2 output328 (.A(net328),
    .X(S4BEG[9]));
 sky130_fd_sc_hd__buf_2 output329 (.A(net329),
    .X(SS4BEG[0]));
 sky130_fd_sc_hd__buf_2 output330 (.A(net330),
    .X(SS4BEG[10]));
 sky130_fd_sc_hd__buf_2 output331 (.A(net331),
    .X(SS4BEG[11]));
 sky130_fd_sc_hd__buf_2 output332 (.A(net332),
    .X(SS4BEG[12]));
 sky130_fd_sc_hd__buf_8 output333 (.A(\Inst_RegFile_switch_matrix.SS4BEG1 ),
    .X(SS4BEG[13]));
 sky130_fd_sc_hd__buf_8 output334 (.A(net334),
    .X(SS4BEG[14]));
 sky130_fd_sc_hd__buf_4 output335 (.A(net335),
    .X(SS4BEG[15]));
 sky130_fd_sc_hd__buf_2 output336 (.A(net336),
    .X(SS4BEG[1]));
 sky130_fd_sc_hd__buf_2 output337 (.A(net337),
    .X(SS4BEG[2]));
 sky130_fd_sc_hd__buf_2 output338 (.A(net338),
    .X(SS4BEG[3]));
 sky130_fd_sc_hd__buf_2 output339 (.A(net339),
    .X(SS4BEG[4]));
 sky130_fd_sc_hd__buf_2 output340 (.A(net340),
    .X(SS4BEG[5]));
 sky130_fd_sc_hd__buf_2 output341 (.A(net341),
    .X(SS4BEG[6]));
 sky130_fd_sc_hd__buf_2 output342 (.A(net342),
    .X(SS4BEG[7]));
 sky130_fd_sc_hd__buf_2 output343 (.A(net343),
    .X(SS4BEG[8]));
 sky130_fd_sc_hd__buf_2 output344 (.A(net344),
    .X(SS4BEG[9]));
 sky130_fd_sc_hd__buf_1 output345 (.A(net345),
    .X(UserCLKo));
 sky130_fd_sc_hd__buf_4 output346 (.A(net346),
    .X(W1BEG[0]));
 sky130_fd_sc_hd__buf_4 output347 (.A(net347),
    .X(W1BEG[1]));
 sky130_fd_sc_hd__buf_6 output348 (.A(\Inst_RegFile_switch_matrix.W1BEG2 ),
    .X(W1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output349 (.A(net349),
    .X(W1BEG[3]));
 sky130_fd_sc_hd__buf_4 output350 (.A(net350),
    .X(W2BEG[0]));
 sky130_fd_sc_hd__buf_4 output351 (.A(net351),
    .X(W2BEG[1]));
 sky130_fd_sc_hd__buf_4 output352 (.A(net352),
    .X(W2BEG[2]));
 sky130_fd_sc_hd__buf_2 output353 (.A(net353),
    .X(W2BEG[3]));
 sky130_fd_sc_hd__buf_4 output354 (.A(net354),
    .X(W2BEG[4]));
 sky130_fd_sc_hd__buf_8 output355 (.A(\Inst_RegFile_switch_matrix.JW2BEG5 ),
    .X(W2BEG[5]));
 sky130_fd_sc_hd__buf_4 output356 (.A(net356),
    .X(W2BEG[6]));
 sky130_fd_sc_hd__buf_4 output357 (.A(net357),
    .X(W2BEG[7]));
 sky130_fd_sc_hd__buf_2 output358 (.A(net358),
    .X(W2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output359 (.A(net359),
    .X(W2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output360 (.A(net360),
    .X(W2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output361 (.A(net361),
    .X(W2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output362 (.A(net362),
    .X(W2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output363 (.A(net363),
    .X(W2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output364 (.A(net364),
    .X(W2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output365 (.A(net365),
    .X(W2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output366 (.A(net366),
    .X(W6BEG[0]));
 sky130_fd_sc_hd__buf_4 output367 (.A(net367),
    .X(W6BEG[10]));
 sky130_fd_sc_hd__buf_4 output368 (.A(net368),
    .X(W6BEG[11]));
 sky130_fd_sc_hd__buf_2 output369 (.A(net369),
    .X(W6BEG[1]));
 sky130_fd_sc_hd__buf_2 output370 (.A(net370),
    .X(W6BEG[2]));
 sky130_fd_sc_hd__buf_2 output371 (.A(net371),
    .X(W6BEG[3]));
 sky130_fd_sc_hd__buf_2 output372 (.A(net372),
    .X(W6BEG[4]));
 sky130_fd_sc_hd__buf_2 output373 (.A(net373),
    .X(W6BEG[5]));
 sky130_fd_sc_hd__buf_2 output374 (.A(net374),
    .X(W6BEG[6]));
 sky130_fd_sc_hd__buf_2 output375 (.A(net375),
    .X(W6BEG[7]));
 sky130_fd_sc_hd__buf_2 output376 (.A(net376),
    .X(W6BEG[8]));
 sky130_fd_sc_hd__buf_2 output377 (.A(net377),
    .X(W6BEG[9]));
 sky130_fd_sc_hd__buf_2 output378 (.A(net378),
    .X(WW4BEG[0]));
 sky130_fd_sc_hd__buf_2 output379 (.A(net379),
    .X(WW4BEG[10]));
 sky130_fd_sc_hd__buf_2 output380 (.A(net380),
    .X(WW4BEG[11]));
 sky130_fd_sc_hd__buf_2 output381 (.A(net381),
    .X(WW4BEG[12]));
 sky130_fd_sc_hd__buf_8 output382 (.A(net382),
    .X(WW4BEG[13]));
 sky130_fd_sc_hd__buf_6 output383 (.A(net383),
    .X(WW4BEG[14]));
 sky130_fd_sc_hd__buf_8 output384 (.A(net384),
    .X(WW4BEG[15]));
 sky130_fd_sc_hd__buf_2 output385 (.A(net385),
    .X(WW4BEG[1]));
 sky130_fd_sc_hd__buf_2 output386 (.A(net386),
    .X(WW4BEG[2]));
 sky130_fd_sc_hd__buf_2 output387 (.A(net387),
    .X(WW4BEG[3]));
 sky130_fd_sc_hd__buf_2 output388 (.A(net388),
    .X(WW4BEG[4]));
 sky130_fd_sc_hd__buf_2 output389 (.A(net389),
    .X(WW4BEG[5]));
 sky130_fd_sc_hd__buf_2 output390 (.A(net390),
    .X(WW4BEG[6]));
 sky130_fd_sc_hd__buf_2 output391 (.A(net391),
    .X(WW4BEG[7]));
 sky130_fd_sc_hd__buf_2 output392 (.A(net392),
    .X(WW4BEG[8]));
 sky130_fd_sc_hd__buf_2 output393 (.A(net393),
    .X(WW4BEG[9]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_regs_0_UserCLK (.A(UserCLK),
    .X(UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_UserCLK (.A(UserCLK),
    .X(clknet_0_UserCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_UserCLK (.A(clknet_0_UserCLK),
    .X(clknet_1_0__leaf_UserCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_UserCLK_regs (.A(UserCLK_regs),
    .X(clknet_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_0_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_1_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_2_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_3_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_4_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_5_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_6_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_7_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_8_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_9_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_10_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_11_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_12_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_13_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_14_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_15_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinv_2 clkload0 (.A(clknet_4_0_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload1 (.A(clknet_4_1_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_4 clkload2 (.A(clknet_4_2_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinv_2 clkload3 (.A(clknet_4_3_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload4 (.A(clknet_4_4_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinv_2 clkload5 (.A(clknet_4_5_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload6 (.A(clknet_4_6_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinv_2 clkload7 (.A(clknet_4_7_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinv_2 clkload8 (.A(clknet_4_9_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_4 clkload9 (.A(clknet_4_10_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinv_2 clkload10 (.A(clknet_4_12_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload11 (.A(clknet_4_13_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinv_2 clkload12 (.A(clknet_4_14_0_UserCLK_regs));
 sky130_fd_sc_hd__buf_6 rebuffer1 (.A(_0400_),
    .X(net394));
 sky130_fd_sc_hd__a31o_4 clone2 (.A1(_0178_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q ),
    .A3(_0180_),
    .B1(_0191_),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_1 clone3 (.A(_0135_),
    .X(net396));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer4 (.A(_0400_),
    .X(net397));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer5 (.A(AD3),
    .X(net398));
 sky130_fd_sc_hd__buf_6 clone15 (.A(_0163_),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_1 clone16 (.A(BD3),
    .X(net409));
 sky130_fd_sc_hd__buf_6 clone17 (.A(B_ADR0),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_1 clone19 (.A(net684),
    .X(net412));
 sky130_fd_sc_hd__buf_6 clone20 (.A(_0363_),
    .X(net413));
 sky130_fd_sc_hd__buf_6 rebuffer21 (.A(_1036_),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_1 clone22 (.A(net634),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(_0436_),
    .X(net420));
 sky130_fd_sc_hd__buf_6 clone28 (.A(AD3),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_1 clone29 (.A(net647),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_1 clone30 (.A(net655),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\Inst_RegFile_32x4.mem[6][1] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\Inst_RegFile_32x4.mem[4][0] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\Inst_RegFile_32x4.mem[4][3] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\Inst_RegFile_32x4.mem[30][3] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\Inst_RegFile_32x4.mem[6][0] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\Inst_RegFile_32x4.mem[12][2] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\Inst_RegFile_32x4.mem[6][2] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\Inst_RegFile_32x4.mem[4][2] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\Inst_RegFile_32x4.mem[26][0] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\Inst_RegFile_32x4.mem[20][1] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\Inst_RegFile_32x4.mem[4][1] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\Inst_RegFile_32x4.mem[25][0] ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\Inst_RegFile_32x4.mem[1][0] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\Inst_RegFile_32x4.mem[15][0] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\Inst_RegFile_32x4.mem[30][1] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\Inst_RegFile_32x4.mem[24][1] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\Inst_RegFile_32x4.mem[27][2] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\Inst_RegFile_32x4.mem[20][0] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\Inst_RegFile_32x4.mem[13][2] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\Inst_RegFile_32x4.mem[5][0] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\Inst_RegFile_32x4.mem[29][0] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\Inst_RegFile_32x4.mem[11][3] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\Inst_RegFile_32x4.mem[17][1] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\Inst_RegFile_32x4.mem[2][0] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\Inst_RegFile_32x4.mem[19][2] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\Inst_RegFile_32x4.mem[30][0] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\Inst_RegFile_32x4.mem[17][0] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\Inst_RegFile_32x4.mem[19][3] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\Inst_RegFile_32x4.mem[13][1] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\Inst_RegFile_32x4.mem[13][0] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\Inst_RegFile_32x4.mem[3][0] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\Inst_RegFile_32x4.mem[20][3] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\Inst_RegFile_32x4.mem[30][2] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\Inst_RegFile_32x4.mem[12][1] ),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\Inst_RegFile_32x4.mem[31][0] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\Inst_RegFile_32x4.mem[9][1] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\Inst_RegFile_32x4.mem[6][3] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\Inst_RegFile_32x4.mem[21][0] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\Inst_RegFile_32x4.mem[5][2] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\Inst_RegFile_32x4.mem[15][1] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\Inst_RegFile_32x4.mem[31][2] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\Inst_RegFile_32x4.mem[15][2] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\Inst_RegFile_32x4.mem[29][1] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\Inst_RegFile_32x4.mem[19][0] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\Inst_RegFile_32x4.mem[22][0] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\Inst_RegFile_32x4.mem[23][2] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\Inst_RegFile_32x4.mem[9][2] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\Inst_RegFile_32x4.mem[21][3] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\Inst_RegFile_32x4.mem[24][3] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\Inst_RegFile_32x4.mem[13][3] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\Inst_RegFile_32x4.mem[27][0] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\Inst_RegFile_32x4.mem[23][0] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\Inst_RegFile_32x4.mem[11][1] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\Inst_RegFile_32x4.mem[1][3] ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\Inst_RegFile_32x4.mem[9][3] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\Inst_RegFile_32x4.mem[1][1] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\Inst_RegFile_32x4.mem[11][2] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\Inst_RegFile_32x4.mem[5][1] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\Inst_RegFile_32x4.mem[29][3] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\Inst_RegFile_32x4.mem[27][1] ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\Inst_RegFile_32x4.mem[29][2] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\Inst_RegFile_32x4.mem[9][0] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\Inst_RegFile_32x4.mem[10][0] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\Inst_RegFile_32x4.mem[5][3] ),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\Inst_RegFile_32x4.mem[21][1] ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\Inst_RegFile_32x4.mem[27][3] ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\Inst_RegFile_32x4.mem[14][2] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\Inst_RegFile_32x4.mem[2][3] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\Inst_RegFile_32x4.mem[19][1] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\Inst_RegFile_32x4.mem[17][3] ),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\Inst_RegFile_32x4.mem[12][3] ),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\Inst_RegFile_32x4.mem[17][2] ),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\Inst_RegFile_32x4.mem[0][3] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\Inst_RegFile_32x4.mem[14][0] ),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\Inst_RegFile_32x4.mem[23][3] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\Inst_RegFile_32x4.mem[11][0] ),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\Inst_RegFile_32x4.mem[18][2] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\Inst_RegFile_32x4.mem[14][3] ),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\Inst_RegFile_32x4.mem[8][1] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\Inst_RegFile_32x4.mem[20][2] ),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\Inst_RegFile_32x4.mem[0][1] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\Inst_RegFile_32x4.mem[10][1] ),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\Inst_RegFile_32x4.mem[28][3] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\Inst_RegFile_32x4.mem[2][2] ),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\Inst_RegFile_32x4.mem[28][0] ),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\Inst_RegFile_32x4.mem[16][0] ),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\Inst_RegFile_32x4.mem[14][1] ),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\Inst_RegFile_32x4.mem[28][2] ),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\Inst_RegFile_32x4.mem[16][2] ),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\Inst_RegFile_32x4.mem[26][1] ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\Inst_RegFile_32x4.mem[1][2] ),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\Inst_RegFile_32x4.mem[24][2] ),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\Inst_RegFile_32x4.mem[18][3] ),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\Inst_RegFile_32x4.mem[16][1] ),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\Inst_RegFile_32x4.mem[31][3] ),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\Inst_RegFile_32x4.mem[3][2] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\Inst_RegFile_32x4.mem[8][2] ),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\Inst_RegFile_32x4.mem[7][2] ),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\Inst_RegFile_32x4.mem[0][2] ),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\Inst_RegFile_32x4.mem[28][1] ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\Inst_RegFile_32x4.mem[10][2] ),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\Inst_RegFile_32x4.mem[22][1] ),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\Inst_RegFile_32x4.mem[8][3] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\Inst_RegFile_32x4.mem[3][3] ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\Inst_RegFile_32x4.mem[10][3] ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\Inst_RegFile_32x4.mem[2][1] ),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\Inst_RegFile_32x4.mem[3][1] ),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\Inst_RegFile_32x4.mem[7][1] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\Inst_RegFile_32x4.mem[21][2] ),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\Inst_RegFile_32x4.mem[22][3] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\Inst_RegFile_32x4.mem[31][1] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\Inst_RegFile_32x4.mem[18][1] ),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\Inst_RegFile_32x4.mem[12][0] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\Inst_RegFile_32x4.mem[25][1] ),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\Inst_RegFile_32x4.mem[25][2] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\Inst_RegFile_32x4.mem[7][0] ),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\Inst_RegFile_32x4.mem[16][3] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\Inst_RegFile_32x4.mem[22][2] ),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\Inst_RegFile_32x4.mem[7][3] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\Inst_RegFile_32x4.mem[23][1] ),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\Inst_RegFile_32x4.mem[25][3] ),
    .X(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(E6END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(E6END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(E6END[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(E6END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(E6END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(E6END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(E6END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(E6END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(E6END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(E6END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(E6END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(E6END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(EE4END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(EE4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(EE4END[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(EE4END[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(EE4END[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(EE4END[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(EE4END[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(EE4END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(EE4END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(EE4END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(EE4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(FrameData[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(FrameStrobe[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(FrameStrobe[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(FrameStrobe[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(FrameStrobe[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(FrameStrobe[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(FrameStrobe[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(FrameStrobe[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(FrameStrobe[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(FrameStrobe[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(FrameStrobe[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(FrameStrobe[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(FrameStrobe[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(FrameStrobe[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(\Inst_RegFile_switch_matrix.JW2BEG6 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(\Inst_RegFile_switch_matrix.JW2BEG6 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(N4END[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(N4END[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(N4END[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(N4END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(S4END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(S4END[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(S4END[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(S4END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(S4END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(S4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(SS4END[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(W6END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(W6END[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(W6END[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(W6END[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(W6END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(W6END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(W6END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(W6END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(W6END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(W6END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(WW4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(WW4END[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(WW4END[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(WW4END[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(WW4END[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(WW4END[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(WW4END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(WW4END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(WW4END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(WW4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(_0129_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(_0133_));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(_0213_));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(_0213_));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(_0213_));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(E6END[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(E6END[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(EE4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(EE4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(FrameStrobe[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(FrameStrobe[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(N4END[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(N4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(NN4END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(SS4END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(WW4END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(WW4END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(_0264_));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(net777));
 sky130_fd_sc_hd__fill_1 FILLER_0_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_473 ();
endmodule
