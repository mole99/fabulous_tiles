* NGSPICE file created from S_CPU_IF.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt S_CPU_IF Co FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] I_top0 I_top1 I_top10 I_top11
+ I_top12 I_top13 I_top14 I_top15 I_top2 I_top3 I_top4 I_top5 I_top6 I_top7 I_top8
+ I_top9 N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3] N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4]
+ N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5]
+ N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15]
+ N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9]
+ NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1]
+ NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9]
+ O_top0 O_top1 O_top10 O_top11 O_top12 O_top13 O_top14 O_top15 O_top2 O_top3 O_top4
+ O_top5 O_top6 O_top7 O_top8 O_top9 S1END[0] S1END[1] S1END[2] S1END[3] S2END[0]
+ S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1]
+ S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10] S4END[11]
+ S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5]
+ S4END[6] S4END[7] S4END[8] S4END[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13]
+ SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6]
+ SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR
XFILLER_5_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput220 net231 VGND VGND VPWR VPWR NN4BEG[9] sky130_fd_sc_hd__buf_2
X_062_ net78 net56 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit17.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N2BEG1 sky130_fd_sc_hd__mux2_1
X_131_ net30 net43 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_200_ FrameStrobe[11] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_114_ net15 net40 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_045_ net84 net49 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit2.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N4BEG2 sky130_fd_sc_hd__mux2_1
X_028_ net99 net48 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit19.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.NN4BEG3 sky130_fd_sc_hd__mux2_1
XFILLER_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput210 net221 VGND VGND VPWR VPWR NN4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput221 net232 VGND VGND VPWR VPWR UserCLKo sky130_fd_sc_hd__buf_1
X_130_ net29 net43 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_9_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_259_ Inst_S_CPU_IF_switch_matrix.NN4BEG14 VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__buf_1
X_061_ net77 net55 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit18.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N2BEG2 sky130_fd_sc_hd__mux2_1
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_044_ net83 net48 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit3.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N4BEG3 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_113_ net14 net41 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_027_ net98 net47 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit20.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.NN4BEG4 sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput211 net222 VGND VGND VPWR VPWR NN4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput200 net211 VGND VGND VPWR VPWR N4BEG[5] sky130_fd_sc_hd__buf_2
X_060_ net76 net54 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit19.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N2BEG3 sky130_fd_sc_hd__mux2_1
XFILLER_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_189_ net44 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_1
X_258_ Inst_S_CPU_IF_switch_matrix.NN4BEG13 VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__buf_1
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_043_ net82 net47 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit4.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N4BEG4 sky130_fd_sc_hd__mux2_1
X_112_ net13 net41 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_026_ net97 net46 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit21.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.NN4BEG5 sky130_fd_sc_hd__mux2_1
Xinput100 SS4END[9] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_1
XFILLER_0_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_009_ net62 net66 net92 net108 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit12.Q Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit13.Q
+ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__mux4_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput201 net212 VGND VGND VPWR VPWR N4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput212 net223 VGND VGND VPWR VPWR NN4BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_257_ Inst_S_CPU_IF_switch_matrix.NN4BEG12 VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_188_ net25 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
X_111_ net11 net38 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_042_ net81 net46 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit5.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N4BEG5 sky130_fd_sc_hd__mux2_1
XFILLER_3_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_025_ net111 net59 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit22.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.NN4BEG6 sky130_fd_sc_hd__mux2_1
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_008_ net63 net67 net93 net109 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit14.Q Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit15.Q
+ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__mux4_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput213 net224 VGND VGND VPWR VPWR NN4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput202 net213 VGND VGND VPWR VPWR N4BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_256_ Inst_S_CPU_IF_switch_matrix.NN4BEG11 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_1
X_187_ net24 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
X_041_ net95 net59 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit6.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N4BEG6 sky130_fd_sc_hd__mux2_1
X_110_ net10 net38 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_239_ Inst_S_CPU_IF_switch_matrix.N4BEG10 VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__buf_1
X_024_ net110 net58 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit23.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.NN4BEG7 sky130_fd_sc_hd__mux2_1
XFILLER_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_007_ net60 net68 net94 net110 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit16.Q Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit17.Q
+ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__mux4_1
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput214 net225 VGND VGND VPWR VPWR NN4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput203 net214 VGND VGND VPWR VPWR N4BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_186_ net22 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
X_255_ Inst_S_CPU_IF_switch_matrix.NN4BEG10 VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__buf_1
X_040_ net94 net58 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit7.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N4BEG7 sky130_fd_sc_hd__mux2_1
X_238_ Inst_S_CPU_IF_switch_matrix.N4BEG9 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__buf_1
XFILLER_6_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_169_ net4 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_1
X_023_ net109 net57 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit24.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.NN4BEG8 sky130_fd_sc_hd__mux2_1
XFILLER_8_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_006_ net61 net69 net95 net111 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit18.Q Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit19.Q
+ VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__mux4_1
XFILLER_7_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput215 net226 VGND VGND VPWR VPWR NN4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput204 net215 VGND VGND VPWR VPWR N4BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_185_ net21 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__buf_1
X_254_ Inst_S_CPU_IF_switch_matrix.NN4BEG9 VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__buf_1
XFILLER_6_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_099_ net30 net41 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_237_ Inst_S_CPU_IF_switch_matrix.N4BEG8 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_1
X_168_ net3 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_022_ net108 net56 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit25.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.NN4BEG9 sky130_fd_sc_hd__mux2_1
XFILLER_3_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_005_ net62 net70 net81 net97 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit20.Q Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit21.Q
+ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__mux4_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput216 net227 VGND VGND VPWR VPWR NN4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput205 net216 VGND VGND VPWR VPWR NN4BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_4_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_253_ Inst_S_CPU_IF_switch_matrix.NN4BEG8 VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_1
X_184_ net20 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_0_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_236_ Inst_S_CPU_IF_switch_matrix.N4BEG7 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_1
X_098_ net29 net40 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_167_ net2 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_1
X_021_ net107 net55 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit26.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.NN4BEG10 sky130_fd_sc_hd__mux2_1
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_219_ Inst_S_CPU_IF_switch_matrix.N2BEG6 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_1
X_004_ net63 net71 net82 net98 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit22.Q Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit23.Q
+ VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__mux4_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput206 net217 VGND VGND VPWR VPWR NN4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput217 net228 VGND VGND VPWR VPWR NN4BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_252_ Inst_S_CPU_IF_switch_matrix.NN4BEG7 VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_183_ net19 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_0_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout40 net41 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
XFILLER_9_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_235_ Inst_S_CPU_IF_switch_matrix.N4BEG6 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__buf_1
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_166_ net32 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_097_ net28 net41 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_020_ net106 net54 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit27.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.NN4BEG11 sky130_fd_sc_hd__mux2_1
XFILLER_3_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_149_ net18 net44 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_6_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_218_ Inst_S_CPU_IF_switch_matrix.N2BEG5 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
X_003_ net60 net76 net83 net99 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit24.Q Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit25.Q
+ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__mux4_1
XFILLER_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput218 net229 VGND VGND VPWR VPWR NN4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput207 net218 VGND VGND VPWR VPWR NN4BEG[11] sky130_fd_sc_hd__buf_2
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_182_ net18 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_0_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout41 FrameStrobe[1] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
X_251_ Inst_S_CPU_IF_switch_matrix.NN4BEG6 VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_165_ net31 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
X_234_ Inst_S_CPU_IF_switch_matrix.N4BEG5 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__buf_1
XFILLER_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_096_ net27 net41 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_148_ net17 net44 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_217_ Inst_S_CPU_IF_switch_matrix.N2BEG4 VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_079_ net11 net36 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_002_ net61 net77 net84 net100 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit26.Q Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit27.Q
+ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__mux4_1
XFILLER_7_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput208 net219 VGND VGND VPWR VPWR NN4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput219 net230 VGND VGND VPWR VPWR NN4BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_4_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_181_ net17 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__buf_1
XFILLER_6_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout42 net43 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_250_ Inst_S_CPU_IF_switch_matrix.NN4BEG5 VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__buf_1
XFILLER_9_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_164_ net30 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__buf_1
X_095_ net26 net38 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_233_ Inst_S_CPU_IF_switch_matrix.N4BEG4 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_216_ Inst_S_CPU_IF_switch_matrix.N2BEG3 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_1
X_147_ net16 net42 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_078_ net10 net36 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_001_ net62 net78 net85 net101 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit28.Q Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit29.Q
+ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__mux4_1
XFILLER_7_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput90 SS4END[14] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput209 net220 VGND VGND VPWR VPWR NN4BEG[13] sky130_fd_sc_hd__buf_2
XFILLER_4_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout43 net45 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
X_180_ net16 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_9_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_232_ Inst_S_CPU_IF_switch_matrix.N4BEG3 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__buf_1
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_094_ net23 net38 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_163_ net29 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__buf_1
XFILLER_10_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_077_ net9 net36 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_6_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_215_ Inst_S_CPU_IF_switch_matrix.N2BEG2 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_146_ net15 net44 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_000_ net63 net79 net86 net102 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit30.Q Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit31.Q
+ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__mux4_1
Xinput80 S4END[5] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_1
Xinput91 SS4END[15] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_1
X_129_ net28 net42 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout44 net45 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_9_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_093_ net12 net38 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_231_ Inst_S_CPU_IF_switch_matrix.N4BEG2 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_1
X_162_ net28 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput1 FrameData[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
X_214_ Inst_S_CPU_IF_switch_matrix.N2BEG1 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_076_ net8 net35 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_145_ net14 net44 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput190 net201 VGND VGND VPWR VPWR N4BEG[10] sky130_fd_sc_hd__buf_2
X_059_ net75 net53 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit20.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N2BEG4 sky130_fd_sc_hd__mux2_1
X_128_ net27 net42 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput92 SS4END[1] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__buf_1
Xinput70 S4END[10] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_1
Xinput81 S4END[6] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_3_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout45 FrameStrobe[0] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_230_ Inst_S_CPU_IF_switch_matrix.N4BEG1 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__buf_1
XFILLER_6_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_161_ net27 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_1
X_092_ net1 net38 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit0.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_5_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 FrameData[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
X_213_ Inst_S_CPU_IF_switch_matrix.N2BEG0 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_144_ net13 net44 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_075_ net7 net37 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput191 net202 VGND VGND VPWR VPWR N4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput180 net191 VGND VGND VPWR VPWR N2BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_127_ net26 net43 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_058_ net74 net52 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit21.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N2BEG5 sky130_fd_sc_hd__mux2_1
Xinput71 S4END[11] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_1
Xinput82 S4END[7] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_1
Xinput60 S2END[7] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_1
Xinput93 SS4END[2] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout35 net36 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_0_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_091_ net25 net35 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_160_ net26 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_7_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput3 FrameData[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
X_212_ Inst_S_CPU_IF_switch_matrix.N1BEG3 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__buf_1
X_074_ net6 net37 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_143_ net11 net42 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput192 net203 VGND VGND VPWR VPWR N4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput181 net192 VGND VGND VPWR VPWR N2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput170 net181 VGND VGND VPWR VPWR N1BEG[1] sky130_fd_sc_hd__buf_2
X_057_ net73 net34 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit22.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N2BEG6 sky130_fd_sc_hd__mux2_1
X_126_ net23 net43 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput94 SS4END[3] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__buf_1
Xinput83 S4END[8] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_1
Xinput50 S1END[1] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput72 S4END[12] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_1
Xinput61 S2MID[0] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_109_ net9 net39 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout36 net37 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_090_ net24 net37 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput4 FrameData[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
X_142_ net10 net42 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_211_ Inst_S_CPU_IF_switch_matrix.N1BEG2 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_073_ net5 net35 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_11_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput182 net193 VGND VGND VPWR VPWR N2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput171 net182 VGND VGND VPWR VPWR N1BEG[2] sky130_fd_sc_hd__buf_2
Xoutput193 net204 VGND VGND VPWR VPWR N4BEG[13] sky130_fd_sc_hd__buf_2
XFILLER_7_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput160 net171 VGND VGND VPWR VPWR I_top15 sky130_fd_sc_hd__buf_2
X_056_ net72 net33 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit23.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N2BEG7 sky130_fd_sc_hd__mux2_1
X_125_ net12 net43 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput95 SS4END[4] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_1
Xinput84 S4END[9] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_1
Xinput73 S4END[13] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_1
Xinput51 S1END[2] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_10_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput62 S2MID[1] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_7_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput40 O_top15 VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_1
X_039_ net93 net57 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit8.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N4BEG8 sky130_fd_sc_hd__mux2_1
XFILLER_7_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_108_ net8 net38 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_10_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout37 FrameStrobe[2] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput5 FrameData[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_141_ net9 net44 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_210_ Inst_S_CPU_IF_switch_matrix.N1BEG1 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_072_ net4 net35 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput150 net161 VGND VGND VPWR VPWR FrameStrobe_O[7] sky130_fd_sc_hd__buf_2
Xoutput172 net183 VGND VGND VPWR VPWR N1BEG[3] sky130_fd_sc_hd__buf_2
X_055_ net71 net51 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit24.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N2BEGb0 sky130_fd_sc_hd__mux2_1
Xoutput194 net205 VGND VGND VPWR VPWR N4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput183 net194 VGND VGND VPWR VPWR N2BEGb[2] sky130_fd_sc_hd__buf_2
XFILLER_7_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput161 net172 VGND VGND VPWR VPWR I_top2 sky130_fd_sc_hd__buf_2
X_124_ net1 net43 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit0.Q sky130_fd_sc_hd__dlxtp_1
Xinput96 SS4END[5] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput85 SS4END[0] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_1
Xinput74 S4END[14] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_1
Xinput52 S1END[3] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput63 S2MID[2] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_7_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput41 O_top2 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_2
Xinput30 FrameData[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlymetal6s2s_1
X_038_ net92 net56 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit9.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N4BEG9 sky130_fd_sc_hd__mux2_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_107_ net7 net40 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout38 net39 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_4_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput6 FrameData[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
X_071_ net3 net35 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_140_ net8 net44 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput140 net151 VGND VGND VPWR VPWR FrameStrobe_O[16] sky130_fd_sc_hd__buf_2
Xoutput151 net162 VGND VGND VPWR VPWR FrameStrobe_O[8] sky130_fd_sc_hd__buf_2
Xoutput195 net206 VGND VGND VPWR VPWR N4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput173 net184 VGND VGND VPWR VPWR N2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput184 net195 VGND VGND VPWR VPWR N2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput162 net173 VGND VGND VPWR VPWR I_top3 sky130_fd_sc_hd__buf_2
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput20 FrameData[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
X_054_ net70 net50 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit25.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N2BEGb1 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_123_ net25 net40 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput31 FrameData[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_1
Xinput97 SS4END[6] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_1
Xinput75 S4END[15] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_1
Xinput53 S2END[0] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_1
Xinput86 SS4END[10] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
Xinput64 S2MID[3] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput42 O_top3 VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_2
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_106_ net6 net40 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_037_ net91 net55 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit10.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N4BEG10 sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout39 net40 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
XFILLER_1_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput7 FrameData[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
XFILLER_5_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_070_ net2 net35 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_199_ FrameStrobe[10] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_1
Xoutput141 net152 VGND VGND VPWR VPWR FrameStrobe_O[17] sky130_fd_sc_hd__buf_2
Xoutput152 net163 VGND VGND VPWR VPWR FrameStrobe_O[9] sky130_fd_sc_hd__buf_2
Xoutput196 net207 VGND VGND VPWR VPWR N4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput185 net196 VGND VGND VPWR VPWR N2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput174 net185 VGND VGND VPWR VPWR N2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput163 net174 VGND VGND VPWR VPWR I_top4 sky130_fd_sc_hd__buf_2
Xoutput130 net141 VGND VGND VPWR VPWR FrameData_O[7] sky130_fd_sc_hd__buf_2
XFILLER_7_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_122_ net24 net40 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_053_ net69 net49 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit26.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N2BEGb2 sky130_fd_sc_hd__mux2_1
Xinput98 SS4END[7] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_1
Xinput76 S4END[1] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_1
Xinput54 S2END[1] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_1
Xinput65 S2MID[4] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
Xinput21 FrameData[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
Xinput87 SS4END[11] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_1
XFILLER_6_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput10 FrameData[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
Xinput43 O_top4 VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput32 FrameData[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
X_105_ net5 net40 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_4_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_036_ net90 net54 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit11.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N4BEG11 sky130_fd_sc_hd__mux2_1
XFILLER_8_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_019_ net105 net53 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit28.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.NN4BEG12 sky130_fd_sc_hd__mux2_1
XFILLER_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 FrameData[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
XFILLER_5_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_198_ FrameStrobe[9] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_1
Xoutput142 net153 VGND VGND VPWR VPWR FrameStrobe_O[18] sky130_fd_sc_hd__buf_2
Xoutput186 net197 VGND VGND VPWR VPWR N2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput175 net186 VGND VGND VPWR VPWR N2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput120 net131 VGND VGND VPWR VPWR FrameData_O[27] sky130_fd_sc_hd__buf_2
Xoutput197 net208 VGND VGND VPWR VPWR N4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput164 net175 VGND VGND VPWR VPWR I_top5 sky130_fd_sc_hd__buf_2
Xoutput153 net164 VGND VGND VPWR VPWR I_top0 sky130_fd_sc_hd__buf_2
Xoutput131 net142 VGND VGND VPWR VPWR FrameData_O[8] sky130_fd_sc_hd__buf_2
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_052_ net68 net48 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit27.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N2BEGb3 sky130_fd_sc_hd__mux2_1
X_121_ net22 net41 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput99 SS4END[8] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__buf_1
Xinput55 S2END[2] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_1
Xinput88 SS4END[12] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_1
Xinput77 S4END[2] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_1
Xinput66 S2MID[5] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_1
Xinput22 FrameData[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
Xinput11 FrameData[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_7_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput44 O_top5 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_1
Xinput33 O_top0 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlymetal6s2s_1
X_035_ net89 net53 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit12.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N4BEG12 sky130_fd_sc_hd__mux2_1
XFILLER_8_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_104_ net4 net39 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_018_ net104 net52 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit29.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.NN4BEG13 sky130_fd_sc_hd__mux2_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 FrameData[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_197_ FrameStrobe[8] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput143 net154 VGND VGND VPWR VPWR FrameStrobe_O[19] sky130_fd_sc_hd__buf_2
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput110 net121 VGND VGND VPWR VPWR FrameData_O[18] sky130_fd_sc_hd__buf_2
Xoutput121 net132 VGND VGND VPWR VPWR FrameData_O[28] sky130_fd_sc_hd__buf_2
XFILLER_2_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput132 net143 VGND VGND VPWR VPWR FrameData_O[9] sky130_fd_sc_hd__buf_2
X_120_ net21 net39 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput187 net198 VGND VGND VPWR VPWR N2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput176 net187 VGND VGND VPWR VPWR N2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput198 net209 VGND VGND VPWR VPWR N4BEG[3] sky130_fd_sc_hd__buf_2
X_051_ net67 net47 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit28.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N2BEGb4 sky130_fd_sc_hd__mux2_1
Xoutput165 net176 VGND VGND VPWR VPWR I_top6 sky130_fd_sc_hd__buf_2
Xoutput154 net165 VGND VGND VPWR VPWR I_top1 sky130_fd_sc_hd__buf_2
Xinput89 SS4END[13] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput56 S2END[3] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_1
Xinput78 S4END[3] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_1
Xinput67 S2MID[6] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_7_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_249_ Inst_S_CPU_IF_switch_matrix.NN4BEG4 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__buf_1
Xinput45 O_top6 VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_2
Xinput23 FrameData[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_1
Xinput12 FrameData[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput34 O_top1 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_103_ net3 net39 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_034_ net88 net52 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit13.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N4BEG13 sky130_fd_sc_hd__mux2_1
XFILLER_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_017_ net103 net34 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit30.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.NN4BEG14 sky130_fd_sc_hd__mux2_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_196_ FrameStrobe[7] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput144 net155 VGND VGND VPWR VPWR FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput133 net144 VGND VGND VPWR VPWR FrameStrobe_O[0] sky130_fd_sc_hd__buf_2
Xoutput188 net199 VGND VGND VPWR VPWR N2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput177 net188 VGND VGND VPWR VPWR N2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput122 net133 VGND VGND VPWR VPWR FrameData_O[29] sky130_fd_sc_hd__buf_2
Xoutput199 net210 VGND VGND VPWR VPWR N4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput111 net122 VGND VGND VPWR VPWR FrameData_O[19] sky130_fd_sc_hd__buf_2
X_050_ net66 net46 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit29.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N2BEGb5 sky130_fd_sc_hd__mux2_1
Xoutput155 net166 VGND VGND VPWR VPWR I_top10 sky130_fd_sc_hd__buf_2
Xoutput166 net177 VGND VGND VPWR VPWR I_top7 sky130_fd_sc_hd__buf_2
Xinput79 S4END[4] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_1
Xinput57 S2END[4] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
Xinput68 S2MID[7] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_1
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput24 FrameData[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput13 FrameData[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_7_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_248_ Inst_S_CPU_IF_switch_matrix.NN4BEG3 VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_1
Xinput35 O_top10 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_2
Xinput46 O_top7 VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_1
X_179_ net15 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__buf_1
X_102_ net2 net39 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_033_ net87 net34 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit14.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N4BEG14 sky130_fd_sc_hd__mux2_1
XFILLER_8_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_016_ net96 net33 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit31.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.NN4BEG15 sky130_fd_sc_hd__mux2_1
XFILLER_3_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_195_ FrameStrobe[6] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_1
Xoutput134 net145 VGND VGND VPWR VPWR FrameStrobe_O[10] sky130_fd_sc_hd__buf_2
Xoutput145 net156 VGND VGND VPWR VPWR FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
Xoutput178 net189 VGND VGND VPWR VPWR N2BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput189 net200 VGND VGND VPWR VPWR N4BEG[0] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_6_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput167 net178 VGND VGND VPWR VPWR I_top8 sky130_fd_sc_hd__buf_2
Xoutput156 net167 VGND VGND VPWR VPWR I_top11 sky130_fd_sc_hd__buf_2
Xoutput123 net134 VGND VGND VPWR VPWR FrameData_O[2] sky130_fd_sc_hd__buf_2
Xoutput112 net123 VGND VGND VPWR VPWR FrameData_O[1] sky130_fd_sc_hd__buf_2
Xoutput101 net112 VGND VGND VPWR VPWR FrameData_O[0] sky130_fd_sc_hd__buf_2
Xinput25 FrameData[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput14 FrameData[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
Xinput36 O_top11 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_1
X_247_ Inst_S_CPU_IF_switch_matrix.NN4BEG2 VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__buf_1
Xinput69 S4END[0] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
Xinput58 S2END[5] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_1
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput47 O_top8 VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_1
X_178_ net14 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_1
X_101_ net32 net38 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_032_ net80 net33 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit15.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N4BEG15 sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_9_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_015_ net60 net72 net80 net96 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit0.Q Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit1.Q
+ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__mux4_1
XFILLER_8_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_194_ FrameStrobe[5] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput146 net157 VGND VGND VPWR VPWR FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
Xoutput179 net190 VGND VGND VPWR VPWR N2BEG[6] sky130_fd_sc_hd__buf_2
Xoutput135 net146 VGND VGND VPWR VPWR FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
Xoutput113 net124 VGND VGND VPWR VPWR FrameData_O[20] sky130_fd_sc_hd__buf_2
Xoutput124 net135 VGND VGND VPWR VPWR FrameData_O[30] sky130_fd_sc_hd__buf_2
Xoutput168 net179 VGND VGND VPWR VPWR I_top9 sky130_fd_sc_hd__buf_2
Xoutput157 net168 VGND VGND VPWR VPWR I_top12 sky130_fd_sc_hd__buf_2
Xoutput102 net113 VGND VGND VPWR VPWR FrameData_O[10] sky130_fd_sc_hd__buf_2
Xinput59 S2END[6] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_1
X_246_ Inst_S_CPU_IF_switch_matrix.NN4BEG1 VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__buf_1
Xinput15 FrameData[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
Xinput37 O_top12 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_1
Xinput48 O_top9 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_1
Xinput26 FrameData[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_1
X_177_ net13 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__buf_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_100_ net31 net38 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_031_ net102 net51 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit16.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.NN4BEG0 sky130_fd_sc_hd__mux2_1
X_229_ Inst_S_CPU_IF_switch_matrix.N4BEG0 VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_014_ net61 net73 net87 net103 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit2.Q Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit3.Q
+ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__mux4_1
XS_CPU_IF_222 VGND VGND VPWR VPWR S_CPU_IF_222/HI Co sky130_fd_sc_hd__conb_1
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_193_ FrameStrobe[4] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput136 net147 VGND VGND VPWR VPWR FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
Xoutput147 net158 VGND VGND VPWR VPWR FrameStrobe_O[4] sky130_fd_sc_hd__buf_2
Xoutput169 net180 VGND VGND VPWR VPWR N1BEG[0] sky130_fd_sc_hd__buf_2
Xoutput125 net136 VGND VGND VPWR VPWR FrameData_O[31] sky130_fd_sc_hd__buf_2
Xoutput114 net125 VGND VGND VPWR VPWR FrameData_O[21] sky130_fd_sc_hd__buf_2
Xoutput103 net114 VGND VGND VPWR VPWR FrameData_O[11] sky130_fd_sc_hd__buf_2
Xoutput158 net169 VGND VGND VPWR VPWR I_top13 sky130_fd_sc_hd__buf_2
Xinput49 S1END[0] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_1
Xinput16 FrameData[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_245_ Inst_S_CPU_IF_switch_matrix.NN4BEG0 VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_1
X_176_ net11 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
Xinput38 O_top13 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_1
Xinput27 FrameData[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlymetal6s2s_1
X_030_ net101 net50 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit17.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.NN4BEG1 sky130_fd_sc_hd__mux2_1
XFILLER_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_228_ Inst_S_CPU_IF_switch_matrix.N2BEGb7 VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_159_ net23 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_013_ net62 net74 net88 net104 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit4.Q Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit5.Q
+ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__mux4_1
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_192_ FrameStrobe[3] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_1
X_261_ UserCLK VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__buf_2
Xoutput148 net159 VGND VGND VPWR VPWR FrameStrobe_O[5] sky130_fd_sc_hd__buf_2
Xoutput115 net126 VGND VGND VPWR VPWR FrameData_O[22] sky130_fd_sc_hd__buf_2
Xoutput137 net148 VGND VGND VPWR VPWR FrameStrobe_O[13] sky130_fd_sc_hd__buf_2
XFILLER_1_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput159 net170 VGND VGND VPWR VPWR I_top14 sky130_fd_sc_hd__buf_2
XFILLER_1_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput126 net137 VGND VGND VPWR VPWR FrameData_O[3] sky130_fd_sc_hd__buf_2
Xoutput104 net115 VGND VGND VPWR VPWR FrameData_O[12] sky130_fd_sc_hd__buf_2
XFILLER_11_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput17 FrameData[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput39 O_top14 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
X_175_ net10 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
Xinput28 FrameData[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_2
X_244_ Inst_S_CPU_IF_switch_matrix.N4BEG15 VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_089_ net22 net37 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_158_ net12 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__buf_1
X_227_ Inst_S_CPU_IF_switch_matrix.N2BEGb6 VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__buf_1
X_012_ net63 net75 net89 net105 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit6.Q Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit7.Q
+ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_260_ Inst_S_CPU_IF_switch_matrix.NN4BEG15 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_191_ net37 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_1
Xoutput138 net149 VGND VGND VPWR VPWR FrameStrobe_O[14] sky130_fd_sc_hd__buf_2
Xoutput149 net160 VGND VGND VPWR VPWR FrameStrobe_O[6] sky130_fd_sc_hd__buf_2
Xoutput116 net127 VGND VGND VPWR VPWR FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput105 net116 VGND VGND VPWR VPWR FrameData_O[13] sky130_fd_sc_hd__buf_2
Xoutput127 net138 VGND VGND VPWR VPWR FrameData_O[4] sky130_fd_sc_hd__buf_2
XFILLER_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput18 FrameData[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
X_174_ net9 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_1
Xinput29 FrameData[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_1
X_243_ Inst_S_CPU_IF_switch_matrix.N4BEG14 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_226_ Inst_S_CPU_IF_switch_matrix.N2BEGb5 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_2
X_088_ net21 net37 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_157_ net1 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_8_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_011_ net60 net64 net90 net106 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit8.Q Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit9.Q
+ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__mux4_1
XFILLER_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_209_ Inst_S_CPU_IF_switch_matrix.N1BEG0 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_190_ net41 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_1
Xoutput117 net128 VGND VGND VPWR VPWR FrameData_O[24] sky130_fd_sc_hd__buf_2
Xoutput139 net150 VGND VGND VPWR VPWR FrameStrobe_O[15] sky130_fd_sc_hd__buf_2
XFILLER_9_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput106 net117 VGND VGND VPWR VPWR FrameData_O[14] sky130_fd_sc_hd__buf_2
Xoutput128 net139 VGND VGND VPWR VPWR FrameData_O[5] sky130_fd_sc_hd__buf_2
Xinput19 FrameData[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_1
X_173_ net8 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_1_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_242_ Inst_S_CPU_IF_switch_matrix.N4BEG13 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__buf_1
XFILLER_10_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_225_ Inst_S_CPU_IF_switch_matrix.N2BEGb4 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__buf_1
XFILLER_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_087_ net20 net36 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_010_ net61 net65 net91 net107 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit10.Q Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit11.Q
+ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__mux4_1
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_208_ FrameStrobe[19] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_1
X_139_ net7 net42 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_5_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput118 net129 VGND VGND VPWR VPWR FrameData_O[25] sky130_fd_sc_hd__buf_2
XFILLER_9_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput107 net118 VGND VGND VPWR VPWR FrameData_O[15] sky130_fd_sc_hd__buf_2
Xoutput129 net140 VGND VGND VPWR VPWR FrameData_O[6] sky130_fd_sc_hd__buf_2
X_241_ Inst_S_CPU_IF_switch_matrix.N4BEG12 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_172_ net7 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_1
X_224_ Inst_S_CPU_IF_switch_matrix.N2BEGb3 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__buf_1
XFILLER_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_155_ net25 net42 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_086_ net19 net36 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_8_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_069_ net32 net36 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_138_ net6 net42 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_207_ FrameStrobe[18] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput119 net130 VGND VGND VPWR VPWR FrameData_O[26] sky130_fd_sc_hd__buf_2
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput108 net119 VGND VGND VPWR VPWR FrameData_O[16] sky130_fd_sc_hd__buf_2
XFILLER_1_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_240_ Inst_S_CPU_IF_switch_matrix.N4BEG11 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_171_ net6 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__buf_1
X_223_ Inst_S_CPU_IF_switch_matrix.N2BEGb2 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_085_ net18 net35 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_154_ net24 net45 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_206_ FrameStrobe[17] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_1
X_068_ net31 net36 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_137_ net5 net44 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput109 net120 VGND VGND VPWR VPWR FrameData_O[17] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_170_ net5 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__buf_1
XFILLER_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_084_ net17 net36 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_222_ Inst_S_CPU_IF_switch_matrix.N2BEGb1 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__buf_1
X_153_ net22 net45 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_205_ FrameStrobe[16] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_1
X_136_ net4 net44 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_067_ net63 net53 net57 net51 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit8.Q Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit9.Q
+ VGND VGND VPWR VPWR Inst_S_CPU_IF_switch_matrix.N1BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_2_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_119_ net20 net40 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_4_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_221_ Inst_S_CPU_IF_switch_matrix.N2BEGb0 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_1
X_152_ net21 net45 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_083_ net16 net35 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_204_ FrameStrobe[15] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_1
X_066_ net62 net52 net56 net50 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit10.Q Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit11.Q
+ VGND VGND VPWR VPWR Inst_S_CPU_IF_switch_matrix.N1BEG1 sky130_fd_sc_hd__mux4_1
X_135_ net3 net42 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_049_ net65 net59 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit30.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N2BEGb6 sky130_fd_sc_hd__mux2_1
X_118_ net19 net39 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_1 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_151_ net20 net43 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_082_ net15 net35 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_220_ Inst_S_CPU_IF_switch_matrix.N2BEG7 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__buf_1
X_203_ FrameStrobe[14] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_065_ net61 net34 net55 net49 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit12.Q Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit13.Q
+ VGND VGND VPWR VPWR Inst_S_CPU_IF_switch_matrix.N1BEG2 sky130_fd_sc_hd__mux4_1
X_134_ net2 net42 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_11_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_117_ net18 net39 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_048_ net64 net58 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit31.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N2BEGb7 sky130_fd_sc_hd__mux2_1
XANTENNA_2 FrameStrobe[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_150_ net19 net45 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_081_ net14 net36 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_202_ FrameStrobe[13] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_1
X_133_ net32 net43 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_064_ net60 net33 net54 net48 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit14.Q Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit15.Q
+ VGND VGND VPWR VPWR Inst_S_CPU_IF_switch_matrix.N1BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_116_ net17 net38 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_047_ net86 net51 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit0.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N4BEG0 sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_3 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_080_ net13 net35 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_8_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_132_ net31 net43 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_063_ net79 net57 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit16.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N2BEG0 sky130_fd_sc_hd__mux2_1
X_201_ FrameStrobe[12] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_046_ net85 net50 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit1.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.N4BEG1 sky130_fd_sc_hd__mux2_1
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_115_ net16 net41 VGND VGND VPWR VPWR Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_4 net195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_029_ net100 net49 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit18.Q VGND VGND VPWR VPWR
+ Inst_S_CPU_IF_switch_matrix.NN4BEG2 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

