magic
tech sky130A
magscale 1 2
timestamp 1740383317
<< viali >>
rect 1409 8585 1443 8619
rect 3893 8585 3927 8619
rect 5733 8585 5767 8619
rect 7849 8585 7883 8619
rect 9965 8585 9999 8619
rect 12081 8585 12115 8619
rect 14197 8585 14231 8619
rect 16313 8585 16347 8619
rect 18429 8585 18463 8619
rect 20545 8585 20579 8619
rect 22661 8585 22695 8619
rect 24777 8585 24811 8619
rect 27077 8585 27111 8619
rect 29009 8585 29043 8619
rect 31125 8585 31159 8619
rect 33241 8585 33275 8619
rect 35449 8585 35483 8619
rect 37473 8585 37507 8619
rect 40049 8585 40083 8619
rect 41429 8585 41463 8619
rect 41797 8585 41831 8619
rect 42165 8585 42199 8619
rect 42717 8585 42751 8619
rect 1593 8449 1627 8483
rect 4077 8449 4111 8483
rect 5917 8449 5951 8483
rect 8033 8449 8067 8483
rect 10149 8449 10183 8483
rect 12265 8449 12299 8483
rect 14381 8449 14415 8483
rect 16497 8449 16531 8483
rect 18613 8449 18647 8483
rect 20729 8449 20763 8483
rect 22845 8449 22879 8483
rect 24961 8449 24995 8483
rect 27261 8449 27295 8483
rect 29193 8449 29227 8483
rect 31309 8449 31343 8483
rect 33425 8449 33459 8483
rect 35265 8449 35299 8483
rect 37657 8449 37691 8483
rect 39865 8449 39899 8483
rect 41245 8449 41279 8483
rect 41613 8449 41647 8483
rect 41981 8449 42015 8483
rect 42533 8449 42567 8483
rect 42901 8449 42935 8483
rect 43269 8449 43303 8483
rect 43085 8313 43119 8347
rect 43453 8313 43487 8347
rect 17509 8041 17543 8075
rect 17877 8041 17911 8075
rect 21373 8041 21407 8075
rect 23765 8041 23799 8075
rect 24593 8041 24627 8075
rect 26341 8041 26375 8075
rect 26709 8041 26743 8075
rect 41981 8041 42015 8075
rect 42349 8041 42383 8075
rect 42717 8041 42751 8075
rect 20545 7973 20579 8007
rect 20729 7973 20763 8007
rect 21097 7973 21131 8007
rect 3801 7837 3835 7871
rect 4169 7837 4203 7871
rect 16037 7837 16071 7871
rect 17601 7837 17635 7871
rect 17693 7837 17727 7871
rect 19349 7837 19383 7871
rect 19625 7837 19659 7871
rect 20361 7837 20395 7871
rect 20821 7837 20855 7871
rect 20913 7837 20947 7871
rect 21189 7837 21223 7871
rect 23489 7837 23523 7871
rect 23581 7837 23615 7871
rect 24409 7837 24443 7871
rect 24685 7837 24719 7871
rect 26433 7837 26467 7871
rect 26525 7837 26559 7871
rect 26985 7837 27019 7871
rect 27077 7837 27111 7871
rect 27537 7837 27571 7871
rect 28365 7837 28399 7871
rect 29561 7837 29595 7871
rect 29837 7837 29871 7871
rect 41797 7837 41831 7871
rect 42165 7837 42199 7871
rect 42533 7837 42567 7871
rect 42901 7837 42935 7871
rect 43269 7837 43303 7871
rect 3985 7701 4019 7735
rect 4353 7701 4387 7735
rect 16221 7701 16255 7735
rect 19533 7701 19567 7735
rect 21465 7701 21499 7735
rect 23489 7701 23523 7735
rect 26893 7701 26927 7735
rect 27261 7701 27295 7735
rect 27353 7701 27387 7735
rect 28181 7701 28215 7735
rect 29745 7701 29779 7735
rect 43085 7701 43119 7735
rect 43453 7701 43487 7735
rect 43085 7497 43119 7531
rect 18889 7361 18923 7395
rect 18981 7361 19015 7395
rect 22017 7361 22051 7395
rect 31217 7361 31251 7395
rect 42901 7361 42935 7395
rect 43269 7361 43303 7395
rect 18797 7293 18831 7327
rect 19165 7225 19199 7259
rect 22201 7157 22235 7191
rect 31033 7157 31067 7191
rect 43453 7157 43487 7191
rect 9597 6885 9631 6919
rect 25329 6885 25363 6919
rect 1961 6749 1995 6783
rect 9413 6749 9447 6783
rect 12909 6749 12943 6783
rect 15853 6749 15887 6783
rect 16129 6749 16163 6783
rect 22845 6749 22879 6783
rect 25053 6749 25087 6783
rect 25145 6749 25179 6783
rect 26985 6749 27019 6783
rect 27169 6749 27203 6783
rect 29929 6749 29963 6783
rect 30021 6749 30055 6783
rect 34897 6749 34931 6783
rect 42901 6749 42935 6783
rect 43269 6749 43303 6783
rect 24961 6681 24995 6715
rect 2145 6613 2179 6647
rect 13093 6613 13127 6647
rect 16037 6613 16071 6647
rect 16313 6613 16347 6647
rect 23029 6613 23063 6647
rect 27353 6613 27387 6647
rect 29837 6613 29871 6647
rect 30205 6613 30239 6647
rect 35081 6613 35115 6647
rect 43085 6613 43119 6647
rect 43453 6613 43487 6647
rect 9229 6409 9263 6443
rect 17693 6409 17727 6443
rect 18061 6409 18095 6443
rect 21189 6409 21223 6443
rect 25513 6409 25547 6443
rect 31769 6409 31803 6443
rect 37749 6409 37783 6443
rect 38485 6409 38519 6443
rect 41337 6409 41371 6443
rect 43453 6409 43487 6443
rect 5917 6273 5951 6307
rect 9137 6273 9171 6307
rect 9413 6273 9447 6307
rect 10885 6273 10919 6307
rect 13737 6273 13771 6307
rect 17785 6273 17819 6307
rect 17877 6273 17911 6307
rect 20361 6273 20395 6307
rect 21281 6273 21315 6307
rect 21373 6273 21407 6307
rect 25697 6273 25731 6307
rect 31401 6273 31435 6307
rect 31953 6273 31987 6307
rect 37933 6273 37967 6307
rect 38301 6273 38335 6307
rect 39129 6273 39163 6307
rect 41153 6273 41187 6307
rect 42901 6273 42935 6307
rect 43269 6273 43303 6307
rect 39313 6137 39347 6171
rect 6101 6069 6135 6103
rect 11069 6069 11103 6103
rect 13921 6069 13955 6103
rect 20545 6069 20579 6103
rect 21557 6069 21591 6103
rect 31217 6069 31251 6103
rect 43085 6069 43119 6103
rect 15209 5865 15243 5899
rect 15485 5865 15519 5899
rect 18705 5797 18739 5831
rect 21649 5797 21683 5831
rect 33701 5797 33735 5831
rect 43453 5797 43487 5831
rect 6653 5661 6687 5695
rect 15025 5661 15059 5695
rect 15301 5661 15335 5695
rect 18521 5661 18555 5695
rect 21465 5661 21499 5695
rect 26249 5661 26283 5695
rect 28365 5661 28399 5695
rect 30941 5661 30975 5695
rect 33885 5661 33919 5695
rect 35265 5661 35299 5695
rect 35541 5661 35575 5695
rect 42901 5661 42935 5695
rect 43269 5661 43303 5695
rect 6837 5525 6871 5559
rect 26065 5525 26099 5559
rect 28549 5525 28583 5559
rect 30757 5525 30791 5559
rect 35173 5525 35207 5559
rect 35357 5525 35391 5559
rect 43085 5525 43119 5559
rect 22017 5321 22051 5355
rect 23213 5321 23247 5355
rect 25881 5321 25915 5355
rect 36921 5321 36955 5355
rect 43453 5321 43487 5355
rect 2329 5185 2363 5219
rect 3985 5185 4019 5219
rect 9689 5185 9723 5219
rect 9965 5185 9999 5219
rect 17601 5185 17635 5219
rect 17693 5185 17727 5219
rect 18153 5185 18187 5219
rect 21833 5185 21867 5219
rect 22109 5185 22143 5219
rect 23305 5185 23339 5219
rect 23397 5185 23431 5219
rect 25697 5185 25731 5219
rect 26065 5185 26099 5219
rect 27353 5185 27387 5219
rect 27537 5185 27571 5219
rect 33241 5185 33275 5219
rect 33609 5185 33643 5219
rect 37105 5185 37139 5219
rect 37473 5185 37507 5219
rect 37565 5185 37599 5219
rect 42901 5185 42935 5219
rect 43269 5185 43303 5219
rect 9781 5049 9815 5083
rect 26249 5049 26283 5083
rect 27721 5049 27755 5083
rect 2513 4981 2547 5015
rect 4169 4981 4203 5015
rect 17509 4981 17543 5015
rect 17877 4981 17911 5015
rect 18337 4981 18371 5015
rect 23581 4981 23615 5015
rect 33425 4981 33459 5015
rect 37289 4981 37323 5015
rect 37565 4981 37599 5015
rect 43085 4981 43119 5015
rect 17509 4777 17543 4811
rect 30113 4777 30147 4811
rect 26341 4709 26375 4743
rect 26985 4709 27019 4743
rect 43453 4709 43487 4743
rect 28273 4641 28307 4675
rect 7297 4573 7331 4607
rect 13461 4573 13495 4607
rect 17325 4573 17359 4607
rect 22201 4573 22235 4607
rect 26433 4573 26467 4607
rect 26525 4573 26559 4607
rect 26801 4573 26835 4607
rect 28365 4573 28399 4607
rect 28457 4573 28491 4607
rect 30297 4573 30331 4607
rect 42901 4573 42935 4607
rect 43269 4573 43303 4607
rect 27077 4505 27111 4539
rect 7481 4437 7515 4471
rect 13277 4437 13311 4471
rect 22385 4437 22419 4471
rect 26709 4437 26743 4471
rect 28641 4437 28675 4471
rect 43085 4437 43119 4471
rect 2053 4097 2087 4131
rect 4077 4097 4111 4131
rect 17141 4097 17175 4131
rect 17417 4097 17451 4131
rect 24225 4097 24259 4131
rect 27721 4097 27755 4131
rect 32413 4097 32447 4131
rect 42901 4097 42935 4131
rect 43269 4097 43303 4131
rect 2237 3961 2271 3995
rect 27905 3961 27939 3995
rect 43453 3961 43487 3995
rect 4261 3893 4295 3927
rect 17233 3893 17267 3927
rect 24409 3893 24443 3927
rect 32229 3893 32263 3927
rect 43085 3893 43119 3927
rect 21833 3689 21867 3723
rect 23489 3689 23523 3723
rect 23765 3689 23799 3723
rect 30297 3689 30331 3723
rect 20177 3621 20211 3655
rect 24685 3621 24719 3655
rect 25053 3621 25087 3655
rect 43453 3621 43487 3655
rect 15485 3485 15519 3519
rect 18705 3485 18739 3519
rect 19533 3485 19567 3519
rect 19717 3485 19751 3519
rect 19993 3485 20027 3519
rect 20269 3485 20303 3519
rect 22017 3485 22051 3519
rect 23489 3485 23523 3519
rect 23581 3485 23615 3519
rect 24777 3485 24811 3519
rect 24869 3485 24903 3519
rect 27537 3485 27571 3519
rect 30113 3485 30147 3519
rect 32413 3485 32447 3519
rect 42901 3485 42935 3519
rect 43269 3485 43303 3519
rect 15669 3349 15703 3383
rect 18889 3349 18923 3383
rect 19901 3349 19935 3383
rect 27353 3349 27387 3383
rect 32229 3349 32263 3383
rect 43085 3349 43119 3383
rect 12633 3145 12667 3179
rect 30205 3145 30239 3179
rect 30573 3145 30607 3179
rect 31769 3145 31803 3179
rect 34253 3145 34287 3179
rect 36829 3145 36863 3179
rect 38117 3145 38151 3179
rect 43453 3145 43487 3179
rect 1869 3009 1903 3043
rect 7573 3009 7607 3043
rect 12449 3009 12483 3043
rect 14565 3009 14599 3043
rect 15945 3009 15979 3043
rect 16313 3009 16347 3043
rect 20085 3009 20119 3043
rect 21189 3009 21223 3043
rect 22017 3009 22051 3043
rect 25329 3009 25363 3043
rect 25881 3009 25915 3043
rect 26709 3009 26743 3043
rect 27169 3009 27203 3043
rect 27261 3009 27295 3043
rect 27537 3009 27571 3043
rect 28365 3009 28399 3043
rect 28733 3009 28767 3043
rect 30021 3009 30055 3043
rect 30297 3009 30331 3043
rect 30389 3009 30423 3043
rect 31137 3009 31171 3043
rect 31401 3009 31435 3043
rect 31585 3009 31619 3043
rect 32413 3009 32447 3043
rect 32505 3009 32539 3043
rect 32781 3009 32815 3043
rect 33057 3009 33091 3043
rect 33241 3009 33275 3043
rect 33609 3009 33643 3043
rect 34161 3009 34195 3043
rect 34437 3009 34471 3043
rect 34713 3009 34747 3043
rect 34805 3009 34839 3043
rect 35173 3009 35207 3043
rect 35725 3009 35759 3043
rect 36093 3009 36127 3043
rect 37013 3009 37047 3043
rect 38301 3009 38335 3043
rect 42533 3009 42567 3043
rect 42901 3009 42935 3043
rect 43269 3009 43303 3043
rect 27077 2941 27111 2975
rect 16129 2873 16163 2907
rect 16497 2873 16531 2907
rect 27445 2873 27479 2907
rect 32321 2873 32355 2907
rect 32689 2873 32723 2907
rect 34529 2873 34563 2907
rect 35909 2873 35943 2907
rect 2053 2805 2087 2839
rect 7757 2805 7791 2839
rect 14749 2805 14783 2839
rect 20269 2805 20303 2839
rect 21373 2805 21407 2839
rect 22201 2805 22235 2839
rect 25513 2805 25547 2839
rect 26065 2805 26099 2839
rect 26525 2805 26559 2839
rect 27721 2805 27755 2839
rect 28549 2805 28583 2839
rect 28917 2805 28951 2839
rect 29837 2805 29871 2839
rect 30941 2805 30975 2839
rect 31401 2805 31435 2839
rect 32965 2805 32999 2839
rect 33425 2805 33459 2839
rect 33793 2805 33827 2839
rect 34069 2805 34103 2839
rect 34989 2805 35023 2839
rect 42717 2805 42751 2839
rect 43085 2805 43119 2839
rect 24961 2601 24995 2635
rect 25329 2601 25363 2635
rect 28273 2601 28307 2635
rect 31677 2601 31711 2635
rect 33793 2601 33827 2635
rect 26433 2533 26467 2567
rect 27537 2533 27571 2567
rect 28641 2533 28675 2567
rect 29745 2533 29779 2567
rect 30757 2533 30791 2567
rect 32597 2533 32631 2567
rect 43453 2533 43487 2567
rect 19533 2397 19567 2431
rect 19901 2397 19935 2431
rect 20269 2397 20303 2431
rect 20637 2397 20671 2431
rect 21005 2397 21039 2431
rect 21373 2397 21407 2431
rect 21833 2397 21867 2431
rect 22201 2397 22235 2431
rect 22569 2397 22603 2431
rect 22937 2397 22971 2431
rect 23305 2397 23339 2431
rect 23673 2397 23707 2431
rect 24409 2397 24443 2431
rect 24777 2397 24811 2431
rect 25145 2397 25179 2431
rect 25513 2397 25547 2431
rect 25881 2397 25915 2431
rect 26249 2397 26283 2431
rect 27261 2397 27295 2431
rect 27353 2397 27387 2431
rect 27721 2397 27755 2431
rect 28089 2397 28123 2431
rect 28457 2397 28491 2431
rect 28825 2397 28859 2431
rect 29561 2397 29595 2431
rect 29929 2397 29963 2431
rect 30297 2397 30331 2431
rect 30941 2397 30975 2431
rect 31493 2397 31527 2431
rect 31861 2397 31895 2431
rect 32413 2397 32447 2431
rect 32781 2397 32815 2431
rect 33149 2397 33183 2431
rect 33241 2397 33275 2431
rect 33609 2397 33643 2431
rect 33977 2397 34011 2431
rect 34713 2397 34747 2431
rect 35081 2397 35115 2431
rect 41981 2397 42015 2431
rect 42533 2397 42567 2431
rect 42901 2397 42935 2431
rect 43269 2397 43303 2431
rect 19717 2261 19751 2295
rect 20085 2261 20119 2295
rect 20453 2261 20487 2295
rect 20821 2261 20855 2295
rect 21189 2261 21223 2295
rect 21557 2261 21591 2295
rect 22017 2261 22051 2295
rect 22385 2261 22419 2295
rect 22753 2261 22787 2295
rect 23121 2261 23155 2295
rect 23489 2261 23523 2295
rect 23857 2261 23891 2295
rect 24593 2261 24627 2295
rect 25697 2261 25731 2295
rect 26065 2261 26099 2295
rect 27077 2261 27111 2295
rect 27905 2261 27939 2295
rect 29009 2261 29043 2295
rect 30113 2261 30147 2295
rect 30481 2261 30515 2295
rect 31309 2261 31343 2295
rect 32229 2261 32263 2295
rect 32965 2261 32999 2295
rect 33425 2261 33459 2295
rect 34161 2261 34195 2295
rect 34897 2261 34931 2295
rect 35265 2261 35299 2295
rect 42165 2261 42199 2295
rect 42717 2261 42751 2295
rect 43085 2261 43119 2295
<< metal1 >>
rect 25866 9160 25872 9172
rect 22066 9132 25872 9160
rect 16482 9052 16488 9104
rect 16540 9092 16546 9104
rect 22066 9092 22094 9132
rect 25866 9120 25872 9132
rect 25924 9120 25930 9172
rect 25498 9092 25504 9104
rect 16540 9064 22094 9092
rect 24780 9064 25504 9092
rect 16540 9052 16546 9064
rect 18598 8984 18604 9036
rect 18656 9024 18662 9036
rect 24780 9024 24808 9064
rect 25498 9052 25504 9064
rect 25556 9052 25562 9104
rect 18656 8996 24808 9024
rect 18656 8984 18662 8996
rect 24854 8984 24860 9036
rect 24912 9024 24918 9036
rect 24912 8996 31754 9024
rect 24912 8984 24918 8996
rect 22066 8928 22876 8956
rect 22066 8888 22094 8928
rect 12406 8860 22094 8888
rect 22848 8888 22876 8928
rect 22922 8916 22928 8968
rect 22980 8956 22986 8968
rect 26142 8956 26148 8968
rect 22980 8928 26148 8956
rect 22980 8916 22986 8928
rect 26142 8916 26148 8928
rect 26200 8916 26206 8968
rect 31726 8956 31754 8996
rect 31726 8928 43944 8956
rect 31846 8888 31852 8900
rect 22848 8860 31852 8888
rect 12250 8780 12256 8832
rect 12308 8820 12314 8832
rect 12406 8820 12434 8860
rect 31846 8848 31852 8860
rect 31904 8848 31910 8900
rect 12308 8792 12434 8820
rect 12308 8780 12314 8792
rect 20714 8780 20720 8832
rect 20772 8820 20778 8832
rect 22738 8820 22744 8832
rect 20772 8792 22744 8820
rect 20772 8780 20778 8792
rect 22738 8780 22744 8792
rect 22796 8780 22802 8832
rect 22830 8780 22836 8832
rect 22888 8820 22894 8832
rect 31018 8820 31024 8832
rect 22888 8792 31024 8820
rect 22888 8780 22894 8792
rect 31018 8780 31024 8792
rect 31076 8780 31082 8832
rect 41414 8780 41420 8832
rect 41472 8820 41478 8832
rect 43622 8820 43628 8832
rect 41472 8792 43628 8820
rect 41472 8780 41478 8792
rect 43622 8780 43628 8792
rect 43680 8780 43686 8832
rect 1104 8730 43884 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 39010 8730
rect 39062 8678 39074 8730
rect 39126 8678 39138 8730
rect 39190 8678 39202 8730
rect 39254 8678 39266 8730
rect 39318 8678 43884 8730
rect 1104 8656 43884 8678
rect 1302 8576 1308 8628
rect 1360 8616 1366 8628
rect 1397 8619 1455 8625
rect 1397 8616 1409 8619
rect 1360 8588 1409 8616
rect 1360 8576 1366 8588
rect 1397 8585 1409 8588
rect 1443 8585 1455 8619
rect 1397 8579 1455 8585
rect 3418 8576 3424 8628
rect 3476 8616 3482 8628
rect 3881 8619 3939 8625
rect 3881 8616 3893 8619
rect 3476 8588 3893 8616
rect 3476 8576 3482 8588
rect 3881 8585 3893 8588
rect 3927 8585 3939 8619
rect 3881 8579 3939 8585
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 5721 8619 5779 8625
rect 5721 8616 5733 8619
rect 5592 8588 5733 8616
rect 5592 8576 5598 8588
rect 5721 8585 5733 8588
rect 5767 8585 5779 8619
rect 5721 8579 5779 8585
rect 7650 8576 7656 8628
rect 7708 8616 7714 8628
rect 7837 8619 7895 8625
rect 7837 8616 7849 8619
rect 7708 8588 7849 8616
rect 7708 8576 7714 8588
rect 7837 8585 7849 8588
rect 7883 8585 7895 8619
rect 7837 8579 7895 8585
rect 9766 8576 9772 8628
rect 9824 8616 9830 8628
rect 9953 8619 10011 8625
rect 9953 8616 9965 8619
rect 9824 8588 9965 8616
rect 9824 8576 9830 8588
rect 9953 8585 9965 8588
rect 9999 8585 10011 8619
rect 9953 8579 10011 8585
rect 11882 8576 11888 8628
rect 11940 8616 11946 8628
rect 12069 8619 12127 8625
rect 12069 8616 12081 8619
rect 11940 8588 12081 8616
rect 11940 8576 11946 8588
rect 12069 8585 12081 8588
rect 12115 8585 12127 8619
rect 12069 8579 12127 8585
rect 12250 8576 12256 8628
rect 12308 8576 12314 8628
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 14185 8619 14243 8625
rect 14185 8616 14197 8619
rect 14056 8588 14197 8616
rect 14056 8576 14062 8588
rect 14185 8585 14197 8588
rect 14231 8585 14243 8619
rect 14185 8579 14243 8585
rect 16114 8576 16120 8628
rect 16172 8616 16178 8628
rect 16301 8619 16359 8625
rect 16301 8616 16313 8619
rect 16172 8588 16313 8616
rect 16172 8576 16178 8588
rect 16301 8585 16313 8588
rect 16347 8585 16359 8619
rect 16301 8579 16359 8585
rect 18230 8576 18236 8628
rect 18288 8616 18294 8628
rect 18417 8619 18475 8625
rect 18417 8616 18429 8619
rect 18288 8588 18429 8616
rect 18288 8576 18294 8588
rect 18417 8585 18429 8588
rect 18463 8585 18475 8619
rect 18417 8579 18475 8585
rect 20346 8576 20352 8628
rect 20404 8616 20410 8628
rect 20533 8619 20591 8625
rect 20533 8616 20545 8619
rect 20404 8588 20545 8616
rect 20404 8576 20410 8588
rect 20533 8585 20545 8588
rect 20579 8585 20591 8619
rect 20533 8579 20591 8585
rect 22462 8576 22468 8628
rect 22520 8616 22526 8628
rect 22649 8619 22707 8625
rect 22649 8616 22661 8619
rect 22520 8588 22661 8616
rect 22520 8576 22526 8588
rect 22649 8585 22661 8588
rect 22695 8585 22707 8619
rect 22649 8579 22707 8585
rect 24578 8576 24584 8628
rect 24636 8616 24642 8628
rect 24765 8619 24823 8625
rect 24765 8616 24777 8619
rect 24636 8588 24777 8616
rect 24636 8576 24642 8588
rect 24765 8585 24777 8588
rect 24811 8585 24823 8619
rect 24765 8579 24823 8585
rect 26694 8576 26700 8628
rect 26752 8616 26758 8628
rect 27065 8619 27123 8625
rect 27065 8616 27077 8619
rect 26752 8588 27077 8616
rect 26752 8576 26758 8588
rect 27065 8585 27077 8588
rect 27111 8585 27123 8619
rect 27065 8579 27123 8585
rect 27154 8576 27160 8628
rect 27212 8616 27218 8628
rect 28718 8616 28724 8628
rect 27212 8588 28724 8616
rect 27212 8576 27218 8588
rect 28718 8576 28724 8588
rect 28776 8576 28782 8628
rect 28810 8576 28816 8628
rect 28868 8616 28874 8628
rect 28997 8619 29055 8625
rect 28997 8616 29009 8619
rect 28868 8588 29009 8616
rect 28868 8576 28874 8588
rect 28997 8585 29009 8588
rect 29043 8585 29055 8619
rect 28997 8579 29055 8585
rect 30926 8576 30932 8628
rect 30984 8616 30990 8628
rect 31113 8619 31171 8625
rect 31113 8616 31125 8619
rect 30984 8588 31125 8616
rect 30984 8576 30990 8588
rect 31113 8585 31125 8588
rect 31159 8585 31171 8619
rect 31113 8579 31171 8585
rect 32858 8576 32864 8628
rect 32916 8616 32922 8628
rect 33229 8619 33287 8625
rect 33229 8616 33241 8619
rect 32916 8588 33241 8616
rect 32916 8576 32922 8588
rect 33229 8585 33241 8588
rect 33275 8585 33287 8619
rect 33229 8579 33287 8585
rect 35158 8576 35164 8628
rect 35216 8616 35222 8628
rect 35437 8619 35495 8625
rect 35437 8616 35449 8619
rect 35216 8588 35449 8616
rect 35216 8576 35222 8588
rect 35437 8585 35449 8588
rect 35483 8585 35495 8619
rect 35437 8579 35495 8585
rect 37274 8576 37280 8628
rect 37332 8616 37338 8628
rect 37461 8619 37519 8625
rect 37461 8616 37473 8619
rect 37332 8588 37473 8616
rect 37332 8576 37338 8588
rect 37461 8585 37473 8588
rect 37507 8585 37519 8619
rect 37461 8579 37519 8585
rect 39390 8576 39396 8628
rect 39448 8616 39454 8628
rect 40037 8619 40095 8625
rect 40037 8616 40049 8619
rect 39448 8588 40049 8616
rect 39448 8576 39454 8588
rect 40037 8585 40049 8588
rect 40083 8585 40095 8619
rect 40037 8579 40095 8585
rect 41414 8576 41420 8628
rect 41472 8576 41478 8628
rect 41506 8576 41512 8628
rect 41564 8616 41570 8628
rect 41785 8619 41843 8625
rect 41785 8616 41797 8619
rect 41564 8588 41797 8616
rect 41564 8576 41570 8588
rect 41785 8585 41797 8588
rect 41831 8585 41843 8619
rect 41785 8579 41843 8585
rect 42150 8576 42156 8628
rect 42208 8576 42214 8628
rect 42702 8576 42708 8628
rect 42760 8576 42766 8628
rect 8036 8520 12204 8548
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8449 1639 8483
rect 1581 8443 1639 8449
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8480 4123 8483
rect 5810 8480 5816 8492
rect 4111 8452 5816 8480
rect 4111 8449 4123 8452
rect 4065 8443 4123 8449
rect 1596 8412 1624 8443
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 6822 8480 6828 8492
rect 5951 8452 6828 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 6822 8440 6828 8452
rect 6880 8440 6886 8492
rect 8036 8489 8064 8520
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8449 8079 8483
rect 8021 8443 8079 8449
rect 10137 8483 10195 8489
rect 10137 8449 10149 8483
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 5442 8412 5448 8424
rect 1596 8384 5448 8412
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 10152 8344 10180 8443
rect 12176 8412 12204 8520
rect 12268 8489 12296 8576
rect 14384 8520 22094 8548
rect 14384 8489 14412 8520
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8449 12311 8483
rect 12253 8443 12311 8449
rect 14369 8483 14427 8489
rect 14369 8449 14381 8483
rect 14415 8449 14427 8483
rect 14369 8443 14427 8449
rect 16482 8440 16488 8492
rect 16540 8440 16546 8492
rect 18598 8440 18604 8492
rect 18656 8440 18662 8492
rect 20714 8440 20720 8492
rect 20772 8440 20778 8492
rect 17126 8412 17132 8424
rect 12176 8384 17132 8412
rect 17126 8372 17132 8384
rect 17184 8372 17190 8424
rect 22066 8412 22094 8520
rect 23750 8508 23756 8560
rect 23808 8548 23814 8560
rect 23808 8520 27384 8548
rect 23808 8508 23814 8520
rect 22830 8440 22836 8492
rect 22888 8440 22894 8492
rect 24949 8483 25007 8489
rect 24949 8449 24961 8483
rect 24995 8480 25007 8483
rect 27154 8480 27160 8492
rect 24995 8452 27160 8480
rect 24995 8449 25007 8452
rect 24949 8443 25007 8449
rect 27154 8440 27160 8452
rect 27212 8440 27218 8492
rect 27249 8483 27307 8489
rect 27249 8449 27261 8483
rect 27295 8449 27307 8483
rect 27356 8480 27384 8520
rect 29104 8520 29316 8548
rect 29104 8480 29132 8520
rect 27356 8452 29132 8480
rect 27249 8443 27307 8449
rect 26786 8412 26792 8424
rect 22066 8384 26792 8412
rect 26786 8372 26792 8384
rect 26844 8372 26850 8424
rect 27264 8412 27292 8443
rect 29178 8440 29184 8492
rect 29236 8440 29242 8492
rect 29288 8480 29316 8520
rect 29362 8508 29368 8560
rect 29420 8548 29426 8560
rect 29420 8520 42564 8548
rect 29420 8508 29426 8520
rect 31297 8483 31355 8489
rect 29288 8452 30420 8480
rect 29086 8412 29092 8424
rect 27264 8384 29092 8412
rect 29086 8372 29092 8384
rect 29144 8372 29150 8424
rect 30392 8412 30420 8452
rect 31297 8449 31309 8483
rect 31343 8480 31355 8483
rect 33318 8480 33324 8492
rect 31343 8452 33324 8480
rect 31343 8449 31355 8452
rect 31297 8443 31355 8449
rect 33318 8440 33324 8452
rect 33376 8440 33382 8492
rect 33413 8483 33471 8489
rect 33413 8449 33425 8483
rect 33459 8480 33471 8483
rect 34974 8480 34980 8492
rect 33459 8452 34980 8480
rect 33459 8449 33471 8452
rect 33413 8443 33471 8449
rect 34974 8440 34980 8452
rect 35032 8440 35038 8492
rect 35066 8440 35072 8492
rect 35124 8480 35130 8492
rect 35253 8483 35311 8489
rect 35253 8480 35265 8483
rect 35124 8452 35265 8480
rect 35124 8440 35130 8452
rect 35253 8449 35265 8452
rect 35299 8449 35311 8483
rect 35253 8443 35311 8449
rect 37642 8440 37648 8492
rect 37700 8440 37706 8492
rect 39850 8440 39856 8492
rect 39908 8440 39914 8492
rect 41230 8440 41236 8492
rect 41288 8440 41294 8492
rect 41598 8440 41604 8492
rect 41656 8440 41662 8492
rect 42536 8489 42564 8520
rect 41969 8483 42027 8489
rect 41969 8480 41981 8483
rect 41892 8452 41981 8480
rect 40034 8412 40040 8424
rect 30392 8384 40040 8412
rect 40034 8372 40040 8384
rect 40092 8372 40098 8424
rect 20438 8344 20444 8356
rect 10152 8316 20444 8344
rect 20438 8304 20444 8316
rect 20496 8304 20502 8356
rect 23382 8304 23388 8356
rect 23440 8344 23446 8356
rect 41892 8344 41920 8452
rect 41969 8449 41981 8452
rect 42015 8449 42027 8483
rect 41969 8443 42027 8449
rect 42521 8483 42579 8489
rect 42521 8449 42533 8483
rect 42567 8449 42579 8483
rect 42521 8443 42579 8449
rect 42889 8483 42947 8489
rect 42889 8449 42901 8483
rect 42935 8449 42947 8483
rect 42889 8443 42947 8449
rect 43257 8483 43315 8489
rect 43257 8449 43269 8483
rect 43303 8480 43315 8483
rect 43916 8480 43944 8928
rect 43303 8452 43944 8480
rect 43303 8449 43315 8452
rect 43257 8443 43315 8449
rect 23440 8316 29132 8344
rect 23440 8304 23446 8316
rect 21358 8236 21364 8288
rect 21416 8276 21422 8288
rect 23198 8276 23204 8288
rect 21416 8248 23204 8276
rect 21416 8236 21422 8248
rect 23198 8236 23204 8248
rect 23256 8236 23262 8288
rect 26142 8236 26148 8288
rect 26200 8276 26206 8288
rect 28166 8276 28172 8288
rect 26200 8248 28172 8276
rect 26200 8236 26206 8248
rect 28166 8236 28172 8248
rect 28224 8236 28230 8288
rect 29104 8276 29132 8316
rect 34486 8316 41920 8344
rect 34486 8276 34514 8316
rect 29104 8248 34514 8276
rect 40034 8236 40040 8288
rect 40092 8276 40098 8288
rect 42904 8276 42932 8443
rect 43070 8304 43076 8356
rect 43128 8304 43134 8356
rect 43438 8304 43444 8356
rect 43496 8304 43502 8356
rect 40092 8248 42932 8276
rect 40092 8236 40098 8248
rect 1104 8186 43884 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 37950 8186
rect 38002 8134 38014 8186
rect 38066 8134 38078 8186
rect 38130 8134 38142 8186
rect 38194 8134 38206 8186
rect 38258 8134 43884 8186
rect 1104 8112 43884 8134
rect 14918 8032 14924 8084
rect 14976 8072 14982 8084
rect 17497 8075 17555 8081
rect 17497 8072 17509 8075
rect 14976 8044 17509 8072
rect 14976 8032 14982 8044
rect 17497 8041 17509 8044
rect 17543 8041 17555 8075
rect 17497 8035 17555 8041
rect 17865 8075 17923 8081
rect 17865 8041 17877 8075
rect 17911 8072 17923 8075
rect 21266 8072 21272 8084
rect 17911 8044 21272 8072
rect 17911 8041 17923 8044
rect 17865 8035 17923 8041
rect 21266 8032 21272 8044
rect 21324 8032 21330 8084
rect 21358 8032 21364 8084
rect 21416 8032 21422 8084
rect 23382 8072 23388 8084
rect 21652 8044 23388 8072
rect 20533 8007 20591 8013
rect 20533 7973 20545 8007
rect 20579 7973 20591 8007
rect 20533 7967 20591 7973
rect 20548 7936 20576 7967
rect 20714 7964 20720 8016
rect 20772 7964 20778 8016
rect 21085 8007 21143 8013
rect 21085 7973 21097 8007
rect 21131 8004 21143 8007
rect 21652 8004 21680 8044
rect 23382 8032 23388 8044
rect 23440 8032 23446 8084
rect 23750 8032 23756 8084
rect 23808 8032 23814 8084
rect 24581 8075 24639 8081
rect 24581 8041 24593 8075
rect 24627 8072 24639 8075
rect 24854 8072 24860 8084
rect 24627 8044 24860 8072
rect 24627 8041 24639 8044
rect 24581 8035 24639 8041
rect 24854 8032 24860 8044
rect 24912 8032 24918 8084
rect 26326 8032 26332 8084
rect 26384 8032 26390 8084
rect 26697 8075 26755 8081
rect 26697 8041 26709 8075
rect 26743 8072 26755 8075
rect 29362 8072 29368 8084
rect 26743 8044 29368 8072
rect 26743 8041 26755 8044
rect 26697 8035 26755 8041
rect 29362 8032 29368 8044
rect 29420 8032 29426 8084
rect 41966 8032 41972 8084
rect 42024 8032 42030 8084
rect 42334 8032 42340 8084
rect 42392 8032 42398 8084
rect 42610 8032 42616 8084
rect 42668 8072 42674 8084
rect 42705 8075 42763 8081
rect 42705 8072 42717 8075
rect 42668 8044 42717 8072
rect 42668 8032 42674 8044
rect 42705 8041 42717 8044
rect 42751 8041 42763 8075
rect 42705 8035 42763 8041
rect 23106 8004 23112 8016
rect 21131 7976 21680 8004
rect 21744 7976 23112 8004
rect 21131 7973 21143 7976
rect 21085 7967 21143 7973
rect 21744 7936 21772 7976
rect 23106 7964 23112 7976
rect 23164 7964 23170 8016
rect 23198 7964 23204 8016
rect 23256 8004 23262 8016
rect 23256 7976 42564 8004
rect 23256 7964 23262 7976
rect 36538 7936 36544 7948
rect 20548 7908 21772 7936
rect 22066 7908 36544 7936
rect 3789 7871 3847 7877
rect 3789 7837 3801 7871
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7868 4215 7871
rect 7834 7868 7840 7880
rect 4203 7840 7840 7868
rect 4203 7837 4215 7840
rect 4157 7831 4215 7837
rect 3804 7800 3832 7831
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 10870 7828 10876 7880
rect 10928 7868 10934 7880
rect 16025 7871 16083 7877
rect 16025 7868 16037 7871
rect 10928 7840 16037 7868
rect 10928 7828 10934 7840
rect 16025 7837 16037 7840
rect 16071 7837 16083 7871
rect 16025 7831 16083 7837
rect 17589 7871 17647 7877
rect 17589 7837 17601 7871
rect 17635 7868 17647 7871
rect 17681 7871 17739 7877
rect 17681 7868 17693 7871
rect 17635 7840 17693 7868
rect 17635 7837 17647 7840
rect 17589 7831 17647 7837
rect 17681 7837 17693 7840
rect 17727 7837 17739 7871
rect 17681 7831 17739 7837
rect 19334 7828 19340 7880
rect 19392 7868 19398 7880
rect 19613 7871 19671 7877
rect 19613 7868 19625 7871
rect 19392 7840 19625 7868
rect 19392 7828 19398 7840
rect 19613 7837 19625 7840
rect 19659 7837 19671 7871
rect 19613 7831 19671 7837
rect 20346 7828 20352 7880
rect 20404 7828 20410 7880
rect 20809 7871 20867 7877
rect 20809 7837 20821 7871
rect 20855 7868 20867 7871
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 20855 7840 20913 7868
rect 20855 7837 20867 7840
rect 20809 7831 20867 7837
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 20990 7828 20996 7880
rect 21048 7868 21054 7880
rect 21177 7871 21235 7877
rect 21177 7868 21189 7871
rect 21048 7840 21189 7868
rect 21048 7828 21054 7840
rect 21177 7837 21189 7840
rect 21223 7837 21235 7871
rect 21177 7831 21235 7837
rect 21266 7828 21272 7880
rect 21324 7868 21330 7880
rect 22066 7868 22094 7908
rect 36538 7896 36544 7908
rect 36596 7896 36602 7948
rect 21324 7840 22094 7868
rect 23477 7871 23535 7877
rect 21324 7828 21330 7840
rect 23477 7837 23489 7871
rect 23523 7868 23535 7871
rect 23569 7871 23627 7877
rect 23569 7868 23581 7871
rect 23523 7840 23581 7868
rect 23523 7837 23535 7840
rect 23477 7831 23535 7837
rect 23569 7837 23581 7840
rect 23615 7837 23627 7871
rect 23569 7831 23627 7837
rect 23658 7828 23664 7880
rect 23716 7868 23722 7880
rect 24397 7871 24455 7877
rect 24397 7868 24409 7871
rect 23716 7840 24409 7868
rect 23716 7828 23722 7840
rect 24397 7837 24409 7840
rect 24443 7868 24455 7871
rect 24673 7871 24731 7877
rect 24673 7868 24685 7871
rect 24443 7840 24685 7868
rect 24443 7837 24455 7840
rect 24397 7831 24455 7837
rect 24673 7837 24685 7840
rect 24719 7837 24731 7871
rect 24673 7831 24731 7837
rect 26421 7871 26479 7877
rect 26421 7837 26433 7871
rect 26467 7868 26479 7871
rect 26513 7871 26571 7877
rect 26513 7868 26525 7871
rect 26467 7840 26525 7868
rect 26467 7837 26479 7840
rect 26421 7831 26479 7837
rect 26513 7837 26525 7840
rect 26559 7837 26571 7871
rect 26513 7831 26571 7837
rect 26973 7871 27031 7877
rect 26973 7837 26985 7871
rect 27019 7868 27031 7871
rect 27065 7871 27123 7877
rect 27065 7868 27077 7871
rect 27019 7840 27077 7868
rect 27019 7837 27031 7840
rect 26973 7831 27031 7837
rect 27065 7837 27077 7840
rect 27111 7837 27123 7871
rect 27065 7831 27123 7837
rect 27522 7828 27528 7880
rect 27580 7828 27586 7880
rect 28350 7828 28356 7880
rect 28408 7828 28414 7880
rect 29546 7828 29552 7880
rect 29604 7868 29610 7880
rect 29825 7871 29883 7877
rect 29825 7868 29837 7871
rect 29604 7840 29837 7868
rect 29604 7828 29610 7840
rect 29825 7837 29837 7840
rect 29871 7837 29883 7871
rect 29825 7831 29883 7837
rect 41782 7828 41788 7880
rect 41840 7828 41846 7880
rect 42536 7877 42564 7976
rect 42153 7871 42211 7877
rect 42153 7837 42165 7871
rect 42199 7837 42211 7871
rect 42153 7831 42211 7837
rect 42521 7871 42579 7877
rect 42521 7837 42533 7871
rect 42567 7837 42579 7871
rect 42521 7831 42579 7837
rect 7558 7800 7564 7812
rect 3804 7772 7564 7800
rect 7558 7760 7564 7772
rect 7616 7760 7622 7812
rect 42168 7800 42196 7831
rect 42610 7828 42616 7880
rect 42668 7868 42674 7880
rect 42889 7871 42947 7877
rect 42889 7868 42901 7871
rect 42668 7840 42901 7868
rect 42668 7828 42674 7840
rect 42889 7837 42901 7840
rect 42935 7837 42947 7871
rect 42889 7831 42947 7837
rect 43254 7828 43260 7880
rect 43312 7828 43318 7880
rect 19536 7772 42196 7800
rect 3970 7692 3976 7744
rect 4028 7692 4034 7744
rect 4338 7692 4344 7744
rect 4396 7692 4402 7744
rect 8846 7692 8852 7744
rect 8904 7732 8910 7744
rect 9398 7732 9404 7744
rect 8904 7704 9404 7732
rect 8904 7692 8910 7704
rect 9398 7692 9404 7704
rect 9456 7692 9462 7744
rect 16209 7735 16267 7741
rect 16209 7701 16221 7735
rect 16255 7732 16267 7735
rect 19058 7732 19064 7744
rect 16255 7704 19064 7732
rect 16255 7701 16267 7704
rect 16209 7695 16267 7701
rect 19058 7692 19064 7704
rect 19116 7692 19122 7744
rect 19536 7741 19564 7772
rect 19521 7735 19579 7741
rect 19521 7701 19533 7735
rect 19567 7701 19579 7735
rect 19521 7695 19579 7701
rect 20990 7692 20996 7744
rect 21048 7732 21054 7744
rect 21453 7735 21511 7741
rect 21453 7732 21465 7735
rect 21048 7704 21465 7732
rect 21048 7692 21054 7704
rect 21453 7701 21465 7704
rect 21499 7701 21511 7735
rect 21453 7695 21511 7701
rect 23474 7692 23480 7744
rect 23532 7692 23538 7744
rect 26878 7692 26884 7744
rect 26936 7692 26942 7744
rect 27246 7692 27252 7744
rect 27304 7692 27310 7744
rect 27341 7735 27399 7741
rect 27341 7701 27353 7735
rect 27387 7732 27399 7735
rect 27430 7732 27436 7744
rect 27387 7704 27436 7732
rect 27387 7701 27399 7704
rect 27341 7695 27399 7701
rect 27430 7692 27436 7704
rect 27488 7692 27494 7744
rect 28166 7692 28172 7744
rect 28224 7692 28230 7744
rect 29730 7692 29736 7744
rect 29788 7692 29794 7744
rect 43070 7692 43076 7744
rect 43128 7692 43134 7744
rect 43438 7692 43444 7744
rect 43496 7692 43502 7744
rect 1104 7642 43884 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 39010 7642
rect 39062 7590 39074 7642
rect 39126 7590 39138 7642
rect 39190 7590 39202 7642
rect 39254 7590 39266 7642
rect 39318 7590 43884 7642
rect 1104 7568 43884 7590
rect 4338 7488 4344 7540
rect 4396 7528 4402 7540
rect 20714 7528 20720 7540
rect 4396 7500 20720 7528
rect 4396 7488 4402 7500
rect 20714 7488 20720 7500
rect 20772 7488 20778 7540
rect 20806 7488 20812 7540
rect 20864 7528 20870 7540
rect 27522 7528 27528 7540
rect 20864 7500 27528 7528
rect 20864 7488 20870 7500
rect 27522 7488 27528 7500
rect 27580 7488 27586 7540
rect 29730 7488 29736 7540
rect 29788 7528 29794 7540
rect 41782 7528 41788 7540
rect 29788 7500 41788 7528
rect 29788 7488 29794 7500
rect 41782 7488 41788 7500
rect 41840 7488 41846 7540
rect 43073 7531 43131 7537
rect 43073 7497 43085 7531
rect 43119 7528 43131 7531
rect 43162 7528 43168 7540
rect 43119 7500 43168 7528
rect 43119 7497 43131 7500
rect 43073 7491 43131 7497
rect 43162 7488 43168 7500
rect 43220 7488 43226 7540
rect 18046 7420 18052 7472
rect 18104 7460 18110 7472
rect 18104 7432 26924 7460
rect 18104 7420 18110 7432
rect 18877 7395 18935 7401
rect 18877 7361 18889 7395
rect 18923 7392 18935 7395
rect 18969 7395 19027 7401
rect 18969 7392 18981 7395
rect 18923 7364 18981 7392
rect 18923 7361 18935 7364
rect 18877 7355 18935 7361
rect 18969 7361 18981 7364
rect 19015 7361 19027 7395
rect 20346 7392 20352 7404
rect 18969 7355 19027 7361
rect 19076 7364 20352 7392
rect 18782 7284 18788 7336
rect 18840 7284 18846 7336
rect 11146 7216 11152 7268
rect 11204 7256 11210 7268
rect 19076 7256 19104 7364
rect 20346 7352 20352 7364
rect 20404 7352 20410 7404
rect 22002 7352 22008 7404
rect 22060 7352 22066 7404
rect 23106 7352 23112 7404
rect 23164 7392 23170 7404
rect 25130 7392 25136 7404
rect 23164 7364 25136 7392
rect 23164 7352 23170 7364
rect 25130 7352 25136 7364
rect 25188 7352 25194 7404
rect 20622 7324 20628 7336
rect 19168 7296 20628 7324
rect 19168 7265 19196 7296
rect 20622 7284 20628 7296
rect 20680 7284 20686 7336
rect 11204 7228 19104 7256
rect 19153 7259 19211 7265
rect 11204 7216 11210 7228
rect 19153 7225 19165 7259
rect 19199 7225 19211 7259
rect 26896 7256 26924 7432
rect 27338 7420 27344 7472
rect 27396 7460 27402 7472
rect 29454 7460 29460 7472
rect 27396 7432 29460 7460
rect 27396 7420 27402 7432
rect 29454 7420 29460 7432
rect 29512 7420 29518 7472
rect 36814 7460 36820 7472
rect 31726 7432 36820 7460
rect 31205 7395 31263 7401
rect 31205 7361 31217 7395
rect 31251 7392 31263 7395
rect 31726 7392 31754 7432
rect 36814 7420 36820 7432
rect 36872 7420 36878 7472
rect 31251 7364 31754 7392
rect 31251 7361 31263 7364
rect 31205 7355 31263 7361
rect 36538 7352 36544 7404
rect 36596 7392 36602 7404
rect 42889 7395 42947 7401
rect 42889 7392 42901 7395
rect 36596 7364 42901 7392
rect 36596 7352 36602 7364
rect 42889 7361 42901 7364
rect 42935 7361 42947 7395
rect 42889 7355 42947 7361
rect 43257 7395 43315 7401
rect 43257 7361 43269 7395
rect 43303 7361 43315 7395
rect 43257 7355 43315 7361
rect 28350 7284 28356 7336
rect 28408 7324 28414 7336
rect 36446 7324 36452 7336
rect 28408 7296 36452 7324
rect 28408 7284 28414 7296
rect 36446 7284 36452 7296
rect 36504 7284 36510 7336
rect 43272 7256 43300 7355
rect 26896 7228 43300 7256
rect 19153 7219 19211 7225
rect 13722 7148 13728 7200
rect 13780 7188 13786 7200
rect 21818 7188 21824 7200
rect 13780 7160 21824 7188
rect 13780 7148 13786 7160
rect 21818 7148 21824 7160
rect 21876 7148 21882 7200
rect 22186 7148 22192 7200
rect 22244 7148 22250 7200
rect 31018 7148 31024 7200
rect 31076 7148 31082 7200
rect 43438 7148 43444 7200
rect 43496 7148 43502 7200
rect 1104 7098 43884 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 37950 7098
rect 38002 7046 38014 7098
rect 38066 7046 38078 7098
rect 38130 7046 38142 7098
rect 38194 7046 38206 7098
rect 38258 7046 43884 7098
rect 1104 7024 43884 7046
rect 3970 6944 3976 6996
rect 4028 6984 4034 6996
rect 13722 6984 13728 6996
rect 4028 6956 13728 6984
rect 4028 6944 4034 6956
rect 13722 6944 13728 6956
rect 13780 6944 13786 6996
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 20806 6984 20812 6996
rect 13872 6956 20812 6984
rect 13872 6944 13878 6956
rect 20806 6944 20812 6956
rect 20864 6944 20870 6996
rect 22186 6944 22192 6996
rect 22244 6984 22250 6996
rect 35618 6984 35624 6996
rect 22244 6956 35624 6984
rect 22244 6944 22250 6956
rect 35618 6944 35624 6956
rect 35676 6944 35682 6996
rect 9582 6876 9588 6928
rect 9640 6876 9646 6928
rect 20622 6876 20628 6928
rect 20680 6916 20686 6928
rect 25222 6916 25228 6928
rect 20680 6888 25228 6916
rect 20680 6876 20686 6888
rect 25222 6876 25228 6888
rect 25280 6876 25286 6928
rect 25317 6919 25375 6925
rect 25317 6885 25329 6919
rect 25363 6885 25375 6919
rect 25317 6879 25375 6885
rect 12526 6808 12532 6860
rect 12584 6848 12590 6860
rect 12584 6820 16160 6848
rect 12584 6808 12590 6820
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6780 2007 6783
rect 6178 6780 6184 6792
rect 1995 6752 6184 6780
rect 1995 6749 2007 6752
rect 1949 6743 2007 6749
rect 6178 6740 6184 6752
rect 6236 6740 6242 6792
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6780 9459 6783
rect 10042 6780 10048 6792
rect 9447 6752 10048 6780
rect 9447 6749 9459 6752
rect 9401 6743 9459 6749
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 10594 6740 10600 6792
rect 10652 6780 10658 6792
rect 16132 6789 16160 6820
rect 16482 6808 16488 6860
rect 16540 6848 16546 6860
rect 25332 6848 25360 6879
rect 25406 6876 25412 6928
rect 25464 6916 25470 6928
rect 43254 6916 43260 6928
rect 25464 6888 43260 6916
rect 25464 6876 25470 6888
rect 43254 6876 43260 6888
rect 43312 6876 43318 6928
rect 16540 6820 25268 6848
rect 25332 6820 41414 6848
rect 16540 6808 16546 6820
rect 12897 6783 12955 6789
rect 12897 6780 12909 6783
rect 10652 6752 12909 6780
rect 10652 6740 10658 6752
rect 12897 6749 12909 6752
rect 12943 6749 12955 6783
rect 12897 6743 12955 6749
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 16117 6783 16175 6789
rect 16117 6749 16129 6783
rect 16163 6749 16175 6783
rect 16117 6743 16175 6749
rect 10226 6712 10232 6724
rect 2148 6684 10232 6712
rect 2148 6653 2176 6684
rect 10226 6672 10232 6684
rect 10284 6672 10290 6724
rect 12250 6672 12256 6724
rect 12308 6712 12314 6724
rect 15856 6712 15884 6743
rect 18690 6740 18696 6792
rect 18748 6780 18754 6792
rect 22833 6783 22891 6789
rect 22833 6780 22845 6783
rect 18748 6752 22845 6780
rect 18748 6740 18754 6752
rect 22833 6749 22845 6752
rect 22879 6749 22891 6783
rect 22833 6743 22891 6749
rect 25041 6783 25099 6789
rect 25041 6749 25053 6783
rect 25087 6780 25099 6783
rect 25133 6783 25191 6789
rect 25133 6780 25145 6783
rect 25087 6752 25145 6780
rect 25087 6749 25099 6752
rect 25041 6743 25099 6749
rect 25133 6749 25145 6752
rect 25179 6749 25191 6783
rect 25240 6780 25268 6820
rect 26973 6783 27031 6789
rect 26973 6780 26985 6783
rect 25240 6752 26985 6780
rect 25133 6743 25191 6749
rect 26973 6749 26985 6752
rect 27019 6780 27031 6783
rect 27157 6783 27215 6789
rect 27157 6780 27169 6783
rect 27019 6752 27169 6780
rect 27019 6749 27031 6752
rect 26973 6743 27031 6749
rect 27157 6749 27169 6752
rect 27203 6749 27215 6783
rect 27157 6743 27215 6749
rect 29917 6783 29975 6789
rect 29917 6749 29929 6783
rect 29963 6780 29975 6783
rect 30009 6783 30067 6789
rect 30009 6780 30021 6783
rect 29963 6752 30021 6780
rect 29963 6749 29975 6752
rect 29917 6743 29975 6749
rect 30009 6749 30021 6752
rect 30055 6749 30067 6783
rect 30009 6743 30067 6749
rect 34885 6783 34943 6789
rect 34885 6749 34897 6783
rect 34931 6780 34943 6783
rect 38470 6780 38476 6792
rect 34931 6752 38476 6780
rect 34931 6749 34943 6752
rect 34885 6743 34943 6749
rect 38470 6740 38476 6752
rect 38528 6740 38534 6792
rect 41386 6780 41414 6820
rect 42889 6783 42947 6789
rect 42889 6780 42901 6783
rect 41386 6752 42901 6780
rect 42889 6749 42901 6752
rect 42935 6749 42947 6783
rect 42889 6743 42947 6749
rect 42978 6740 42984 6792
rect 43036 6780 43042 6792
rect 43257 6783 43315 6789
rect 43257 6780 43269 6783
rect 43036 6752 43269 6780
rect 43036 6740 43042 6752
rect 43257 6749 43269 6752
rect 43303 6749 43315 6783
rect 43257 6743 43315 6749
rect 22002 6712 22008 6724
rect 12308 6684 15884 6712
rect 15948 6684 22008 6712
rect 12308 6672 12314 6684
rect 2133 6647 2191 6653
rect 2133 6613 2145 6647
rect 2179 6613 2191 6647
rect 2133 6607 2191 6613
rect 9582 6604 9588 6656
rect 9640 6644 9646 6656
rect 12894 6644 12900 6656
rect 9640 6616 12900 6644
rect 9640 6604 9646 6616
rect 12894 6604 12900 6616
rect 12952 6604 12958 6656
rect 13081 6647 13139 6653
rect 13081 6613 13093 6647
rect 13127 6644 13139 6647
rect 13170 6644 13176 6656
rect 13127 6616 13176 6644
rect 13127 6613 13139 6616
rect 13081 6607 13139 6613
rect 13170 6604 13176 6616
rect 13228 6604 13234 6656
rect 14918 6604 14924 6656
rect 14976 6644 14982 6656
rect 15948 6644 15976 6684
rect 22002 6672 22008 6684
rect 22060 6672 22066 6724
rect 24946 6672 24952 6724
rect 25004 6672 25010 6724
rect 29362 6712 29368 6724
rect 27264 6684 29368 6712
rect 14976 6616 15976 6644
rect 14976 6604 14982 6616
rect 16022 6604 16028 6656
rect 16080 6604 16086 6656
rect 16298 6604 16304 6656
rect 16356 6604 16362 6656
rect 23017 6647 23075 6653
rect 23017 6613 23029 6647
rect 23063 6644 23075 6647
rect 27264 6644 27292 6684
rect 29362 6672 29368 6684
rect 29420 6672 29426 6724
rect 23063 6616 27292 6644
rect 27341 6647 27399 6653
rect 23063 6613 23075 6616
rect 23017 6607 23075 6613
rect 27341 6613 27353 6647
rect 27387 6644 27399 6647
rect 29546 6644 29552 6656
rect 27387 6616 29552 6644
rect 27387 6613 27399 6616
rect 27341 6607 27399 6613
rect 29546 6604 29552 6616
rect 29604 6604 29610 6656
rect 29822 6604 29828 6656
rect 29880 6604 29886 6656
rect 30193 6647 30251 6653
rect 30193 6613 30205 6647
rect 30239 6644 30251 6647
rect 34422 6644 34428 6656
rect 30239 6616 34428 6644
rect 30239 6613 30251 6616
rect 30193 6607 30251 6613
rect 34422 6604 34428 6616
rect 34480 6604 34486 6656
rect 35066 6604 35072 6656
rect 35124 6604 35130 6656
rect 43070 6604 43076 6656
rect 43128 6604 43134 6656
rect 43438 6604 43444 6656
rect 43496 6604 43502 6656
rect 1104 6554 43884 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 39010 6554
rect 39062 6502 39074 6554
rect 39126 6502 39138 6554
rect 39190 6502 39202 6554
rect 39254 6502 39266 6554
rect 39318 6502 43884 6554
rect 1104 6480 43884 6502
rect 5810 6400 5816 6452
rect 5868 6440 5874 6452
rect 9217 6443 9275 6449
rect 9217 6440 9229 6443
rect 5868 6412 9229 6440
rect 5868 6400 5874 6412
rect 9217 6409 9229 6412
rect 9263 6409 9275 6443
rect 9217 6403 9275 6409
rect 12342 6400 12348 6452
rect 12400 6440 12406 6452
rect 17681 6443 17739 6449
rect 17681 6440 17693 6443
rect 12400 6412 17693 6440
rect 12400 6400 12406 6412
rect 17681 6409 17693 6412
rect 17727 6409 17739 6443
rect 17681 6403 17739 6409
rect 18046 6400 18052 6452
rect 18104 6400 18110 6452
rect 20898 6400 20904 6452
rect 20956 6440 20962 6452
rect 21177 6443 21235 6449
rect 21177 6440 21189 6443
rect 20956 6412 21189 6440
rect 20956 6400 20962 6412
rect 21177 6409 21189 6412
rect 21223 6409 21235 6443
rect 21177 6403 21235 6409
rect 25498 6400 25504 6452
rect 25556 6400 25562 6452
rect 27522 6440 27528 6452
rect 25608 6412 27528 6440
rect 10226 6332 10232 6384
rect 10284 6372 10290 6384
rect 12986 6372 12992 6384
rect 10284 6344 12992 6372
rect 10284 6332 10290 6344
rect 12986 6332 12992 6344
rect 13044 6332 13050 6384
rect 15194 6332 15200 6384
rect 15252 6372 15258 6384
rect 24670 6372 24676 6384
rect 15252 6344 24676 6372
rect 15252 6332 15258 6344
rect 24670 6332 24676 6344
rect 24728 6332 24734 6384
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6304 5963 6307
rect 7282 6304 7288 6316
rect 5951 6276 7288 6304
rect 5951 6273 5963 6276
rect 5905 6267 5963 6273
rect 7282 6264 7288 6276
rect 7340 6264 7346 6316
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6304 9183 6307
rect 9398 6304 9404 6316
rect 9171 6276 9404 6304
rect 9171 6273 9183 6276
rect 9125 6267 9183 6273
rect 9398 6264 9404 6276
rect 9456 6264 9462 6316
rect 10873 6307 10931 6313
rect 10873 6273 10885 6307
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 10888 6236 10916 6267
rect 13630 6264 13636 6316
rect 13688 6304 13694 6316
rect 13725 6307 13783 6313
rect 13725 6304 13737 6307
rect 13688 6276 13737 6304
rect 13688 6264 13694 6276
rect 13725 6273 13737 6276
rect 13771 6273 13783 6307
rect 13725 6267 13783 6273
rect 17773 6307 17831 6313
rect 17773 6273 17785 6307
rect 17819 6304 17831 6307
rect 17865 6307 17923 6313
rect 17865 6304 17877 6307
rect 17819 6276 17877 6304
rect 17819 6273 17831 6276
rect 17773 6267 17831 6273
rect 17865 6273 17877 6276
rect 17911 6273 17923 6307
rect 17865 6267 17923 6273
rect 20349 6307 20407 6313
rect 20349 6273 20361 6307
rect 20395 6273 20407 6307
rect 20349 6267 20407 6273
rect 21269 6307 21327 6313
rect 21269 6273 21281 6307
rect 21315 6304 21327 6307
rect 21361 6307 21419 6313
rect 21361 6304 21373 6307
rect 21315 6276 21373 6304
rect 21315 6273 21327 6276
rect 21269 6267 21327 6273
rect 21361 6273 21373 6276
rect 21407 6273 21419 6307
rect 21361 6267 21419 6273
rect 14734 6236 14740 6248
rect 10888 6208 14740 6236
rect 14734 6196 14740 6208
rect 14792 6196 14798 6248
rect 17678 6196 17684 6248
rect 17736 6236 17742 6248
rect 20364 6236 20392 6267
rect 21450 6264 21456 6316
rect 21508 6304 21514 6316
rect 25608 6304 25636 6412
rect 27522 6400 27528 6412
rect 27580 6400 27586 6452
rect 29178 6400 29184 6452
rect 29236 6440 29242 6452
rect 31757 6443 31815 6449
rect 31757 6440 31769 6443
rect 29236 6412 31769 6440
rect 29236 6400 29242 6412
rect 31757 6409 31769 6412
rect 31803 6409 31815 6443
rect 36262 6440 36268 6452
rect 31757 6403 31815 6409
rect 33980 6412 36268 6440
rect 33980 6372 34008 6412
rect 36262 6400 36268 6412
rect 36320 6400 36326 6452
rect 37642 6400 37648 6452
rect 37700 6440 37706 6452
rect 37737 6443 37795 6449
rect 37737 6440 37749 6443
rect 37700 6412 37749 6440
rect 37700 6400 37706 6412
rect 37737 6409 37749 6412
rect 37783 6409 37795 6443
rect 37737 6403 37795 6409
rect 38473 6443 38531 6449
rect 38473 6409 38485 6443
rect 38519 6440 38531 6443
rect 39850 6440 39856 6452
rect 38519 6412 39856 6440
rect 38519 6409 38531 6412
rect 38473 6403 38531 6409
rect 39850 6400 39856 6412
rect 39908 6400 39914 6452
rect 41230 6400 41236 6452
rect 41288 6440 41294 6452
rect 41325 6443 41383 6449
rect 41325 6440 41337 6443
rect 41288 6412 41337 6440
rect 41288 6400 41294 6412
rect 41325 6409 41337 6412
rect 41371 6409 41383 6443
rect 41325 6403 41383 6409
rect 43438 6400 43444 6452
rect 43496 6400 43502 6452
rect 25700 6344 34008 6372
rect 25700 6313 25728 6344
rect 35618 6332 35624 6384
rect 35676 6372 35682 6384
rect 43162 6372 43168 6384
rect 35676 6344 43168 6372
rect 35676 6332 35682 6344
rect 43162 6332 43168 6344
rect 43220 6332 43226 6384
rect 21508 6276 25636 6304
rect 25685 6307 25743 6313
rect 21508 6264 21514 6276
rect 25685 6273 25697 6307
rect 25731 6273 25743 6307
rect 25685 6267 25743 6273
rect 31389 6307 31447 6313
rect 31389 6273 31401 6307
rect 31435 6304 31447 6307
rect 31941 6307 31999 6313
rect 31435 6276 31754 6304
rect 31435 6273 31447 6276
rect 31389 6267 31447 6273
rect 29822 6236 29828 6248
rect 17736 6208 20392 6236
rect 20456 6208 29828 6236
rect 17736 6196 17742 6208
rect 1302 6128 1308 6180
rect 1360 6168 1366 6180
rect 18782 6168 18788 6180
rect 1360 6140 18788 6168
rect 1360 6128 1366 6140
rect 18782 6128 18788 6140
rect 18840 6128 18846 6180
rect 6089 6103 6147 6109
rect 6089 6069 6101 6103
rect 6135 6100 6147 6103
rect 9582 6100 9588 6112
rect 6135 6072 9588 6100
rect 6135 6069 6147 6072
rect 6089 6063 6147 6069
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 11054 6060 11060 6112
rect 11112 6060 11118 6112
rect 13909 6103 13967 6109
rect 13909 6069 13921 6103
rect 13955 6100 13967 6103
rect 14826 6100 14832 6112
rect 13955 6072 14832 6100
rect 13955 6069 13967 6072
rect 13909 6063 13967 6069
rect 14826 6060 14832 6072
rect 14884 6060 14890 6112
rect 15010 6060 15016 6112
rect 15068 6100 15074 6112
rect 20456 6100 20484 6208
rect 29822 6196 29828 6208
rect 29880 6196 29886 6248
rect 31726 6236 31754 6276
rect 31941 6273 31953 6307
rect 31987 6304 31999 6307
rect 37642 6304 37648 6316
rect 31987 6276 37648 6304
rect 31987 6273 31999 6276
rect 31941 6267 31999 6273
rect 37642 6264 37648 6276
rect 37700 6264 37706 6316
rect 37921 6307 37979 6313
rect 37921 6273 37933 6307
rect 37967 6273 37979 6307
rect 37921 6267 37979 6273
rect 38289 6307 38347 6313
rect 38289 6273 38301 6307
rect 38335 6304 38347 6307
rect 38930 6304 38936 6316
rect 38335 6276 38936 6304
rect 38335 6273 38347 6276
rect 38289 6267 38347 6273
rect 37182 6236 37188 6248
rect 31726 6208 37188 6236
rect 37182 6196 37188 6208
rect 37240 6196 37246 6248
rect 37936 6236 37964 6267
rect 38930 6264 38936 6276
rect 38988 6264 38994 6316
rect 39117 6307 39175 6313
rect 39117 6273 39129 6307
rect 39163 6304 39175 6307
rect 39390 6304 39396 6316
rect 39163 6276 39396 6304
rect 39163 6273 39175 6276
rect 39117 6267 39175 6273
rect 39390 6264 39396 6276
rect 39448 6264 39454 6316
rect 39574 6264 39580 6316
rect 39632 6304 39638 6316
rect 41141 6307 41199 6313
rect 41141 6304 41153 6307
rect 39632 6276 41153 6304
rect 39632 6264 39638 6276
rect 41141 6273 41153 6276
rect 41187 6273 41199 6307
rect 41141 6267 41199 6273
rect 42886 6264 42892 6316
rect 42944 6264 42950 6316
rect 43254 6264 43260 6316
rect 43312 6264 43318 6316
rect 38746 6236 38752 6248
rect 37936 6208 38752 6236
rect 38746 6196 38752 6208
rect 38804 6196 38810 6248
rect 29454 6128 29460 6180
rect 29512 6168 29518 6180
rect 29512 6140 31892 6168
rect 29512 6128 29518 6140
rect 15068 6072 20484 6100
rect 15068 6060 15074 6072
rect 20530 6060 20536 6112
rect 20588 6060 20594 6112
rect 21545 6103 21603 6109
rect 21545 6069 21557 6103
rect 21591 6100 21603 6103
rect 25406 6100 25412 6112
rect 21591 6072 25412 6100
rect 21591 6069 21603 6072
rect 21545 6063 21603 6069
rect 25406 6060 25412 6072
rect 25464 6060 25470 6112
rect 28718 6060 28724 6112
rect 28776 6100 28782 6112
rect 31205 6103 31263 6109
rect 31205 6100 31217 6103
rect 28776 6072 31217 6100
rect 28776 6060 28782 6072
rect 31205 6069 31217 6072
rect 31251 6069 31263 6103
rect 31864 6100 31892 6140
rect 33226 6128 33232 6180
rect 33284 6168 33290 6180
rect 37366 6168 37372 6180
rect 33284 6140 37372 6168
rect 33284 6128 33290 6140
rect 37366 6128 37372 6140
rect 37424 6128 37430 6180
rect 39301 6171 39359 6177
rect 39301 6137 39313 6171
rect 39347 6168 39359 6171
rect 41598 6168 41604 6180
rect 39347 6140 41604 6168
rect 39347 6137 39359 6140
rect 39301 6131 39359 6137
rect 41598 6128 41604 6140
rect 41656 6128 41662 6180
rect 42334 6100 42340 6112
rect 31864 6072 42340 6100
rect 31205 6063 31263 6069
rect 42334 6060 42340 6072
rect 42392 6060 42398 6112
rect 43070 6060 43076 6112
rect 43128 6060 43134 6112
rect 1104 6010 43884 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 37950 6010
rect 38002 5958 38014 6010
rect 38066 5958 38078 6010
rect 38130 5958 38142 6010
rect 38194 5958 38206 6010
rect 38258 5958 43884 6010
rect 1104 5936 43884 5958
rect 11606 5856 11612 5908
rect 11664 5896 11670 5908
rect 14918 5896 14924 5908
rect 11664 5868 14924 5896
rect 11664 5856 11670 5868
rect 14918 5856 14924 5868
rect 14976 5856 14982 5908
rect 15194 5856 15200 5908
rect 15252 5856 15258 5908
rect 15473 5899 15531 5905
rect 15473 5865 15485 5899
rect 15519 5896 15531 5899
rect 21450 5896 21456 5908
rect 15519 5868 21456 5896
rect 15519 5865 15531 5868
rect 15473 5859 15531 5865
rect 21450 5856 21456 5868
rect 21508 5856 21514 5908
rect 21560 5868 22094 5896
rect 934 5788 940 5840
rect 992 5828 998 5840
rect 18693 5831 18751 5837
rect 992 5800 18644 5828
rect 992 5788 998 5800
rect 11974 5720 11980 5772
rect 12032 5760 12038 5772
rect 12032 5732 18552 5760
rect 12032 5720 12038 5732
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5692 6699 5695
rect 7006 5692 7012 5704
rect 6687 5664 7012 5692
rect 6687 5661 6699 5664
rect 6641 5655 6699 5661
rect 7006 5652 7012 5664
rect 7064 5652 7070 5704
rect 9490 5652 9496 5704
rect 9548 5692 9554 5704
rect 15013 5695 15071 5701
rect 15013 5692 15025 5695
rect 9548 5664 15025 5692
rect 9548 5652 9554 5664
rect 15013 5661 15025 5664
rect 15059 5661 15071 5695
rect 15013 5655 15071 5661
rect 15286 5652 15292 5704
rect 15344 5652 15350 5704
rect 18524 5701 18552 5732
rect 18509 5695 18567 5701
rect 18509 5661 18521 5695
rect 18555 5661 18567 5695
rect 18616 5692 18644 5800
rect 18693 5797 18705 5831
rect 18739 5797 18751 5831
rect 18693 5791 18751 5797
rect 18708 5760 18736 5791
rect 18782 5788 18788 5840
rect 18840 5828 18846 5840
rect 21560 5828 21588 5868
rect 18840 5800 21588 5828
rect 18840 5788 18846 5800
rect 21634 5788 21640 5840
rect 21692 5788 21698 5840
rect 22066 5828 22094 5868
rect 25406 5856 25412 5908
rect 25464 5896 25470 5908
rect 42978 5896 42984 5908
rect 25464 5868 42984 5896
rect 25464 5856 25470 5868
rect 42978 5856 42984 5868
rect 43036 5856 43042 5908
rect 26050 5828 26056 5840
rect 22066 5800 26056 5828
rect 26050 5788 26056 5800
rect 26108 5788 26114 5840
rect 26252 5800 33364 5828
rect 18708 5732 21680 5760
rect 21453 5695 21511 5701
rect 21453 5692 21465 5695
rect 18616 5664 21465 5692
rect 18509 5655 18567 5661
rect 21453 5661 21465 5664
rect 21499 5661 21511 5695
rect 21652 5692 21680 5732
rect 25774 5692 25780 5704
rect 21652 5664 25780 5692
rect 21453 5655 21511 5661
rect 25774 5652 25780 5664
rect 25832 5652 25838 5704
rect 26252 5701 26280 5800
rect 33226 5760 33232 5772
rect 30944 5732 33232 5760
rect 26237 5695 26295 5701
rect 26237 5661 26249 5695
rect 26283 5661 26295 5695
rect 26237 5655 26295 5661
rect 28350 5652 28356 5704
rect 28408 5652 28414 5704
rect 29086 5652 29092 5704
rect 29144 5692 29150 5704
rect 30944 5701 30972 5732
rect 33226 5720 33232 5732
rect 33284 5720 33290 5772
rect 33336 5760 33364 5800
rect 33410 5788 33416 5840
rect 33468 5828 33474 5840
rect 33689 5831 33747 5837
rect 33689 5828 33701 5831
rect 33468 5800 33701 5828
rect 33468 5788 33474 5800
rect 33689 5797 33701 5800
rect 33735 5797 33747 5831
rect 35802 5828 35808 5840
rect 33689 5791 33747 5797
rect 33796 5800 35808 5828
rect 33796 5760 33824 5800
rect 35802 5788 35808 5800
rect 35860 5788 35866 5840
rect 43438 5788 43444 5840
rect 43496 5788 43502 5840
rect 33336 5732 33824 5760
rect 33962 5720 33968 5772
rect 34020 5760 34026 5772
rect 34020 5732 43300 5760
rect 34020 5720 34026 5732
rect 30929 5695 30987 5701
rect 29144 5664 30788 5692
rect 29144 5652 29150 5664
rect 7374 5584 7380 5636
rect 7432 5624 7438 5636
rect 23198 5624 23204 5636
rect 7432 5596 23204 5624
rect 7432 5584 7438 5596
rect 23198 5584 23204 5596
rect 23256 5584 23262 5636
rect 6825 5559 6883 5565
rect 6825 5525 6837 5559
rect 6871 5556 6883 5559
rect 8478 5556 8484 5568
rect 6871 5528 8484 5556
rect 6871 5525 6883 5528
rect 6825 5519 6883 5525
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 12802 5516 12808 5568
rect 12860 5556 12866 5568
rect 15286 5556 15292 5568
rect 12860 5528 15292 5556
rect 12860 5516 12866 5528
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 20530 5516 20536 5568
rect 20588 5556 20594 5568
rect 25406 5556 25412 5568
rect 20588 5528 25412 5556
rect 20588 5516 20594 5528
rect 25406 5516 25412 5528
rect 25464 5516 25470 5568
rect 25866 5516 25872 5568
rect 25924 5556 25930 5568
rect 26053 5559 26111 5565
rect 26053 5556 26065 5559
rect 25924 5528 26065 5556
rect 25924 5516 25930 5528
rect 26053 5525 26065 5528
rect 26099 5525 26111 5559
rect 26053 5519 26111 5525
rect 28537 5559 28595 5565
rect 28537 5525 28549 5559
rect 28583 5556 28595 5559
rect 30374 5556 30380 5568
rect 28583 5528 30380 5556
rect 28583 5525 28595 5528
rect 28537 5519 28595 5525
rect 30374 5516 30380 5528
rect 30432 5516 30438 5568
rect 30760 5565 30788 5664
rect 30929 5661 30941 5695
rect 30975 5661 30987 5695
rect 30929 5655 30987 5661
rect 33873 5695 33931 5701
rect 33873 5661 33885 5695
rect 33919 5692 33931 5695
rect 35253 5695 35311 5701
rect 33919 5664 35112 5692
rect 33919 5661 33931 5664
rect 33873 5655 33931 5661
rect 31110 5584 31116 5636
rect 31168 5624 31174 5636
rect 35084 5624 35112 5664
rect 35253 5661 35265 5695
rect 35299 5692 35311 5695
rect 35529 5695 35587 5701
rect 35529 5692 35541 5695
rect 35299 5664 35541 5692
rect 35299 5661 35311 5664
rect 35253 5655 35311 5661
rect 35529 5661 35541 5664
rect 35575 5661 35587 5695
rect 35529 5655 35587 5661
rect 38654 5652 38660 5704
rect 38712 5692 38718 5704
rect 43272 5701 43300 5732
rect 42889 5695 42947 5701
rect 42889 5692 42901 5695
rect 38712 5664 42901 5692
rect 38712 5652 38718 5664
rect 42889 5661 42901 5664
rect 42935 5661 42947 5695
rect 42889 5655 42947 5661
rect 43257 5695 43315 5701
rect 43257 5661 43269 5695
rect 43303 5661 43315 5695
rect 43257 5655 43315 5661
rect 37826 5624 37832 5636
rect 31168 5596 33824 5624
rect 35084 5596 37832 5624
rect 31168 5584 31174 5596
rect 30745 5559 30803 5565
rect 30745 5525 30757 5559
rect 30791 5525 30803 5559
rect 33796 5556 33824 5596
rect 37826 5584 37832 5596
rect 37884 5584 37890 5636
rect 35161 5559 35219 5565
rect 35161 5556 35173 5559
rect 33796 5528 35173 5556
rect 30745 5519 30803 5525
rect 35161 5525 35173 5528
rect 35207 5525 35219 5559
rect 35161 5519 35219 5525
rect 35342 5516 35348 5568
rect 35400 5516 35406 5568
rect 43070 5516 43076 5568
rect 43128 5516 43134 5568
rect 1104 5466 43884 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 39010 5466
rect 39062 5414 39074 5466
rect 39126 5414 39138 5466
rect 39190 5414 39202 5466
rect 39254 5414 39266 5466
rect 39318 5414 43884 5466
rect 1104 5392 43884 5414
rect 8846 5312 8852 5364
rect 8904 5352 8910 5364
rect 22005 5355 22063 5361
rect 8904 5324 17908 5352
rect 8904 5312 8910 5324
rect 17880 5284 17908 5324
rect 22005 5321 22017 5355
rect 22051 5321 22063 5355
rect 22005 5315 22063 5321
rect 22020 5284 22048 5315
rect 23198 5312 23204 5364
rect 23256 5312 23262 5364
rect 25869 5355 25927 5361
rect 25869 5321 25881 5355
rect 25915 5352 25927 5355
rect 25915 5324 31754 5352
rect 25915 5321 25927 5324
rect 25869 5315 25927 5321
rect 29638 5284 29644 5296
rect 9968 5256 12434 5284
rect 17880 5256 18828 5284
rect 22020 5256 29644 5284
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5185 2375 5219
rect 2317 5179 2375 5185
rect 3973 5219 4031 5225
rect 3973 5185 3985 5219
rect 4019 5216 4031 5219
rect 7742 5216 7748 5228
rect 4019 5188 7748 5216
rect 4019 5185 4031 5188
rect 3973 5179 4031 5185
rect 2332 5148 2360 5179
rect 7742 5176 7748 5188
rect 7800 5176 7806 5228
rect 9968 5225 9996 5256
rect 9677 5219 9735 5225
rect 9677 5185 9689 5219
rect 9723 5216 9735 5219
rect 9953 5219 10011 5225
rect 9953 5216 9965 5219
rect 9723 5188 9965 5216
rect 9723 5185 9735 5188
rect 9677 5179 9735 5185
rect 9953 5185 9965 5188
rect 9999 5185 10011 5219
rect 12406 5216 12434 5256
rect 17494 5216 17500 5228
rect 12406 5188 17500 5216
rect 9953 5179 10011 5185
rect 17494 5176 17500 5188
rect 17552 5176 17558 5228
rect 17604 5225 17724 5240
rect 17589 5219 17739 5225
rect 17589 5185 17601 5219
rect 17635 5212 17693 5219
rect 17635 5185 17647 5212
rect 17589 5179 17647 5185
rect 17681 5185 17693 5212
rect 17727 5185 17739 5219
rect 17681 5179 17739 5185
rect 17862 5176 17868 5228
rect 17920 5216 17926 5228
rect 18141 5219 18199 5225
rect 18141 5216 18153 5219
rect 17920 5188 18153 5216
rect 17920 5176 17926 5188
rect 18141 5185 18153 5188
rect 18187 5185 18199 5219
rect 18800 5216 18828 5256
rect 29638 5244 29644 5256
rect 29696 5244 29702 5296
rect 31726 5284 31754 5324
rect 34974 5312 34980 5364
rect 35032 5352 35038 5364
rect 36909 5355 36967 5361
rect 36909 5352 36921 5355
rect 35032 5324 36921 5352
rect 35032 5312 35038 5324
rect 36909 5321 36921 5324
rect 36955 5321 36967 5355
rect 36909 5315 36967 5321
rect 43438 5312 43444 5364
rect 43496 5312 43502 5364
rect 33502 5284 33508 5296
rect 31726 5256 33508 5284
rect 33502 5244 33508 5256
rect 33560 5244 33566 5296
rect 42610 5284 42616 5296
rect 33704 5256 42616 5284
rect 21821 5219 21879 5225
rect 21821 5216 21833 5219
rect 18800 5188 21833 5216
rect 18141 5179 18199 5185
rect 21821 5185 21833 5188
rect 21867 5216 21879 5219
rect 22097 5219 22155 5225
rect 22097 5216 22109 5219
rect 21867 5188 22109 5216
rect 21867 5185 21879 5188
rect 21821 5179 21879 5185
rect 22097 5185 22109 5188
rect 22143 5185 22155 5219
rect 22097 5179 22155 5185
rect 23293 5219 23351 5225
rect 23293 5185 23305 5219
rect 23339 5216 23351 5219
rect 23385 5219 23443 5225
rect 23385 5216 23397 5219
rect 23339 5188 23397 5216
rect 23339 5185 23351 5188
rect 23293 5179 23351 5185
rect 23385 5185 23397 5188
rect 23431 5185 23443 5219
rect 23385 5179 23443 5185
rect 25685 5219 25743 5225
rect 25685 5185 25697 5219
rect 25731 5185 25743 5219
rect 25685 5179 25743 5185
rect 5902 5148 5908 5160
rect 2332 5120 5908 5148
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 7190 5108 7196 5160
rect 7248 5148 7254 5160
rect 25700 5148 25728 5179
rect 26050 5176 26056 5228
rect 26108 5176 26114 5228
rect 27338 5176 27344 5228
rect 27396 5216 27402 5228
rect 27525 5219 27583 5225
rect 27525 5216 27537 5219
rect 27396 5188 27537 5216
rect 27396 5176 27402 5188
rect 27525 5185 27537 5188
rect 27571 5185 27583 5219
rect 27525 5179 27583 5185
rect 31202 5176 31208 5228
rect 31260 5216 31266 5228
rect 33229 5219 33287 5225
rect 33229 5216 33241 5219
rect 31260 5188 33241 5216
rect 31260 5176 31266 5188
rect 33229 5185 33241 5188
rect 33275 5216 33287 5219
rect 33597 5219 33655 5225
rect 33597 5216 33609 5219
rect 33275 5188 33609 5216
rect 33275 5185 33287 5188
rect 33229 5179 33287 5185
rect 33597 5185 33609 5188
rect 33643 5185 33655 5219
rect 33597 5179 33655 5185
rect 33134 5148 33140 5160
rect 7248 5120 17908 5148
rect 7248 5108 7254 5120
rect 6822 5040 6828 5092
rect 6880 5080 6886 5092
rect 9769 5083 9827 5089
rect 9769 5080 9781 5083
rect 6880 5052 9781 5080
rect 6880 5040 6886 5052
rect 9769 5049 9781 5052
rect 9815 5049 9827 5083
rect 17880 5080 17908 5120
rect 18248 5120 25728 5148
rect 31726 5120 33140 5148
rect 18248 5080 18276 5120
rect 17880 5052 18276 5080
rect 26237 5083 26295 5089
rect 9769 5043 9827 5049
rect 26237 5049 26249 5083
rect 26283 5080 26295 5083
rect 27709 5083 27767 5089
rect 26283 5052 27660 5080
rect 26283 5049 26295 5052
rect 26237 5043 26295 5049
rect 2498 4972 2504 5024
rect 2556 4972 2562 5024
rect 4157 5015 4215 5021
rect 4157 4981 4169 5015
rect 4203 5012 4215 5015
rect 7466 5012 7472 5024
rect 4203 4984 7472 5012
rect 4203 4981 4215 4984
rect 4157 4975 4215 4981
rect 7466 4972 7472 4984
rect 7524 4972 7530 5024
rect 8754 4972 8760 5024
rect 8812 5012 8818 5024
rect 17497 5015 17555 5021
rect 17497 5012 17509 5015
rect 8812 4984 17509 5012
rect 8812 4972 8818 4984
rect 17497 4981 17509 4984
rect 17543 4981 17555 5015
rect 17497 4975 17555 4981
rect 17770 4972 17776 5024
rect 17828 5012 17834 5024
rect 17865 5015 17923 5021
rect 17865 5012 17877 5015
rect 17828 4984 17877 5012
rect 17828 4972 17834 4984
rect 17865 4981 17877 4984
rect 17911 4981 17923 5015
rect 17865 4975 17923 4981
rect 18325 5015 18383 5021
rect 18325 4981 18337 5015
rect 18371 5012 18383 5015
rect 20622 5012 20628 5024
rect 18371 4984 20628 5012
rect 18371 4981 18383 4984
rect 18325 4975 18383 4981
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 23569 5015 23627 5021
rect 23569 4981 23581 5015
rect 23615 5012 23627 5015
rect 26418 5012 26424 5024
rect 23615 4984 26424 5012
rect 23615 4981 23627 4984
rect 23569 4975 23627 4981
rect 26418 4972 26424 4984
rect 26476 4972 26482 5024
rect 27632 5012 27660 5052
rect 27709 5049 27721 5083
rect 27755 5080 27767 5083
rect 31726 5080 31754 5120
rect 33134 5108 33140 5120
rect 33192 5108 33198 5160
rect 33704 5148 33732 5256
rect 42610 5244 42616 5256
rect 42668 5244 42674 5296
rect 37093 5219 37151 5225
rect 37093 5185 37105 5219
rect 37139 5185 37151 5219
rect 37093 5179 37151 5185
rect 37461 5219 37519 5225
rect 37461 5185 37473 5219
rect 37507 5216 37519 5219
rect 37553 5219 37611 5225
rect 37553 5216 37565 5219
rect 37507 5188 37565 5216
rect 37507 5185 37519 5188
rect 37461 5179 37519 5185
rect 37553 5185 37565 5188
rect 37599 5185 37611 5219
rect 37553 5179 37611 5185
rect 33244 5120 33732 5148
rect 37108 5148 37136 5179
rect 42794 5176 42800 5228
rect 42852 5216 42858 5228
rect 42889 5219 42947 5225
rect 42889 5216 42901 5219
rect 42852 5188 42901 5216
rect 42852 5176 42858 5188
rect 42889 5185 42901 5188
rect 42935 5185 42947 5219
rect 42889 5179 42947 5185
rect 43254 5176 43260 5228
rect 43312 5176 43318 5228
rect 38286 5148 38292 5160
rect 37108 5120 38292 5148
rect 27755 5052 31754 5080
rect 27755 5049 27767 5052
rect 27709 5043 27767 5049
rect 33244 5012 33272 5120
rect 38286 5108 38292 5120
rect 38344 5108 38350 5160
rect 33318 5040 33324 5092
rect 33376 5080 33382 5092
rect 42886 5080 42892 5092
rect 33376 5052 42892 5080
rect 33376 5040 33382 5052
rect 42886 5040 42892 5052
rect 42944 5040 42950 5092
rect 27632 4984 33272 5012
rect 33410 4972 33416 5024
rect 33468 4972 33474 5024
rect 37274 4972 37280 5024
rect 37332 4972 37338 5024
rect 37550 4972 37556 5024
rect 37608 4972 37614 5024
rect 43070 4972 43076 5024
rect 43128 4972 43134 5024
rect 1104 4922 43884 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 37950 4922
rect 38002 4870 38014 4922
rect 38066 4870 38078 4922
rect 38130 4870 38142 4922
rect 38194 4870 38206 4922
rect 38258 4870 43884 4922
rect 1104 4848 43884 4870
rect 2498 4768 2504 4820
rect 2556 4808 2562 4820
rect 13722 4808 13728 4820
rect 2556 4780 13728 4808
rect 2556 4768 2562 4780
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 17497 4811 17555 4817
rect 17497 4777 17509 4811
rect 17543 4808 17555 4811
rect 23842 4808 23848 4820
rect 17543 4780 23848 4808
rect 17543 4777 17555 4780
rect 17497 4771 17555 4777
rect 23842 4768 23848 4780
rect 23900 4768 23906 4820
rect 26786 4768 26792 4820
rect 26844 4808 26850 4820
rect 30101 4811 30159 4817
rect 30101 4808 30113 4811
rect 26844 4780 30113 4808
rect 26844 4768 26850 4780
rect 30101 4777 30113 4780
rect 30147 4777 30159 4811
rect 30101 4771 30159 4777
rect 30374 4768 30380 4820
rect 30432 4808 30438 4820
rect 36538 4808 36544 4820
rect 30432 4780 36544 4808
rect 30432 4768 30438 4780
rect 36538 4768 36544 4780
rect 36596 4768 36602 4820
rect 26329 4743 26387 4749
rect 26329 4740 26341 4743
rect 6886 4712 26341 4740
rect 5534 4632 5540 4684
rect 5592 4672 5598 4684
rect 6886 4672 6914 4712
rect 26329 4709 26341 4712
rect 26375 4709 26387 4743
rect 26329 4703 26387 4709
rect 26973 4743 27031 4749
rect 26973 4709 26985 4743
rect 27019 4740 27031 4743
rect 29914 4740 29920 4752
rect 27019 4712 29920 4740
rect 27019 4709 27031 4712
rect 26973 4703 27031 4709
rect 29914 4700 29920 4712
rect 29972 4700 29978 4752
rect 33502 4700 33508 4752
rect 33560 4740 33566 4752
rect 41966 4740 41972 4752
rect 33560 4712 41972 4740
rect 33560 4700 33566 4712
rect 41966 4700 41972 4712
rect 42024 4700 42030 4752
rect 43438 4700 43444 4752
rect 43496 4700 43502 4752
rect 5592 4644 6914 4672
rect 5592 4632 5598 4644
rect 11698 4632 11704 4684
rect 11756 4672 11762 4684
rect 11756 4644 17448 4672
rect 11756 4632 11762 4644
rect 6730 4564 6736 4616
rect 6788 4604 6794 4616
rect 7285 4607 7343 4613
rect 7285 4604 7297 4607
rect 6788 4576 7297 4604
rect 6788 4564 6794 4576
rect 7285 4573 7297 4576
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 8662 4564 8668 4616
rect 8720 4604 8726 4616
rect 8720 4576 13400 4604
rect 8720 4564 8726 4576
rect 13372 4536 13400 4576
rect 13446 4564 13452 4616
rect 13504 4564 13510 4616
rect 17313 4607 17371 4613
rect 17313 4573 17325 4607
rect 17359 4573 17371 4607
rect 17313 4567 17371 4573
rect 17328 4536 17356 4567
rect 6886 4508 12434 4536
rect 13372 4508 17356 4536
rect 17420 4536 17448 4644
rect 17494 4632 17500 4684
rect 17552 4672 17558 4684
rect 21818 4672 21824 4684
rect 17552 4644 21824 4672
rect 17552 4632 17558 4644
rect 21818 4632 21824 4644
rect 21876 4632 21882 4684
rect 24762 4632 24768 4684
rect 24820 4672 24826 4684
rect 28261 4675 28319 4681
rect 28261 4672 28273 4675
rect 24820 4644 28273 4672
rect 24820 4632 24826 4644
rect 28261 4641 28273 4644
rect 28307 4641 28319 4675
rect 28261 4635 28319 4641
rect 28718 4632 28724 4684
rect 28776 4672 28782 4684
rect 28776 4644 41414 4672
rect 28776 4632 28782 4644
rect 21450 4564 21456 4616
rect 21508 4604 21514 4616
rect 22189 4607 22247 4613
rect 22189 4604 22201 4607
rect 21508 4576 22201 4604
rect 21508 4564 21514 4576
rect 22189 4573 22201 4576
rect 22235 4573 22247 4607
rect 22189 4567 22247 4573
rect 26421 4607 26479 4613
rect 26421 4573 26433 4607
rect 26467 4604 26479 4607
rect 26513 4607 26571 4613
rect 26513 4604 26525 4607
rect 26467 4576 26525 4604
rect 26467 4573 26479 4576
rect 26421 4567 26479 4573
rect 26513 4573 26525 4576
rect 26559 4573 26571 4607
rect 26513 4567 26571 4573
rect 26789 4607 26847 4613
rect 26789 4573 26801 4607
rect 26835 4573 26847 4607
rect 26789 4567 26847 4573
rect 28353 4607 28411 4613
rect 28353 4573 28365 4607
rect 28399 4604 28411 4607
rect 28445 4607 28503 4613
rect 28445 4604 28457 4607
rect 28399 4576 28457 4604
rect 28399 4573 28411 4576
rect 28353 4567 28411 4573
rect 28445 4573 28457 4576
rect 28491 4573 28503 4607
rect 28445 4567 28503 4573
rect 30285 4607 30343 4613
rect 30285 4573 30297 4607
rect 30331 4604 30343 4607
rect 35618 4604 35624 4616
rect 30331 4576 35624 4604
rect 30331 4573 30343 4576
rect 30285 4567 30343 4573
rect 26804 4536 26832 4567
rect 35618 4564 35624 4576
rect 35676 4564 35682 4616
rect 41386 4604 41414 4644
rect 42889 4607 42947 4613
rect 42889 4604 42901 4607
rect 41386 4576 42901 4604
rect 42889 4573 42901 4576
rect 42935 4573 42947 4607
rect 42889 4567 42947 4573
rect 42978 4564 42984 4616
rect 43036 4604 43042 4616
rect 43257 4607 43315 4613
rect 43257 4604 43269 4607
rect 43036 4576 43269 4604
rect 43036 4564 43042 4576
rect 43257 4573 43269 4576
rect 43303 4573 43315 4607
rect 43257 4567 43315 4573
rect 27065 4539 27123 4545
rect 27065 4536 27077 4539
rect 17420 4508 27077 4536
rect 5442 4428 5448 4480
rect 5500 4468 5506 4480
rect 6886 4468 6914 4508
rect 5500 4440 6914 4468
rect 7469 4471 7527 4477
rect 5500 4428 5506 4440
rect 7469 4437 7481 4471
rect 7515 4468 7527 4471
rect 10962 4468 10968 4480
rect 7515 4440 10968 4468
rect 7515 4437 7527 4440
rect 7469 4431 7527 4437
rect 10962 4428 10968 4440
rect 11020 4428 11026 4480
rect 12406 4468 12434 4508
rect 27065 4505 27077 4508
rect 27111 4505 27123 4539
rect 27065 4499 27123 4505
rect 28644 4508 31754 4536
rect 13265 4471 13323 4477
rect 13265 4468 13277 4471
rect 12406 4440 13277 4468
rect 13265 4437 13277 4440
rect 13311 4437 13323 4471
rect 13265 4431 13323 4437
rect 13354 4428 13360 4480
rect 13412 4468 13418 4480
rect 17862 4468 17868 4480
rect 13412 4440 17868 4468
rect 13412 4428 13418 4440
rect 17862 4428 17868 4440
rect 17920 4428 17926 4480
rect 22373 4471 22431 4477
rect 22373 4437 22385 4471
rect 22419 4468 22431 4471
rect 25866 4468 25872 4480
rect 22419 4440 25872 4468
rect 22419 4437 22431 4440
rect 22373 4431 22431 4437
rect 25866 4428 25872 4440
rect 25924 4428 25930 4480
rect 26694 4428 26700 4480
rect 26752 4428 26758 4480
rect 28644 4477 28672 4508
rect 28629 4471 28687 4477
rect 28629 4437 28641 4471
rect 28675 4437 28687 4471
rect 31726 4468 31754 4508
rect 42886 4468 42892 4480
rect 31726 4440 42892 4468
rect 28629 4431 28687 4437
rect 42886 4428 42892 4440
rect 42944 4428 42950 4480
rect 43070 4428 43076 4480
rect 43128 4428 43134 4480
rect 1104 4378 43884 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 39010 4378
rect 39062 4326 39074 4378
rect 39126 4326 39138 4378
rect 39190 4326 39202 4378
rect 39254 4326 39266 4378
rect 39318 4326 43884 4378
rect 1104 4304 43884 4326
rect 1302 4224 1308 4276
rect 1360 4264 1366 4276
rect 26602 4264 26608 4276
rect 1360 4236 26608 4264
rect 1360 4224 1366 4236
rect 26602 4224 26608 4236
rect 26660 4224 26666 4276
rect 26694 4224 26700 4276
rect 26752 4264 26758 4276
rect 40034 4264 40040 4276
rect 26752 4236 40040 4264
rect 26752 4224 26758 4236
rect 40034 4224 40040 4236
rect 40092 4224 40098 4276
rect 1210 4156 1216 4208
rect 1268 4196 1274 4208
rect 28350 4196 28356 4208
rect 1268 4168 28356 4196
rect 1268 4156 1274 4168
rect 28350 4156 28356 4168
rect 28408 4156 28414 4208
rect 36538 4156 36544 4208
rect 36596 4196 36602 4208
rect 36596 4168 43300 4196
rect 36596 4156 36602 4168
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4097 2099 4131
rect 2041 4091 2099 4097
rect 4065 4131 4123 4137
rect 4065 4097 4077 4131
rect 4111 4128 4123 4131
rect 8386 4128 8392 4140
rect 4111 4100 8392 4128
rect 4111 4097 4123 4100
rect 4065 4091 4123 4097
rect 2056 4060 2084 4091
rect 8386 4088 8392 4100
rect 8444 4088 8450 4140
rect 17129 4131 17187 4137
rect 17129 4097 17141 4131
rect 17175 4128 17187 4131
rect 17402 4128 17408 4140
rect 17175 4100 17408 4128
rect 17175 4097 17187 4100
rect 17129 4091 17187 4097
rect 17402 4088 17408 4100
rect 17460 4088 17466 4140
rect 22094 4088 22100 4140
rect 22152 4128 22158 4140
rect 24213 4131 24271 4137
rect 24213 4128 24225 4131
rect 22152 4100 24225 4128
rect 22152 4088 22158 4100
rect 24213 4097 24225 4100
rect 24259 4097 24271 4131
rect 24213 4091 24271 4097
rect 27709 4131 27767 4137
rect 27709 4097 27721 4131
rect 27755 4128 27767 4131
rect 27798 4128 27804 4140
rect 27755 4100 27804 4128
rect 27755 4097 27767 4100
rect 27709 4091 27767 4097
rect 27798 4088 27804 4100
rect 27856 4088 27862 4140
rect 32401 4131 32459 4137
rect 32401 4097 32413 4131
rect 32447 4128 32459 4131
rect 32858 4128 32864 4140
rect 32447 4100 32864 4128
rect 32447 4097 32459 4100
rect 32401 4091 32459 4097
rect 32858 4088 32864 4100
rect 32916 4088 32922 4140
rect 43272 4137 43300 4168
rect 42889 4131 42947 4137
rect 42889 4128 42901 4131
rect 41386 4100 42901 4128
rect 5626 4060 5632 4072
rect 2056 4032 5632 4060
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 16114 4020 16120 4072
rect 16172 4060 16178 4072
rect 23750 4060 23756 4072
rect 16172 4032 23756 4060
rect 16172 4020 16178 4032
rect 23750 4020 23756 4032
rect 23808 4020 23814 4072
rect 29546 4020 29552 4072
rect 29604 4060 29610 4072
rect 41386 4060 41414 4100
rect 42889 4097 42901 4100
rect 42935 4097 42947 4131
rect 42889 4091 42947 4097
rect 43257 4131 43315 4137
rect 43257 4097 43269 4131
rect 43303 4097 43315 4131
rect 43257 4091 43315 4097
rect 29604 4032 41414 4060
rect 29604 4020 29610 4032
rect 2225 3995 2283 4001
rect 2225 3961 2237 3995
rect 2271 3992 2283 3995
rect 19702 3992 19708 4004
rect 2271 3964 19708 3992
rect 2271 3961 2283 3964
rect 2225 3955 2283 3961
rect 19702 3952 19708 3964
rect 19760 3952 19766 4004
rect 23842 3952 23848 4004
rect 23900 3992 23906 4004
rect 25682 3992 25688 4004
rect 23900 3964 25688 3992
rect 23900 3952 23906 3964
rect 25682 3952 25688 3964
rect 25740 3952 25746 4004
rect 25774 3952 25780 4004
rect 25832 3992 25838 4004
rect 27614 3992 27620 4004
rect 25832 3964 27620 3992
rect 25832 3952 25838 3964
rect 27614 3952 27620 3964
rect 27672 3952 27678 4004
rect 27893 3995 27951 4001
rect 27893 3961 27905 3995
rect 27939 3992 27951 3995
rect 33594 3992 33600 4004
rect 27939 3964 33600 3992
rect 27939 3961 27951 3964
rect 27893 3955 27951 3961
rect 33594 3952 33600 3964
rect 33652 3952 33658 4004
rect 43438 3952 43444 4004
rect 43496 3952 43502 4004
rect 4246 3884 4252 3936
rect 4304 3884 4310 3936
rect 17126 3884 17132 3936
rect 17184 3924 17190 3936
rect 17221 3927 17279 3933
rect 17221 3924 17233 3927
rect 17184 3896 17233 3924
rect 17184 3884 17190 3896
rect 17221 3893 17233 3896
rect 17267 3893 17279 3927
rect 17221 3887 17279 3893
rect 24397 3927 24455 3933
rect 24397 3893 24409 3927
rect 24443 3924 24455 3927
rect 30650 3924 30656 3936
rect 24443 3896 30656 3924
rect 24443 3893 24455 3896
rect 24397 3887 24455 3893
rect 30650 3884 30656 3896
rect 30708 3884 30714 3936
rect 31846 3884 31852 3936
rect 31904 3924 31910 3936
rect 32217 3927 32275 3933
rect 32217 3924 32229 3927
rect 31904 3896 32229 3924
rect 31904 3884 31910 3896
rect 32217 3893 32229 3896
rect 32263 3893 32275 3927
rect 32217 3887 32275 3893
rect 43070 3884 43076 3936
rect 43128 3884 43134 3936
rect 1104 3834 43884 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 37950 3834
rect 38002 3782 38014 3834
rect 38066 3782 38078 3834
rect 38130 3782 38142 3834
rect 38194 3782 38206 3834
rect 38258 3782 43884 3834
rect 1104 3760 43884 3782
rect 4246 3680 4252 3732
rect 4304 3720 4310 3732
rect 20346 3720 20352 3732
rect 4304 3692 20352 3720
rect 4304 3680 4310 3692
rect 20346 3680 20352 3692
rect 20404 3680 20410 3732
rect 20438 3680 20444 3732
rect 20496 3720 20502 3732
rect 21821 3723 21879 3729
rect 21821 3720 21833 3723
rect 20496 3692 21833 3720
rect 20496 3680 20502 3692
rect 21821 3689 21833 3692
rect 21867 3689 21879 3723
rect 21821 3683 21879 3689
rect 22020 3692 23336 3720
rect 13722 3612 13728 3664
rect 13780 3652 13786 3664
rect 20070 3652 20076 3664
rect 13780 3624 20076 3652
rect 13780 3612 13786 3624
rect 20070 3612 20076 3624
rect 20128 3612 20134 3664
rect 20162 3612 20168 3664
rect 20220 3612 20226 3664
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 21358 3584 21364 3596
rect 9640 3556 21364 3584
rect 9640 3544 9646 3556
rect 21358 3544 21364 3556
rect 21416 3544 21422 3596
rect 9398 3476 9404 3528
rect 9456 3516 9462 3528
rect 15473 3519 15531 3525
rect 15473 3516 15485 3519
rect 9456 3488 15485 3516
rect 9456 3476 9462 3488
rect 15473 3485 15485 3488
rect 15519 3485 15531 3519
rect 15473 3479 15531 3485
rect 18693 3519 18751 3525
rect 18693 3485 18705 3519
rect 18739 3485 18751 3519
rect 18693 3479 18751 3485
rect 13078 3408 13084 3460
rect 13136 3448 13142 3460
rect 18708 3448 18736 3479
rect 19518 3476 19524 3528
rect 19576 3516 19582 3528
rect 19705 3519 19763 3525
rect 19705 3516 19717 3519
rect 19576 3488 19717 3516
rect 19576 3476 19582 3488
rect 19705 3485 19717 3488
rect 19751 3485 19763 3519
rect 19705 3479 19763 3485
rect 19794 3476 19800 3528
rect 19852 3516 19858 3528
rect 22020 3525 22048 3692
rect 23308 3584 23336 3692
rect 23474 3680 23480 3732
rect 23532 3680 23538 3732
rect 23753 3723 23811 3729
rect 23753 3689 23765 3723
rect 23799 3720 23811 3723
rect 26326 3720 26332 3732
rect 23799 3692 26332 3720
rect 23799 3689 23811 3692
rect 23753 3683 23811 3689
rect 26326 3680 26332 3692
rect 26384 3680 26390 3732
rect 30285 3723 30343 3729
rect 30285 3689 30297 3723
rect 30331 3720 30343 3723
rect 34698 3720 34704 3732
rect 30331 3692 34704 3720
rect 30331 3689 30343 3692
rect 30285 3683 30343 3689
rect 34698 3680 34704 3692
rect 34756 3680 34762 3732
rect 23382 3612 23388 3664
rect 23440 3652 23446 3664
rect 24673 3655 24731 3661
rect 24673 3652 24685 3655
rect 23440 3624 24685 3652
rect 23440 3612 23446 3624
rect 24673 3621 24685 3624
rect 24719 3621 24731 3655
rect 24673 3615 24731 3621
rect 25041 3655 25099 3661
rect 25041 3621 25053 3655
rect 25087 3652 25099 3655
rect 25087 3624 31754 3652
rect 25087 3621 25099 3624
rect 25041 3615 25099 3621
rect 30374 3584 30380 3596
rect 23308 3556 30380 3584
rect 30374 3544 30380 3556
rect 30432 3544 30438 3596
rect 31726 3584 31754 3624
rect 34422 3612 34428 3664
rect 34480 3652 34486 3664
rect 34480 3624 43300 3652
rect 34480 3612 34486 3624
rect 42978 3584 42984 3596
rect 31726 3556 42984 3584
rect 42978 3544 42984 3556
rect 43036 3544 43042 3596
rect 19981 3519 20039 3525
rect 19981 3516 19993 3519
rect 19852 3488 19993 3516
rect 19852 3476 19858 3488
rect 19981 3485 19993 3488
rect 20027 3516 20039 3519
rect 20257 3519 20315 3525
rect 20257 3516 20269 3519
rect 20027 3488 20269 3516
rect 20027 3485 20039 3488
rect 19981 3479 20039 3485
rect 20257 3485 20269 3488
rect 20303 3485 20315 3519
rect 20257 3479 20315 3485
rect 22005 3519 22063 3525
rect 22005 3485 22017 3519
rect 22051 3485 22063 3519
rect 22005 3479 22063 3485
rect 23477 3519 23535 3525
rect 23477 3485 23489 3519
rect 23523 3516 23535 3519
rect 23569 3519 23627 3525
rect 23569 3516 23581 3519
rect 23523 3488 23581 3516
rect 23523 3485 23535 3488
rect 23477 3479 23535 3485
rect 23569 3485 23581 3488
rect 23615 3485 23627 3519
rect 23569 3479 23627 3485
rect 24765 3519 24823 3525
rect 24765 3485 24777 3519
rect 24811 3516 24823 3519
rect 24857 3519 24915 3525
rect 24857 3516 24869 3519
rect 24811 3488 24869 3516
rect 24811 3485 24823 3488
rect 24765 3479 24823 3485
rect 24857 3485 24869 3488
rect 24903 3485 24915 3519
rect 24857 3479 24915 3485
rect 26694 3476 26700 3528
rect 26752 3516 26758 3528
rect 27525 3519 27583 3525
rect 27525 3516 27537 3519
rect 26752 3488 27537 3516
rect 26752 3476 26758 3488
rect 27525 3485 27537 3488
rect 27571 3485 27583 3519
rect 30101 3519 30159 3525
rect 30101 3516 30113 3519
rect 27525 3479 27583 3485
rect 27632 3488 30113 3516
rect 23290 3448 23296 3460
rect 13136 3420 18736 3448
rect 18800 3420 23296 3448
rect 13136 3408 13142 3420
rect 15654 3340 15660 3392
rect 15712 3340 15718 3392
rect 15746 3340 15752 3392
rect 15804 3380 15810 3392
rect 18800 3380 18828 3420
rect 23290 3408 23296 3420
rect 23348 3408 23354 3460
rect 26234 3408 26240 3460
rect 26292 3448 26298 3460
rect 27632 3448 27660 3488
rect 30101 3485 30113 3488
rect 30147 3485 30159 3519
rect 30101 3479 30159 3485
rect 32401 3519 32459 3525
rect 32401 3485 32413 3519
rect 32447 3516 32459 3519
rect 34238 3516 34244 3528
rect 32447 3488 34244 3516
rect 32447 3485 32459 3488
rect 32401 3479 32459 3485
rect 34238 3476 34244 3488
rect 34296 3476 34302 3528
rect 42886 3476 42892 3528
rect 42944 3476 42950 3528
rect 43272 3525 43300 3624
rect 43438 3612 43444 3664
rect 43496 3612 43502 3664
rect 43257 3519 43315 3525
rect 43257 3485 43269 3519
rect 43303 3485 43315 3519
rect 43257 3479 43315 3485
rect 26292 3420 27660 3448
rect 26292 3408 26298 3420
rect 30006 3408 30012 3460
rect 30064 3448 30070 3460
rect 38102 3448 38108 3460
rect 30064 3420 38108 3448
rect 30064 3408 30070 3420
rect 38102 3408 38108 3420
rect 38160 3408 38166 3460
rect 15804 3352 18828 3380
rect 15804 3340 15810 3352
rect 18874 3340 18880 3392
rect 18932 3340 18938 3392
rect 19886 3340 19892 3392
rect 19944 3340 19950 3392
rect 27338 3340 27344 3392
rect 27396 3340 27402 3392
rect 31846 3340 31852 3392
rect 31904 3380 31910 3392
rect 32217 3383 32275 3389
rect 32217 3380 32229 3383
rect 31904 3352 32229 3380
rect 31904 3340 31910 3352
rect 32217 3349 32229 3352
rect 32263 3349 32275 3383
rect 32217 3343 32275 3349
rect 43070 3340 43076 3392
rect 43128 3340 43134 3392
rect 1104 3290 43884 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 39010 3290
rect 39062 3238 39074 3290
rect 39126 3238 39138 3290
rect 39190 3238 39202 3290
rect 39254 3238 39266 3290
rect 39318 3238 43884 3290
rect 1104 3216 43884 3238
rect 12621 3179 12679 3185
rect 12621 3145 12633 3179
rect 12667 3176 12679 3179
rect 12667 3148 14872 3176
rect 12667 3145 12679 3148
rect 12621 3139 12679 3145
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 5350 3040 5356 3052
rect 1903 3012 5356 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 7561 3043 7619 3049
rect 7561 3040 7573 3043
rect 6512 3012 7573 3040
rect 6512 3000 6518 3012
rect 7561 3009 7573 3012
rect 7607 3009 7619 3043
rect 7561 3003 7619 3009
rect 10318 3000 10324 3052
rect 10376 3040 10382 3052
rect 12437 3043 12495 3049
rect 12437 3040 12449 3043
rect 10376 3012 12449 3040
rect 10376 3000 10382 3012
rect 12437 3009 12449 3012
rect 12483 3009 12495 3043
rect 12437 3003 12495 3009
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3009 14611 3043
rect 14844 3040 14872 3148
rect 15654 3136 15660 3188
rect 15712 3176 15718 3188
rect 24486 3176 24492 3188
rect 15712 3148 24492 3176
rect 15712 3136 15718 3148
rect 24486 3136 24492 3148
rect 24544 3136 24550 3188
rect 25958 3136 25964 3188
rect 26016 3176 26022 3188
rect 30193 3179 30251 3185
rect 30193 3176 30205 3179
rect 26016 3148 30205 3176
rect 26016 3136 26022 3148
rect 30193 3145 30205 3148
rect 30239 3145 30251 3179
rect 30193 3139 30251 3145
rect 30561 3179 30619 3185
rect 30561 3145 30573 3179
rect 30607 3176 30619 3179
rect 31662 3176 31668 3188
rect 30607 3148 31668 3176
rect 30607 3145 30619 3148
rect 30561 3139 30619 3145
rect 31662 3136 31668 3148
rect 31720 3136 31726 3188
rect 31757 3179 31815 3185
rect 31757 3145 31769 3179
rect 31803 3176 31815 3179
rect 33042 3176 33048 3188
rect 31803 3148 33048 3176
rect 31803 3145 31815 3148
rect 31757 3139 31815 3145
rect 33042 3136 33048 3148
rect 33100 3136 33106 3188
rect 34238 3136 34244 3188
rect 34296 3136 34302 3188
rect 34422 3136 34428 3188
rect 34480 3176 34486 3188
rect 36817 3179 36875 3185
rect 36817 3176 36829 3179
rect 34480 3148 36829 3176
rect 34480 3136 34486 3148
rect 36817 3145 36829 3148
rect 36863 3145 36875 3179
rect 36817 3139 36875 3145
rect 38102 3136 38108 3188
rect 38160 3136 38166 3188
rect 43438 3136 43444 3188
rect 43496 3136 43502 3188
rect 14918 3068 14924 3120
rect 14976 3108 14982 3120
rect 14976 3080 16344 3108
rect 14976 3068 14982 3080
rect 15746 3040 15752 3052
rect 14844 3012 15752 3040
rect 14553 3003 14611 3009
rect 9766 2932 9772 2984
rect 9824 2972 9830 2984
rect 14568 2972 14596 3003
rect 15746 3000 15752 3012
rect 15804 3000 15810 3052
rect 16316 3049 16344 3080
rect 18874 3068 18880 3120
rect 18932 3108 18938 3120
rect 25590 3108 25596 3120
rect 18932 3080 25596 3108
rect 18932 3068 18938 3080
rect 25590 3068 25596 3080
rect 25648 3068 25654 3120
rect 27430 3108 27436 3120
rect 26712 3080 27436 3108
rect 15933 3043 15991 3049
rect 15933 3009 15945 3043
rect 15979 3009 15991 3043
rect 15933 3003 15991 3009
rect 16301 3043 16359 3049
rect 16301 3009 16313 3043
rect 16347 3009 16359 3043
rect 16301 3003 16359 3009
rect 9824 2944 14596 2972
rect 9824 2932 9830 2944
rect 8846 2864 8852 2916
rect 8904 2904 8910 2916
rect 15948 2904 15976 3003
rect 20070 3000 20076 3052
rect 20128 3000 20134 3052
rect 20714 3000 20720 3052
rect 20772 3040 20778 3052
rect 21177 3043 21235 3049
rect 21177 3040 21189 3043
rect 20772 3012 21189 3040
rect 20772 3000 20778 3012
rect 21177 3009 21189 3012
rect 21223 3009 21235 3043
rect 21177 3003 21235 3009
rect 21358 3000 21364 3052
rect 21416 3040 21422 3052
rect 22005 3043 22063 3049
rect 22005 3040 22017 3043
rect 21416 3012 22017 3040
rect 21416 3000 21422 3012
rect 22005 3009 22017 3012
rect 22051 3009 22063 3043
rect 22005 3003 22063 3009
rect 25317 3043 25375 3049
rect 25317 3009 25329 3043
rect 25363 3009 25375 3043
rect 25317 3003 25375 3009
rect 22370 2972 22376 2984
rect 8904 2876 15976 2904
rect 16040 2944 22376 2972
rect 8904 2864 8910 2876
rect 2041 2839 2099 2845
rect 2041 2805 2053 2839
rect 2087 2836 2099 2839
rect 7650 2836 7656 2848
rect 2087 2808 7656 2836
rect 2087 2805 2099 2808
rect 2041 2799 2099 2805
rect 7650 2796 7656 2808
rect 7708 2796 7714 2848
rect 7745 2839 7803 2845
rect 7745 2805 7757 2839
rect 7791 2836 7803 2839
rect 14274 2836 14280 2848
rect 7791 2808 14280 2836
rect 7791 2805 7803 2808
rect 7745 2799 7803 2805
rect 14274 2796 14280 2808
rect 14332 2796 14338 2848
rect 14737 2839 14795 2845
rect 14737 2805 14749 2839
rect 14783 2836 14795 2839
rect 16040 2836 16068 2944
rect 22370 2932 22376 2944
rect 22428 2932 22434 2984
rect 16114 2864 16120 2916
rect 16172 2864 16178 2916
rect 16485 2907 16543 2913
rect 16485 2873 16497 2907
rect 16531 2904 16543 2907
rect 25332 2904 25360 3003
rect 25866 3000 25872 3052
rect 25924 3000 25930 3052
rect 26712 3049 26740 3080
rect 27430 3068 27436 3080
rect 27488 3068 27494 3120
rect 33410 3108 33416 3120
rect 31312 3080 33416 3108
rect 26697 3043 26755 3049
rect 26697 3009 26709 3043
rect 26743 3009 26755 3043
rect 26697 3003 26755 3009
rect 27157 3043 27215 3049
rect 27157 3009 27169 3043
rect 27203 3040 27215 3043
rect 27249 3043 27307 3049
rect 27249 3040 27261 3043
rect 27203 3012 27261 3040
rect 27203 3009 27215 3012
rect 27157 3003 27215 3009
rect 27249 3009 27261 3012
rect 27295 3009 27307 3043
rect 27249 3003 27307 3009
rect 27522 3000 27528 3052
rect 27580 3000 27586 3052
rect 27614 3000 27620 3052
rect 27672 3040 27678 3052
rect 28353 3043 28411 3049
rect 28353 3040 28365 3043
rect 27672 3012 28365 3040
rect 27672 3000 27678 3012
rect 28353 3009 28365 3012
rect 28399 3009 28411 3043
rect 28353 3003 28411 3009
rect 28721 3043 28779 3049
rect 28721 3009 28733 3043
rect 28767 3009 28779 3043
rect 28721 3003 28779 3009
rect 26602 2932 26608 2984
rect 26660 2972 26666 2984
rect 27065 2975 27123 2981
rect 27065 2972 27077 2975
rect 26660 2944 27077 2972
rect 26660 2932 26666 2944
rect 27065 2941 27077 2944
rect 27111 2941 27123 2975
rect 28736 2972 28764 3003
rect 30006 3000 30012 3052
rect 30064 3000 30070 3052
rect 30285 3043 30343 3049
rect 30285 3009 30297 3043
rect 30331 3040 30343 3043
rect 30377 3043 30435 3049
rect 30377 3040 30389 3043
rect 30331 3012 30389 3040
rect 30331 3009 30343 3012
rect 30285 3003 30343 3009
rect 30377 3009 30389 3012
rect 30423 3009 30435 3043
rect 31018 3040 31024 3052
rect 30377 3003 30435 3009
rect 30760 3012 31024 3040
rect 27065 2935 27123 2941
rect 27172 2944 28764 2972
rect 16531 2876 25360 2904
rect 16531 2873 16543 2876
rect 16485 2867 16543 2873
rect 25406 2864 25412 2916
rect 25464 2904 25470 2916
rect 27172 2904 27200 2944
rect 30098 2932 30104 2984
rect 30156 2972 30162 2984
rect 30760 2972 30788 3012
rect 31018 3000 31024 3012
rect 31076 3000 31082 3052
rect 31125 3043 31183 3049
rect 31125 3009 31137 3043
rect 31171 3040 31183 3043
rect 31312 3040 31340 3080
rect 33410 3068 33416 3080
rect 33468 3068 33474 3120
rect 42334 3068 42340 3120
rect 42392 3108 42398 3120
rect 42392 3080 43300 3108
rect 42392 3068 42398 3080
rect 31171 3012 31340 3040
rect 31389 3043 31447 3049
rect 31171 3009 31183 3012
rect 31125 3003 31183 3009
rect 31389 3009 31401 3043
rect 31435 3040 31447 3043
rect 31573 3043 31631 3049
rect 31573 3040 31585 3043
rect 31435 3012 31585 3040
rect 31435 3009 31447 3012
rect 31389 3003 31447 3009
rect 31573 3009 31585 3012
rect 31619 3009 31631 3043
rect 31573 3003 31631 3009
rect 32401 3043 32459 3049
rect 32401 3009 32413 3043
rect 32447 3040 32459 3043
rect 32493 3043 32551 3049
rect 32493 3040 32505 3043
rect 32447 3012 32505 3040
rect 32447 3009 32459 3012
rect 32401 3003 32459 3009
rect 32493 3009 32505 3012
rect 32539 3009 32551 3043
rect 32493 3003 32551 3009
rect 32766 3000 32772 3052
rect 32824 3040 32830 3052
rect 33045 3043 33103 3049
rect 33045 3040 33057 3043
rect 32824 3012 33057 3040
rect 32824 3000 32830 3012
rect 33045 3009 33057 3012
rect 33091 3009 33103 3043
rect 33045 3003 33103 3009
rect 33229 3043 33287 3049
rect 33229 3009 33241 3043
rect 33275 3009 33287 3043
rect 33229 3003 33287 3009
rect 30156 2944 30788 2972
rect 30156 2932 30162 2944
rect 30834 2932 30840 2984
rect 30892 2972 30898 2984
rect 31478 2972 31484 2984
rect 30892 2944 31484 2972
rect 30892 2932 30898 2944
rect 31478 2932 31484 2944
rect 31536 2932 31542 2984
rect 31662 2932 31668 2984
rect 31720 2972 31726 2984
rect 33244 2972 33272 3003
rect 33594 3000 33600 3052
rect 33652 3000 33658 3052
rect 34149 3043 34207 3049
rect 34149 3009 34161 3043
rect 34195 3040 34207 3043
rect 34425 3043 34483 3049
rect 34425 3040 34437 3043
rect 34195 3012 34437 3040
rect 34195 3009 34207 3012
rect 34149 3003 34207 3009
rect 34425 3009 34437 3012
rect 34471 3009 34483 3043
rect 34425 3003 34483 3009
rect 34701 3043 34759 3049
rect 34701 3009 34713 3043
rect 34747 3040 34759 3043
rect 34790 3040 34796 3052
rect 34747 3012 34796 3040
rect 34747 3009 34759 3012
rect 34701 3003 34759 3009
rect 34790 3000 34796 3012
rect 34848 3000 34854 3052
rect 35161 3043 35219 3049
rect 35161 3009 35173 3043
rect 35207 3009 35219 3043
rect 35161 3003 35219 3009
rect 31720 2944 33272 2972
rect 31720 2932 31726 2944
rect 33686 2932 33692 2984
rect 33744 2972 33750 2984
rect 35176 2972 35204 3003
rect 35710 3000 35716 3052
rect 35768 3040 35774 3052
rect 36081 3043 36139 3049
rect 36081 3040 36093 3043
rect 35768 3012 36093 3040
rect 35768 3000 35774 3012
rect 36081 3009 36093 3012
rect 36127 3009 36139 3043
rect 36081 3003 36139 3009
rect 36998 3000 37004 3052
rect 37056 3000 37062 3052
rect 37090 3000 37096 3052
rect 37148 3040 37154 3052
rect 38289 3043 38347 3049
rect 38289 3040 38301 3043
rect 37148 3012 38301 3040
rect 37148 3000 37154 3012
rect 38289 3009 38301 3012
rect 38335 3009 38347 3043
rect 38289 3003 38347 3009
rect 40034 3000 40040 3052
rect 40092 3040 40098 3052
rect 42521 3043 42579 3049
rect 42521 3040 42533 3043
rect 40092 3012 42533 3040
rect 40092 3000 40098 3012
rect 42521 3009 42533 3012
rect 42567 3009 42579 3043
rect 42521 3003 42579 3009
rect 42889 3043 42947 3049
rect 42889 3009 42901 3043
rect 42935 3040 42947 3043
rect 43162 3040 43168 3052
rect 42935 3012 43168 3040
rect 42935 3009 42947 3012
rect 42889 3003 42947 3009
rect 43162 3000 43168 3012
rect 43220 3000 43226 3052
rect 43272 3049 43300 3080
rect 43257 3043 43315 3049
rect 43257 3009 43269 3043
rect 43303 3009 43315 3043
rect 43257 3003 43315 3009
rect 33744 2944 35204 2972
rect 33744 2932 33750 2944
rect 25464 2876 27200 2904
rect 27433 2907 27491 2913
rect 25464 2864 25470 2876
rect 27433 2873 27445 2907
rect 27479 2904 27491 2907
rect 28718 2904 28724 2916
rect 27479 2876 28724 2904
rect 27479 2873 27491 2876
rect 27433 2867 27491 2873
rect 28718 2864 28724 2876
rect 28776 2864 28782 2916
rect 28994 2864 29000 2916
rect 29052 2904 29058 2916
rect 32309 2907 32367 2913
rect 32309 2904 32321 2907
rect 29052 2876 32321 2904
rect 29052 2864 29058 2876
rect 32309 2873 32321 2876
rect 32355 2873 32367 2907
rect 32309 2867 32367 2873
rect 32677 2907 32735 2913
rect 32677 2873 32689 2907
rect 32723 2904 32735 2907
rect 33594 2904 33600 2916
rect 32723 2876 33600 2904
rect 32723 2873 32735 2876
rect 32677 2867 32735 2873
rect 33594 2864 33600 2876
rect 33652 2864 33658 2916
rect 33870 2864 33876 2916
rect 33928 2904 33934 2916
rect 34517 2907 34575 2913
rect 34517 2904 34529 2907
rect 33928 2876 34529 2904
rect 33928 2864 33934 2876
rect 34517 2873 34529 2876
rect 34563 2873 34575 2907
rect 35897 2907 35955 2913
rect 35897 2904 35909 2907
rect 34517 2867 34575 2873
rect 34624 2876 35909 2904
rect 14783 2808 16068 2836
rect 14783 2805 14795 2808
rect 14737 2799 14795 2805
rect 19794 2796 19800 2848
rect 19852 2836 19858 2848
rect 20257 2839 20315 2845
rect 20257 2836 20269 2839
rect 19852 2808 20269 2836
rect 19852 2796 19858 2808
rect 20257 2805 20269 2808
rect 20303 2805 20315 2839
rect 20257 2799 20315 2805
rect 20898 2796 20904 2848
rect 20956 2836 20962 2848
rect 21361 2839 21419 2845
rect 21361 2836 21373 2839
rect 20956 2808 21373 2836
rect 20956 2796 20962 2808
rect 21361 2805 21373 2808
rect 21407 2805 21419 2839
rect 21361 2799 21419 2805
rect 21910 2796 21916 2848
rect 21968 2836 21974 2848
rect 22189 2839 22247 2845
rect 22189 2836 22201 2839
rect 21968 2808 22201 2836
rect 21968 2796 21974 2808
rect 22189 2805 22201 2808
rect 22235 2805 22247 2839
rect 22189 2799 22247 2805
rect 25222 2796 25228 2848
rect 25280 2836 25286 2848
rect 25501 2839 25559 2845
rect 25501 2836 25513 2839
rect 25280 2808 25513 2836
rect 25280 2796 25286 2808
rect 25501 2805 25513 2808
rect 25547 2805 25559 2839
rect 25501 2799 25559 2805
rect 25774 2796 25780 2848
rect 25832 2836 25838 2848
rect 26053 2839 26111 2845
rect 26053 2836 26065 2839
rect 25832 2808 26065 2836
rect 25832 2796 25838 2808
rect 26053 2805 26065 2808
rect 26099 2805 26111 2839
rect 26053 2799 26111 2805
rect 26326 2796 26332 2848
rect 26384 2836 26390 2848
rect 26513 2839 26571 2845
rect 26513 2836 26525 2839
rect 26384 2808 26525 2836
rect 26384 2796 26390 2808
rect 26513 2805 26525 2808
rect 26559 2805 26571 2839
rect 26513 2799 26571 2805
rect 27522 2796 27528 2848
rect 27580 2836 27586 2848
rect 27709 2839 27767 2845
rect 27709 2836 27721 2839
rect 27580 2808 27721 2836
rect 27580 2796 27586 2808
rect 27709 2805 27721 2808
rect 27755 2805 27767 2839
rect 27709 2799 27767 2805
rect 28258 2796 28264 2848
rect 28316 2836 28322 2848
rect 28537 2839 28595 2845
rect 28537 2836 28549 2839
rect 28316 2808 28549 2836
rect 28316 2796 28322 2808
rect 28537 2805 28549 2808
rect 28583 2805 28595 2839
rect 28537 2799 28595 2805
rect 28626 2796 28632 2848
rect 28684 2836 28690 2848
rect 28905 2839 28963 2845
rect 28905 2836 28917 2839
rect 28684 2808 28917 2836
rect 28684 2796 28690 2808
rect 28905 2805 28917 2808
rect 28951 2805 28963 2839
rect 28905 2799 28963 2805
rect 29638 2796 29644 2848
rect 29696 2836 29702 2848
rect 29825 2839 29883 2845
rect 29825 2836 29837 2839
rect 29696 2808 29837 2836
rect 29696 2796 29702 2808
rect 29825 2805 29837 2808
rect 29871 2805 29883 2839
rect 29825 2799 29883 2805
rect 30742 2796 30748 2848
rect 30800 2836 30806 2848
rect 30929 2839 30987 2845
rect 30929 2836 30941 2839
rect 30800 2808 30941 2836
rect 30800 2796 30806 2808
rect 30929 2805 30941 2808
rect 30975 2805 30987 2839
rect 30929 2799 30987 2805
rect 31018 2796 31024 2848
rect 31076 2836 31082 2848
rect 31389 2839 31447 2845
rect 31389 2836 31401 2839
rect 31076 2808 31401 2836
rect 31076 2796 31082 2808
rect 31389 2805 31401 2808
rect 31435 2805 31447 2839
rect 31389 2799 31447 2805
rect 31478 2796 31484 2848
rect 31536 2836 31542 2848
rect 32766 2836 32772 2848
rect 31536 2808 32772 2836
rect 31536 2796 31542 2808
rect 32766 2796 32772 2808
rect 32824 2796 32830 2848
rect 32950 2796 32956 2848
rect 33008 2796 33014 2848
rect 33410 2796 33416 2848
rect 33468 2796 33474 2848
rect 33502 2796 33508 2848
rect 33560 2836 33566 2848
rect 33781 2839 33839 2845
rect 33781 2836 33793 2839
rect 33560 2808 33793 2836
rect 33560 2796 33566 2808
rect 33781 2805 33793 2808
rect 33827 2805 33839 2839
rect 33781 2799 33839 2805
rect 33962 2796 33968 2848
rect 34020 2836 34026 2848
rect 34057 2839 34115 2845
rect 34057 2836 34069 2839
rect 34020 2808 34069 2836
rect 34020 2796 34026 2808
rect 34057 2805 34069 2808
rect 34103 2805 34115 2839
rect 34057 2799 34115 2805
rect 34330 2796 34336 2848
rect 34388 2836 34394 2848
rect 34624 2836 34652 2876
rect 35897 2873 35909 2876
rect 35943 2873 35955 2907
rect 35897 2867 35955 2873
rect 34388 2808 34652 2836
rect 34388 2796 34394 2808
rect 34974 2796 34980 2848
rect 35032 2796 35038 2848
rect 42705 2839 42763 2845
rect 42705 2805 42717 2839
rect 42751 2836 42763 2839
rect 42978 2836 42984 2848
rect 42751 2808 42984 2836
rect 42751 2805 42763 2808
rect 42705 2799 42763 2805
rect 42978 2796 42984 2808
rect 43036 2796 43042 2848
rect 43070 2796 43076 2848
rect 43128 2796 43134 2848
rect 1104 2746 43884 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 37950 2746
rect 38002 2694 38014 2746
rect 38066 2694 38078 2746
rect 38130 2694 38142 2746
rect 38194 2694 38206 2746
rect 38258 2694 43884 2746
rect 1104 2672 43884 2694
rect 10962 2592 10968 2644
rect 11020 2632 11026 2644
rect 24949 2635 25007 2641
rect 24949 2632 24961 2635
rect 11020 2604 22094 2632
rect 11020 2592 11026 2604
rect 8266 2536 20300 2564
rect 7650 2456 7656 2508
rect 7708 2496 7714 2508
rect 8266 2496 8294 2536
rect 7708 2468 8294 2496
rect 7708 2456 7714 2468
rect 7466 2388 7472 2440
rect 7524 2428 7530 2440
rect 7524 2400 12434 2428
rect 7524 2388 7530 2400
rect 12406 2360 12434 2400
rect 12986 2388 12992 2440
rect 13044 2428 13050 2440
rect 19521 2431 19579 2437
rect 19521 2428 19533 2431
rect 13044 2400 19533 2428
rect 13044 2388 13050 2400
rect 19521 2397 19533 2400
rect 19567 2397 19579 2431
rect 19521 2391 19579 2397
rect 19702 2388 19708 2440
rect 19760 2428 19766 2440
rect 20272 2437 20300 2536
rect 20714 2524 20720 2576
rect 20772 2564 20778 2576
rect 21450 2564 21456 2576
rect 20772 2536 21456 2564
rect 20772 2524 20778 2536
rect 21450 2524 21456 2536
rect 21508 2524 21514 2576
rect 21726 2496 21732 2508
rect 21376 2468 21732 2496
rect 19889 2431 19947 2437
rect 19889 2428 19901 2431
rect 19760 2400 19901 2428
rect 19760 2388 19766 2400
rect 19889 2397 19901 2400
rect 19935 2397 19947 2431
rect 19889 2391 19947 2397
rect 20257 2431 20315 2437
rect 20257 2397 20269 2431
rect 20303 2397 20315 2431
rect 20257 2391 20315 2397
rect 20346 2388 20352 2440
rect 20404 2428 20410 2440
rect 21376 2437 21404 2468
rect 21726 2456 21732 2468
rect 21784 2456 21790 2508
rect 20625 2431 20683 2437
rect 20625 2428 20637 2431
rect 20404 2400 20637 2428
rect 20404 2388 20410 2400
rect 20625 2397 20637 2400
rect 20671 2397 20683 2431
rect 20625 2391 20683 2397
rect 20993 2431 21051 2437
rect 20993 2397 21005 2431
rect 21039 2397 21051 2431
rect 20993 2391 21051 2397
rect 21361 2431 21419 2437
rect 21361 2397 21373 2431
rect 21407 2397 21419 2431
rect 21361 2391 21419 2397
rect 21008 2360 21036 2391
rect 21542 2388 21548 2440
rect 21600 2428 21606 2440
rect 21821 2431 21879 2437
rect 21821 2428 21833 2431
rect 21600 2400 21833 2428
rect 21600 2388 21606 2400
rect 21821 2397 21833 2400
rect 21867 2397 21879 2431
rect 22066 2428 22094 2604
rect 24780 2604 24961 2632
rect 24118 2524 24124 2576
rect 24176 2564 24182 2576
rect 24780 2564 24808 2604
rect 24949 2601 24961 2604
rect 24995 2601 25007 2635
rect 24949 2595 25007 2601
rect 25038 2592 25044 2644
rect 25096 2632 25102 2644
rect 25317 2635 25375 2641
rect 25317 2632 25329 2635
rect 25096 2604 25329 2632
rect 25096 2592 25102 2604
rect 25317 2601 25329 2604
rect 25363 2601 25375 2635
rect 25317 2595 25375 2601
rect 27338 2592 27344 2644
rect 27396 2632 27402 2644
rect 28261 2635 28319 2641
rect 28261 2632 28273 2635
rect 27396 2604 28273 2632
rect 27396 2592 27402 2604
rect 28261 2601 28273 2604
rect 28307 2601 28319 2635
rect 28261 2595 28319 2601
rect 30190 2592 30196 2644
rect 30248 2632 30254 2644
rect 31665 2635 31723 2641
rect 31665 2632 31677 2635
rect 30248 2604 31677 2632
rect 30248 2592 30254 2604
rect 31665 2601 31677 2604
rect 31711 2601 31723 2635
rect 31665 2595 31723 2601
rect 32398 2592 32404 2644
rect 32456 2632 32462 2644
rect 33781 2635 33839 2641
rect 33781 2632 33793 2635
rect 32456 2604 33793 2632
rect 32456 2592 32462 2604
rect 33781 2601 33793 2604
rect 33827 2601 33839 2635
rect 33781 2595 33839 2601
rect 41386 2604 42932 2632
rect 24176 2536 24808 2564
rect 24176 2524 24182 2536
rect 25498 2524 25504 2576
rect 25556 2564 25562 2576
rect 26421 2567 26479 2573
rect 26421 2564 26433 2567
rect 25556 2536 26433 2564
rect 25556 2524 25562 2536
rect 26421 2533 26433 2536
rect 26467 2533 26479 2567
rect 26421 2527 26479 2533
rect 26602 2524 26608 2576
rect 26660 2564 26666 2576
rect 27525 2567 27583 2573
rect 27525 2564 27537 2567
rect 26660 2536 27537 2564
rect 26660 2524 26666 2536
rect 27525 2533 27537 2536
rect 27571 2533 27583 2567
rect 27525 2527 27583 2533
rect 27706 2524 27712 2576
rect 27764 2564 27770 2576
rect 28629 2567 28687 2573
rect 28629 2564 28641 2567
rect 27764 2536 28641 2564
rect 27764 2524 27770 2536
rect 28629 2533 28641 2536
rect 28675 2533 28687 2567
rect 28629 2527 28687 2533
rect 28810 2524 28816 2576
rect 28868 2564 28874 2576
rect 29733 2567 29791 2573
rect 29733 2564 29745 2567
rect 28868 2536 29745 2564
rect 28868 2524 28874 2536
rect 29733 2533 29745 2536
rect 29779 2533 29791 2567
rect 29733 2527 29791 2533
rect 29914 2524 29920 2576
rect 29972 2564 29978 2576
rect 30745 2567 30803 2573
rect 30745 2564 30757 2567
rect 29972 2536 30757 2564
rect 29972 2524 29978 2536
rect 30745 2533 30757 2536
rect 30791 2533 30803 2567
rect 30745 2527 30803 2533
rect 31294 2524 31300 2576
rect 31352 2564 31358 2576
rect 32585 2567 32643 2573
rect 32585 2564 32597 2567
rect 31352 2536 32597 2564
rect 31352 2524 31358 2536
rect 32585 2533 32597 2536
rect 32631 2533 32643 2567
rect 41386 2564 41414 2604
rect 32585 2527 32643 2533
rect 32876 2536 41414 2564
rect 22370 2456 22376 2508
rect 22428 2496 22434 2508
rect 22428 2468 24440 2496
rect 22428 2456 22434 2468
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 22066 2400 22201 2428
rect 21821 2391 21879 2397
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 22554 2388 22560 2440
rect 22612 2388 22618 2440
rect 22922 2388 22928 2440
rect 22980 2388 22986 2440
rect 23290 2388 23296 2440
rect 23348 2388 23354 2440
rect 23382 2388 23388 2440
rect 23440 2428 23446 2440
rect 24412 2437 24440 2468
rect 24964 2468 25544 2496
rect 23661 2431 23719 2437
rect 23661 2428 23673 2431
rect 23440 2400 23673 2428
rect 23440 2388 23446 2400
rect 23661 2397 23673 2400
rect 23707 2397 23719 2431
rect 23661 2391 23719 2397
rect 24397 2431 24455 2437
rect 24397 2397 24409 2431
rect 24443 2397 24455 2431
rect 24397 2391 24455 2397
rect 24762 2388 24768 2440
rect 24820 2388 24826 2440
rect 24964 2428 24992 2468
rect 24872 2400 24992 2428
rect 25133 2431 25191 2437
rect 12406 2332 21036 2360
rect 21450 2320 21456 2372
rect 21508 2360 21514 2372
rect 23198 2360 23204 2372
rect 21508 2332 23204 2360
rect 21508 2320 21514 2332
rect 23198 2320 23204 2332
rect 23256 2320 23262 2372
rect 23750 2320 23756 2372
rect 23808 2360 23814 2372
rect 24872 2360 24900 2400
rect 25133 2397 25145 2431
rect 25179 2428 25191 2431
rect 25314 2428 25320 2440
rect 25179 2400 25320 2428
rect 25179 2397 25191 2400
rect 25133 2391 25191 2397
rect 25314 2388 25320 2400
rect 25372 2388 25378 2440
rect 25516 2437 25544 2468
rect 25590 2456 25596 2508
rect 25648 2496 25654 2508
rect 25648 2468 28120 2496
rect 25648 2456 25654 2468
rect 25501 2431 25559 2437
rect 25501 2397 25513 2431
rect 25547 2397 25559 2431
rect 25501 2391 25559 2397
rect 25682 2388 25688 2440
rect 25740 2428 25746 2440
rect 25869 2431 25927 2437
rect 25869 2428 25881 2431
rect 25740 2400 25881 2428
rect 25740 2388 25746 2400
rect 25869 2397 25881 2400
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 25958 2388 25964 2440
rect 26016 2428 26022 2440
rect 26237 2431 26295 2437
rect 26237 2428 26249 2431
rect 26016 2400 26249 2428
rect 26016 2388 26022 2400
rect 26237 2397 26249 2400
rect 26283 2397 26295 2431
rect 26237 2391 26295 2397
rect 27246 2388 27252 2440
rect 27304 2388 27310 2440
rect 27341 2431 27399 2437
rect 27341 2397 27353 2431
rect 27387 2428 27399 2431
rect 27522 2428 27528 2440
rect 27387 2400 27528 2428
rect 27387 2397 27399 2400
rect 27341 2391 27399 2397
rect 27522 2388 27528 2400
rect 27580 2388 27586 2440
rect 27614 2388 27620 2440
rect 27672 2428 27678 2440
rect 28092 2437 28120 2468
rect 30006 2456 30012 2508
rect 30064 2496 30070 2508
rect 32876 2496 32904 2536
rect 30064 2468 32904 2496
rect 30064 2456 30070 2468
rect 32950 2456 32956 2508
rect 33008 2496 33014 2508
rect 33008 2468 33272 2496
rect 33008 2456 33014 2468
rect 27709 2431 27767 2437
rect 27709 2428 27721 2431
rect 27672 2400 27721 2428
rect 27672 2388 27678 2400
rect 27709 2397 27721 2400
rect 27755 2397 27767 2431
rect 27709 2391 27767 2397
rect 28077 2431 28135 2437
rect 28077 2397 28089 2431
rect 28123 2397 28135 2431
rect 28077 2391 28135 2397
rect 28442 2388 28448 2440
rect 28500 2388 28506 2440
rect 28626 2388 28632 2440
rect 28684 2428 28690 2440
rect 28813 2431 28871 2437
rect 28813 2428 28825 2431
rect 28684 2400 28825 2428
rect 28684 2388 28690 2400
rect 28813 2397 28825 2400
rect 28859 2397 28871 2431
rect 28813 2391 28871 2397
rect 29546 2388 29552 2440
rect 29604 2388 29610 2440
rect 29730 2388 29736 2440
rect 29788 2428 29794 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29788 2400 29929 2428
rect 29788 2388 29794 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 30282 2388 30288 2440
rect 30340 2388 30346 2440
rect 30926 2388 30932 2440
rect 30984 2388 30990 2440
rect 31478 2388 31484 2440
rect 31536 2388 31542 2440
rect 31849 2431 31907 2437
rect 31849 2397 31861 2431
rect 31895 2428 31907 2431
rect 32306 2428 32312 2440
rect 31895 2400 32312 2428
rect 31895 2397 31907 2400
rect 31849 2391 31907 2397
rect 32306 2388 32312 2400
rect 32364 2388 32370 2440
rect 32401 2431 32459 2437
rect 32401 2397 32413 2431
rect 32447 2428 32459 2431
rect 32674 2428 32680 2440
rect 32447 2400 32680 2428
rect 32447 2397 32459 2400
rect 32401 2391 32459 2397
rect 32674 2388 32680 2400
rect 32732 2388 32738 2440
rect 32766 2388 32772 2440
rect 32824 2388 32830 2440
rect 33244 2437 33272 2468
rect 33318 2456 33324 2508
rect 33376 2496 33382 2508
rect 33376 2468 34008 2496
rect 33376 2456 33382 2468
rect 33137 2431 33195 2437
rect 33137 2397 33149 2431
rect 33183 2397 33195 2431
rect 33137 2391 33195 2397
rect 33229 2431 33287 2437
rect 33229 2397 33241 2431
rect 33275 2397 33287 2431
rect 33229 2391 33287 2397
rect 23808 2332 24900 2360
rect 23808 2320 23814 2332
rect 24946 2320 24952 2372
rect 25004 2360 25010 2372
rect 25004 2332 26096 2360
rect 25004 2320 25010 2332
rect 19702 2252 19708 2304
rect 19760 2252 19766 2304
rect 20073 2295 20131 2301
rect 20073 2261 20085 2295
rect 20119 2292 20131 2295
rect 20254 2292 20260 2304
rect 20119 2264 20260 2292
rect 20119 2261 20131 2264
rect 20073 2255 20131 2261
rect 20254 2252 20260 2264
rect 20312 2252 20318 2304
rect 20441 2295 20499 2301
rect 20441 2261 20453 2295
rect 20487 2292 20499 2295
rect 20530 2292 20536 2304
rect 20487 2264 20536 2292
rect 20487 2261 20499 2264
rect 20441 2255 20499 2261
rect 20530 2252 20536 2264
rect 20588 2252 20594 2304
rect 20806 2252 20812 2304
rect 20864 2252 20870 2304
rect 21177 2295 21235 2301
rect 21177 2261 21189 2295
rect 21223 2292 21235 2295
rect 21358 2292 21364 2304
rect 21223 2264 21364 2292
rect 21223 2261 21235 2264
rect 21177 2255 21235 2261
rect 21358 2252 21364 2264
rect 21416 2252 21422 2304
rect 21545 2295 21603 2301
rect 21545 2261 21557 2295
rect 21591 2292 21603 2295
rect 21634 2292 21640 2304
rect 21591 2264 21640 2292
rect 21591 2261 21603 2264
rect 21545 2255 21603 2261
rect 21634 2252 21640 2264
rect 21692 2252 21698 2304
rect 22005 2295 22063 2301
rect 22005 2261 22017 2295
rect 22051 2292 22063 2295
rect 22186 2292 22192 2304
rect 22051 2264 22192 2292
rect 22051 2261 22063 2264
rect 22005 2255 22063 2261
rect 22186 2252 22192 2264
rect 22244 2252 22250 2304
rect 22373 2295 22431 2301
rect 22373 2261 22385 2295
rect 22419 2292 22431 2295
rect 22462 2292 22468 2304
rect 22419 2264 22468 2292
rect 22419 2261 22431 2264
rect 22373 2255 22431 2261
rect 22462 2252 22468 2264
rect 22520 2252 22526 2304
rect 22738 2252 22744 2304
rect 22796 2252 22802 2304
rect 23014 2252 23020 2304
rect 23072 2292 23078 2304
rect 23109 2295 23167 2301
rect 23109 2292 23121 2295
rect 23072 2264 23121 2292
rect 23072 2252 23078 2264
rect 23109 2261 23121 2264
rect 23155 2261 23167 2295
rect 23109 2255 23167 2261
rect 23290 2252 23296 2304
rect 23348 2292 23354 2304
rect 23477 2295 23535 2301
rect 23477 2292 23489 2295
rect 23348 2264 23489 2292
rect 23348 2252 23354 2264
rect 23477 2261 23489 2264
rect 23523 2261 23535 2295
rect 23477 2255 23535 2261
rect 23566 2252 23572 2304
rect 23624 2292 23630 2304
rect 23845 2295 23903 2301
rect 23845 2292 23857 2295
rect 23624 2264 23857 2292
rect 23624 2252 23630 2264
rect 23845 2261 23857 2264
rect 23891 2261 23903 2295
rect 23845 2255 23903 2261
rect 23934 2252 23940 2304
rect 23992 2292 23998 2304
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 23992 2264 24593 2292
rect 23992 2252 23998 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 24670 2252 24676 2304
rect 24728 2292 24734 2304
rect 26068 2301 26096 2332
rect 26878 2320 26884 2372
rect 26936 2360 26942 2372
rect 26936 2332 27936 2360
rect 26936 2320 26942 2332
rect 25685 2295 25743 2301
rect 25685 2292 25697 2295
rect 24728 2264 25697 2292
rect 24728 2252 24734 2264
rect 25685 2261 25697 2264
rect 25731 2261 25743 2295
rect 25685 2255 25743 2261
rect 26053 2295 26111 2301
rect 26053 2261 26065 2295
rect 26099 2261 26111 2295
rect 26053 2255 26111 2261
rect 26142 2252 26148 2304
rect 26200 2292 26206 2304
rect 27908 2301 27936 2332
rect 27982 2320 27988 2372
rect 28040 2360 28046 2372
rect 28040 2332 29040 2360
rect 28040 2320 28046 2332
rect 29012 2301 29040 2332
rect 29362 2320 29368 2372
rect 29420 2360 29426 2372
rect 29420 2332 30512 2360
rect 29420 2320 29426 2332
rect 27065 2295 27123 2301
rect 27065 2292 27077 2295
rect 26200 2264 27077 2292
rect 26200 2252 26206 2264
rect 27065 2261 27077 2264
rect 27111 2261 27123 2295
rect 27065 2255 27123 2261
rect 27893 2295 27951 2301
rect 27893 2261 27905 2295
rect 27939 2261 27951 2295
rect 27893 2255 27951 2261
rect 28997 2295 29055 2301
rect 28997 2261 29009 2295
rect 29043 2261 29055 2295
rect 28997 2255 29055 2261
rect 29086 2252 29092 2304
rect 29144 2292 29150 2304
rect 30484 2301 30512 2332
rect 30558 2320 30564 2372
rect 30616 2360 30622 2372
rect 30616 2332 31432 2360
rect 30616 2320 30622 2332
rect 30101 2295 30159 2301
rect 30101 2292 30113 2295
rect 29144 2264 30113 2292
rect 29144 2252 29150 2264
rect 30101 2261 30113 2264
rect 30147 2261 30159 2295
rect 30101 2255 30159 2261
rect 30469 2295 30527 2301
rect 30469 2261 30481 2295
rect 30515 2261 30527 2295
rect 30469 2255 30527 2261
rect 31018 2252 31024 2304
rect 31076 2292 31082 2304
rect 31297 2295 31355 2301
rect 31297 2292 31309 2295
rect 31076 2264 31309 2292
rect 31076 2252 31082 2264
rect 31297 2261 31309 2264
rect 31343 2261 31355 2295
rect 31404 2292 31432 2332
rect 31570 2320 31576 2372
rect 31628 2360 31634 2372
rect 33152 2360 33180 2391
rect 33594 2388 33600 2440
rect 33652 2388 33658 2440
rect 33778 2388 33784 2440
rect 33836 2388 33842 2440
rect 33980 2437 34008 2468
rect 33965 2431 34023 2437
rect 33965 2397 33977 2431
rect 34011 2397 34023 2431
rect 33965 2391 34023 2397
rect 34698 2388 34704 2440
rect 34756 2388 34762 2440
rect 35066 2388 35072 2440
rect 35124 2388 35130 2440
rect 41966 2388 41972 2440
rect 42024 2388 42030 2440
rect 42518 2388 42524 2440
rect 42576 2388 42582 2440
rect 42904 2437 42932 2604
rect 43438 2524 43444 2576
rect 43496 2524 43502 2576
rect 42889 2431 42947 2437
rect 42889 2397 42901 2431
rect 42935 2397 42947 2431
rect 42889 2391 42947 2397
rect 43257 2431 43315 2437
rect 43257 2397 43269 2431
rect 43303 2428 43315 2431
rect 43303 2400 43944 2428
rect 43303 2397 43315 2400
rect 43257 2391 43315 2397
rect 33796 2360 33824 2388
rect 31628 2332 32996 2360
rect 33152 2332 33824 2360
rect 31628 2320 31634 2332
rect 32968 2301 32996 2332
rect 33870 2320 33876 2372
rect 33928 2360 33934 2372
rect 33928 2332 35296 2360
rect 33928 2320 33934 2332
rect 32217 2295 32275 2301
rect 32217 2292 32229 2295
rect 31404 2264 32229 2292
rect 31297 2255 31355 2261
rect 32217 2261 32229 2264
rect 32263 2261 32275 2295
rect 32217 2255 32275 2261
rect 32953 2295 33011 2301
rect 32953 2261 32965 2295
rect 32999 2261 33011 2295
rect 32953 2255 33011 2261
rect 33134 2252 33140 2304
rect 33192 2292 33198 2304
rect 33413 2295 33471 2301
rect 33413 2292 33425 2295
rect 33192 2264 33425 2292
rect 33192 2252 33198 2264
rect 33413 2261 33425 2264
rect 33459 2261 33471 2295
rect 33413 2255 33471 2261
rect 33594 2252 33600 2304
rect 33652 2292 33658 2304
rect 34149 2295 34207 2301
rect 34149 2292 34161 2295
rect 33652 2264 34161 2292
rect 33652 2252 33658 2264
rect 34149 2261 34161 2264
rect 34195 2261 34207 2295
rect 34149 2255 34207 2261
rect 34238 2252 34244 2304
rect 34296 2292 34302 2304
rect 35268 2301 35296 2332
rect 34885 2295 34943 2301
rect 34885 2292 34897 2295
rect 34296 2264 34897 2292
rect 34296 2252 34302 2264
rect 34885 2261 34897 2264
rect 34931 2261 34943 2295
rect 34885 2255 34943 2261
rect 35253 2295 35311 2301
rect 35253 2261 35265 2295
rect 35299 2261 35311 2295
rect 35253 2255 35311 2261
rect 42150 2252 42156 2304
rect 42208 2252 42214 2304
rect 42702 2252 42708 2304
rect 42760 2252 42766 2304
rect 43070 2252 43076 2304
rect 43128 2252 43134 2304
rect 1104 2202 43884 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 39010 2202
rect 39062 2150 39074 2202
rect 39126 2150 39138 2202
rect 39190 2150 39202 2202
rect 39254 2150 39266 2202
rect 39318 2150 43884 2202
rect 1104 2128 43884 2150
rect 16298 2048 16304 2100
rect 16356 2088 16362 2100
rect 21450 2088 21456 2100
rect 16356 2060 21456 2088
rect 16356 2048 16362 2060
rect 21450 2048 21456 2060
rect 21508 2048 21514 2100
rect 26786 2088 26792 2100
rect 21560 2060 26792 2088
rect 19426 1980 19432 2032
rect 19484 2020 19490 2032
rect 21560 2020 21588 2060
rect 26786 2048 26792 2060
rect 26844 2048 26850 2100
rect 32766 2048 32772 2100
rect 32824 2088 32830 2100
rect 34330 2088 34336 2100
rect 32824 2060 34336 2088
rect 32824 2048 32830 2060
rect 34330 2048 34336 2060
rect 34388 2048 34394 2100
rect 19484 1992 21588 2020
rect 19484 1980 19490 1992
rect 23198 1980 23204 2032
rect 23256 2020 23262 2032
rect 28442 2020 28448 2032
rect 23256 1992 28448 2020
rect 23256 1980 23262 1992
rect 28442 1980 28448 1992
rect 28500 1980 28506 2032
rect 32674 1980 32680 2032
rect 32732 2020 32738 2032
rect 34974 2020 34980 2032
rect 32732 1992 34980 2020
rect 32732 1980 32738 1992
rect 34974 1980 34980 1992
rect 35032 1980 35038 2032
rect 16942 1912 16948 1964
rect 17000 1952 17006 1964
rect 24854 1952 24860 1964
rect 17000 1924 24860 1952
rect 17000 1912 17006 1924
rect 24854 1912 24860 1924
rect 24912 1912 24918 1964
rect 25130 1912 25136 1964
rect 25188 1952 25194 1964
rect 29730 1952 29736 1964
rect 25188 1924 29736 1952
rect 25188 1912 25194 1924
rect 29730 1912 29736 1924
rect 29788 1912 29794 1964
rect 32306 1912 32312 1964
rect 32364 1952 32370 1964
rect 35342 1952 35348 1964
rect 32364 1924 35348 1952
rect 32364 1912 32370 1924
rect 35342 1912 35348 1924
rect 35400 1912 35406 1964
rect 43916 1952 43944 2400
rect 41386 1924 43944 1952
rect 16022 1844 16028 1896
rect 16080 1884 16086 1896
rect 28626 1884 28632 1896
rect 16080 1856 24900 1884
rect 16080 1844 16086 1856
rect 14274 1776 14280 1828
rect 14332 1816 14338 1828
rect 22554 1816 22560 1828
rect 14332 1788 22560 1816
rect 14332 1776 14338 1788
rect 22554 1776 22560 1788
rect 22612 1776 22618 1828
rect 14826 1708 14832 1760
rect 14884 1748 14890 1760
rect 24872 1748 24900 1856
rect 25240 1856 28632 1884
rect 25240 1748 25268 1856
rect 28626 1844 28632 1856
rect 28684 1844 28690 1896
rect 31478 1844 31484 1896
rect 31536 1884 31542 1896
rect 34422 1884 34428 1896
rect 31536 1856 34428 1884
rect 31536 1844 31542 1856
rect 34422 1844 34428 1856
rect 34480 1844 34486 1896
rect 30926 1776 30932 1828
rect 30984 1816 30990 1828
rect 37274 1816 37280 1828
rect 30984 1788 37280 1816
rect 30984 1776 30990 1788
rect 37274 1776 37280 1788
rect 37332 1776 37338 1828
rect 14884 1720 24716 1748
rect 24872 1720 25268 1748
rect 14884 1708 14890 1720
rect 13170 1640 13176 1692
rect 13228 1680 13234 1692
rect 22922 1680 22928 1692
rect 13228 1652 22928 1680
rect 13228 1640 13234 1652
rect 22922 1640 22928 1652
rect 22980 1640 22986 1692
rect 24688 1680 24716 1720
rect 26786 1708 26792 1760
rect 26844 1748 26850 1760
rect 37090 1748 37096 1760
rect 26844 1720 37096 1748
rect 26844 1708 26850 1720
rect 37090 1708 37096 1720
rect 37148 1708 37154 1760
rect 27522 1680 27528 1692
rect 24688 1652 27528 1680
rect 27522 1640 27528 1652
rect 27580 1640 27586 1692
rect 30650 1640 30656 1692
rect 30708 1680 30714 1692
rect 35066 1680 35072 1692
rect 30708 1652 35072 1680
rect 30708 1640 30714 1652
rect 35066 1640 35072 1652
rect 35124 1640 35130 1692
rect 20622 1572 20628 1624
rect 20680 1612 20686 1624
rect 27614 1612 27620 1624
rect 20680 1584 27620 1612
rect 20680 1572 20686 1584
rect 27614 1572 27620 1584
rect 27672 1572 27678 1624
rect 41386 1612 41414 1924
rect 31726 1584 41414 1612
rect 26418 1504 26424 1556
rect 26476 1544 26482 1556
rect 31726 1544 31754 1584
rect 26476 1516 31754 1544
rect 26476 1504 26482 1516
rect 24854 1436 24860 1488
rect 24912 1476 24918 1488
rect 30834 1476 30840 1488
rect 24912 1448 30840 1476
rect 24912 1436 24918 1448
rect 30834 1436 30840 1448
rect 30892 1436 30898 1488
rect 14458 1368 14464 1420
rect 14516 1408 14522 1420
rect 20714 1408 20720 1420
rect 14516 1380 20720 1408
rect 14516 1368 14522 1380
rect 20714 1368 20720 1380
rect 20772 1368 20778 1420
rect 24394 1368 24400 1420
rect 24452 1408 24458 1420
rect 24762 1408 24768 1420
rect 24452 1380 24768 1408
rect 24452 1368 24458 1380
rect 24762 1368 24768 1380
rect 24820 1368 24826 1420
rect 34238 1408 34244 1420
rect 33244 1380 34244 1408
rect 33244 1352 33272 1380
rect 34238 1368 34244 1380
rect 34296 1368 34302 1420
rect 33226 1300 33232 1352
rect 33284 1300 33290 1352
rect 32858 1232 32864 1284
rect 32916 1272 32922 1284
rect 35434 1272 35440 1284
rect 32916 1244 35440 1272
rect 32916 1232 32922 1244
rect 35434 1232 35440 1244
rect 35492 1232 35498 1284
rect 11698 1096 11704 1148
rect 11756 1136 11762 1148
rect 17678 1136 17684 1148
rect 11756 1108 17684 1136
rect 11756 1096 11762 1108
rect 17678 1096 17684 1108
rect 17736 1096 17742 1148
rect 15286 416 15292 468
rect 15344 456 15350 468
rect 22094 456 22100 468
rect 15344 428 22100 456
rect 15344 416 15350 428
rect 22094 416 22100 428
rect 22152 416 22158 468
rect 16114 348 16120 400
rect 16172 388 16178 400
rect 25866 388 25872 400
rect 16172 360 25872 388
rect 16172 348 16178 360
rect 25866 348 25872 360
rect 25924 348 25930 400
rect 15562 280 15568 332
rect 15620 320 15626 332
rect 27798 320 27804 332
rect 15620 292 27804 320
rect 15620 280 15626 292
rect 27798 280 27804 292
rect 27856 280 27862 332
rect 14182 212 14188 264
rect 14240 252 14246 264
rect 26694 252 26700 264
rect 14240 224 26700 252
rect 14240 212 14246 224
rect 26694 212 26700 224
rect 26752 212 26758 264
rect 17218 144 17224 196
rect 17276 184 17282 196
rect 33962 184 33968 196
rect 17276 156 33968 184
rect 17276 144 17282 156
rect 33962 144 33968 156
rect 34020 144 34026 196
rect 19242 76 19248 128
rect 19300 116 19306 128
rect 37550 116 37556 128
rect 19300 88 37556 116
rect 19300 76 19306 88
rect 37550 76 37556 88
rect 37608 76 37614 128
rect 18138 8 18144 60
rect 18196 48 18202 60
rect 36998 48 37004 60
rect 18196 20 37004 48
rect 18196 8 18202 20
rect 36998 8 37004 20
rect 37056 8 37062 60
<< via1 >>
rect 16488 9052 16540 9104
rect 25872 9120 25924 9172
rect 18604 8984 18656 9036
rect 25504 9052 25556 9104
rect 24860 8984 24912 9036
rect 22928 8916 22980 8968
rect 26148 8916 26200 8968
rect 12256 8780 12308 8832
rect 31852 8848 31904 8900
rect 20720 8780 20772 8832
rect 22744 8780 22796 8832
rect 22836 8780 22888 8832
rect 31024 8780 31076 8832
rect 41420 8780 41472 8832
rect 43628 8780 43680 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 39010 8678 39062 8730
rect 39074 8678 39126 8730
rect 39138 8678 39190 8730
rect 39202 8678 39254 8730
rect 39266 8678 39318 8730
rect 1308 8576 1360 8628
rect 3424 8576 3476 8628
rect 5540 8576 5592 8628
rect 7656 8576 7708 8628
rect 9772 8576 9824 8628
rect 11888 8576 11940 8628
rect 12256 8576 12308 8628
rect 14004 8576 14056 8628
rect 16120 8576 16172 8628
rect 18236 8576 18288 8628
rect 20352 8576 20404 8628
rect 22468 8576 22520 8628
rect 24584 8576 24636 8628
rect 26700 8576 26752 8628
rect 27160 8576 27212 8628
rect 28724 8576 28776 8628
rect 28816 8576 28868 8628
rect 30932 8576 30984 8628
rect 32864 8576 32916 8628
rect 35164 8576 35216 8628
rect 37280 8576 37332 8628
rect 39396 8576 39448 8628
rect 41420 8619 41472 8628
rect 41420 8585 41429 8619
rect 41429 8585 41463 8619
rect 41463 8585 41472 8619
rect 41420 8576 41472 8585
rect 41512 8576 41564 8628
rect 42156 8619 42208 8628
rect 42156 8585 42165 8619
rect 42165 8585 42199 8619
rect 42199 8585 42208 8619
rect 42156 8576 42208 8585
rect 42708 8619 42760 8628
rect 42708 8585 42717 8619
rect 42717 8585 42751 8619
rect 42751 8585 42760 8619
rect 42708 8576 42760 8585
rect 5816 8440 5868 8492
rect 6828 8440 6880 8492
rect 5448 8372 5500 8424
rect 16488 8483 16540 8492
rect 16488 8449 16497 8483
rect 16497 8449 16531 8483
rect 16531 8449 16540 8483
rect 16488 8440 16540 8449
rect 18604 8483 18656 8492
rect 18604 8449 18613 8483
rect 18613 8449 18647 8483
rect 18647 8449 18656 8483
rect 18604 8440 18656 8449
rect 20720 8483 20772 8492
rect 20720 8449 20729 8483
rect 20729 8449 20763 8483
rect 20763 8449 20772 8483
rect 20720 8440 20772 8449
rect 17132 8372 17184 8424
rect 23756 8508 23808 8560
rect 22836 8483 22888 8492
rect 22836 8449 22845 8483
rect 22845 8449 22879 8483
rect 22879 8449 22888 8483
rect 22836 8440 22888 8449
rect 27160 8440 27212 8492
rect 26792 8372 26844 8424
rect 29184 8483 29236 8492
rect 29184 8449 29193 8483
rect 29193 8449 29227 8483
rect 29227 8449 29236 8483
rect 29184 8440 29236 8449
rect 29368 8508 29420 8560
rect 29092 8372 29144 8424
rect 33324 8440 33376 8492
rect 34980 8440 35032 8492
rect 35072 8440 35124 8492
rect 37648 8483 37700 8492
rect 37648 8449 37657 8483
rect 37657 8449 37691 8483
rect 37691 8449 37700 8483
rect 37648 8440 37700 8449
rect 39856 8483 39908 8492
rect 39856 8449 39865 8483
rect 39865 8449 39899 8483
rect 39899 8449 39908 8483
rect 39856 8440 39908 8449
rect 41236 8483 41288 8492
rect 41236 8449 41245 8483
rect 41245 8449 41279 8483
rect 41279 8449 41288 8483
rect 41236 8440 41288 8449
rect 41604 8483 41656 8492
rect 41604 8449 41613 8483
rect 41613 8449 41647 8483
rect 41647 8449 41656 8483
rect 41604 8440 41656 8449
rect 40040 8372 40092 8424
rect 20444 8304 20496 8356
rect 23388 8304 23440 8356
rect 21364 8236 21416 8288
rect 23204 8236 23256 8288
rect 26148 8236 26200 8288
rect 28172 8236 28224 8288
rect 40040 8236 40092 8288
rect 43076 8347 43128 8356
rect 43076 8313 43085 8347
rect 43085 8313 43119 8347
rect 43119 8313 43128 8347
rect 43076 8304 43128 8313
rect 43444 8347 43496 8356
rect 43444 8313 43453 8347
rect 43453 8313 43487 8347
rect 43487 8313 43496 8347
rect 43444 8304 43496 8313
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 37950 8134 38002 8186
rect 38014 8134 38066 8186
rect 38078 8134 38130 8186
rect 38142 8134 38194 8186
rect 38206 8134 38258 8186
rect 14924 8032 14976 8084
rect 21272 8032 21324 8084
rect 21364 8075 21416 8084
rect 21364 8041 21373 8075
rect 21373 8041 21407 8075
rect 21407 8041 21416 8075
rect 21364 8032 21416 8041
rect 20720 8007 20772 8016
rect 20720 7973 20729 8007
rect 20729 7973 20763 8007
rect 20763 7973 20772 8007
rect 20720 7964 20772 7973
rect 23388 8032 23440 8084
rect 23756 8075 23808 8084
rect 23756 8041 23765 8075
rect 23765 8041 23799 8075
rect 23799 8041 23808 8075
rect 23756 8032 23808 8041
rect 24860 8032 24912 8084
rect 26332 8075 26384 8084
rect 26332 8041 26341 8075
rect 26341 8041 26375 8075
rect 26375 8041 26384 8075
rect 26332 8032 26384 8041
rect 29368 8032 29420 8084
rect 41972 8075 42024 8084
rect 41972 8041 41981 8075
rect 41981 8041 42015 8075
rect 42015 8041 42024 8075
rect 41972 8032 42024 8041
rect 42340 8075 42392 8084
rect 42340 8041 42349 8075
rect 42349 8041 42383 8075
rect 42383 8041 42392 8075
rect 42340 8032 42392 8041
rect 42616 8032 42668 8084
rect 23112 7964 23164 8016
rect 23204 7964 23256 8016
rect 7840 7828 7892 7880
rect 10876 7828 10928 7880
rect 19340 7871 19392 7880
rect 19340 7837 19349 7871
rect 19349 7837 19383 7871
rect 19383 7837 19392 7871
rect 19340 7828 19392 7837
rect 20352 7871 20404 7880
rect 20352 7837 20361 7871
rect 20361 7837 20395 7871
rect 20395 7837 20404 7871
rect 20352 7828 20404 7837
rect 20996 7828 21048 7880
rect 21272 7828 21324 7880
rect 36544 7896 36596 7948
rect 23664 7828 23716 7880
rect 27528 7871 27580 7880
rect 27528 7837 27537 7871
rect 27537 7837 27571 7871
rect 27571 7837 27580 7871
rect 27528 7828 27580 7837
rect 28356 7871 28408 7880
rect 28356 7837 28365 7871
rect 28365 7837 28399 7871
rect 28399 7837 28408 7871
rect 28356 7828 28408 7837
rect 29552 7871 29604 7880
rect 29552 7837 29561 7871
rect 29561 7837 29595 7871
rect 29595 7837 29604 7871
rect 29552 7828 29604 7837
rect 41788 7871 41840 7880
rect 41788 7837 41797 7871
rect 41797 7837 41831 7871
rect 41831 7837 41840 7871
rect 41788 7828 41840 7837
rect 7564 7760 7616 7812
rect 42616 7828 42668 7880
rect 43260 7871 43312 7880
rect 43260 7837 43269 7871
rect 43269 7837 43303 7871
rect 43303 7837 43312 7871
rect 43260 7828 43312 7837
rect 3976 7735 4028 7744
rect 3976 7701 3985 7735
rect 3985 7701 4019 7735
rect 4019 7701 4028 7735
rect 3976 7692 4028 7701
rect 4344 7735 4396 7744
rect 4344 7701 4353 7735
rect 4353 7701 4387 7735
rect 4387 7701 4396 7735
rect 4344 7692 4396 7701
rect 8852 7692 8904 7744
rect 9404 7692 9456 7744
rect 19064 7692 19116 7744
rect 20996 7692 21048 7744
rect 23480 7735 23532 7744
rect 23480 7701 23489 7735
rect 23489 7701 23523 7735
rect 23523 7701 23532 7735
rect 23480 7692 23532 7701
rect 26884 7735 26936 7744
rect 26884 7701 26893 7735
rect 26893 7701 26927 7735
rect 26927 7701 26936 7735
rect 26884 7692 26936 7701
rect 27252 7735 27304 7744
rect 27252 7701 27261 7735
rect 27261 7701 27295 7735
rect 27295 7701 27304 7735
rect 27252 7692 27304 7701
rect 27436 7692 27488 7744
rect 28172 7735 28224 7744
rect 28172 7701 28181 7735
rect 28181 7701 28215 7735
rect 28215 7701 28224 7735
rect 28172 7692 28224 7701
rect 29736 7735 29788 7744
rect 29736 7701 29745 7735
rect 29745 7701 29779 7735
rect 29779 7701 29788 7735
rect 29736 7692 29788 7701
rect 43076 7735 43128 7744
rect 43076 7701 43085 7735
rect 43085 7701 43119 7735
rect 43119 7701 43128 7735
rect 43076 7692 43128 7701
rect 43444 7735 43496 7744
rect 43444 7701 43453 7735
rect 43453 7701 43487 7735
rect 43487 7701 43496 7735
rect 43444 7692 43496 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 39010 7590 39062 7642
rect 39074 7590 39126 7642
rect 39138 7590 39190 7642
rect 39202 7590 39254 7642
rect 39266 7590 39318 7642
rect 4344 7488 4396 7540
rect 20720 7488 20772 7540
rect 20812 7488 20864 7540
rect 27528 7488 27580 7540
rect 29736 7488 29788 7540
rect 41788 7488 41840 7540
rect 43168 7488 43220 7540
rect 18052 7420 18104 7472
rect 18788 7327 18840 7336
rect 18788 7293 18797 7327
rect 18797 7293 18831 7327
rect 18831 7293 18840 7327
rect 18788 7284 18840 7293
rect 11152 7216 11204 7268
rect 20352 7352 20404 7404
rect 22008 7395 22060 7404
rect 22008 7361 22017 7395
rect 22017 7361 22051 7395
rect 22051 7361 22060 7395
rect 22008 7352 22060 7361
rect 23112 7352 23164 7404
rect 25136 7352 25188 7404
rect 20628 7284 20680 7336
rect 27344 7420 27396 7472
rect 29460 7420 29512 7472
rect 36820 7420 36872 7472
rect 36544 7352 36596 7404
rect 28356 7284 28408 7336
rect 36452 7284 36504 7336
rect 13728 7148 13780 7200
rect 21824 7148 21876 7200
rect 22192 7191 22244 7200
rect 22192 7157 22201 7191
rect 22201 7157 22235 7191
rect 22235 7157 22244 7191
rect 22192 7148 22244 7157
rect 31024 7191 31076 7200
rect 31024 7157 31033 7191
rect 31033 7157 31067 7191
rect 31067 7157 31076 7191
rect 31024 7148 31076 7157
rect 43444 7191 43496 7200
rect 43444 7157 43453 7191
rect 43453 7157 43487 7191
rect 43487 7157 43496 7191
rect 43444 7148 43496 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 37950 7046 38002 7098
rect 38014 7046 38066 7098
rect 38078 7046 38130 7098
rect 38142 7046 38194 7098
rect 38206 7046 38258 7098
rect 3976 6944 4028 6996
rect 13728 6944 13780 6996
rect 13820 6944 13872 6996
rect 20812 6944 20864 6996
rect 22192 6944 22244 6996
rect 35624 6944 35676 6996
rect 9588 6919 9640 6928
rect 9588 6885 9597 6919
rect 9597 6885 9631 6919
rect 9631 6885 9640 6919
rect 9588 6876 9640 6885
rect 20628 6876 20680 6928
rect 25228 6876 25280 6928
rect 12532 6808 12584 6860
rect 6184 6740 6236 6792
rect 10048 6740 10100 6792
rect 10600 6740 10652 6792
rect 16488 6808 16540 6860
rect 25412 6876 25464 6928
rect 43260 6876 43312 6928
rect 10232 6672 10284 6724
rect 12256 6672 12308 6724
rect 18696 6740 18748 6792
rect 38476 6740 38528 6792
rect 42984 6740 43036 6792
rect 9588 6604 9640 6656
rect 12900 6604 12952 6656
rect 13176 6604 13228 6656
rect 14924 6604 14976 6656
rect 22008 6672 22060 6724
rect 24952 6715 25004 6724
rect 24952 6681 24961 6715
rect 24961 6681 24995 6715
rect 24995 6681 25004 6715
rect 24952 6672 25004 6681
rect 16028 6647 16080 6656
rect 16028 6613 16037 6647
rect 16037 6613 16071 6647
rect 16071 6613 16080 6647
rect 16028 6604 16080 6613
rect 16304 6647 16356 6656
rect 16304 6613 16313 6647
rect 16313 6613 16347 6647
rect 16347 6613 16356 6647
rect 16304 6604 16356 6613
rect 29368 6672 29420 6724
rect 29552 6604 29604 6656
rect 29828 6647 29880 6656
rect 29828 6613 29837 6647
rect 29837 6613 29871 6647
rect 29871 6613 29880 6647
rect 29828 6604 29880 6613
rect 34428 6604 34480 6656
rect 35072 6647 35124 6656
rect 35072 6613 35081 6647
rect 35081 6613 35115 6647
rect 35115 6613 35124 6647
rect 35072 6604 35124 6613
rect 43076 6647 43128 6656
rect 43076 6613 43085 6647
rect 43085 6613 43119 6647
rect 43119 6613 43128 6647
rect 43076 6604 43128 6613
rect 43444 6647 43496 6656
rect 43444 6613 43453 6647
rect 43453 6613 43487 6647
rect 43487 6613 43496 6647
rect 43444 6604 43496 6613
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 39010 6502 39062 6554
rect 39074 6502 39126 6554
rect 39138 6502 39190 6554
rect 39202 6502 39254 6554
rect 39266 6502 39318 6554
rect 5816 6400 5868 6452
rect 12348 6400 12400 6452
rect 18052 6443 18104 6452
rect 18052 6409 18061 6443
rect 18061 6409 18095 6443
rect 18095 6409 18104 6443
rect 18052 6400 18104 6409
rect 20904 6400 20956 6452
rect 25504 6443 25556 6452
rect 25504 6409 25513 6443
rect 25513 6409 25547 6443
rect 25547 6409 25556 6443
rect 25504 6400 25556 6409
rect 10232 6332 10284 6384
rect 12992 6332 13044 6384
rect 15200 6332 15252 6384
rect 24676 6332 24728 6384
rect 7288 6264 7340 6316
rect 9404 6307 9456 6316
rect 9404 6273 9413 6307
rect 9413 6273 9447 6307
rect 9447 6273 9456 6307
rect 9404 6264 9456 6273
rect 13636 6264 13688 6316
rect 14740 6196 14792 6248
rect 17684 6196 17736 6248
rect 21456 6264 21508 6316
rect 27528 6400 27580 6452
rect 29184 6400 29236 6452
rect 36268 6400 36320 6452
rect 37648 6400 37700 6452
rect 39856 6400 39908 6452
rect 41236 6400 41288 6452
rect 43444 6443 43496 6452
rect 43444 6409 43453 6443
rect 43453 6409 43487 6443
rect 43487 6409 43496 6443
rect 43444 6400 43496 6409
rect 35624 6332 35676 6384
rect 43168 6332 43220 6384
rect 1308 6128 1360 6180
rect 18788 6128 18840 6180
rect 9588 6060 9640 6112
rect 11060 6103 11112 6112
rect 11060 6069 11069 6103
rect 11069 6069 11103 6103
rect 11103 6069 11112 6103
rect 11060 6060 11112 6069
rect 14832 6060 14884 6112
rect 15016 6060 15068 6112
rect 29828 6196 29880 6248
rect 37648 6264 37700 6316
rect 37188 6196 37240 6248
rect 38936 6264 38988 6316
rect 39396 6264 39448 6316
rect 39580 6264 39632 6316
rect 42892 6307 42944 6316
rect 42892 6273 42901 6307
rect 42901 6273 42935 6307
rect 42935 6273 42944 6307
rect 42892 6264 42944 6273
rect 43260 6307 43312 6316
rect 43260 6273 43269 6307
rect 43269 6273 43303 6307
rect 43303 6273 43312 6307
rect 43260 6264 43312 6273
rect 38752 6196 38804 6248
rect 29460 6128 29512 6180
rect 20536 6103 20588 6112
rect 20536 6069 20545 6103
rect 20545 6069 20579 6103
rect 20579 6069 20588 6103
rect 20536 6060 20588 6069
rect 25412 6060 25464 6112
rect 28724 6060 28776 6112
rect 33232 6128 33284 6180
rect 37372 6128 37424 6180
rect 41604 6128 41656 6180
rect 42340 6060 42392 6112
rect 43076 6103 43128 6112
rect 43076 6069 43085 6103
rect 43085 6069 43119 6103
rect 43119 6069 43128 6103
rect 43076 6060 43128 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 37950 5958 38002 6010
rect 38014 5958 38066 6010
rect 38078 5958 38130 6010
rect 38142 5958 38194 6010
rect 38206 5958 38258 6010
rect 11612 5856 11664 5908
rect 14924 5856 14976 5908
rect 15200 5899 15252 5908
rect 15200 5865 15209 5899
rect 15209 5865 15243 5899
rect 15243 5865 15252 5899
rect 15200 5856 15252 5865
rect 21456 5856 21508 5908
rect 940 5788 992 5840
rect 11980 5720 12032 5772
rect 7012 5652 7064 5704
rect 9496 5652 9548 5704
rect 15292 5695 15344 5704
rect 15292 5661 15301 5695
rect 15301 5661 15335 5695
rect 15335 5661 15344 5695
rect 15292 5652 15344 5661
rect 18788 5788 18840 5840
rect 21640 5831 21692 5840
rect 21640 5797 21649 5831
rect 21649 5797 21683 5831
rect 21683 5797 21692 5831
rect 21640 5788 21692 5797
rect 25412 5856 25464 5908
rect 42984 5856 43036 5908
rect 26056 5788 26108 5840
rect 25780 5652 25832 5704
rect 28356 5695 28408 5704
rect 28356 5661 28365 5695
rect 28365 5661 28399 5695
rect 28399 5661 28408 5695
rect 28356 5652 28408 5661
rect 29092 5652 29144 5704
rect 33232 5720 33284 5772
rect 33416 5788 33468 5840
rect 35808 5788 35860 5840
rect 43444 5831 43496 5840
rect 43444 5797 43453 5831
rect 43453 5797 43487 5831
rect 43487 5797 43496 5831
rect 43444 5788 43496 5797
rect 33968 5720 34020 5772
rect 7380 5584 7432 5636
rect 23204 5584 23256 5636
rect 8484 5516 8536 5568
rect 12808 5516 12860 5568
rect 15292 5516 15344 5568
rect 20536 5516 20588 5568
rect 25412 5516 25464 5568
rect 25872 5516 25924 5568
rect 30380 5516 30432 5568
rect 31116 5584 31168 5636
rect 38660 5652 38712 5704
rect 37832 5584 37884 5636
rect 35348 5559 35400 5568
rect 35348 5525 35357 5559
rect 35357 5525 35391 5559
rect 35391 5525 35400 5559
rect 35348 5516 35400 5525
rect 43076 5559 43128 5568
rect 43076 5525 43085 5559
rect 43085 5525 43119 5559
rect 43119 5525 43128 5559
rect 43076 5516 43128 5525
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 39010 5414 39062 5466
rect 39074 5414 39126 5466
rect 39138 5414 39190 5466
rect 39202 5414 39254 5466
rect 39266 5414 39318 5466
rect 8852 5312 8904 5364
rect 23204 5355 23256 5364
rect 23204 5321 23213 5355
rect 23213 5321 23247 5355
rect 23247 5321 23256 5355
rect 23204 5312 23256 5321
rect 7748 5176 7800 5228
rect 17500 5176 17552 5228
rect 17868 5176 17920 5228
rect 29644 5244 29696 5296
rect 34980 5312 35032 5364
rect 43444 5355 43496 5364
rect 43444 5321 43453 5355
rect 43453 5321 43487 5355
rect 43487 5321 43496 5355
rect 43444 5312 43496 5321
rect 33508 5244 33560 5296
rect 5908 5108 5960 5160
rect 7196 5108 7248 5160
rect 26056 5219 26108 5228
rect 26056 5185 26065 5219
rect 26065 5185 26099 5219
rect 26099 5185 26108 5219
rect 26056 5176 26108 5185
rect 27344 5219 27396 5228
rect 27344 5185 27353 5219
rect 27353 5185 27387 5219
rect 27387 5185 27396 5219
rect 27344 5176 27396 5185
rect 31208 5176 31260 5228
rect 6828 5040 6880 5092
rect 2504 5015 2556 5024
rect 2504 4981 2513 5015
rect 2513 4981 2547 5015
rect 2547 4981 2556 5015
rect 2504 4972 2556 4981
rect 7472 4972 7524 5024
rect 8760 4972 8812 5024
rect 17776 4972 17828 5024
rect 20628 4972 20680 5024
rect 26424 4972 26476 5024
rect 33140 5108 33192 5160
rect 42616 5244 42668 5296
rect 42800 5176 42852 5228
rect 43260 5219 43312 5228
rect 43260 5185 43269 5219
rect 43269 5185 43303 5219
rect 43303 5185 43312 5219
rect 43260 5176 43312 5185
rect 38292 5108 38344 5160
rect 33324 5040 33376 5092
rect 42892 5040 42944 5092
rect 33416 5015 33468 5024
rect 33416 4981 33425 5015
rect 33425 4981 33459 5015
rect 33459 4981 33468 5015
rect 33416 4972 33468 4981
rect 37280 5015 37332 5024
rect 37280 4981 37289 5015
rect 37289 4981 37323 5015
rect 37323 4981 37332 5015
rect 37280 4972 37332 4981
rect 37556 5015 37608 5024
rect 37556 4981 37565 5015
rect 37565 4981 37599 5015
rect 37599 4981 37608 5015
rect 37556 4972 37608 4981
rect 43076 5015 43128 5024
rect 43076 4981 43085 5015
rect 43085 4981 43119 5015
rect 43119 4981 43128 5015
rect 43076 4972 43128 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 37950 4870 38002 4922
rect 38014 4870 38066 4922
rect 38078 4870 38130 4922
rect 38142 4870 38194 4922
rect 38206 4870 38258 4922
rect 2504 4768 2556 4820
rect 13728 4768 13780 4820
rect 23848 4768 23900 4820
rect 26792 4768 26844 4820
rect 30380 4768 30432 4820
rect 36544 4768 36596 4820
rect 5540 4632 5592 4684
rect 29920 4700 29972 4752
rect 33508 4700 33560 4752
rect 41972 4700 42024 4752
rect 43444 4743 43496 4752
rect 43444 4709 43453 4743
rect 43453 4709 43487 4743
rect 43487 4709 43496 4743
rect 43444 4700 43496 4709
rect 11704 4632 11756 4684
rect 6736 4564 6788 4616
rect 8668 4564 8720 4616
rect 13452 4607 13504 4616
rect 13452 4573 13461 4607
rect 13461 4573 13495 4607
rect 13495 4573 13504 4607
rect 13452 4564 13504 4573
rect 17500 4632 17552 4684
rect 21824 4632 21876 4684
rect 24768 4632 24820 4684
rect 28724 4632 28776 4684
rect 21456 4564 21508 4616
rect 35624 4564 35676 4616
rect 42984 4564 43036 4616
rect 5448 4428 5500 4480
rect 10968 4428 11020 4480
rect 13360 4428 13412 4480
rect 17868 4428 17920 4480
rect 25872 4428 25924 4480
rect 26700 4471 26752 4480
rect 26700 4437 26709 4471
rect 26709 4437 26743 4471
rect 26743 4437 26752 4471
rect 26700 4428 26752 4437
rect 42892 4428 42944 4480
rect 43076 4471 43128 4480
rect 43076 4437 43085 4471
rect 43085 4437 43119 4471
rect 43119 4437 43128 4471
rect 43076 4428 43128 4437
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 39010 4326 39062 4378
rect 39074 4326 39126 4378
rect 39138 4326 39190 4378
rect 39202 4326 39254 4378
rect 39266 4326 39318 4378
rect 1308 4224 1360 4276
rect 26608 4224 26660 4276
rect 26700 4224 26752 4276
rect 40040 4224 40092 4276
rect 1216 4156 1268 4208
rect 28356 4156 28408 4208
rect 36544 4156 36596 4208
rect 8392 4088 8444 4140
rect 17408 4131 17460 4140
rect 17408 4097 17417 4131
rect 17417 4097 17451 4131
rect 17451 4097 17460 4131
rect 17408 4088 17460 4097
rect 22100 4088 22152 4140
rect 27804 4088 27856 4140
rect 32864 4088 32916 4140
rect 5632 4020 5684 4072
rect 16120 4020 16172 4072
rect 23756 4020 23808 4072
rect 29552 4020 29604 4072
rect 19708 3952 19760 4004
rect 23848 3952 23900 4004
rect 25688 3952 25740 4004
rect 25780 3952 25832 4004
rect 27620 3952 27672 4004
rect 33600 3952 33652 4004
rect 43444 3995 43496 4004
rect 43444 3961 43453 3995
rect 43453 3961 43487 3995
rect 43487 3961 43496 3995
rect 43444 3952 43496 3961
rect 4252 3927 4304 3936
rect 4252 3893 4261 3927
rect 4261 3893 4295 3927
rect 4295 3893 4304 3927
rect 4252 3884 4304 3893
rect 17132 3884 17184 3936
rect 30656 3884 30708 3936
rect 31852 3884 31904 3936
rect 43076 3927 43128 3936
rect 43076 3893 43085 3927
rect 43085 3893 43119 3927
rect 43119 3893 43128 3927
rect 43076 3884 43128 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 37950 3782 38002 3834
rect 38014 3782 38066 3834
rect 38078 3782 38130 3834
rect 38142 3782 38194 3834
rect 38206 3782 38258 3834
rect 4252 3680 4304 3732
rect 20352 3680 20404 3732
rect 20444 3680 20496 3732
rect 13728 3612 13780 3664
rect 20076 3612 20128 3664
rect 20168 3655 20220 3664
rect 20168 3621 20177 3655
rect 20177 3621 20211 3655
rect 20211 3621 20220 3655
rect 20168 3612 20220 3621
rect 9588 3544 9640 3596
rect 21364 3544 21416 3596
rect 9404 3476 9456 3528
rect 13084 3408 13136 3460
rect 19524 3519 19576 3528
rect 19524 3485 19533 3519
rect 19533 3485 19567 3519
rect 19567 3485 19576 3519
rect 19524 3476 19576 3485
rect 19800 3476 19852 3528
rect 23480 3723 23532 3732
rect 23480 3689 23489 3723
rect 23489 3689 23523 3723
rect 23523 3689 23532 3723
rect 23480 3680 23532 3689
rect 26332 3680 26384 3732
rect 34704 3680 34756 3732
rect 23388 3612 23440 3664
rect 30380 3544 30432 3596
rect 34428 3612 34480 3664
rect 42984 3544 43036 3596
rect 26700 3476 26752 3528
rect 15660 3383 15712 3392
rect 15660 3349 15669 3383
rect 15669 3349 15703 3383
rect 15703 3349 15712 3383
rect 15660 3340 15712 3349
rect 15752 3340 15804 3392
rect 23296 3408 23348 3460
rect 26240 3408 26292 3460
rect 34244 3476 34296 3528
rect 42892 3519 42944 3528
rect 42892 3485 42901 3519
rect 42901 3485 42935 3519
rect 42935 3485 42944 3519
rect 42892 3476 42944 3485
rect 43444 3655 43496 3664
rect 43444 3621 43453 3655
rect 43453 3621 43487 3655
rect 43487 3621 43496 3655
rect 43444 3612 43496 3621
rect 30012 3408 30064 3460
rect 38108 3408 38160 3460
rect 18880 3383 18932 3392
rect 18880 3349 18889 3383
rect 18889 3349 18923 3383
rect 18923 3349 18932 3383
rect 18880 3340 18932 3349
rect 19892 3383 19944 3392
rect 19892 3349 19901 3383
rect 19901 3349 19935 3383
rect 19935 3349 19944 3383
rect 19892 3340 19944 3349
rect 27344 3383 27396 3392
rect 27344 3349 27353 3383
rect 27353 3349 27387 3383
rect 27387 3349 27396 3383
rect 27344 3340 27396 3349
rect 31852 3340 31904 3392
rect 43076 3383 43128 3392
rect 43076 3349 43085 3383
rect 43085 3349 43119 3383
rect 43119 3349 43128 3383
rect 43076 3340 43128 3349
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 39010 3238 39062 3290
rect 39074 3238 39126 3290
rect 39138 3238 39190 3290
rect 39202 3238 39254 3290
rect 39266 3238 39318 3290
rect 5356 3000 5408 3052
rect 6460 3000 6512 3052
rect 10324 3000 10376 3052
rect 15660 3136 15712 3188
rect 24492 3136 24544 3188
rect 25964 3136 26016 3188
rect 31668 3136 31720 3188
rect 33048 3136 33100 3188
rect 34244 3179 34296 3188
rect 34244 3145 34253 3179
rect 34253 3145 34287 3179
rect 34287 3145 34296 3179
rect 34244 3136 34296 3145
rect 34428 3136 34480 3188
rect 38108 3179 38160 3188
rect 38108 3145 38117 3179
rect 38117 3145 38151 3179
rect 38151 3145 38160 3179
rect 38108 3136 38160 3145
rect 43444 3179 43496 3188
rect 43444 3145 43453 3179
rect 43453 3145 43487 3179
rect 43487 3145 43496 3179
rect 43444 3136 43496 3145
rect 14924 3068 14976 3120
rect 9772 2932 9824 2984
rect 15752 3000 15804 3052
rect 18880 3068 18932 3120
rect 25596 3068 25648 3120
rect 8852 2864 8904 2916
rect 20076 3043 20128 3052
rect 20076 3009 20085 3043
rect 20085 3009 20119 3043
rect 20119 3009 20128 3043
rect 20076 3000 20128 3009
rect 20720 3000 20772 3052
rect 21364 3000 21416 3052
rect 7656 2796 7708 2848
rect 14280 2796 14332 2848
rect 22376 2932 22428 2984
rect 16120 2907 16172 2916
rect 16120 2873 16129 2907
rect 16129 2873 16163 2907
rect 16163 2873 16172 2907
rect 16120 2864 16172 2873
rect 25872 3043 25924 3052
rect 25872 3009 25881 3043
rect 25881 3009 25915 3043
rect 25915 3009 25924 3043
rect 25872 3000 25924 3009
rect 27436 3068 27488 3120
rect 27528 3043 27580 3052
rect 27528 3009 27537 3043
rect 27537 3009 27571 3043
rect 27571 3009 27580 3043
rect 27528 3000 27580 3009
rect 27620 3000 27672 3052
rect 26608 2932 26660 2984
rect 30012 3043 30064 3052
rect 30012 3009 30021 3043
rect 30021 3009 30055 3043
rect 30055 3009 30064 3043
rect 30012 3000 30064 3009
rect 25412 2864 25464 2916
rect 30104 2932 30156 2984
rect 31024 3000 31076 3052
rect 33416 3068 33468 3120
rect 42340 3068 42392 3120
rect 32772 3043 32824 3052
rect 32772 3009 32781 3043
rect 32781 3009 32815 3043
rect 32815 3009 32824 3043
rect 32772 3000 32824 3009
rect 30840 2932 30892 2984
rect 31484 2932 31536 2984
rect 31668 2932 31720 2984
rect 33600 3043 33652 3052
rect 33600 3009 33609 3043
rect 33609 3009 33643 3043
rect 33643 3009 33652 3043
rect 33600 3000 33652 3009
rect 34796 3043 34848 3052
rect 34796 3009 34805 3043
rect 34805 3009 34839 3043
rect 34839 3009 34848 3043
rect 34796 3000 34848 3009
rect 33692 2932 33744 2984
rect 35716 3043 35768 3052
rect 35716 3009 35725 3043
rect 35725 3009 35759 3043
rect 35759 3009 35768 3043
rect 35716 3000 35768 3009
rect 37004 3043 37056 3052
rect 37004 3009 37013 3043
rect 37013 3009 37047 3043
rect 37047 3009 37056 3043
rect 37004 3000 37056 3009
rect 37096 3000 37148 3052
rect 40040 3000 40092 3052
rect 43168 3000 43220 3052
rect 28724 2864 28776 2916
rect 29000 2864 29052 2916
rect 33600 2864 33652 2916
rect 33876 2864 33928 2916
rect 19800 2796 19852 2848
rect 20904 2796 20956 2848
rect 21916 2796 21968 2848
rect 25228 2796 25280 2848
rect 25780 2796 25832 2848
rect 26332 2796 26384 2848
rect 27528 2796 27580 2848
rect 28264 2796 28316 2848
rect 28632 2796 28684 2848
rect 29644 2796 29696 2848
rect 30748 2796 30800 2848
rect 31024 2796 31076 2848
rect 31484 2796 31536 2848
rect 32772 2796 32824 2848
rect 32956 2839 33008 2848
rect 32956 2805 32965 2839
rect 32965 2805 32999 2839
rect 32999 2805 33008 2839
rect 32956 2796 33008 2805
rect 33416 2839 33468 2848
rect 33416 2805 33425 2839
rect 33425 2805 33459 2839
rect 33459 2805 33468 2839
rect 33416 2796 33468 2805
rect 33508 2796 33560 2848
rect 33968 2796 34020 2848
rect 34336 2796 34388 2848
rect 34980 2839 35032 2848
rect 34980 2805 34989 2839
rect 34989 2805 35023 2839
rect 35023 2805 35032 2839
rect 34980 2796 35032 2805
rect 42984 2796 43036 2848
rect 43076 2839 43128 2848
rect 43076 2805 43085 2839
rect 43085 2805 43119 2839
rect 43119 2805 43128 2839
rect 43076 2796 43128 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 37950 2694 38002 2746
rect 38014 2694 38066 2746
rect 38078 2694 38130 2746
rect 38142 2694 38194 2746
rect 38206 2694 38258 2746
rect 10968 2592 11020 2644
rect 7656 2456 7708 2508
rect 7472 2388 7524 2440
rect 12992 2388 13044 2440
rect 19708 2388 19760 2440
rect 20720 2524 20772 2576
rect 21456 2524 21508 2576
rect 20352 2388 20404 2440
rect 21732 2456 21784 2508
rect 21548 2388 21600 2440
rect 24124 2524 24176 2576
rect 25044 2592 25096 2644
rect 27344 2592 27396 2644
rect 30196 2592 30248 2644
rect 32404 2592 32456 2644
rect 25504 2524 25556 2576
rect 26608 2524 26660 2576
rect 27712 2524 27764 2576
rect 28816 2524 28868 2576
rect 29920 2524 29972 2576
rect 31300 2524 31352 2576
rect 22376 2456 22428 2508
rect 22560 2431 22612 2440
rect 22560 2397 22569 2431
rect 22569 2397 22603 2431
rect 22603 2397 22612 2431
rect 22560 2388 22612 2397
rect 22928 2431 22980 2440
rect 22928 2397 22937 2431
rect 22937 2397 22971 2431
rect 22971 2397 22980 2431
rect 22928 2388 22980 2397
rect 23296 2431 23348 2440
rect 23296 2397 23305 2431
rect 23305 2397 23339 2431
rect 23339 2397 23348 2431
rect 23296 2388 23348 2397
rect 23388 2388 23440 2440
rect 24768 2431 24820 2440
rect 24768 2397 24777 2431
rect 24777 2397 24811 2431
rect 24811 2397 24820 2431
rect 24768 2388 24820 2397
rect 21456 2320 21508 2372
rect 23204 2320 23256 2372
rect 23756 2320 23808 2372
rect 25320 2388 25372 2440
rect 25596 2456 25648 2508
rect 25688 2388 25740 2440
rect 25964 2388 26016 2440
rect 27252 2431 27304 2440
rect 27252 2397 27261 2431
rect 27261 2397 27295 2431
rect 27295 2397 27304 2431
rect 27252 2388 27304 2397
rect 27528 2388 27580 2440
rect 27620 2388 27672 2440
rect 30012 2456 30064 2508
rect 32956 2456 33008 2508
rect 28448 2431 28500 2440
rect 28448 2397 28457 2431
rect 28457 2397 28491 2431
rect 28491 2397 28500 2431
rect 28448 2388 28500 2397
rect 28632 2388 28684 2440
rect 29552 2431 29604 2440
rect 29552 2397 29561 2431
rect 29561 2397 29595 2431
rect 29595 2397 29604 2431
rect 29552 2388 29604 2397
rect 29736 2388 29788 2440
rect 30288 2431 30340 2440
rect 30288 2397 30297 2431
rect 30297 2397 30331 2431
rect 30331 2397 30340 2431
rect 30288 2388 30340 2397
rect 30932 2431 30984 2440
rect 30932 2397 30941 2431
rect 30941 2397 30975 2431
rect 30975 2397 30984 2431
rect 30932 2388 30984 2397
rect 31484 2431 31536 2440
rect 31484 2397 31493 2431
rect 31493 2397 31527 2431
rect 31527 2397 31536 2431
rect 31484 2388 31536 2397
rect 32312 2388 32364 2440
rect 32680 2388 32732 2440
rect 32772 2431 32824 2440
rect 32772 2397 32781 2431
rect 32781 2397 32815 2431
rect 32815 2397 32824 2431
rect 32772 2388 32824 2397
rect 33324 2456 33376 2508
rect 24952 2320 25004 2372
rect 19708 2295 19760 2304
rect 19708 2261 19717 2295
rect 19717 2261 19751 2295
rect 19751 2261 19760 2295
rect 19708 2252 19760 2261
rect 20260 2252 20312 2304
rect 20536 2252 20588 2304
rect 20812 2295 20864 2304
rect 20812 2261 20821 2295
rect 20821 2261 20855 2295
rect 20855 2261 20864 2295
rect 20812 2252 20864 2261
rect 21364 2252 21416 2304
rect 21640 2252 21692 2304
rect 22192 2252 22244 2304
rect 22468 2252 22520 2304
rect 22744 2295 22796 2304
rect 22744 2261 22753 2295
rect 22753 2261 22787 2295
rect 22787 2261 22796 2295
rect 22744 2252 22796 2261
rect 23020 2252 23072 2304
rect 23296 2252 23348 2304
rect 23572 2252 23624 2304
rect 23940 2252 23992 2304
rect 24676 2252 24728 2304
rect 26884 2320 26936 2372
rect 26148 2252 26200 2304
rect 27988 2320 28040 2372
rect 29368 2320 29420 2372
rect 29092 2252 29144 2304
rect 30564 2320 30616 2372
rect 31024 2252 31076 2304
rect 31576 2320 31628 2372
rect 33600 2431 33652 2440
rect 33600 2397 33609 2431
rect 33609 2397 33643 2431
rect 33643 2397 33652 2431
rect 33600 2388 33652 2397
rect 33784 2388 33836 2440
rect 34704 2431 34756 2440
rect 34704 2397 34713 2431
rect 34713 2397 34747 2431
rect 34747 2397 34756 2431
rect 34704 2388 34756 2397
rect 35072 2431 35124 2440
rect 35072 2397 35081 2431
rect 35081 2397 35115 2431
rect 35115 2397 35124 2431
rect 35072 2388 35124 2397
rect 41972 2431 42024 2440
rect 41972 2397 41981 2431
rect 41981 2397 42015 2431
rect 42015 2397 42024 2431
rect 41972 2388 42024 2397
rect 42524 2431 42576 2440
rect 42524 2397 42533 2431
rect 42533 2397 42567 2431
rect 42567 2397 42576 2431
rect 42524 2388 42576 2397
rect 43444 2567 43496 2576
rect 43444 2533 43453 2567
rect 43453 2533 43487 2567
rect 43487 2533 43496 2567
rect 43444 2524 43496 2533
rect 33876 2320 33928 2372
rect 33140 2252 33192 2304
rect 33600 2252 33652 2304
rect 34244 2252 34296 2304
rect 42156 2295 42208 2304
rect 42156 2261 42165 2295
rect 42165 2261 42199 2295
rect 42199 2261 42208 2295
rect 42156 2252 42208 2261
rect 42708 2295 42760 2304
rect 42708 2261 42717 2295
rect 42717 2261 42751 2295
rect 42751 2261 42760 2295
rect 42708 2252 42760 2261
rect 43076 2295 43128 2304
rect 43076 2261 43085 2295
rect 43085 2261 43119 2295
rect 43119 2261 43128 2295
rect 43076 2252 43128 2261
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 39010 2150 39062 2202
rect 39074 2150 39126 2202
rect 39138 2150 39190 2202
rect 39202 2150 39254 2202
rect 39266 2150 39318 2202
rect 16304 2048 16356 2100
rect 21456 2048 21508 2100
rect 19432 1980 19484 2032
rect 26792 2048 26844 2100
rect 32772 2048 32824 2100
rect 34336 2048 34388 2100
rect 23204 1980 23256 2032
rect 28448 1980 28500 2032
rect 32680 1980 32732 2032
rect 34980 1980 35032 2032
rect 16948 1912 17000 1964
rect 24860 1912 24912 1964
rect 25136 1912 25188 1964
rect 29736 1912 29788 1964
rect 32312 1912 32364 1964
rect 35348 1912 35400 1964
rect 16028 1844 16080 1896
rect 14280 1776 14332 1828
rect 22560 1776 22612 1828
rect 14832 1708 14884 1760
rect 28632 1844 28684 1896
rect 31484 1844 31536 1896
rect 34428 1844 34480 1896
rect 30932 1776 30984 1828
rect 37280 1776 37332 1828
rect 13176 1640 13228 1692
rect 22928 1640 22980 1692
rect 26792 1708 26844 1760
rect 37096 1708 37148 1760
rect 27528 1640 27580 1692
rect 30656 1640 30708 1692
rect 35072 1640 35124 1692
rect 20628 1572 20680 1624
rect 27620 1572 27672 1624
rect 26424 1504 26476 1556
rect 24860 1436 24912 1488
rect 30840 1436 30892 1488
rect 14464 1368 14516 1420
rect 20720 1368 20772 1420
rect 24400 1368 24452 1420
rect 24768 1368 24820 1420
rect 34244 1368 34296 1420
rect 33232 1300 33284 1352
rect 32864 1232 32916 1284
rect 35440 1232 35492 1284
rect 11704 1096 11756 1148
rect 17684 1096 17736 1148
rect 15292 416 15344 468
rect 22100 416 22152 468
rect 16120 348 16172 400
rect 25872 348 25924 400
rect 15568 280 15620 332
rect 27804 280 27856 332
rect 14188 212 14240 264
rect 26700 212 26752 264
rect 17224 144 17276 196
rect 33968 144 34020 196
rect 19248 76 19300 128
rect 37556 76 37608 128
rect 18144 8 18196 60
rect 37004 8 37056 60
<< metal2 >>
rect 1306 11194 1362 11250
rect 3422 11194 3478 11250
rect 5538 11194 5594 11250
rect 7654 11194 7710 11250
rect 9770 11194 9826 11250
rect 11886 11194 11942 11250
rect 14002 11194 14058 11250
rect 16118 11194 16174 11250
rect 18234 11194 18290 11250
rect 20350 11194 20406 11250
rect 22466 11194 22522 11250
rect 24582 11194 24638 11250
rect 26698 11194 26754 11250
rect 28814 11194 28870 11250
rect 30930 11194 30986 11250
rect 33046 11194 33102 11250
rect 35162 11194 35218 11250
rect 37278 11194 37334 11250
rect 39394 11194 39450 11250
rect 41510 11194 41566 11250
rect 43626 11194 43682 11250
rect 1214 9888 1270 9897
rect 1214 9823 1270 9832
rect 1228 8401 1256 9823
rect 1320 8634 1348 11194
rect 2870 8800 2926 8809
rect 2870 8735 2926 8744
rect 1308 8628 1360 8634
rect 1308 8570 1360 8576
rect 2884 8401 2912 8735
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 3436 8634 3464 11194
rect 5552 8634 5580 11194
rect 7668 8634 7696 11194
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 9784 8634 9812 11194
rect 11900 8634 11928 11194
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12268 8634 12296 8774
rect 14016 8634 14044 11194
rect 14922 9344 14978 9353
rect 14922 9279 14978 9288
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 5448 8424 5500 8430
rect 1214 8392 1270 8401
rect 1214 8327 1270 8336
rect 2870 8392 2926 8401
rect 5448 8366 5500 8372
rect 2870 8327 2926 8336
rect 1766 8256 1822 8265
rect 1766 8191 1822 8200
rect 1780 7449 1808 8191
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 1306 7440 1362 7449
rect 1306 7375 1362 7384
rect 1766 7440 1822 7449
rect 1766 7375 1822 7384
rect 1320 6186 1348 7375
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 3988 7002 4016 7686
rect 4356 7546 4384 7686
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 1308 6180 1360 6186
rect 1308 6122 1360 6128
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 940 5840 992 5846
rect 940 5782 992 5788
rect 952 1465 980 5782
rect 2870 5536 2926 5545
rect 2870 5471 2926 5480
rect 2884 5137 2912 5471
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 2870 5128 2926 5137
rect 2870 5063 2926 5072
rect 2504 5024 2556 5030
rect 1766 4992 1822 5001
rect 2504 4966 2556 4972
rect 1766 4927 1822 4936
rect 1306 4448 1362 4457
rect 1306 4383 1362 4392
rect 1320 4282 1348 4383
rect 1308 4276 1360 4282
rect 1308 4218 1360 4224
rect 1216 4208 1268 4214
rect 1214 4176 1216 4185
rect 1780 4185 1808 4927
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2516 4826 2544 4966
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 5460 4486 5488 8366
rect 5828 6458 5856 8434
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 1268 4176 1270 4185
rect 1214 4111 1270 4120
rect 1766 4176 1822 4185
rect 1766 4111 1822 4120
rect 2870 4040 2926 4049
rect 2870 3975 2926 3984
rect 1766 3904 1822 3913
rect 1766 3839 1822 3848
rect 1780 3505 1808 3839
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1766 3496 1822 3505
rect 1766 3431 1822 3440
rect 2884 3369 2912 3975
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4264 3738 4292 3878
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 2870 3360 2926 3369
rect 2870 3295 2926 3304
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 938 1456 994 1465
rect 938 1391 994 1400
rect 5368 56 5396 2994
rect 5552 2009 5580 4626
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5538 2000 5594 2009
rect 5538 1935 5594 1944
rect 5644 56 5672 4014
rect 5920 56 5948 5102
rect 6196 56 6224 6734
rect 6840 5098 6868 8434
rect 7746 8256 7802 8265
rect 7746 8191 7802 8200
rect 7760 7857 7788 8191
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 14936 8090 14964 9279
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 16132 8634 16160 11194
rect 16488 9104 16540 9110
rect 16488 9046 16540 9052
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16500 8498 16528 9046
rect 18248 8634 18276 11194
rect 19338 9616 19394 9625
rect 19338 9551 19394 9560
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18616 8498 18644 8978
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 7840 7880 7892 7886
rect 7746 7848 7802 7857
rect 7564 7812 7616 7818
rect 7840 7822 7892 7828
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 7746 7783 7802 7792
rect 7564 7754 7616 7760
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6472 56 6500 2994
rect 6748 56 6776 4558
rect 7024 56 7052 5646
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 7208 1737 7236 5102
rect 7194 1728 7250 1737
rect 7194 1663 7250 1672
rect 7300 56 7328 6258
rect 7380 5636 7432 5642
rect 7380 5578 7432 5584
rect 7392 2553 7420 5578
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7378 2544 7434 2553
rect 7378 2479 7434 2488
rect 7484 2446 7512 4966
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7576 56 7604 7754
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7656 2848 7708 2854
rect 7656 2790 7708 2796
rect 7668 2514 7696 2790
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 7760 82 7788 5170
rect 7852 218 7880 7822
rect 8852 7744 8904 7750
rect 8850 7712 8852 7721
rect 9404 7744 9456 7750
rect 8904 7712 8906 7721
rect 9404 7686 9456 7692
rect 8850 7647 8906 7656
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 9416 7585 9444 7686
rect 9402 7576 9458 7585
rect 9402 7511 9458 7520
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 9600 6662 9628 6870
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 8758 6352 8814 6361
rect 8758 6287 8814 6296
rect 9404 6316 9456 6322
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 8482 5672 8538 5681
rect 8482 5607 8538 5616
rect 8496 5574 8524 5607
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8772 5030 8800 6287
rect 9404 6258 9456 6264
rect 9416 6225 9444 6258
rect 9402 6216 9458 6225
rect 9402 6151 9458 6160
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 8850 5808 8906 5817
rect 8850 5743 8906 5752
rect 8864 5370 8892 5743
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 7852 190 7972 218
rect 7760 56 7880 82
rect 5354 0 5410 56
rect 5630 0 5686 56
rect 5906 0 5962 56
rect 6182 0 6238 56
rect 6458 0 6514 56
rect 6734 0 6790 56
rect 7010 0 7066 56
rect 7286 0 7342 56
rect 7562 0 7618 56
rect 7760 54 7894 56
rect 7838 0 7894 54
rect 7944 42 7972 190
rect 8036 56 8156 82
rect 8404 56 8432 4082
rect 8680 56 8708 4558
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 8852 2916 8904 2922
rect 8852 2858 8904 2864
rect 8864 1578 8892 2858
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 8864 1550 8984 1578
rect 8956 56 8984 1550
rect 9232 56 9352 82
rect 8036 54 8170 56
rect 8036 42 8064 54
rect 7944 14 8064 42
rect 8114 0 8170 54
rect 8390 0 8446 56
rect 8666 0 8722 56
rect 8942 0 8998 56
rect 9218 54 9352 56
rect 9218 0 9274 54
rect 9324 42 9352 54
rect 9416 42 9444 3470
rect 9508 56 9536 5646
rect 9600 3602 9628 6054
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9784 56 9812 2926
rect 10060 56 10088 6734
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 10244 6390 10272 6666
rect 10232 6384 10284 6390
rect 10232 6326 10284 6332
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10336 56 10364 2994
rect 10612 56 10640 6734
rect 10888 56 10916 7822
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 14830 7576 14886 7585
rect 15010 7579 15318 7588
rect 14830 7511 14886 7520
rect 14844 7313 14872 7511
rect 12346 7304 12402 7313
rect 11152 7268 11204 7274
rect 12346 7239 12402 7248
rect 13266 7304 13322 7313
rect 13266 7239 13322 7248
rect 14830 7304 14886 7313
rect 14830 7239 14886 7248
rect 11152 7210 11204 7216
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 10980 2650 11008 4422
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 11072 2553 11100 6054
rect 11058 2544 11114 2553
rect 11058 2479 11114 2488
rect 11164 56 11192 7210
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11624 2961 11652 5850
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11610 2952 11666 2961
rect 11610 2887 11666 2896
rect 11716 2417 11744 4626
rect 11702 2408 11758 2417
rect 11702 2343 11758 2352
rect 11426 2000 11482 2009
rect 11426 1935 11482 1944
rect 11440 56 11468 1935
rect 11704 1148 11756 1154
rect 11704 1090 11756 1096
rect 11716 56 11744 1090
rect 11992 56 12020 5714
rect 12268 56 12296 6666
rect 12360 6458 12388 7239
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12544 56 12572 6802
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12820 56 12848 5510
rect 12912 2417 12940 6598
rect 12992 6384 13044 6390
rect 12992 6326 13044 6332
rect 13004 2446 13032 6326
rect 13084 3460 13136 3466
rect 13084 3402 13136 3408
rect 12992 2440 13044 2446
rect 12898 2408 12954 2417
rect 12992 2382 13044 2388
rect 12898 2343 12954 2352
rect 13096 56 13124 3402
rect 13188 1698 13216 6598
rect 13280 3097 13308 7239
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13740 7002 13768 7142
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13450 4720 13506 4729
rect 13450 4655 13506 4664
rect 13464 4622 13492 4655
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13266 3088 13322 3097
rect 13266 3023 13322 3032
rect 13176 1692 13228 1698
rect 13176 1634 13228 1640
rect 13372 56 13400 4422
rect 13648 56 13676 6258
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13740 3670 13768 4762
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13832 456 13860 6938
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 14280 2848 14332 2854
rect 14280 2790 14332 2796
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 14292 1834 14320 2790
rect 14280 1828 14332 1834
rect 14280 1770 14332 1776
rect 14464 1420 14516 1426
rect 14464 1362 14516 1368
rect 13832 428 13952 456
rect 13924 56 13952 428
rect 14188 264 14240 270
rect 14188 206 14240 212
rect 14200 56 14228 206
rect 14476 56 14504 1362
rect 14752 56 14780 6190
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 14844 1766 14872 6054
rect 14936 5914 14964 6598
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 15028 5658 15056 6054
rect 15212 5914 15240 6326
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 14936 5630 15056 5658
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 14936 3641 14964 5630
rect 15304 5574 15332 5646
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 14922 3632 14978 3641
rect 14922 3567 14978 3576
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 15010 3227 15318 3236
rect 15672 3194 15700 3334
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 14832 1760 14884 1766
rect 14832 1702 14884 1708
rect 14936 1442 14964 3062
rect 15764 3058 15792 3334
rect 15842 3224 15898 3233
rect 15842 3159 15898 3168
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 14936 1414 15056 1442
rect 15028 56 15056 1414
rect 15292 468 15344 474
rect 15292 410 15344 416
rect 15304 56 15332 410
rect 15568 332 15620 338
rect 15568 274 15620 280
rect 15580 56 15608 274
rect 15856 56 15884 3159
rect 16040 1902 16068 6598
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 16132 2922 16160 4014
rect 16120 2916 16172 2922
rect 16120 2858 16172 2864
rect 16316 2106 16344 6598
rect 16500 3505 16528 6802
rect 16946 5944 17002 5953
rect 16946 5879 17002 5888
rect 16960 5681 16988 5879
rect 16946 5672 17002 5681
rect 16946 5607 17002 5616
rect 17144 3942 17172 8366
rect 19352 7886 19380 9551
rect 20364 8634 20392 11194
rect 20902 9072 20958 9081
rect 20902 9007 20958 9016
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20732 8498 20760 8774
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20718 8392 20774 8401
rect 20444 8356 20496 8362
rect 20718 8327 20774 8336
rect 20444 8298 20496 8304
rect 19950 8188 20258 8197
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 18052 7472 18104 7478
rect 18052 7414 18104 7420
rect 18064 6458 18092 7414
rect 18788 7336 18840 7342
rect 18786 7304 18788 7313
rect 18840 7304 18842 7313
rect 18786 7239 18842 7248
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 17222 6352 17278 6361
rect 17222 6287 17278 6296
rect 17774 6352 17830 6361
rect 17774 6287 17830 6296
rect 17236 5681 17264 6287
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 17222 5672 17278 5681
rect 17222 5607 17278 5616
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 17512 4690 17540 5170
rect 17500 4684 17552 4690
rect 17500 4626 17552 4632
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 16486 3496 16542 3505
rect 16486 3431 16542 3440
rect 16670 2952 16726 2961
rect 16670 2887 16726 2896
rect 16304 2100 16356 2106
rect 16304 2042 16356 2048
rect 16028 1896 16080 1902
rect 16028 1838 16080 1844
rect 16394 504 16450 513
rect 16394 439 16450 448
rect 16120 400 16172 406
rect 16120 342 16172 348
rect 16132 56 16160 342
rect 16408 56 16436 439
rect 16684 56 16712 2887
rect 16948 1964 17000 1970
rect 16948 1906 17000 1912
rect 16960 56 16988 1906
rect 17224 196 17276 202
rect 17224 138 17276 144
rect 17236 56 17264 138
rect 17420 105 17448 4082
rect 17696 1154 17724 6190
rect 17788 5030 17816 6287
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17880 4486 17908 5170
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17866 3088 17922 3097
rect 17866 3023 17922 3032
rect 17880 1442 17908 3023
rect 18708 2009 18736 6734
rect 18788 6180 18840 6186
rect 18788 6122 18840 6128
rect 18800 5846 18828 6122
rect 18788 5840 18840 5846
rect 18788 5782 18840 5788
rect 19076 5409 19104 7686
rect 20364 7410 20392 7822
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 19062 5400 19118 5409
rect 19062 5335 19118 5344
rect 19522 5264 19578 5273
rect 19522 5199 19578 5208
rect 19536 3534 19564 5199
rect 19798 5128 19854 5137
rect 19798 5063 19854 5072
rect 19708 4004 19760 4010
rect 19708 3946 19760 3952
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 18880 3392 18932 3398
rect 18880 3334 18932 3340
rect 18892 3126 18920 3334
rect 18880 3120 18932 3126
rect 18880 3062 18932 3068
rect 19720 2446 19748 3946
rect 19812 3534 19840 5063
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 19950 3836 20258 3845
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 20456 3738 20484 8298
rect 20732 8022 20760 8327
rect 20720 8016 20772 8022
rect 20720 7958 20772 7964
rect 20916 7970 20944 9007
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 22480 8634 22508 11194
rect 22928 8968 22980 8974
rect 22756 8916 22928 8922
rect 22756 8910 22980 8916
rect 22756 8894 22968 8910
rect 22756 8838 22784 8894
rect 22744 8832 22796 8838
rect 22744 8774 22796 8780
rect 22836 8832 22888 8838
rect 22836 8774 22888 8780
rect 22468 8628 22520 8634
rect 22468 8570 22520 8576
rect 22848 8498 22876 8774
rect 24596 8634 24624 11194
rect 25872 9172 25924 9178
rect 25872 9114 25924 9120
rect 25504 9104 25556 9110
rect 25504 9046 25556 9052
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 24584 8628 24636 8634
rect 24584 8570 24636 8576
rect 23756 8560 23808 8566
rect 23756 8502 23808 8508
rect 22836 8492 22888 8498
rect 22836 8434 22888 8440
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 23204 8288 23256 8294
rect 23204 8230 23256 8236
rect 21376 8090 21404 8230
rect 21272 8084 21324 8090
rect 21272 8026 21324 8032
rect 21364 8084 21416 8090
rect 21364 8026 21416 8032
rect 20916 7942 21036 7970
rect 21008 7886 21036 7942
rect 21284 7886 21312 8026
rect 23216 8022 23244 8230
rect 23400 8090 23428 8298
rect 23768 8090 23796 8502
rect 24872 8090 24900 8978
rect 23388 8084 23440 8090
rect 23388 8026 23440 8032
rect 23756 8084 23808 8090
rect 23756 8026 23808 8032
rect 24860 8084 24912 8090
rect 24860 8026 24912 8032
rect 23112 8016 23164 8022
rect 23112 7958 23164 7964
rect 23204 8016 23256 8022
rect 23204 7958 23256 7964
rect 23662 7984 23718 7993
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21008 7750 21036 7822
rect 20996 7744 21048 7750
rect 20996 7686 21048 7692
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20640 6934 20668 7278
rect 20628 6928 20680 6934
rect 20628 6870 20680 6876
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 20548 5574 20576 6054
rect 20536 5568 20588 5574
rect 20536 5510 20588 5516
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20444 3732 20496 3738
rect 20444 3674 20496 3680
rect 20076 3664 20128 3670
rect 20168 3664 20220 3670
rect 20076 3606 20128 3612
rect 20166 3632 20168 3641
rect 20220 3632 20222 3641
rect 19800 3528 19852 3534
rect 19800 3470 19852 3476
rect 19890 3496 19946 3505
rect 19890 3431 19946 3440
rect 19904 3398 19932 3431
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 20088 3058 20116 3606
rect 20166 3567 20222 3576
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 19708 2440 19760 2446
rect 19708 2382 19760 2388
rect 19708 2304 19760 2310
rect 19708 2246 19760 2252
rect 19432 2032 19484 2038
rect 18694 2000 18750 2009
rect 18694 1935 18750 1944
rect 18878 2000 18934 2009
rect 19432 1974 19484 1980
rect 18878 1935 18934 1944
rect 17788 1414 17908 1442
rect 17684 1148 17736 1154
rect 17684 1090 17736 1096
rect 17498 232 17554 241
rect 17498 167 17554 176
rect 17406 96 17462 105
rect 9324 14 9444 42
rect 9494 0 9550 56
rect 9770 0 9826 56
rect 10046 0 10102 56
rect 10322 0 10378 56
rect 10598 0 10654 56
rect 10874 0 10930 56
rect 11150 0 11206 56
rect 11426 0 11482 56
rect 11702 0 11758 56
rect 11978 0 12034 56
rect 12254 0 12310 56
rect 12530 0 12586 56
rect 12806 0 12862 56
rect 13082 0 13138 56
rect 13358 0 13414 56
rect 13634 0 13690 56
rect 13910 0 13966 56
rect 14186 0 14242 56
rect 14462 0 14518 56
rect 14738 0 14794 56
rect 15014 0 15070 56
rect 15290 0 15346 56
rect 15566 0 15622 56
rect 15842 0 15898 56
rect 16118 0 16174 56
rect 16394 0 16450 56
rect 16670 0 16726 56
rect 16946 0 17002 56
rect 17222 0 17278 56
rect 17512 56 17540 167
rect 17788 56 17816 1414
rect 18326 640 18382 649
rect 18326 575 18382 584
rect 18064 66 18184 82
rect 18064 60 18196 66
rect 18064 56 18144 60
rect 17406 31 17462 40
rect 17498 0 17554 56
rect 17774 0 17830 56
rect 18050 54 18144 56
rect 18050 0 18106 54
rect 18340 56 18368 575
rect 18602 368 18658 377
rect 18602 303 18658 312
rect 18616 56 18644 303
rect 18892 56 18920 1935
rect 19248 128 19300 134
rect 19168 76 19248 82
rect 19168 70 19300 76
rect 19168 56 19288 70
rect 19444 56 19472 1974
rect 19720 56 19748 2246
rect 18144 2 18196 8
rect 18326 0 18382 56
rect 18602 0 18658 56
rect 18878 0 18934 56
rect 19154 54 19288 56
rect 19154 0 19210 54
rect 19430 0 19486 56
rect 19706 0 19762 56
rect 19812 42 19840 2790
rect 19950 2748 20258 2757
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 20364 2446 20392 3674
rect 20442 3224 20498 3233
rect 20442 3159 20498 3168
rect 20456 2825 20484 3159
rect 20442 2816 20498 2825
rect 20442 2751 20498 2760
rect 20352 2440 20404 2446
rect 20352 2382 20404 2388
rect 20260 2304 20312 2310
rect 20260 2246 20312 2252
rect 20536 2304 20588 2310
rect 20536 2246 20588 2252
rect 19904 56 20024 82
rect 20272 56 20300 2246
rect 20548 56 20576 2246
rect 20640 1630 20668 4966
rect 20732 3058 20760 7482
rect 20824 7002 20852 7482
rect 23124 7410 23152 7958
rect 23662 7919 23718 7928
rect 23676 7886 23704 7919
rect 23664 7880 23716 7886
rect 23664 7822 23716 7828
rect 23480 7744 23532 7750
rect 23480 7686 23532 7692
rect 23492 7449 23520 7686
rect 23478 7440 23534 7449
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 23112 7404 23164 7410
rect 23478 7375 23534 7384
rect 25136 7404 25188 7410
rect 23112 7346 23164 7352
rect 25136 7346 25188 7352
rect 21824 7200 21876 7206
rect 21824 7142 21876 7148
rect 20812 6996 20864 7002
rect 20812 6938 20864 6944
rect 20902 6896 20958 6905
rect 20902 6831 20958 6840
rect 20916 6458 20944 6831
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 21456 6316 21508 6322
rect 21456 6258 21508 6264
rect 21468 5914 21496 6258
rect 21456 5908 21508 5914
rect 21456 5850 21508 5856
rect 21640 5840 21692 5846
rect 21454 5808 21510 5817
rect 21638 5808 21640 5817
rect 21692 5808 21694 5817
rect 21510 5766 21588 5794
rect 21454 5743 21510 5752
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 21456 4616 21508 4622
rect 21456 4558 21508 4564
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 21376 3058 21404 3538
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 20904 2848 20956 2854
rect 20904 2790 20956 2796
rect 20720 2576 20772 2582
rect 20720 2518 20772 2524
rect 20628 1624 20680 1630
rect 20628 1566 20680 1572
rect 20732 1426 20760 2518
rect 20812 2304 20864 2310
rect 20812 2246 20864 2252
rect 20720 1420 20772 1426
rect 20720 1362 20772 1368
rect 20824 56 20852 2246
rect 19904 54 20038 56
rect 19904 42 19932 54
rect 19812 14 19932 42
rect 19982 0 20038 54
rect 20258 0 20314 56
rect 20534 0 20590 56
rect 20810 0 20866 56
rect 20916 42 20944 2790
rect 21468 2582 21496 4558
rect 21456 2576 21508 2582
rect 21456 2518 21508 2524
rect 21560 2446 21588 5766
rect 21638 5743 21694 5752
rect 21836 5658 21864 7142
rect 22020 6730 22048 7346
rect 22192 7200 22244 7206
rect 22192 7142 22244 7148
rect 22204 7002 22232 7142
rect 22192 6996 22244 7002
rect 22192 6938 22244 6944
rect 24950 6760 25006 6769
rect 22008 6724 22060 6730
rect 24950 6695 24952 6704
rect 22008 6666 22060 6672
rect 25004 6695 25006 6704
rect 24952 6666 25004 6672
rect 24676 6384 24728 6390
rect 24676 6326 24728 6332
rect 21744 5630 21864 5658
rect 23204 5636 23256 5642
rect 21638 3088 21694 3097
rect 21638 3023 21694 3032
rect 21652 2825 21680 3023
rect 21638 2816 21694 2825
rect 21638 2751 21694 2760
rect 21744 2514 21772 5630
rect 23204 5578 23256 5584
rect 23216 5370 23244 5578
rect 23204 5364 23256 5370
rect 23204 5306 23256 5312
rect 23848 4820 23900 4826
rect 23848 4762 23900 4768
rect 21824 4684 21876 4690
rect 21824 4626 21876 4632
rect 21732 2508 21784 2514
rect 21732 2450 21784 2456
rect 21548 2440 21600 2446
rect 21548 2382 21600 2388
rect 21456 2372 21508 2378
rect 21456 2314 21508 2320
rect 21364 2304 21416 2310
rect 21364 2246 21416 2252
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 21008 56 21128 82
rect 21376 56 21404 2246
rect 21468 2106 21496 2314
rect 21640 2304 21692 2310
rect 21640 2246 21692 2252
rect 21456 2100 21508 2106
rect 21456 2042 21508 2048
rect 21652 56 21680 2246
rect 21836 1737 21864 4626
rect 23386 4584 23442 4593
rect 23386 4519 23442 4528
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 21822 1728 21878 1737
rect 21822 1663 21878 1672
rect 21928 56 21956 2790
rect 22112 474 22140 4082
rect 23400 3670 23428 4519
rect 23478 4176 23534 4185
rect 23478 4111 23534 4120
rect 23492 3738 23520 4111
rect 23756 4072 23808 4078
rect 23756 4014 23808 4020
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23388 3664 23440 3670
rect 23388 3606 23440 3612
rect 23296 3460 23348 3466
rect 23296 3402 23348 3408
rect 22376 2984 22428 2990
rect 22376 2926 22428 2932
rect 22388 2514 22416 2926
rect 22376 2508 22428 2514
rect 22376 2450 22428 2456
rect 23308 2446 23336 3402
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 22928 2440 22980 2446
rect 22928 2382 22980 2388
rect 23296 2440 23348 2446
rect 23388 2440 23440 2446
rect 23296 2382 23348 2388
rect 23386 2408 23388 2417
rect 23440 2408 23442 2417
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 22468 2304 22520 2310
rect 22468 2246 22520 2252
rect 22100 468 22152 474
rect 22100 410 22152 416
rect 22204 56 22232 2246
rect 22480 56 22508 2246
rect 22572 1834 22600 2382
rect 22744 2304 22796 2310
rect 22744 2246 22796 2252
rect 22560 1828 22612 1834
rect 22560 1770 22612 1776
rect 22756 56 22784 2246
rect 22940 1698 22968 2382
rect 23204 2372 23256 2378
rect 23768 2378 23796 4014
rect 23860 4010 23888 4762
rect 23848 4004 23900 4010
rect 23848 3946 23900 3952
rect 24492 3188 24544 3194
rect 24492 3130 24544 3136
rect 24504 2689 24532 3130
rect 24688 2774 24716 6326
rect 24768 4684 24820 4690
rect 24768 4626 24820 4632
rect 24780 4049 24808 4626
rect 24766 4040 24822 4049
rect 24766 3975 24822 3984
rect 24688 2746 24808 2774
rect 24490 2680 24546 2689
rect 24490 2615 24546 2624
rect 24124 2576 24176 2582
rect 24124 2518 24176 2524
rect 23386 2343 23442 2352
rect 23756 2372 23808 2378
rect 23204 2314 23256 2320
rect 23756 2314 23808 2320
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 22928 1692 22980 1698
rect 22928 1634 22980 1640
rect 23032 56 23060 2246
rect 23216 2038 23244 2314
rect 23296 2304 23348 2310
rect 23296 2246 23348 2252
rect 23572 2304 23624 2310
rect 23940 2304 23992 2310
rect 23572 2246 23624 2252
rect 23860 2264 23940 2292
rect 23204 2032 23256 2038
rect 23204 1974 23256 1980
rect 23308 56 23336 2246
rect 23584 56 23612 2246
rect 23860 56 23888 2264
rect 23940 2246 23992 2252
rect 24136 56 24164 2518
rect 24780 2446 24808 2746
rect 25044 2644 25096 2650
rect 25044 2586 25096 2592
rect 25056 2496 25084 2586
rect 24872 2468 25084 2496
rect 24768 2440 24820 2446
rect 24768 2382 24820 2388
rect 24676 2304 24728 2310
rect 24872 2292 24900 2468
rect 24952 2372 25004 2378
rect 24952 2314 25004 2320
rect 24676 2246 24728 2252
rect 24780 2264 24900 2292
rect 24400 1420 24452 1426
rect 24400 1362 24452 1368
rect 24412 56 24440 1362
rect 24688 56 24716 2246
rect 24780 1426 24808 2264
rect 24860 1964 24912 1970
rect 24860 1906 24912 1912
rect 24872 1494 24900 1906
rect 24860 1488 24912 1494
rect 24860 1430 24912 1436
rect 24768 1420 24820 1426
rect 24768 1362 24820 1368
rect 24964 56 24992 2314
rect 25148 1970 25176 7346
rect 25228 6928 25280 6934
rect 25412 6928 25464 6934
rect 25280 6876 25412 6882
rect 25228 6870 25464 6876
rect 25240 6854 25452 6870
rect 25516 6458 25544 9046
rect 25504 6452 25556 6458
rect 25504 6394 25556 6400
rect 25412 6112 25464 6118
rect 25412 6054 25464 6060
rect 25424 5914 25452 6054
rect 25412 5908 25464 5914
rect 25412 5850 25464 5856
rect 25780 5704 25832 5710
rect 25780 5646 25832 5652
rect 25412 5568 25464 5574
rect 25412 5510 25464 5516
rect 25424 2922 25452 5510
rect 25792 4010 25820 5646
rect 25884 5574 25912 9114
rect 26148 8968 26200 8974
rect 26148 8910 26200 8916
rect 26160 8294 26188 8910
rect 26712 8634 26740 11194
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 28828 8634 28856 11194
rect 30944 8634 30972 11194
rect 31852 8900 31904 8906
rect 31852 8842 31904 8848
rect 31024 8832 31076 8838
rect 31024 8774 31076 8780
rect 26700 8628 26752 8634
rect 26700 8570 26752 8576
rect 27160 8628 27212 8634
rect 27160 8570 27212 8576
rect 28724 8628 28776 8634
rect 28724 8570 28776 8576
rect 28816 8628 28868 8634
rect 28816 8570 28868 8576
rect 30932 8628 30984 8634
rect 30932 8570 30984 8576
rect 26330 8528 26386 8537
rect 27172 8498 27200 8570
rect 26330 8463 26386 8472
rect 27160 8492 27212 8498
rect 26148 8288 26200 8294
rect 26148 8230 26200 8236
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 26344 8090 26372 8463
rect 27160 8434 27212 8440
rect 26792 8424 26844 8430
rect 26792 8366 26844 8372
rect 26332 8084 26384 8090
rect 26332 8026 26384 8032
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 26056 5840 26108 5846
rect 26056 5782 26108 5788
rect 25872 5568 25924 5574
rect 25872 5510 25924 5516
rect 26068 5234 26096 5782
rect 26056 5228 26108 5234
rect 26056 5170 26108 5176
rect 26424 5024 26476 5030
rect 26424 4966 26476 4972
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 25872 4480 25924 4486
rect 25872 4422 25924 4428
rect 25688 4004 25740 4010
rect 25688 3946 25740 3952
rect 25780 4004 25832 4010
rect 25780 3946 25832 3952
rect 25596 3120 25648 3126
rect 25596 3062 25648 3068
rect 25412 2916 25464 2922
rect 25412 2858 25464 2864
rect 25228 2848 25280 2854
rect 25228 2790 25280 2796
rect 25136 1964 25188 1970
rect 25136 1906 25188 1912
rect 25240 56 25268 2790
rect 25318 2680 25374 2689
rect 25318 2615 25374 2624
rect 25332 2446 25360 2615
rect 25504 2576 25556 2582
rect 25504 2518 25556 2524
rect 25320 2440 25372 2446
rect 25320 2382 25372 2388
rect 25516 56 25544 2518
rect 25608 2514 25636 3062
rect 25596 2508 25648 2514
rect 25596 2450 25648 2456
rect 25700 2446 25728 3946
rect 25884 3058 25912 4422
rect 26330 4040 26386 4049
rect 26330 3975 26386 3984
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 26344 3738 26372 3975
rect 26332 3732 26384 3738
rect 26332 3674 26384 3680
rect 26240 3460 26292 3466
rect 26240 3402 26292 3408
rect 25964 3188 26016 3194
rect 25964 3130 26016 3136
rect 25872 3052 25924 3058
rect 25872 2994 25924 3000
rect 25780 2848 25832 2854
rect 25976 2836 26004 3130
rect 26252 3097 26280 3402
rect 26238 3088 26294 3097
rect 26238 3023 26294 3032
rect 25780 2790 25832 2796
rect 25884 2808 26004 2836
rect 26332 2848 26384 2854
rect 25688 2440 25740 2446
rect 25688 2382 25740 2388
rect 25792 56 25820 2790
rect 25884 406 25912 2808
rect 26332 2790 26384 2796
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 25962 2544 26018 2553
rect 25962 2479 26018 2488
rect 25976 2446 26004 2479
rect 25964 2440 26016 2446
rect 25964 2382 26016 2388
rect 26148 2304 26200 2310
rect 26068 2264 26148 2292
rect 25872 400 25924 406
rect 25872 342 25924 348
rect 26068 56 26096 2264
rect 26148 2246 26200 2252
rect 26344 56 26372 2790
rect 26436 1562 26464 4966
rect 26804 4826 26832 8366
rect 28172 8288 28224 8294
rect 28172 8230 28224 8236
rect 27528 7880 27580 7886
rect 27264 7806 27384 7834
rect 27528 7822 27580 7828
rect 27264 7750 27292 7806
rect 26884 7744 26936 7750
rect 26884 7686 26936 7692
rect 27252 7744 27304 7750
rect 27252 7686 27304 7692
rect 26896 7313 26924 7686
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 27356 7478 27384 7806
rect 27436 7744 27488 7750
rect 27436 7686 27488 7692
rect 27344 7472 27396 7478
rect 27344 7414 27396 7420
rect 26882 7304 26938 7313
rect 26882 7239 26938 7248
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 27342 5672 27398 5681
rect 27342 5607 27398 5616
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 27356 5234 27384 5607
rect 27344 5228 27396 5234
rect 27344 5170 27396 5176
rect 26792 4820 26844 4826
rect 26792 4762 26844 4768
rect 26700 4480 26752 4486
rect 26700 4422 26752 4428
rect 26712 4282 26740 4422
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 26608 4276 26660 4282
rect 26608 4218 26660 4224
rect 26700 4276 26752 4282
rect 26700 4218 26752 4224
rect 26620 2990 26648 4218
rect 26700 3528 26752 3534
rect 26700 3470 26752 3476
rect 26608 2984 26660 2990
rect 26608 2926 26660 2932
rect 26608 2576 26660 2582
rect 26608 2518 26660 2524
rect 26424 1556 26476 1562
rect 26424 1498 26476 1504
rect 26620 56 26648 2518
rect 26712 270 26740 3470
rect 27344 3392 27396 3398
rect 27344 3334 27396 3340
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 27356 2774 27384 3334
rect 27448 3126 27476 7686
rect 27540 7546 27568 7822
rect 28184 7750 28212 8230
rect 28356 7880 28408 7886
rect 28356 7822 28408 7828
rect 28172 7744 28224 7750
rect 28172 7686 28224 7692
rect 27528 7540 27580 7546
rect 27528 7482 27580 7488
rect 28368 7342 28396 7822
rect 28356 7336 28408 7342
rect 28356 7278 28408 7284
rect 27528 6452 27580 6458
rect 27528 6394 27580 6400
rect 27436 3120 27488 3126
rect 27436 3062 27488 3068
rect 27540 3058 27568 6394
rect 28736 6118 28764 8570
rect 29368 8560 29420 8566
rect 29368 8502 29420 8508
rect 29184 8492 29236 8498
rect 29184 8434 29236 8440
rect 29092 8424 29144 8430
rect 29092 8366 29144 8372
rect 28724 6112 28776 6118
rect 28724 6054 28776 6060
rect 29104 5710 29132 8366
rect 29196 6458 29224 8434
rect 29380 8090 29408 8502
rect 29368 8084 29420 8090
rect 29368 8026 29420 8032
rect 29552 7880 29604 7886
rect 29550 7848 29552 7857
rect 29604 7848 29606 7857
rect 29550 7783 29606 7792
rect 29736 7744 29788 7750
rect 29736 7686 29788 7692
rect 29748 7546 29776 7686
rect 29736 7540 29788 7546
rect 29736 7482 29788 7488
rect 29460 7472 29512 7478
rect 29460 7414 29512 7420
rect 29368 6724 29420 6730
rect 29368 6666 29420 6672
rect 29184 6452 29236 6458
rect 29184 6394 29236 6400
rect 28356 5704 28408 5710
rect 28356 5646 28408 5652
rect 29092 5704 29144 5710
rect 29092 5646 29144 5652
rect 28368 4214 28396 5646
rect 28724 4684 28776 4690
rect 28724 4626 28776 4632
rect 28356 4208 28408 4214
rect 28356 4150 28408 4156
rect 27804 4140 27856 4146
rect 27804 4082 27856 4088
rect 27620 4004 27672 4010
rect 27620 3946 27672 3952
rect 27632 3058 27660 3946
rect 27528 3052 27580 3058
rect 27528 2994 27580 3000
rect 27620 3052 27672 3058
rect 27620 2994 27672 3000
rect 27528 2848 27580 2854
rect 27264 2746 27384 2774
rect 27448 2808 27528 2836
rect 27264 2446 27292 2746
rect 27344 2644 27396 2650
rect 27344 2586 27396 2592
rect 27252 2440 27304 2446
rect 27252 2382 27304 2388
rect 26884 2372 26936 2378
rect 26884 2314 26936 2320
rect 26792 2100 26844 2106
rect 26792 2042 26844 2048
rect 26804 1766 26832 2042
rect 26792 1760 26844 1766
rect 26792 1702 26844 1708
rect 26700 264 26752 270
rect 26700 206 26752 212
rect 26896 56 26924 2314
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 27172 56 27292 82
rect 21008 54 21142 56
rect 21008 42 21036 54
rect 20916 14 21036 42
rect 21086 0 21142 54
rect 21362 0 21418 56
rect 21638 0 21694 56
rect 21914 0 21970 56
rect 22190 0 22246 56
rect 22466 0 22522 56
rect 22742 0 22798 56
rect 23018 0 23074 56
rect 23294 0 23350 56
rect 23570 0 23626 56
rect 23846 0 23902 56
rect 24122 0 24178 56
rect 24398 0 24454 56
rect 24674 0 24730 56
rect 24950 0 25006 56
rect 25226 0 25282 56
rect 25502 0 25558 56
rect 25778 0 25834 56
rect 26054 0 26110 56
rect 26330 0 26386 56
rect 26606 0 26662 56
rect 26882 0 26938 56
rect 27158 54 27292 56
rect 27158 0 27214 54
rect 27264 42 27292 54
rect 27356 42 27384 2586
rect 27448 56 27476 2808
rect 27528 2790 27580 2796
rect 27712 2576 27764 2582
rect 27712 2518 27764 2524
rect 27528 2440 27580 2446
rect 27528 2382 27580 2388
rect 27620 2440 27672 2446
rect 27620 2382 27672 2388
rect 27540 1698 27568 2382
rect 27528 1692 27580 1698
rect 27528 1634 27580 1640
rect 27632 1630 27660 2382
rect 27620 1624 27672 1630
rect 27620 1566 27672 1572
rect 27724 56 27752 2518
rect 27816 338 27844 4082
rect 28736 2922 28764 4626
rect 28998 2952 29054 2961
rect 28724 2916 28776 2922
rect 28998 2887 29000 2896
rect 28724 2858 28776 2864
rect 29052 2887 29054 2896
rect 29000 2858 29052 2864
rect 28264 2848 28316 2854
rect 28632 2848 28684 2854
rect 28264 2790 28316 2796
rect 28552 2808 28632 2836
rect 27988 2372 28040 2378
rect 27988 2314 28040 2320
rect 27804 332 27856 338
rect 27804 274 27856 280
rect 28000 56 28028 2314
rect 28276 56 28304 2790
rect 28448 2440 28500 2446
rect 28448 2382 28500 2388
rect 28460 2038 28488 2382
rect 28448 2032 28500 2038
rect 28448 1974 28500 1980
rect 28552 56 28580 2808
rect 28632 2790 28684 2796
rect 29380 2774 29408 6666
rect 29472 6186 29500 7414
rect 31036 7206 31064 8774
rect 31024 7200 31076 7206
rect 31024 7142 31076 7148
rect 29552 6656 29604 6662
rect 29552 6598 29604 6604
rect 29828 6656 29880 6662
rect 29828 6598 29880 6604
rect 29460 6180 29512 6186
rect 29460 6122 29512 6128
rect 29564 4078 29592 6598
rect 29840 6254 29868 6598
rect 29828 6248 29880 6254
rect 29828 6190 29880 6196
rect 29642 5672 29698 5681
rect 29642 5607 29698 5616
rect 31116 5636 31168 5642
rect 29656 5302 29684 5607
rect 31116 5578 31168 5584
rect 30380 5568 30432 5574
rect 30380 5510 30432 5516
rect 29644 5296 29696 5302
rect 29644 5238 29696 5244
rect 30286 5264 30342 5273
rect 30286 5199 30342 5208
rect 29920 4752 29972 4758
rect 29920 4694 29972 4700
rect 29552 4072 29604 4078
rect 29552 4014 29604 4020
rect 29644 2848 29696 2854
rect 29644 2790 29696 2796
rect 29380 2746 29592 2774
rect 28816 2576 28868 2582
rect 28816 2518 28868 2524
rect 28632 2440 28684 2446
rect 28632 2382 28684 2388
rect 28644 1902 28672 2382
rect 28632 1896 28684 1902
rect 28632 1838 28684 1844
rect 28828 56 28856 2518
rect 29564 2446 29592 2746
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 29368 2372 29420 2378
rect 29368 2314 29420 2320
rect 29092 2304 29144 2310
rect 29092 2246 29144 2252
rect 29104 56 29132 2246
rect 29380 56 29408 2314
rect 29656 56 29684 2790
rect 29932 2774 29960 4694
rect 30012 3460 30064 3466
rect 30012 3402 30064 3408
rect 30024 3058 30052 3402
rect 30012 3052 30064 3058
rect 30012 2994 30064 3000
rect 30104 2984 30156 2990
rect 30104 2926 30156 2932
rect 29932 2746 30052 2774
rect 29920 2576 29972 2582
rect 29920 2518 29972 2524
rect 29736 2440 29788 2446
rect 29736 2382 29788 2388
rect 29748 1970 29776 2382
rect 29736 1964 29788 1970
rect 29736 1906 29788 1912
rect 29932 56 29960 2518
rect 30024 2514 30052 2746
rect 30012 2508 30064 2514
rect 30012 2450 30064 2456
rect 30116 513 30144 2926
rect 30300 2774 30328 5199
rect 30392 4826 30420 5510
rect 30380 4820 30432 4826
rect 30380 4762 30432 4768
rect 30656 3936 30708 3942
rect 30656 3878 30708 3884
rect 30380 3596 30432 3602
rect 30380 3538 30432 3544
rect 30392 2961 30420 3538
rect 30378 2952 30434 2961
rect 30378 2887 30434 2896
rect 30300 2746 30420 2774
rect 30392 2666 30420 2746
rect 30196 2644 30248 2650
rect 30196 2586 30248 2592
rect 30300 2638 30420 2666
rect 30102 504 30158 513
rect 30102 439 30158 448
rect 30208 56 30236 2586
rect 30300 2446 30328 2638
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 30564 2372 30616 2378
rect 30564 2314 30616 2320
rect 30576 1170 30604 2314
rect 30668 1698 30696 3878
rect 31024 3052 31076 3058
rect 31024 2994 31076 3000
rect 30840 2984 30892 2990
rect 30840 2926 30892 2932
rect 30748 2848 30800 2854
rect 30748 2790 30800 2796
rect 30656 1692 30708 1698
rect 30656 1634 30708 1640
rect 30484 1142 30604 1170
rect 30484 56 30512 1142
rect 30760 56 30788 2790
rect 30852 1494 30880 2926
rect 31036 2854 31064 2994
rect 31024 2848 31076 2854
rect 31024 2790 31076 2796
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 30944 1834 30972 2382
rect 31024 2304 31076 2310
rect 31024 2246 31076 2252
rect 30932 1828 30984 1834
rect 30932 1770 30984 1776
rect 30840 1488 30892 1494
rect 30840 1430 30892 1436
rect 31036 56 31064 2246
rect 31128 2009 31156 5578
rect 31208 5228 31260 5234
rect 31208 5170 31260 5176
rect 31114 2000 31170 2009
rect 31114 1935 31170 1944
rect 31220 649 31248 5170
rect 31864 3942 31892 8842
rect 33060 8820 33088 11194
rect 32876 8792 33088 8820
rect 32876 8634 32904 8792
rect 33010 8732 33318 8741
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 33010 8667 33318 8676
rect 35176 8634 35204 11194
rect 37292 8634 37320 11194
rect 39010 8732 39318 8741
rect 39010 8730 39016 8732
rect 39072 8730 39096 8732
rect 39152 8730 39176 8732
rect 39232 8730 39256 8732
rect 39312 8730 39318 8732
rect 39072 8678 39074 8730
rect 39254 8678 39256 8730
rect 39010 8676 39016 8678
rect 39072 8676 39096 8678
rect 39152 8676 39176 8678
rect 39232 8676 39256 8678
rect 39312 8676 39318 8678
rect 39010 8667 39318 8676
rect 39408 8634 39436 11194
rect 41420 8832 41472 8838
rect 41420 8774 41472 8780
rect 41432 8634 41460 8774
rect 41524 8634 41552 11194
rect 41970 9888 42026 9897
rect 41970 9823 42026 9832
rect 32864 8628 32916 8634
rect 32864 8570 32916 8576
rect 35164 8628 35216 8634
rect 35164 8570 35216 8576
rect 37280 8628 37332 8634
rect 37280 8570 37332 8576
rect 39396 8628 39448 8634
rect 39396 8570 39448 8576
rect 41420 8628 41472 8634
rect 41420 8570 41472 8576
rect 41512 8628 41564 8634
rect 41512 8570 41564 8576
rect 33324 8492 33376 8498
rect 34980 8492 35032 8498
rect 33376 8452 33456 8480
rect 33324 8434 33376 8440
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 33010 7644 33318 7653
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 33010 6556 33318 6565
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 33232 6180 33284 6186
rect 33232 6122 33284 6128
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 33244 5778 33272 6122
rect 33428 5846 33456 8452
rect 34980 8434 35032 8440
rect 35072 8492 35124 8498
rect 35072 8434 35124 8440
rect 37648 8492 37700 8498
rect 37648 8434 37700 8440
rect 39856 8492 39908 8498
rect 39856 8434 39908 8440
rect 41236 8492 41288 8498
rect 41236 8434 41288 8440
rect 41604 8492 41656 8498
rect 41604 8434 41656 8440
rect 34428 6656 34480 6662
rect 34428 6598 34480 6604
rect 34150 6216 34206 6225
rect 34150 6151 34206 6160
rect 33416 5840 33468 5846
rect 33416 5782 33468 5788
rect 33232 5772 33284 5778
rect 33232 5714 33284 5720
rect 33968 5772 34020 5778
rect 33968 5714 34020 5720
rect 33980 5681 34008 5714
rect 33966 5672 34022 5681
rect 33966 5607 34022 5616
rect 33010 5468 33318 5477
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 33010 5403 33318 5412
rect 33508 5296 33560 5302
rect 33508 5238 33560 5244
rect 33140 5160 33192 5166
rect 33192 5108 33364 5114
rect 33140 5102 33364 5108
rect 33152 5098 33364 5102
rect 33152 5092 33376 5098
rect 33152 5086 33324 5092
rect 33324 5034 33376 5040
rect 33416 5024 33468 5030
rect 33416 4966 33468 4972
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 33010 4380 33318 4389
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 32864 4140 32916 4146
rect 32864 4082 32916 4088
rect 31852 3936 31904 3942
rect 31852 3878 31904 3884
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 31852 3392 31904 3398
rect 31852 3334 31904 3340
rect 31668 3188 31720 3194
rect 31668 3130 31720 3136
rect 31680 2990 31708 3130
rect 31484 2984 31536 2990
rect 31484 2926 31536 2932
rect 31668 2984 31720 2990
rect 31668 2926 31720 2932
rect 31496 2854 31524 2926
rect 31484 2848 31536 2854
rect 31484 2790 31536 2796
rect 31300 2576 31352 2582
rect 31300 2518 31352 2524
rect 31206 640 31262 649
rect 31206 575 31262 584
rect 31312 56 31340 2518
rect 31484 2440 31536 2446
rect 31484 2382 31536 2388
rect 31496 1902 31524 2382
rect 31576 2372 31628 2378
rect 31576 2314 31628 2320
rect 31484 1896 31536 1902
rect 31484 1838 31536 1844
rect 31588 56 31616 2314
rect 31864 56 31892 3334
rect 32772 3052 32824 3058
rect 32772 2994 32824 3000
rect 32784 2854 32812 2994
rect 32772 2848 32824 2854
rect 32772 2790 32824 2796
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 32404 2644 32456 2650
rect 32404 2586 32456 2592
rect 32312 2440 32364 2446
rect 32126 2408 32182 2417
rect 32312 2382 32364 2388
rect 32126 2343 32182 2352
rect 32140 56 32168 2343
rect 32324 1970 32352 2382
rect 32312 1964 32364 1970
rect 32312 1906 32364 1912
rect 32416 56 32444 2586
rect 32680 2440 32732 2446
rect 32680 2382 32732 2388
rect 32772 2440 32824 2446
rect 32772 2382 32824 2388
rect 32692 2038 32720 2382
rect 32784 2106 32812 2382
rect 32772 2100 32824 2106
rect 32772 2042 32824 2048
rect 32680 2032 32732 2038
rect 32680 1974 32732 1980
rect 32678 1456 32734 1465
rect 32678 1391 32734 1400
rect 32692 56 32720 1391
rect 32876 1290 32904 4082
rect 33010 3292 33318 3301
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 33048 3188 33100 3194
rect 33048 3130 33100 3136
rect 32956 2848 33008 2854
rect 32956 2790 33008 2796
rect 32968 2514 32996 2790
rect 33060 2530 33088 3130
rect 33428 3126 33456 4966
rect 33520 4758 33548 5238
rect 33508 4752 33560 4758
rect 33508 4694 33560 4700
rect 34058 4720 34114 4729
rect 34058 4655 34114 4664
rect 33600 4004 33652 4010
rect 33600 3946 33652 3952
rect 33416 3120 33468 3126
rect 33416 3062 33468 3068
rect 33612 3058 33640 3946
rect 33600 3052 33652 3058
rect 33600 2994 33652 3000
rect 33692 2984 33744 2990
rect 33692 2926 33744 2932
rect 33600 2916 33652 2922
rect 33600 2858 33652 2864
rect 33416 2848 33468 2854
rect 33416 2790 33468 2796
rect 33508 2848 33560 2854
rect 33508 2790 33560 2796
rect 33060 2514 33364 2530
rect 32956 2508 33008 2514
rect 33060 2508 33376 2514
rect 33060 2502 33324 2508
rect 32956 2450 33008 2456
rect 33324 2450 33376 2456
rect 33138 2408 33194 2417
rect 33138 2343 33194 2352
rect 33152 2310 33180 2343
rect 33140 2304 33192 2310
rect 33140 2246 33192 2252
rect 33010 2204 33318 2213
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 33428 1442 33456 2790
rect 32968 1414 33456 1442
rect 32864 1284 32916 1290
rect 32864 1226 32916 1232
rect 32968 56 32996 1414
rect 33232 1352 33284 1358
rect 33232 1294 33284 1300
rect 33244 56 33272 1294
rect 33520 56 33548 2790
rect 33612 2446 33640 2858
rect 33600 2440 33652 2446
rect 33600 2382 33652 2388
rect 33600 2304 33652 2310
rect 33600 2246 33652 2252
rect 33612 1465 33640 2246
rect 33598 1456 33654 1465
rect 33598 1391 33654 1400
rect 33704 377 33732 2926
rect 33876 2916 33928 2922
rect 33876 2858 33928 2864
rect 33888 2774 33916 2858
rect 33968 2848 34020 2854
rect 33968 2790 34020 2796
rect 33796 2746 33916 2774
rect 33796 2446 33824 2746
rect 33784 2440 33836 2446
rect 33784 2382 33836 2388
rect 33876 2372 33928 2378
rect 33876 2314 33928 2320
rect 33888 1170 33916 2314
rect 33796 1142 33916 1170
rect 33690 368 33746 377
rect 33690 303 33746 312
rect 33796 56 33824 1142
rect 33980 202 34008 2790
rect 33968 196 34020 202
rect 33968 138 34020 144
rect 34072 56 34100 4655
rect 27264 14 27384 42
rect 27434 0 27490 56
rect 27710 0 27766 56
rect 27986 0 28042 56
rect 28262 0 28318 56
rect 28538 0 28594 56
rect 28814 0 28870 56
rect 29090 0 29146 56
rect 29366 0 29422 56
rect 29642 0 29698 56
rect 29918 0 29974 56
rect 30194 0 30250 56
rect 30470 0 30526 56
rect 30746 0 30802 56
rect 31022 0 31078 56
rect 31298 0 31354 56
rect 31574 0 31630 56
rect 31850 0 31906 56
rect 32126 0 32182 56
rect 32402 0 32458 56
rect 32678 0 32734 56
rect 32954 0 33010 56
rect 33230 0 33286 56
rect 33506 0 33562 56
rect 33782 0 33838 56
rect 34058 0 34114 56
rect 34164 42 34192 6151
rect 34440 3670 34468 6598
rect 34992 5370 35020 8434
rect 35084 6662 35112 8434
rect 36544 7948 36596 7954
rect 36544 7890 36596 7896
rect 36556 7410 36584 7890
rect 36820 7472 36872 7478
rect 36820 7414 36872 7420
rect 36544 7404 36596 7410
rect 36544 7346 36596 7352
rect 36452 7336 36504 7342
rect 36452 7278 36504 7284
rect 35624 6996 35676 7002
rect 35624 6938 35676 6944
rect 35072 6656 35124 6662
rect 35072 6598 35124 6604
rect 35636 6390 35664 6938
rect 36268 6452 36320 6458
rect 36268 6394 36320 6400
rect 35624 6384 35676 6390
rect 35624 6326 35676 6332
rect 35808 5840 35860 5846
rect 35808 5782 35860 5788
rect 35348 5568 35400 5574
rect 35348 5510 35400 5516
rect 34980 5364 35032 5370
rect 34980 5306 35032 5312
rect 34704 3732 34756 3738
rect 34704 3674 34756 3680
rect 34428 3664 34480 3670
rect 34428 3606 34480 3612
rect 34244 3528 34296 3534
rect 34244 3470 34296 3476
rect 34256 3194 34284 3470
rect 34244 3188 34296 3194
rect 34244 3130 34296 3136
rect 34428 3188 34480 3194
rect 34428 3130 34480 3136
rect 34336 2848 34388 2854
rect 34336 2790 34388 2796
rect 34244 2304 34296 2310
rect 34244 2246 34296 2252
rect 34256 1426 34284 2246
rect 34348 2106 34376 2790
rect 34336 2100 34388 2106
rect 34336 2042 34388 2048
rect 34440 1902 34468 3130
rect 34716 2446 34744 3674
rect 34796 3052 34848 3058
rect 34796 2994 34848 3000
rect 34704 2440 34756 2446
rect 34704 2382 34756 2388
rect 34428 1896 34480 1902
rect 34428 1838 34480 1844
rect 34610 1728 34666 1737
rect 34610 1663 34666 1672
rect 34244 1420 34296 1426
rect 34244 1362 34296 1368
rect 34256 56 34376 82
rect 34624 56 34652 1663
rect 34808 241 34836 2994
rect 35162 2952 35218 2961
rect 35162 2887 35218 2896
rect 34980 2848 35032 2854
rect 34980 2790 35032 2796
rect 34992 2038 35020 2790
rect 35072 2440 35124 2446
rect 35072 2382 35124 2388
rect 34980 2032 35032 2038
rect 34980 1974 35032 1980
rect 35084 1698 35112 2382
rect 35072 1692 35124 1698
rect 35072 1634 35124 1640
rect 34794 232 34850 241
rect 34794 167 34850 176
rect 34886 96 34942 105
rect 34256 54 34390 56
rect 34256 42 34284 54
rect 34164 14 34284 42
rect 34334 0 34390 54
rect 34610 0 34666 56
rect 35176 56 35204 2887
rect 35360 1970 35388 5510
rect 35624 4616 35676 4622
rect 35624 4558 35676 4564
rect 35636 2774 35664 4558
rect 35714 3088 35770 3097
rect 35714 3023 35716 3032
rect 35768 3023 35770 3032
rect 35716 2994 35768 3000
rect 35820 2774 35848 5782
rect 35636 2746 35756 2774
rect 35820 2746 36032 2774
rect 35348 1964 35400 1970
rect 35348 1906 35400 1912
rect 35440 1284 35492 1290
rect 35440 1226 35492 1232
rect 35452 56 35480 1226
rect 35728 56 35756 2746
rect 36004 56 36032 2746
rect 36280 56 36308 6394
rect 36464 2774 36492 7278
rect 36544 4820 36596 4826
rect 36544 4762 36596 4768
rect 36556 4214 36584 4762
rect 36544 4208 36596 4214
rect 36544 4150 36596 4156
rect 36464 2746 36584 2774
rect 36556 56 36584 2746
rect 36832 56 36860 7414
rect 37660 6458 37688 8434
rect 37950 8188 38258 8197
rect 37950 8186 37956 8188
rect 38012 8186 38036 8188
rect 38092 8186 38116 8188
rect 38172 8186 38196 8188
rect 38252 8186 38258 8188
rect 38012 8134 38014 8186
rect 38194 8134 38196 8186
rect 37950 8132 37956 8134
rect 38012 8132 38036 8134
rect 38092 8132 38116 8134
rect 38172 8132 38196 8134
rect 38252 8132 38258 8134
rect 37950 8123 38258 8132
rect 39010 7644 39318 7653
rect 39010 7642 39016 7644
rect 39072 7642 39096 7644
rect 39152 7642 39176 7644
rect 39232 7642 39256 7644
rect 39312 7642 39318 7644
rect 39072 7590 39074 7642
rect 39254 7590 39256 7642
rect 39010 7588 39016 7590
rect 39072 7588 39096 7590
rect 39152 7588 39176 7590
rect 39232 7588 39256 7590
rect 39312 7588 39318 7590
rect 39010 7579 39318 7588
rect 37950 7100 38258 7109
rect 37950 7098 37956 7100
rect 38012 7098 38036 7100
rect 38092 7098 38116 7100
rect 38172 7098 38196 7100
rect 38252 7098 38258 7100
rect 38012 7046 38014 7098
rect 38194 7046 38196 7098
rect 37950 7044 37956 7046
rect 38012 7044 38036 7046
rect 38092 7044 38116 7046
rect 38172 7044 38196 7046
rect 38252 7044 38258 7046
rect 37950 7035 38258 7044
rect 38476 6792 38528 6798
rect 38476 6734 38528 6740
rect 37648 6452 37700 6458
rect 37648 6394 37700 6400
rect 37648 6316 37700 6322
rect 37648 6258 37700 6264
rect 37188 6248 37240 6254
rect 37188 6190 37240 6196
rect 37004 3052 37056 3058
rect 37004 2994 37056 3000
rect 37096 3052 37148 3058
rect 37096 2994 37148 3000
rect 37016 66 37044 2994
rect 37108 1766 37136 2994
rect 37096 1760 37148 1766
rect 37096 1702 37148 1708
rect 37200 1442 37228 6190
rect 37372 6180 37424 6186
rect 37372 6122 37424 6128
rect 37280 5024 37332 5030
rect 37280 4966 37332 4972
rect 37292 1834 37320 4966
rect 37280 1828 37332 1834
rect 37280 1770 37332 1776
rect 37108 1414 37228 1442
rect 37004 60 37056 66
rect 34886 0 34942 40
rect 35162 0 35218 56
rect 35438 0 35494 56
rect 35714 0 35770 56
rect 35990 0 36046 56
rect 36266 0 36322 56
rect 36542 0 36598 56
rect 36818 0 36874 56
rect 37108 56 37136 1414
rect 37384 56 37412 6122
rect 37556 5024 37608 5030
rect 37556 4966 37608 4972
rect 37568 134 37596 4966
rect 37556 128 37608 134
rect 37556 70 37608 76
rect 37660 56 37688 6258
rect 37950 6012 38258 6021
rect 37950 6010 37956 6012
rect 38012 6010 38036 6012
rect 38092 6010 38116 6012
rect 38172 6010 38196 6012
rect 38252 6010 38258 6012
rect 38012 5958 38014 6010
rect 38194 5958 38196 6010
rect 37950 5956 37956 5958
rect 38012 5956 38036 5958
rect 38092 5956 38116 5958
rect 38172 5956 38196 5958
rect 38252 5956 38258 5958
rect 37950 5947 38258 5956
rect 37832 5636 37884 5642
rect 37832 5578 37884 5584
rect 37844 1442 37872 5578
rect 38292 5160 38344 5166
rect 38292 5102 38344 5108
rect 37950 4924 38258 4933
rect 37950 4922 37956 4924
rect 38012 4922 38036 4924
rect 38092 4922 38116 4924
rect 38172 4922 38196 4924
rect 38252 4922 38258 4924
rect 38012 4870 38014 4922
rect 38194 4870 38196 4922
rect 37950 4868 37956 4870
rect 38012 4868 38036 4870
rect 38092 4868 38116 4870
rect 38172 4868 38196 4870
rect 38252 4868 38258 4870
rect 37950 4859 38258 4868
rect 37950 3836 38258 3845
rect 37950 3834 37956 3836
rect 38012 3834 38036 3836
rect 38092 3834 38116 3836
rect 38172 3834 38196 3836
rect 38252 3834 38258 3836
rect 38012 3782 38014 3834
rect 38194 3782 38196 3834
rect 37950 3780 37956 3782
rect 38012 3780 38036 3782
rect 38092 3780 38116 3782
rect 38172 3780 38196 3782
rect 38252 3780 38258 3782
rect 37950 3771 38258 3780
rect 38108 3460 38160 3466
rect 38108 3402 38160 3408
rect 38120 3194 38148 3402
rect 38108 3188 38160 3194
rect 38108 3130 38160 3136
rect 37950 2748 38258 2757
rect 37950 2746 37956 2748
rect 38012 2746 38036 2748
rect 38092 2746 38116 2748
rect 38172 2746 38196 2748
rect 38252 2746 38258 2748
rect 38012 2694 38014 2746
rect 38194 2694 38196 2746
rect 37950 2692 37956 2694
rect 38012 2692 38036 2694
rect 38092 2692 38116 2694
rect 38172 2692 38196 2694
rect 38252 2692 38258 2694
rect 37950 2683 38258 2692
rect 38304 1442 38332 5102
rect 37844 1414 37964 1442
rect 37936 56 37964 1414
rect 38212 1414 38332 1442
rect 38212 56 38240 1414
rect 38488 56 38516 6734
rect 39010 6556 39318 6565
rect 39010 6554 39016 6556
rect 39072 6554 39096 6556
rect 39152 6554 39176 6556
rect 39232 6554 39256 6556
rect 39312 6554 39318 6556
rect 39072 6502 39074 6554
rect 39254 6502 39256 6554
rect 39010 6500 39016 6502
rect 39072 6500 39096 6502
rect 39152 6500 39176 6502
rect 39232 6500 39256 6502
rect 39312 6500 39318 6502
rect 39010 6491 39318 6500
rect 39868 6458 39896 8434
rect 40040 8424 40092 8430
rect 40040 8366 40092 8372
rect 40052 8294 40080 8366
rect 40040 8288 40092 8294
rect 40040 8230 40092 8236
rect 41248 6458 41276 8434
rect 39856 6452 39908 6458
rect 39856 6394 39908 6400
rect 41236 6452 41288 6458
rect 41236 6394 41288 6400
rect 38936 6316 38988 6322
rect 38936 6258 38988 6264
rect 39396 6316 39448 6322
rect 39396 6258 39448 6264
rect 39580 6316 39632 6322
rect 39580 6258 39632 6264
rect 38752 6248 38804 6254
rect 38752 6190 38804 6196
rect 38660 5704 38712 5710
rect 38660 5646 38712 5652
rect 38672 3641 38700 5646
rect 38658 3632 38714 3641
rect 38658 3567 38714 3576
rect 38764 56 38792 6190
rect 38948 1442 38976 6258
rect 39010 5468 39318 5477
rect 39010 5466 39016 5468
rect 39072 5466 39096 5468
rect 39152 5466 39176 5468
rect 39232 5466 39256 5468
rect 39312 5466 39318 5468
rect 39072 5414 39074 5466
rect 39254 5414 39256 5466
rect 39010 5412 39016 5414
rect 39072 5412 39096 5414
rect 39152 5412 39176 5414
rect 39232 5412 39256 5414
rect 39312 5412 39318 5414
rect 39010 5403 39318 5412
rect 39010 4380 39318 4389
rect 39010 4378 39016 4380
rect 39072 4378 39096 4380
rect 39152 4378 39176 4380
rect 39232 4378 39256 4380
rect 39312 4378 39318 4380
rect 39072 4326 39074 4378
rect 39254 4326 39256 4378
rect 39010 4324 39016 4326
rect 39072 4324 39096 4326
rect 39152 4324 39176 4326
rect 39232 4324 39256 4326
rect 39312 4324 39318 4326
rect 39010 4315 39318 4324
rect 39010 3292 39318 3301
rect 39010 3290 39016 3292
rect 39072 3290 39096 3292
rect 39152 3290 39176 3292
rect 39232 3290 39256 3292
rect 39312 3290 39318 3292
rect 39072 3238 39074 3290
rect 39254 3238 39256 3290
rect 39010 3236 39016 3238
rect 39072 3236 39096 3238
rect 39152 3236 39176 3238
rect 39232 3236 39256 3238
rect 39312 3236 39318 3238
rect 39010 3227 39318 3236
rect 39010 2204 39318 2213
rect 39010 2202 39016 2204
rect 39072 2202 39096 2204
rect 39152 2202 39176 2204
rect 39232 2202 39256 2204
rect 39312 2202 39318 2204
rect 39072 2150 39074 2202
rect 39254 2150 39256 2202
rect 39010 2148 39016 2150
rect 39072 2148 39096 2150
rect 39152 2148 39176 2150
rect 39232 2148 39256 2150
rect 39312 2148 39318 2150
rect 39010 2139 39318 2148
rect 39408 1442 39436 6258
rect 38948 1414 39068 1442
rect 39040 56 39068 1414
rect 39316 1414 39436 1442
rect 39316 56 39344 1414
rect 39592 56 39620 6258
rect 41616 6186 41644 8434
rect 41984 8090 42012 9823
rect 42338 9616 42394 9625
rect 42338 9551 42394 9560
rect 42154 8800 42210 8809
rect 42154 8735 42210 8744
rect 42168 8634 42196 8735
rect 42156 8628 42208 8634
rect 42156 8570 42208 8576
rect 42352 8090 42380 9551
rect 43166 9344 43222 9353
rect 43166 9279 43222 9288
rect 42614 9072 42670 9081
rect 42614 9007 42670 9016
rect 42628 8090 42656 9007
rect 42708 8628 42760 8634
rect 42708 8570 42760 8576
rect 42720 8537 42748 8570
rect 42706 8528 42762 8537
rect 42706 8463 42762 8472
rect 43076 8356 43128 8362
rect 43076 8298 43128 8304
rect 43088 8265 43116 8298
rect 43074 8256 43130 8265
rect 43074 8191 43130 8200
rect 41972 8084 42024 8090
rect 41972 8026 42024 8032
rect 42340 8084 42392 8090
rect 42340 8026 42392 8032
rect 42616 8084 42668 8090
rect 42616 8026 42668 8032
rect 41788 7880 41840 7886
rect 41788 7822 41840 7828
rect 42616 7880 42668 7886
rect 42616 7822 42668 7828
rect 41800 7546 41828 7822
rect 41788 7540 41840 7546
rect 41788 7482 41840 7488
rect 41604 6180 41656 6186
rect 41604 6122 41656 6128
rect 42340 6112 42392 6118
rect 42340 6054 42392 6060
rect 41972 4752 42024 4758
rect 41972 4694 42024 4700
rect 40040 4276 40092 4282
rect 40040 4218 40092 4224
rect 40052 3058 40080 4218
rect 40040 3052 40092 3058
rect 40040 2994 40092 3000
rect 41984 2446 42012 4694
rect 42352 3126 42380 6054
rect 42628 5302 42656 7822
rect 43076 7744 43128 7750
rect 43076 7686 43128 7692
rect 43088 7449 43116 7686
rect 43180 7546 43208 9279
rect 43640 8838 43668 11194
rect 43628 8832 43680 8838
rect 43628 8774 43680 8780
rect 43444 8356 43496 8362
rect 43444 8298 43496 8304
rect 43456 7993 43484 8298
rect 43442 7984 43498 7993
rect 43442 7919 43498 7928
rect 43260 7880 43312 7886
rect 43260 7822 43312 7828
rect 43168 7540 43220 7546
rect 43168 7482 43220 7488
rect 43074 7440 43130 7449
rect 43074 7375 43130 7384
rect 43272 6934 43300 7822
rect 43444 7744 43496 7750
rect 43442 7712 43444 7721
rect 43496 7712 43498 7721
rect 43442 7647 43498 7656
rect 43444 7200 43496 7206
rect 43442 7168 43444 7177
rect 43496 7168 43498 7177
rect 43442 7103 43498 7112
rect 43260 6928 43312 6934
rect 43260 6870 43312 6876
rect 43442 6896 43498 6905
rect 43442 6831 43498 6840
rect 42984 6792 43036 6798
rect 42984 6734 43036 6740
rect 42892 6316 42944 6322
rect 42892 6258 42944 6264
rect 42616 5296 42668 5302
rect 42616 5238 42668 5244
rect 42800 5228 42852 5234
rect 42800 5170 42852 5176
rect 42812 4049 42840 5170
rect 42904 5098 42932 6258
rect 42996 5914 43024 6734
rect 43456 6662 43484 6831
rect 43076 6656 43128 6662
rect 43074 6624 43076 6633
rect 43444 6656 43496 6662
rect 43128 6624 43130 6633
rect 43444 6598 43496 6604
rect 43074 6559 43130 6568
rect 43444 6452 43496 6458
rect 43444 6394 43496 6400
rect 43168 6384 43220 6390
rect 43456 6361 43484 6394
rect 43168 6326 43220 6332
rect 43258 6352 43314 6361
rect 43076 6112 43128 6118
rect 43074 6080 43076 6089
rect 43128 6080 43130 6089
rect 43074 6015 43130 6024
rect 42984 5908 43036 5914
rect 42984 5850 43036 5856
rect 43076 5568 43128 5574
rect 43074 5536 43076 5545
rect 43128 5536 43130 5545
rect 43074 5471 43130 5480
rect 42892 5092 42944 5098
rect 42892 5034 42944 5040
rect 43076 5024 43128 5030
rect 43074 4992 43076 5001
rect 43128 4992 43130 5001
rect 43074 4927 43130 4936
rect 42984 4616 43036 4622
rect 42984 4558 43036 4564
rect 42892 4480 42944 4486
rect 42892 4422 42944 4428
rect 42798 4040 42854 4049
rect 42798 3975 42854 3984
rect 42904 3534 42932 4422
rect 42996 3602 43024 4558
rect 43076 4480 43128 4486
rect 43074 4448 43076 4457
rect 43128 4448 43130 4457
rect 43074 4383 43130 4392
rect 43076 3936 43128 3942
rect 43074 3904 43076 3913
rect 43128 3904 43130 3913
rect 43074 3839 43130 3848
rect 42984 3596 43036 3602
rect 42984 3538 43036 3544
rect 42892 3528 42944 3534
rect 42892 3470 42944 3476
rect 43076 3392 43128 3398
rect 43074 3360 43076 3369
rect 43128 3360 43130 3369
rect 43074 3295 43130 3304
rect 42340 3120 42392 3126
rect 42340 3062 42392 3068
rect 43180 3058 43208 6326
rect 43258 6287 43260 6296
rect 43312 6287 43314 6296
rect 43442 6352 43498 6361
rect 43442 6287 43498 6296
rect 43260 6258 43312 6264
rect 43444 5840 43496 5846
rect 43442 5808 43444 5817
rect 43496 5808 43498 5817
rect 43442 5743 43498 5752
rect 43444 5364 43496 5370
rect 43444 5306 43496 5312
rect 43456 5273 43484 5306
rect 43442 5264 43498 5273
rect 43260 5228 43312 5234
rect 43442 5199 43498 5208
rect 43260 5170 43312 5176
rect 43272 3505 43300 5170
rect 43444 4752 43496 4758
rect 43442 4720 43444 4729
rect 43496 4720 43498 4729
rect 43442 4655 43498 4664
rect 43442 4176 43498 4185
rect 43442 4111 43498 4120
rect 43456 4010 43484 4111
rect 43444 4004 43496 4010
rect 43444 3946 43496 3952
rect 43444 3664 43496 3670
rect 43442 3632 43444 3641
rect 43496 3632 43498 3641
rect 43442 3567 43498 3576
rect 43258 3496 43314 3505
rect 43258 3431 43314 3440
rect 43444 3188 43496 3194
rect 43444 3130 43496 3136
rect 43456 3097 43484 3130
rect 43442 3088 43498 3097
rect 43168 3052 43220 3058
rect 43442 3023 43498 3032
rect 43168 2994 43220 3000
rect 42984 2848 43036 2854
rect 43076 2848 43128 2854
rect 42984 2790 43036 2796
rect 43074 2816 43076 2825
rect 43128 2816 43130 2825
rect 42522 2544 42578 2553
rect 42522 2479 42578 2488
rect 42536 2446 42564 2479
rect 41972 2440 42024 2446
rect 41972 2382 42024 2388
rect 42524 2440 42576 2446
rect 42524 2382 42576 2388
rect 42156 2304 42208 2310
rect 42156 2246 42208 2252
rect 42708 2304 42760 2310
rect 42708 2246 42760 2252
rect 42168 1737 42196 2246
rect 42154 1728 42210 1737
rect 42154 1663 42210 1672
rect 42720 1465 42748 2246
rect 42996 2009 43024 2790
rect 43074 2751 43130 2760
rect 43444 2576 43496 2582
rect 43442 2544 43444 2553
rect 43496 2544 43498 2553
rect 43442 2479 43498 2488
rect 43076 2304 43128 2310
rect 43074 2272 43076 2281
rect 43128 2272 43130 2281
rect 43074 2207 43130 2216
rect 42982 2000 43038 2009
rect 42982 1935 43038 1944
rect 42706 1456 42762 1465
rect 42706 1391 42762 1400
rect 37004 2 37056 8
rect 37094 0 37150 56
rect 37370 0 37426 56
rect 37646 0 37702 56
rect 37922 0 37978 56
rect 38198 0 38254 56
rect 38474 0 38530 56
rect 38750 0 38806 56
rect 39026 0 39082 56
rect 39302 0 39358 56
rect 39578 0 39634 56
<< via2 >>
rect 1214 9832 1270 9888
rect 2870 8744 2926 8800
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 14922 9288 14978 9344
rect 1214 8336 1270 8392
rect 2870 8336 2926 8392
rect 1766 8200 1822 8256
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 1306 7384 1362 7440
rect 1766 7384 1822 7440
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 2870 5480 2926 5536
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 2870 5072 2926 5128
rect 1766 4936 1822 4992
rect 1306 4392 1362 4448
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 1214 4156 1216 4176
rect 1216 4156 1268 4176
rect 1268 4156 1270 4176
rect 1214 4120 1270 4156
rect 1766 4120 1822 4176
rect 2870 3984 2926 4040
rect 1766 3848 1822 3904
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 1766 3440 1822 3496
rect 2870 3304 2926 3360
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 938 1400 994 1456
rect 5538 1944 5594 2000
rect 7746 8200 7802 8256
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 19338 9560 19394 9616
rect 7746 7792 7802 7848
rect 7194 1672 7250 1728
rect 7378 2488 7434 2544
rect 8850 7692 8852 7712
rect 8852 7692 8904 7712
rect 8904 7692 8906 7712
rect 8850 7656 8906 7692
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 9402 7520 9458 7576
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 8758 6296 8814 6352
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 8482 5616 8538 5672
rect 9402 6160 9458 6216
rect 8850 5752 8906 5808
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 14830 7520 14886 7576
rect 12346 7248 12402 7304
rect 13266 7248 13322 7304
rect 14830 7248 14886 7304
rect 11058 2488 11114 2544
rect 11610 2896 11666 2952
rect 11702 2352 11758 2408
rect 11426 1944 11482 2000
rect 12898 2352 12954 2408
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 13450 4664 13506 4720
rect 13266 3032 13322 3088
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 14922 3576 14978 3632
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 15842 3168 15898 3224
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 16946 5888 17002 5944
rect 16946 5616 17002 5672
rect 20902 9016 20958 9072
rect 20718 8336 20774 8392
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 18786 7284 18788 7304
rect 18788 7284 18840 7304
rect 18840 7284 18842 7304
rect 18786 7248 18842 7284
rect 17222 6296 17278 6352
rect 17774 6296 17830 6352
rect 17222 5616 17278 5672
rect 16486 3440 16542 3496
rect 16670 2896 16726 2952
rect 16394 448 16450 504
rect 17866 3032 17922 3088
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 19062 5344 19118 5400
rect 19522 5208 19578 5264
rect 19798 5072 19854 5128
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 20166 3612 20168 3632
rect 20168 3612 20220 3632
rect 20220 3612 20222 3632
rect 19890 3440 19946 3496
rect 20166 3576 20222 3612
rect 18694 1944 18750 2000
rect 18878 1944 18934 2000
rect 17498 176 17554 232
rect 17406 40 17462 96
rect 18326 584 18382 640
rect 18602 312 18658 368
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 20442 3168 20498 3224
rect 20442 2760 20498 2816
rect 23662 7928 23718 7984
rect 23478 7384 23534 7440
rect 20902 6840 20958 6896
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 21454 5752 21510 5808
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 21638 5788 21640 5808
rect 21640 5788 21692 5808
rect 21692 5788 21694 5808
rect 21638 5752 21694 5788
rect 24950 6724 25006 6760
rect 24950 6704 24952 6724
rect 24952 6704 25004 6724
rect 25004 6704 25006 6724
rect 21638 3032 21694 3088
rect 21638 2760 21694 2816
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 23386 4528 23442 4584
rect 21822 1672 21878 1728
rect 23478 4120 23534 4176
rect 23386 2388 23388 2408
rect 23388 2388 23440 2408
rect 23440 2388 23442 2408
rect 23386 2352 23442 2388
rect 24766 3984 24822 4040
rect 24490 2624 24546 2680
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 26330 8472 26386 8528
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 25318 2624 25374 2680
rect 26330 3984 26386 4040
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 26238 3032 26294 3088
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 25962 2488 26018 2544
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 26882 7248 26938 7304
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 27342 5616 27398 5672
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 29550 7828 29552 7848
rect 29552 7828 29604 7848
rect 29604 7828 29606 7848
rect 29550 7792 29606 7828
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 28998 2916 29054 2952
rect 28998 2896 29000 2916
rect 29000 2896 29052 2916
rect 29052 2896 29054 2916
rect 29642 5616 29698 5672
rect 30286 5208 30342 5264
rect 30378 2896 30434 2952
rect 30102 448 30158 504
rect 31114 1944 31170 2000
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 39016 8730 39072 8732
rect 39096 8730 39152 8732
rect 39176 8730 39232 8732
rect 39256 8730 39312 8732
rect 39016 8678 39062 8730
rect 39062 8678 39072 8730
rect 39096 8678 39126 8730
rect 39126 8678 39138 8730
rect 39138 8678 39152 8730
rect 39176 8678 39190 8730
rect 39190 8678 39202 8730
rect 39202 8678 39232 8730
rect 39256 8678 39266 8730
rect 39266 8678 39312 8730
rect 39016 8676 39072 8678
rect 39096 8676 39152 8678
rect 39176 8676 39232 8678
rect 39256 8676 39312 8678
rect 41970 9832 42026 9888
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 34150 6160 34206 6216
rect 33966 5616 34022 5672
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 31206 584 31262 640
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 32126 2352 32182 2408
rect 32678 1400 32734 1456
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 34058 4664 34114 4720
rect 33138 2352 33194 2408
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
rect 33598 1400 33654 1456
rect 33690 312 33746 368
rect 34610 1672 34666 1728
rect 35162 2896 35218 2952
rect 34794 176 34850 232
rect 34886 40 34942 96
rect 35714 3052 35770 3088
rect 35714 3032 35716 3052
rect 35716 3032 35768 3052
rect 35768 3032 35770 3052
rect 37956 8186 38012 8188
rect 38036 8186 38092 8188
rect 38116 8186 38172 8188
rect 38196 8186 38252 8188
rect 37956 8134 38002 8186
rect 38002 8134 38012 8186
rect 38036 8134 38066 8186
rect 38066 8134 38078 8186
rect 38078 8134 38092 8186
rect 38116 8134 38130 8186
rect 38130 8134 38142 8186
rect 38142 8134 38172 8186
rect 38196 8134 38206 8186
rect 38206 8134 38252 8186
rect 37956 8132 38012 8134
rect 38036 8132 38092 8134
rect 38116 8132 38172 8134
rect 38196 8132 38252 8134
rect 39016 7642 39072 7644
rect 39096 7642 39152 7644
rect 39176 7642 39232 7644
rect 39256 7642 39312 7644
rect 39016 7590 39062 7642
rect 39062 7590 39072 7642
rect 39096 7590 39126 7642
rect 39126 7590 39138 7642
rect 39138 7590 39152 7642
rect 39176 7590 39190 7642
rect 39190 7590 39202 7642
rect 39202 7590 39232 7642
rect 39256 7590 39266 7642
rect 39266 7590 39312 7642
rect 39016 7588 39072 7590
rect 39096 7588 39152 7590
rect 39176 7588 39232 7590
rect 39256 7588 39312 7590
rect 37956 7098 38012 7100
rect 38036 7098 38092 7100
rect 38116 7098 38172 7100
rect 38196 7098 38252 7100
rect 37956 7046 38002 7098
rect 38002 7046 38012 7098
rect 38036 7046 38066 7098
rect 38066 7046 38078 7098
rect 38078 7046 38092 7098
rect 38116 7046 38130 7098
rect 38130 7046 38142 7098
rect 38142 7046 38172 7098
rect 38196 7046 38206 7098
rect 38206 7046 38252 7098
rect 37956 7044 38012 7046
rect 38036 7044 38092 7046
rect 38116 7044 38172 7046
rect 38196 7044 38252 7046
rect 37956 6010 38012 6012
rect 38036 6010 38092 6012
rect 38116 6010 38172 6012
rect 38196 6010 38252 6012
rect 37956 5958 38002 6010
rect 38002 5958 38012 6010
rect 38036 5958 38066 6010
rect 38066 5958 38078 6010
rect 38078 5958 38092 6010
rect 38116 5958 38130 6010
rect 38130 5958 38142 6010
rect 38142 5958 38172 6010
rect 38196 5958 38206 6010
rect 38206 5958 38252 6010
rect 37956 5956 38012 5958
rect 38036 5956 38092 5958
rect 38116 5956 38172 5958
rect 38196 5956 38252 5958
rect 37956 4922 38012 4924
rect 38036 4922 38092 4924
rect 38116 4922 38172 4924
rect 38196 4922 38252 4924
rect 37956 4870 38002 4922
rect 38002 4870 38012 4922
rect 38036 4870 38066 4922
rect 38066 4870 38078 4922
rect 38078 4870 38092 4922
rect 38116 4870 38130 4922
rect 38130 4870 38142 4922
rect 38142 4870 38172 4922
rect 38196 4870 38206 4922
rect 38206 4870 38252 4922
rect 37956 4868 38012 4870
rect 38036 4868 38092 4870
rect 38116 4868 38172 4870
rect 38196 4868 38252 4870
rect 37956 3834 38012 3836
rect 38036 3834 38092 3836
rect 38116 3834 38172 3836
rect 38196 3834 38252 3836
rect 37956 3782 38002 3834
rect 38002 3782 38012 3834
rect 38036 3782 38066 3834
rect 38066 3782 38078 3834
rect 38078 3782 38092 3834
rect 38116 3782 38130 3834
rect 38130 3782 38142 3834
rect 38142 3782 38172 3834
rect 38196 3782 38206 3834
rect 38206 3782 38252 3834
rect 37956 3780 38012 3782
rect 38036 3780 38092 3782
rect 38116 3780 38172 3782
rect 38196 3780 38252 3782
rect 37956 2746 38012 2748
rect 38036 2746 38092 2748
rect 38116 2746 38172 2748
rect 38196 2746 38252 2748
rect 37956 2694 38002 2746
rect 38002 2694 38012 2746
rect 38036 2694 38066 2746
rect 38066 2694 38078 2746
rect 38078 2694 38092 2746
rect 38116 2694 38130 2746
rect 38130 2694 38142 2746
rect 38142 2694 38172 2746
rect 38196 2694 38206 2746
rect 38206 2694 38252 2746
rect 37956 2692 38012 2694
rect 38036 2692 38092 2694
rect 38116 2692 38172 2694
rect 38196 2692 38252 2694
rect 39016 6554 39072 6556
rect 39096 6554 39152 6556
rect 39176 6554 39232 6556
rect 39256 6554 39312 6556
rect 39016 6502 39062 6554
rect 39062 6502 39072 6554
rect 39096 6502 39126 6554
rect 39126 6502 39138 6554
rect 39138 6502 39152 6554
rect 39176 6502 39190 6554
rect 39190 6502 39202 6554
rect 39202 6502 39232 6554
rect 39256 6502 39266 6554
rect 39266 6502 39312 6554
rect 39016 6500 39072 6502
rect 39096 6500 39152 6502
rect 39176 6500 39232 6502
rect 39256 6500 39312 6502
rect 38658 3576 38714 3632
rect 39016 5466 39072 5468
rect 39096 5466 39152 5468
rect 39176 5466 39232 5468
rect 39256 5466 39312 5468
rect 39016 5414 39062 5466
rect 39062 5414 39072 5466
rect 39096 5414 39126 5466
rect 39126 5414 39138 5466
rect 39138 5414 39152 5466
rect 39176 5414 39190 5466
rect 39190 5414 39202 5466
rect 39202 5414 39232 5466
rect 39256 5414 39266 5466
rect 39266 5414 39312 5466
rect 39016 5412 39072 5414
rect 39096 5412 39152 5414
rect 39176 5412 39232 5414
rect 39256 5412 39312 5414
rect 39016 4378 39072 4380
rect 39096 4378 39152 4380
rect 39176 4378 39232 4380
rect 39256 4378 39312 4380
rect 39016 4326 39062 4378
rect 39062 4326 39072 4378
rect 39096 4326 39126 4378
rect 39126 4326 39138 4378
rect 39138 4326 39152 4378
rect 39176 4326 39190 4378
rect 39190 4326 39202 4378
rect 39202 4326 39232 4378
rect 39256 4326 39266 4378
rect 39266 4326 39312 4378
rect 39016 4324 39072 4326
rect 39096 4324 39152 4326
rect 39176 4324 39232 4326
rect 39256 4324 39312 4326
rect 39016 3290 39072 3292
rect 39096 3290 39152 3292
rect 39176 3290 39232 3292
rect 39256 3290 39312 3292
rect 39016 3238 39062 3290
rect 39062 3238 39072 3290
rect 39096 3238 39126 3290
rect 39126 3238 39138 3290
rect 39138 3238 39152 3290
rect 39176 3238 39190 3290
rect 39190 3238 39202 3290
rect 39202 3238 39232 3290
rect 39256 3238 39266 3290
rect 39266 3238 39312 3290
rect 39016 3236 39072 3238
rect 39096 3236 39152 3238
rect 39176 3236 39232 3238
rect 39256 3236 39312 3238
rect 39016 2202 39072 2204
rect 39096 2202 39152 2204
rect 39176 2202 39232 2204
rect 39256 2202 39312 2204
rect 39016 2150 39062 2202
rect 39062 2150 39072 2202
rect 39096 2150 39126 2202
rect 39126 2150 39138 2202
rect 39138 2150 39152 2202
rect 39176 2150 39190 2202
rect 39190 2150 39202 2202
rect 39202 2150 39232 2202
rect 39256 2150 39266 2202
rect 39266 2150 39312 2202
rect 39016 2148 39072 2150
rect 39096 2148 39152 2150
rect 39176 2148 39232 2150
rect 39256 2148 39312 2150
rect 42338 9560 42394 9616
rect 42154 8744 42210 8800
rect 43166 9288 43222 9344
rect 42614 9016 42670 9072
rect 42706 8472 42762 8528
rect 43074 8200 43130 8256
rect 43442 7928 43498 7984
rect 43074 7384 43130 7440
rect 43442 7692 43444 7712
rect 43444 7692 43496 7712
rect 43496 7692 43498 7712
rect 43442 7656 43498 7692
rect 43442 7148 43444 7168
rect 43444 7148 43496 7168
rect 43496 7148 43498 7168
rect 43442 7112 43498 7148
rect 43442 6840 43498 6896
rect 43074 6604 43076 6624
rect 43076 6604 43128 6624
rect 43128 6604 43130 6624
rect 43074 6568 43130 6604
rect 43074 6060 43076 6080
rect 43076 6060 43128 6080
rect 43128 6060 43130 6080
rect 43074 6024 43130 6060
rect 43074 5516 43076 5536
rect 43076 5516 43128 5536
rect 43128 5516 43130 5536
rect 43074 5480 43130 5516
rect 43074 4972 43076 4992
rect 43076 4972 43128 4992
rect 43128 4972 43130 4992
rect 43074 4936 43130 4972
rect 42798 3984 42854 4040
rect 43074 4428 43076 4448
rect 43076 4428 43128 4448
rect 43128 4428 43130 4448
rect 43074 4392 43130 4428
rect 43074 3884 43076 3904
rect 43076 3884 43128 3904
rect 43128 3884 43130 3904
rect 43074 3848 43130 3884
rect 43074 3340 43076 3360
rect 43076 3340 43128 3360
rect 43128 3340 43130 3360
rect 43074 3304 43130 3340
rect 43258 6316 43314 6352
rect 43258 6296 43260 6316
rect 43260 6296 43312 6316
rect 43312 6296 43314 6316
rect 43442 6296 43498 6352
rect 43442 5788 43444 5808
rect 43444 5788 43496 5808
rect 43496 5788 43498 5808
rect 43442 5752 43498 5788
rect 43442 5208 43498 5264
rect 43442 4700 43444 4720
rect 43444 4700 43496 4720
rect 43496 4700 43498 4720
rect 43442 4664 43498 4700
rect 43442 4120 43498 4176
rect 43442 3612 43444 3632
rect 43444 3612 43496 3632
rect 43496 3612 43498 3632
rect 43442 3576 43498 3612
rect 43258 3440 43314 3496
rect 43442 3032 43498 3088
rect 43074 2796 43076 2816
rect 43076 2796 43128 2816
rect 43128 2796 43130 2816
rect 42522 2488 42578 2544
rect 42154 1672 42210 1728
rect 43074 2760 43130 2796
rect 43442 2524 43444 2544
rect 43444 2524 43496 2544
rect 43496 2524 43498 2544
rect 43442 2488 43498 2524
rect 43074 2252 43076 2272
rect 43076 2252 43128 2272
rect 43128 2252 43130 2272
rect 43074 2216 43130 2252
rect 42982 1944 43038 2000
rect 42706 1400 42762 1456
<< metal3 >>
rect 0 9890 120 9920
rect 1209 9890 1275 9893
rect 0 9888 1275 9890
rect 0 9832 1214 9888
rect 1270 9832 1275 9888
rect 0 9830 1275 9832
rect 0 9800 120 9830
rect 1209 9827 1275 9830
rect 41965 9890 42031 9893
rect 44880 9890 45000 9920
rect 41965 9888 45000 9890
rect 41965 9832 41970 9888
rect 42026 9832 45000 9888
rect 41965 9830 45000 9832
rect 41965 9827 42031 9830
rect 44880 9800 45000 9830
rect 0 9618 120 9648
rect 19333 9618 19399 9621
rect 0 9616 19399 9618
rect 0 9560 19338 9616
rect 19394 9560 19399 9616
rect 0 9558 19399 9560
rect 0 9528 120 9558
rect 19333 9555 19399 9558
rect 42333 9618 42399 9621
rect 44880 9618 45000 9648
rect 42333 9616 45000 9618
rect 42333 9560 42338 9616
rect 42394 9560 45000 9616
rect 42333 9558 45000 9560
rect 42333 9555 42399 9558
rect 44880 9528 45000 9558
rect 0 9346 120 9376
rect 14917 9346 14983 9349
rect 0 9344 14983 9346
rect 0 9288 14922 9344
rect 14978 9288 14983 9344
rect 0 9286 14983 9288
rect 0 9256 120 9286
rect 14917 9283 14983 9286
rect 43161 9346 43227 9349
rect 44880 9346 45000 9376
rect 43161 9344 45000 9346
rect 43161 9288 43166 9344
rect 43222 9288 45000 9344
rect 43161 9286 45000 9288
rect 43161 9283 43227 9286
rect 44880 9256 45000 9286
rect 0 9074 120 9104
rect 20897 9074 20963 9077
rect 0 9072 20963 9074
rect 0 9016 20902 9072
rect 20958 9016 20963 9072
rect 0 9014 20963 9016
rect 0 8984 120 9014
rect 20897 9011 20963 9014
rect 42609 9074 42675 9077
rect 44880 9074 45000 9104
rect 42609 9072 45000 9074
rect 42609 9016 42614 9072
rect 42670 9016 45000 9072
rect 42609 9014 45000 9016
rect 42609 9011 42675 9014
rect 44880 8984 45000 9014
rect 0 8802 120 8832
rect 2865 8802 2931 8805
rect 0 8800 2931 8802
rect 0 8744 2870 8800
rect 2926 8744 2931 8800
rect 0 8742 2931 8744
rect 0 8712 120 8742
rect 2865 8739 2931 8742
rect 42149 8802 42215 8805
rect 44880 8802 45000 8832
rect 42149 8800 45000 8802
rect 42149 8744 42154 8800
rect 42210 8744 45000 8800
rect 42149 8742 45000 8744
rect 42149 8739 42215 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 33006 8671 33322 8672
rect 39006 8736 39322 8737
rect 39006 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39322 8736
rect 44880 8712 45000 8742
rect 39006 8671 39322 8672
rect 0 8530 120 8560
rect 26325 8530 26391 8533
rect 0 8528 26391 8530
rect 0 8472 26330 8528
rect 26386 8472 26391 8528
rect 0 8470 26391 8472
rect 0 8440 120 8470
rect 26325 8467 26391 8470
rect 42701 8530 42767 8533
rect 44880 8530 45000 8560
rect 42701 8528 45000 8530
rect 42701 8472 42706 8528
rect 42762 8472 45000 8528
rect 42701 8470 45000 8472
rect 42701 8467 42767 8470
rect 44880 8440 45000 8470
rect 1209 8394 1275 8397
rect 2865 8394 2931 8397
rect 20713 8394 20779 8397
rect 1209 8392 2514 8394
rect 1209 8336 1214 8392
rect 1270 8336 2514 8392
rect 1209 8334 2514 8336
rect 1209 8331 1275 8334
rect 0 8258 120 8288
rect 1761 8258 1827 8261
rect 0 8256 1827 8258
rect 0 8200 1766 8256
rect 1822 8200 1827 8256
rect 0 8198 1827 8200
rect 2454 8258 2514 8334
rect 2865 8392 20779 8394
rect 2865 8336 2870 8392
rect 2926 8336 20718 8392
rect 20774 8336 20779 8392
rect 2865 8334 20779 8336
rect 2865 8331 2931 8334
rect 20713 8331 20779 8334
rect 7741 8258 7807 8261
rect 2454 8256 7807 8258
rect 2454 8200 7746 8256
rect 7802 8200 7807 8256
rect 2454 8198 7807 8200
rect 0 8168 120 8198
rect 1761 8195 1827 8198
rect 7741 8195 7807 8198
rect 43069 8258 43135 8261
rect 44880 8258 45000 8288
rect 43069 8256 45000 8258
rect 43069 8200 43074 8256
rect 43130 8200 45000 8256
rect 43069 8198 45000 8200
rect 43069 8195 43135 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 37946 8192 38262 8193
rect 37946 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38262 8192
rect 44880 8168 45000 8198
rect 37946 8127 38262 8128
rect 0 7986 120 8016
rect 23657 7986 23723 7989
rect 0 7984 23723 7986
rect 0 7928 23662 7984
rect 23718 7928 23723 7984
rect 0 7926 23723 7928
rect 0 7896 120 7926
rect 23657 7923 23723 7926
rect 43437 7986 43503 7989
rect 44880 7986 45000 8016
rect 43437 7984 45000 7986
rect 43437 7928 43442 7984
rect 43498 7928 45000 7984
rect 43437 7926 45000 7928
rect 43437 7923 43503 7926
rect 44880 7896 45000 7926
rect 7741 7850 7807 7853
rect 29545 7850 29611 7853
rect 2822 7790 6930 7850
rect 0 7714 120 7744
rect 2822 7714 2882 7790
rect 0 7654 2882 7714
rect 6870 7714 6930 7790
rect 7741 7848 29611 7850
rect 7741 7792 7746 7848
rect 7802 7792 29550 7848
rect 29606 7792 29611 7848
rect 7741 7790 29611 7792
rect 7741 7787 7807 7790
rect 29545 7787 29611 7790
rect 8845 7714 8911 7717
rect 6870 7712 8911 7714
rect 6870 7656 8850 7712
rect 8906 7656 8911 7712
rect 6870 7654 8911 7656
rect 0 7624 120 7654
rect 8845 7651 8911 7654
rect 43437 7714 43503 7717
rect 44880 7714 45000 7744
rect 43437 7712 45000 7714
rect 43437 7656 43442 7712
rect 43498 7656 45000 7712
rect 43437 7654 45000 7656
rect 43437 7651 43503 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 33006 7583 33322 7584
rect 39006 7648 39322 7649
rect 39006 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39322 7648
rect 44880 7624 45000 7654
rect 39006 7583 39322 7584
rect 9397 7578 9463 7581
rect 14825 7578 14891 7581
rect 9397 7576 14891 7578
rect 9397 7520 9402 7576
rect 9458 7520 14830 7576
rect 14886 7520 14891 7576
rect 9397 7518 14891 7520
rect 9397 7515 9463 7518
rect 14825 7515 14891 7518
rect 0 7442 120 7472
rect 1301 7442 1367 7445
rect 0 7440 1367 7442
rect 0 7384 1306 7440
rect 1362 7384 1367 7440
rect 0 7382 1367 7384
rect 0 7352 120 7382
rect 1301 7379 1367 7382
rect 1761 7442 1827 7445
rect 23473 7442 23539 7445
rect 1761 7440 23539 7442
rect 1761 7384 1766 7440
rect 1822 7384 23478 7440
rect 23534 7384 23539 7440
rect 1761 7382 23539 7384
rect 1761 7379 1827 7382
rect 23473 7379 23539 7382
rect 43069 7442 43135 7445
rect 44880 7442 45000 7472
rect 43069 7440 45000 7442
rect 43069 7384 43074 7440
rect 43130 7384 45000 7440
rect 43069 7382 45000 7384
rect 43069 7379 43135 7382
rect 44880 7352 45000 7382
rect 12341 7306 12407 7309
rect 1718 7304 12407 7306
rect 1718 7248 12346 7304
rect 12402 7248 12407 7304
rect 1718 7246 12407 7248
rect 0 7170 120 7200
rect 1718 7170 1778 7246
rect 12341 7243 12407 7246
rect 13261 7306 13327 7309
rect 14825 7306 14891 7309
rect 18781 7306 18847 7309
rect 26877 7306 26943 7309
rect 13261 7304 14474 7306
rect 13261 7248 13266 7304
rect 13322 7248 14474 7304
rect 13261 7246 14474 7248
rect 13261 7243 13327 7246
rect 0 7110 1778 7170
rect 14414 7170 14474 7246
rect 14825 7304 18847 7306
rect 14825 7248 14830 7304
rect 14886 7248 18786 7304
rect 18842 7248 18847 7304
rect 14825 7246 18847 7248
rect 14825 7243 14891 7246
rect 18781 7243 18847 7246
rect 19014 7304 26943 7306
rect 19014 7248 26882 7304
rect 26938 7248 26943 7304
rect 19014 7246 26943 7248
rect 19014 7170 19074 7246
rect 26877 7243 26943 7246
rect 14414 7110 19074 7170
rect 43437 7170 43503 7173
rect 44880 7170 45000 7200
rect 43437 7168 45000 7170
rect 43437 7112 43442 7168
rect 43498 7112 45000 7168
rect 43437 7110 45000 7112
rect 0 7080 120 7110
rect 43437 7107 43503 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 37946 7104 38262 7105
rect 37946 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38262 7104
rect 44880 7080 45000 7110
rect 37946 7039 38262 7040
rect 0 6898 120 6928
rect 20897 6898 20963 6901
rect 0 6896 20963 6898
rect 0 6840 20902 6896
rect 20958 6840 20963 6896
rect 0 6838 20963 6840
rect 0 6808 120 6838
rect 20897 6835 20963 6838
rect 43437 6898 43503 6901
rect 44880 6898 45000 6928
rect 43437 6896 45000 6898
rect 43437 6840 43442 6896
rect 43498 6840 45000 6896
rect 43437 6838 45000 6840
rect 43437 6835 43503 6838
rect 44880 6808 45000 6838
rect 24945 6762 25011 6765
rect 2822 6760 25011 6762
rect 2822 6704 24950 6760
rect 25006 6704 25011 6760
rect 2822 6702 25011 6704
rect 0 6626 120 6656
rect 2822 6626 2882 6702
rect 24945 6699 25011 6702
rect 0 6566 2882 6626
rect 43069 6626 43135 6629
rect 44880 6626 45000 6656
rect 43069 6624 45000 6626
rect 43069 6568 43074 6624
rect 43130 6568 45000 6624
rect 43069 6566 45000 6568
rect 0 6536 120 6566
rect 43069 6563 43135 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 33006 6495 33322 6496
rect 39006 6560 39322 6561
rect 39006 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39322 6560
rect 44880 6536 45000 6566
rect 39006 6495 39322 6496
rect 0 6354 120 6384
rect 8753 6354 8819 6357
rect 17217 6354 17283 6357
rect 0 6352 8819 6354
rect 0 6296 8758 6352
rect 8814 6296 8819 6352
rect 0 6294 8819 6296
rect 0 6264 120 6294
rect 8753 6291 8819 6294
rect 9262 6352 17283 6354
rect 9262 6296 17222 6352
rect 17278 6296 17283 6352
rect 9262 6294 17283 6296
rect 9262 6218 9322 6294
rect 17217 6291 17283 6294
rect 17769 6354 17835 6357
rect 43253 6354 43319 6357
rect 17769 6352 43319 6354
rect 17769 6296 17774 6352
rect 17830 6296 43258 6352
rect 43314 6296 43319 6352
rect 17769 6294 43319 6296
rect 17769 6291 17835 6294
rect 43253 6291 43319 6294
rect 43437 6354 43503 6357
rect 44880 6354 45000 6384
rect 43437 6352 45000 6354
rect 43437 6296 43442 6352
rect 43498 6296 45000 6352
rect 43437 6294 45000 6296
rect 43437 6291 43503 6294
rect 44880 6264 45000 6294
rect 1718 6158 9322 6218
rect 9397 6218 9463 6221
rect 34145 6218 34211 6221
rect 9397 6216 34211 6218
rect 9397 6160 9402 6216
rect 9458 6160 34150 6216
rect 34206 6160 34211 6216
rect 9397 6158 34211 6160
rect 0 6082 120 6112
rect 1718 6082 1778 6158
rect 9397 6155 9463 6158
rect 34145 6155 34211 6158
rect 0 6022 1778 6082
rect 43069 6082 43135 6085
rect 44880 6082 45000 6112
rect 43069 6080 45000 6082
rect 43069 6024 43074 6080
rect 43130 6024 45000 6080
rect 43069 6022 45000 6024
rect 0 5992 120 6022
rect 43069 6019 43135 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 37946 6016 38262 6017
rect 37946 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38262 6016
rect 44880 5992 45000 6022
rect 37946 5951 38262 5952
rect 16941 5946 17007 5949
rect 16941 5944 17786 5946
rect 16941 5888 16946 5944
rect 17002 5888 17786 5944
rect 16941 5886 17786 5888
rect 16941 5883 17007 5886
rect 0 5810 120 5840
rect 8845 5810 8911 5813
rect 0 5808 8911 5810
rect 0 5752 8850 5808
rect 8906 5752 8911 5808
rect 0 5750 8911 5752
rect 17726 5810 17786 5886
rect 21449 5810 21515 5813
rect 17726 5808 21515 5810
rect 17726 5752 21454 5808
rect 21510 5752 21515 5808
rect 17726 5750 21515 5752
rect 0 5720 120 5750
rect 8845 5747 8911 5750
rect 21449 5747 21515 5750
rect 21633 5810 21699 5813
rect 34462 5810 34468 5812
rect 21633 5808 34468 5810
rect 21633 5752 21638 5808
rect 21694 5752 34468 5808
rect 21633 5750 34468 5752
rect 21633 5747 21699 5750
rect 34462 5748 34468 5750
rect 34532 5748 34538 5812
rect 43437 5810 43503 5813
rect 44880 5810 45000 5840
rect 43437 5808 45000 5810
rect 43437 5752 43442 5808
rect 43498 5752 45000 5808
rect 43437 5750 45000 5752
rect 43437 5747 43503 5750
rect 44880 5720 45000 5750
rect 8477 5674 8543 5677
rect 16941 5674 17007 5677
rect 8477 5672 17007 5674
rect 8477 5616 8482 5672
rect 8538 5616 16946 5672
rect 17002 5616 17007 5672
rect 8477 5614 17007 5616
rect 8477 5611 8543 5614
rect 16941 5611 17007 5614
rect 17217 5674 17283 5677
rect 27337 5674 27403 5677
rect 17217 5672 27403 5674
rect 17217 5616 17222 5672
rect 17278 5616 27342 5672
rect 27398 5616 27403 5672
rect 17217 5614 27403 5616
rect 17217 5611 17283 5614
rect 27337 5611 27403 5614
rect 29637 5674 29703 5677
rect 33961 5674 34027 5677
rect 29637 5672 34027 5674
rect 29637 5616 29642 5672
rect 29698 5616 33966 5672
rect 34022 5616 34027 5672
rect 29637 5614 34027 5616
rect 29637 5611 29703 5614
rect 33961 5611 34027 5614
rect 0 5538 120 5568
rect 2865 5538 2931 5541
rect 0 5536 2931 5538
rect 0 5480 2870 5536
rect 2926 5480 2931 5536
rect 0 5478 2931 5480
rect 0 5448 120 5478
rect 2865 5475 2931 5478
rect 43069 5538 43135 5541
rect 44880 5538 45000 5568
rect 43069 5536 45000 5538
rect 43069 5480 43074 5536
rect 43130 5480 45000 5536
rect 43069 5478 45000 5480
rect 43069 5475 43135 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 33006 5407 33322 5408
rect 39006 5472 39322 5473
rect 39006 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39322 5472
rect 44880 5448 45000 5478
rect 39006 5407 39322 5408
rect 19057 5402 19123 5405
rect 19057 5400 19810 5402
rect 19057 5344 19062 5400
rect 19118 5344 19810 5400
rect 19057 5342 19810 5344
rect 19057 5339 19123 5342
rect 0 5266 120 5296
rect 19517 5266 19583 5269
rect 0 5264 19583 5266
rect 0 5208 19522 5264
rect 19578 5208 19583 5264
rect 0 5206 19583 5208
rect 19750 5266 19810 5342
rect 30281 5266 30347 5269
rect 19750 5264 30347 5266
rect 19750 5208 30286 5264
rect 30342 5208 30347 5264
rect 19750 5206 30347 5208
rect 0 5176 120 5206
rect 19517 5203 19583 5206
rect 30281 5203 30347 5206
rect 43437 5266 43503 5269
rect 44880 5266 45000 5296
rect 43437 5264 45000 5266
rect 43437 5208 43442 5264
rect 43498 5208 45000 5264
rect 43437 5206 45000 5208
rect 43437 5203 43503 5206
rect 44880 5176 45000 5206
rect 2865 5130 2931 5133
rect 19793 5130 19859 5133
rect 2865 5128 19859 5130
rect 2865 5072 2870 5128
rect 2926 5072 19798 5128
rect 19854 5072 19859 5128
rect 2865 5070 19859 5072
rect 2865 5067 2931 5070
rect 19793 5067 19859 5070
rect 0 4994 120 5024
rect 1761 4994 1827 4997
rect 0 4992 1827 4994
rect 0 4936 1766 4992
rect 1822 4936 1827 4992
rect 0 4934 1827 4936
rect 0 4904 120 4934
rect 1761 4931 1827 4934
rect 43069 4994 43135 4997
rect 44880 4994 45000 5024
rect 43069 4992 45000 4994
rect 43069 4936 43074 4992
rect 43130 4936 45000 4992
rect 43069 4934 45000 4936
rect 43069 4931 43135 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 37946 4928 38262 4929
rect 37946 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38262 4928
rect 44880 4904 45000 4934
rect 37946 4863 38262 4864
rect 0 4722 120 4752
rect 13445 4722 13511 4725
rect 34053 4722 34119 4725
rect 0 4662 6930 4722
rect 0 4632 120 4662
rect 6870 4586 6930 4662
rect 13445 4720 34119 4722
rect 13445 4664 13450 4720
rect 13506 4664 34058 4720
rect 34114 4664 34119 4720
rect 13445 4662 34119 4664
rect 13445 4659 13511 4662
rect 34053 4659 34119 4662
rect 43437 4722 43503 4725
rect 44880 4722 45000 4752
rect 43437 4720 45000 4722
rect 43437 4664 43442 4720
rect 43498 4664 45000 4720
rect 43437 4662 45000 4664
rect 43437 4659 43503 4662
rect 44880 4632 45000 4662
rect 23381 4586 23447 4589
rect 6870 4584 23447 4586
rect 6870 4528 23386 4584
rect 23442 4528 23447 4584
rect 6870 4526 23447 4528
rect 23381 4523 23447 4526
rect 0 4450 120 4480
rect 1301 4450 1367 4453
rect 0 4448 1367 4450
rect 0 4392 1306 4448
rect 1362 4392 1367 4448
rect 0 4390 1367 4392
rect 0 4360 120 4390
rect 1301 4387 1367 4390
rect 43069 4450 43135 4453
rect 44880 4450 45000 4480
rect 43069 4448 45000 4450
rect 43069 4392 43074 4448
rect 43130 4392 45000 4448
rect 43069 4390 45000 4392
rect 43069 4387 43135 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 33006 4319 33322 4320
rect 39006 4384 39322 4385
rect 39006 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39322 4384
rect 44880 4360 45000 4390
rect 39006 4319 39322 4320
rect 0 4178 120 4208
rect 1209 4178 1275 4181
rect 0 4176 1275 4178
rect 0 4120 1214 4176
rect 1270 4120 1275 4176
rect 0 4118 1275 4120
rect 0 4088 120 4118
rect 1209 4115 1275 4118
rect 1761 4178 1827 4181
rect 23473 4178 23539 4181
rect 1761 4176 23539 4178
rect 1761 4120 1766 4176
rect 1822 4120 23478 4176
rect 23534 4120 23539 4176
rect 1761 4118 23539 4120
rect 1761 4115 1827 4118
rect 23473 4115 23539 4118
rect 43437 4178 43503 4181
rect 44880 4178 45000 4208
rect 43437 4176 45000 4178
rect 43437 4120 43442 4176
rect 43498 4120 45000 4176
rect 43437 4118 45000 4120
rect 43437 4115 43503 4118
rect 44880 4088 45000 4118
rect 2865 4042 2931 4045
rect 24761 4042 24827 4045
rect 2865 4040 24827 4042
rect 2865 3984 2870 4040
rect 2926 3984 24766 4040
rect 24822 3984 24827 4040
rect 2865 3982 24827 3984
rect 2865 3979 2931 3982
rect 24761 3979 24827 3982
rect 26325 4042 26391 4045
rect 42793 4042 42859 4045
rect 26325 4040 42859 4042
rect 26325 3984 26330 4040
rect 26386 3984 42798 4040
rect 42854 3984 42859 4040
rect 26325 3982 42859 3984
rect 26325 3979 26391 3982
rect 42793 3979 42859 3982
rect 0 3906 120 3936
rect 1761 3906 1827 3909
rect 0 3904 1827 3906
rect 0 3848 1766 3904
rect 1822 3848 1827 3904
rect 0 3846 1827 3848
rect 0 3816 120 3846
rect 1761 3843 1827 3846
rect 43069 3906 43135 3909
rect 44880 3906 45000 3936
rect 43069 3904 45000 3906
rect 43069 3848 43074 3904
rect 43130 3848 45000 3904
rect 43069 3846 45000 3848
rect 43069 3843 43135 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 37946 3840 38262 3841
rect 37946 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38262 3840
rect 44880 3816 45000 3846
rect 37946 3775 38262 3776
rect 0 3634 120 3664
rect 14917 3634 14983 3637
rect 0 3632 14983 3634
rect 0 3576 14922 3632
rect 14978 3576 14983 3632
rect 0 3574 14983 3576
rect 0 3544 120 3574
rect 14917 3571 14983 3574
rect 20161 3634 20227 3637
rect 38653 3634 38719 3637
rect 20161 3632 38719 3634
rect 20161 3576 20166 3632
rect 20222 3576 38658 3632
rect 38714 3576 38719 3632
rect 20161 3574 38719 3576
rect 20161 3571 20227 3574
rect 38653 3571 38719 3574
rect 43437 3634 43503 3637
rect 44880 3634 45000 3664
rect 43437 3632 45000 3634
rect 43437 3576 43442 3632
rect 43498 3576 45000 3632
rect 43437 3574 45000 3576
rect 43437 3571 43503 3574
rect 44880 3544 45000 3574
rect 1761 3498 1827 3501
rect 16481 3498 16547 3501
rect 1761 3496 16547 3498
rect 1761 3440 1766 3496
rect 1822 3440 16486 3496
rect 16542 3440 16547 3496
rect 1761 3438 16547 3440
rect 1761 3435 1827 3438
rect 16481 3435 16547 3438
rect 19885 3498 19951 3501
rect 43253 3498 43319 3501
rect 19885 3496 43319 3498
rect 19885 3440 19890 3496
rect 19946 3440 43258 3496
rect 43314 3440 43319 3496
rect 19885 3438 43319 3440
rect 19885 3435 19951 3438
rect 43253 3435 43319 3438
rect 0 3362 120 3392
rect 2865 3362 2931 3365
rect 0 3360 2931 3362
rect 0 3304 2870 3360
rect 2926 3304 2931 3360
rect 0 3302 2931 3304
rect 0 3272 120 3302
rect 2865 3299 2931 3302
rect 43069 3362 43135 3365
rect 44880 3362 45000 3392
rect 43069 3360 45000 3362
rect 43069 3304 43074 3360
rect 43130 3304 45000 3360
rect 43069 3302 45000 3304
rect 43069 3299 43135 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 33006 3231 33322 3232
rect 39006 3296 39322 3297
rect 39006 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39322 3296
rect 44880 3272 45000 3302
rect 39006 3231 39322 3232
rect 15837 3226 15903 3229
rect 20437 3226 20503 3229
rect 15837 3224 20503 3226
rect 15837 3168 15842 3224
rect 15898 3168 20442 3224
rect 20498 3168 20503 3224
rect 15837 3166 20503 3168
rect 15837 3163 15903 3166
rect 20437 3163 20503 3166
rect 21406 3166 26802 3226
rect 0 3090 120 3120
rect 13261 3090 13327 3093
rect 0 3088 13327 3090
rect 0 3032 13266 3088
rect 13322 3032 13327 3088
rect 0 3030 13327 3032
rect 0 3000 120 3030
rect 13261 3027 13327 3030
rect 17861 3090 17927 3093
rect 21406 3090 21466 3166
rect 17861 3088 21466 3090
rect 17861 3032 17866 3088
rect 17922 3032 21466 3088
rect 17861 3030 21466 3032
rect 21633 3090 21699 3093
rect 26233 3090 26299 3093
rect 21633 3088 26299 3090
rect 21633 3032 21638 3088
rect 21694 3032 26238 3088
rect 26294 3032 26299 3088
rect 21633 3030 26299 3032
rect 26742 3090 26802 3166
rect 35709 3090 35775 3093
rect 26742 3088 35775 3090
rect 26742 3032 35714 3088
rect 35770 3032 35775 3088
rect 26742 3030 35775 3032
rect 17861 3027 17927 3030
rect 21633 3027 21699 3030
rect 26233 3027 26299 3030
rect 35709 3027 35775 3030
rect 43437 3090 43503 3093
rect 44880 3090 45000 3120
rect 43437 3088 45000 3090
rect 43437 3032 43442 3088
rect 43498 3032 45000 3088
rect 43437 3030 45000 3032
rect 43437 3027 43503 3030
rect 44880 3000 45000 3030
rect 11605 2954 11671 2957
rect 1718 2952 11671 2954
rect 1718 2896 11610 2952
rect 11666 2896 11671 2952
rect 1718 2894 11671 2896
rect 0 2818 120 2848
rect 1718 2818 1778 2894
rect 11605 2891 11671 2894
rect 16665 2954 16731 2957
rect 28993 2954 29059 2957
rect 16665 2952 29059 2954
rect 16665 2896 16670 2952
rect 16726 2896 28998 2952
rect 29054 2896 29059 2952
rect 16665 2894 29059 2896
rect 16665 2891 16731 2894
rect 28993 2891 29059 2894
rect 30373 2954 30439 2957
rect 35157 2954 35223 2957
rect 30373 2952 35223 2954
rect 30373 2896 30378 2952
rect 30434 2896 35162 2952
rect 35218 2896 35223 2952
rect 30373 2894 35223 2896
rect 30373 2891 30439 2894
rect 35157 2891 35223 2894
rect 0 2758 1778 2818
rect 20437 2818 20503 2821
rect 21633 2818 21699 2821
rect 20437 2816 21699 2818
rect 20437 2760 20442 2816
rect 20498 2760 21638 2816
rect 21694 2760 21699 2816
rect 20437 2758 21699 2760
rect 0 2728 120 2758
rect 20437 2755 20503 2758
rect 21633 2755 21699 2758
rect 43069 2818 43135 2821
rect 44880 2818 45000 2848
rect 43069 2816 45000 2818
rect 43069 2760 43074 2816
rect 43130 2760 45000 2816
rect 43069 2758 45000 2760
rect 43069 2755 43135 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 37946 2752 38262 2753
rect 37946 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38262 2752
rect 44880 2728 45000 2758
rect 37946 2687 38262 2688
rect 24485 2682 24551 2685
rect 25313 2682 25379 2685
rect 24485 2680 25379 2682
rect 24485 2624 24490 2680
rect 24546 2624 25318 2680
rect 25374 2624 25379 2680
rect 24485 2622 25379 2624
rect 24485 2619 24551 2622
rect 25313 2619 25379 2622
rect 0 2546 120 2576
rect 7373 2546 7439 2549
rect 0 2544 7439 2546
rect 0 2488 7378 2544
rect 7434 2488 7439 2544
rect 0 2486 7439 2488
rect 0 2456 120 2486
rect 7373 2483 7439 2486
rect 11053 2546 11119 2549
rect 25957 2546 26023 2549
rect 11053 2544 26023 2546
rect 11053 2488 11058 2544
rect 11114 2488 25962 2544
rect 26018 2488 26023 2544
rect 11053 2486 26023 2488
rect 11053 2483 11119 2486
rect 25957 2483 26023 2486
rect 34462 2484 34468 2548
rect 34532 2546 34538 2548
rect 42517 2546 42583 2549
rect 34532 2544 42583 2546
rect 34532 2488 42522 2544
rect 42578 2488 42583 2544
rect 34532 2486 42583 2488
rect 34532 2484 34538 2486
rect 42517 2483 42583 2486
rect 43437 2546 43503 2549
rect 44880 2546 45000 2576
rect 43437 2544 45000 2546
rect 43437 2488 43442 2544
rect 43498 2488 45000 2544
rect 43437 2486 45000 2488
rect 43437 2483 43503 2486
rect 44880 2456 45000 2486
rect 11697 2410 11763 2413
rect 2822 2408 11763 2410
rect 2822 2352 11702 2408
rect 11758 2352 11763 2408
rect 2822 2350 11763 2352
rect 0 2274 120 2304
rect 2822 2274 2882 2350
rect 11697 2347 11763 2350
rect 12893 2410 12959 2413
rect 23381 2410 23447 2413
rect 12893 2408 23447 2410
rect 12893 2352 12898 2408
rect 12954 2352 23386 2408
rect 23442 2352 23447 2408
rect 12893 2350 23447 2352
rect 12893 2347 12959 2350
rect 23381 2347 23447 2350
rect 32121 2410 32187 2413
rect 33133 2410 33199 2413
rect 32121 2408 33199 2410
rect 32121 2352 32126 2408
rect 32182 2352 33138 2408
rect 33194 2352 33199 2408
rect 32121 2350 33199 2352
rect 32121 2347 32187 2350
rect 33133 2347 33199 2350
rect 0 2214 2882 2274
rect 43069 2274 43135 2277
rect 44880 2274 45000 2304
rect 43069 2272 45000 2274
rect 43069 2216 43074 2272
rect 43130 2216 45000 2272
rect 43069 2214 45000 2216
rect 0 2184 120 2214
rect 43069 2211 43135 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 33006 2143 33322 2144
rect 39006 2208 39322 2209
rect 39006 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39322 2208
rect 44880 2184 45000 2214
rect 39006 2143 39322 2144
rect 0 2002 120 2032
rect 5533 2002 5599 2005
rect 0 2000 5599 2002
rect 0 1944 5538 2000
rect 5594 1944 5599 2000
rect 0 1942 5599 1944
rect 0 1912 120 1942
rect 5533 1939 5599 1942
rect 11421 2002 11487 2005
rect 18689 2002 18755 2005
rect 11421 2000 18755 2002
rect 11421 1944 11426 2000
rect 11482 1944 18694 2000
rect 18750 1944 18755 2000
rect 11421 1942 18755 1944
rect 11421 1939 11487 1942
rect 18689 1939 18755 1942
rect 18873 2002 18939 2005
rect 31109 2002 31175 2005
rect 18873 2000 31175 2002
rect 18873 1944 18878 2000
rect 18934 1944 31114 2000
rect 31170 1944 31175 2000
rect 18873 1942 31175 1944
rect 18873 1939 18939 1942
rect 31109 1939 31175 1942
rect 42977 2002 43043 2005
rect 44880 2002 45000 2032
rect 42977 2000 45000 2002
rect 42977 1944 42982 2000
rect 43038 1944 45000 2000
rect 42977 1942 45000 1944
rect 42977 1939 43043 1942
rect 44880 1912 45000 1942
rect 0 1730 120 1760
rect 7189 1730 7255 1733
rect 0 1728 7255 1730
rect 0 1672 7194 1728
rect 7250 1672 7255 1728
rect 0 1670 7255 1672
rect 0 1640 120 1670
rect 7189 1667 7255 1670
rect 21817 1730 21883 1733
rect 34605 1730 34671 1733
rect 21817 1728 34671 1730
rect 21817 1672 21822 1728
rect 21878 1672 34610 1728
rect 34666 1672 34671 1728
rect 21817 1670 34671 1672
rect 21817 1667 21883 1670
rect 34605 1667 34671 1670
rect 42149 1730 42215 1733
rect 44880 1730 45000 1760
rect 42149 1728 45000 1730
rect 42149 1672 42154 1728
rect 42210 1672 45000 1728
rect 42149 1670 45000 1672
rect 42149 1667 42215 1670
rect 44880 1640 45000 1670
rect 0 1458 120 1488
rect 933 1458 999 1461
rect 0 1456 999 1458
rect 0 1400 938 1456
rect 994 1400 999 1456
rect 0 1398 999 1400
rect 0 1368 120 1398
rect 933 1395 999 1398
rect 32673 1458 32739 1461
rect 33593 1458 33659 1461
rect 32673 1456 33659 1458
rect 32673 1400 32678 1456
rect 32734 1400 33598 1456
rect 33654 1400 33659 1456
rect 32673 1398 33659 1400
rect 32673 1395 32739 1398
rect 33593 1395 33659 1398
rect 42701 1458 42767 1461
rect 44880 1458 45000 1488
rect 42701 1456 45000 1458
rect 42701 1400 42706 1456
rect 42762 1400 45000 1456
rect 42701 1398 45000 1400
rect 42701 1395 42767 1398
rect 44880 1368 45000 1398
rect 18321 642 18387 645
rect 31201 642 31267 645
rect 18321 640 31267 642
rect 18321 584 18326 640
rect 18382 584 31206 640
rect 31262 584 31267 640
rect 18321 582 31267 584
rect 18321 579 18387 582
rect 31201 579 31267 582
rect 16389 506 16455 509
rect 30097 506 30163 509
rect 16389 504 30163 506
rect 16389 448 16394 504
rect 16450 448 30102 504
rect 30158 448 30163 504
rect 16389 446 30163 448
rect 16389 443 16455 446
rect 30097 443 30163 446
rect 18597 370 18663 373
rect 33685 370 33751 373
rect 18597 368 33751 370
rect 18597 312 18602 368
rect 18658 312 33690 368
rect 33746 312 33751 368
rect 18597 310 33751 312
rect 18597 307 18663 310
rect 33685 307 33751 310
rect 17493 234 17559 237
rect 34789 234 34855 237
rect 17493 232 34855 234
rect 17493 176 17498 232
rect 17554 176 34794 232
rect 34850 176 34855 232
rect 17493 174 34855 176
rect 17493 171 17559 174
rect 34789 171 34855 174
rect 17401 98 17467 101
rect 34881 98 34947 101
rect 17401 96 34947 98
rect 17401 40 17406 96
rect 17462 40 34886 96
rect 34942 40 34947 96
rect 17401 38 34947 40
rect 17401 35 17467 38
rect 34881 35 34947 38
<< via3 >>
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 39012 8732 39076 8736
rect 39012 8676 39016 8732
rect 39016 8676 39072 8732
rect 39072 8676 39076 8732
rect 39012 8672 39076 8676
rect 39092 8732 39156 8736
rect 39092 8676 39096 8732
rect 39096 8676 39152 8732
rect 39152 8676 39156 8732
rect 39092 8672 39156 8676
rect 39172 8732 39236 8736
rect 39172 8676 39176 8732
rect 39176 8676 39232 8732
rect 39232 8676 39236 8732
rect 39172 8672 39236 8676
rect 39252 8732 39316 8736
rect 39252 8676 39256 8732
rect 39256 8676 39312 8732
rect 39312 8676 39316 8732
rect 39252 8672 39316 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 37952 8188 38016 8192
rect 37952 8132 37956 8188
rect 37956 8132 38012 8188
rect 38012 8132 38016 8188
rect 37952 8128 38016 8132
rect 38032 8188 38096 8192
rect 38032 8132 38036 8188
rect 38036 8132 38092 8188
rect 38092 8132 38096 8188
rect 38032 8128 38096 8132
rect 38112 8188 38176 8192
rect 38112 8132 38116 8188
rect 38116 8132 38172 8188
rect 38172 8132 38176 8188
rect 38112 8128 38176 8132
rect 38192 8188 38256 8192
rect 38192 8132 38196 8188
rect 38196 8132 38252 8188
rect 38252 8132 38256 8188
rect 38192 8128 38256 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 39012 7644 39076 7648
rect 39012 7588 39016 7644
rect 39016 7588 39072 7644
rect 39072 7588 39076 7644
rect 39012 7584 39076 7588
rect 39092 7644 39156 7648
rect 39092 7588 39096 7644
rect 39096 7588 39152 7644
rect 39152 7588 39156 7644
rect 39092 7584 39156 7588
rect 39172 7644 39236 7648
rect 39172 7588 39176 7644
rect 39176 7588 39232 7644
rect 39232 7588 39236 7644
rect 39172 7584 39236 7588
rect 39252 7644 39316 7648
rect 39252 7588 39256 7644
rect 39256 7588 39312 7644
rect 39312 7588 39316 7644
rect 39252 7584 39316 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 37952 7100 38016 7104
rect 37952 7044 37956 7100
rect 37956 7044 38012 7100
rect 38012 7044 38016 7100
rect 37952 7040 38016 7044
rect 38032 7100 38096 7104
rect 38032 7044 38036 7100
rect 38036 7044 38092 7100
rect 38092 7044 38096 7100
rect 38032 7040 38096 7044
rect 38112 7100 38176 7104
rect 38112 7044 38116 7100
rect 38116 7044 38172 7100
rect 38172 7044 38176 7100
rect 38112 7040 38176 7044
rect 38192 7100 38256 7104
rect 38192 7044 38196 7100
rect 38196 7044 38252 7100
rect 38252 7044 38256 7100
rect 38192 7040 38256 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 39012 6556 39076 6560
rect 39012 6500 39016 6556
rect 39016 6500 39072 6556
rect 39072 6500 39076 6556
rect 39012 6496 39076 6500
rect 39092 6556 39156 6560
rect 39092 6500 39096 6556
rect 39096 6500 39152 6556
rect 39152 6500 39156 6556
rect 39092 6496 39156 6500
rect 39172 6556 39236 6560
rect 39172 6500 39176 6556
rect 39176 6500 39232 6556
rect 39232 6500 39236 6556
rect 39172 6496 39236 6500
rect 39252 6556 39316 6560
rect 39252 6500 39256 6556
rect 39256 6500 39312 6556
rect 39312 6500 39316 6556
rect 39252 6496 39316 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 37952 6012 38016 6016
rect 37952 5956 37956 6012
rect 37956 5956 38012 6012
rect 38012 5956 38016 6012
rect 37952 5952 38016 5956
rect 38032 6012 38096 6016
rect 38032 5956 38036 6012
rect 38036 5956 38092 6012
rect 38092 5956 38096 6012
rect 38032 5952 38096 5956
rect 38112 6012 38176 6016
rect 38112 5956 38116 6012
rect 38116 5956 38172 6012
rect 38172 5956 38176 6012
rect 38112 5952 38176 5956
rect 38192 6012 38256 6016
rect 38192 5956 38196 6012
rect 38196 5956 38252 6012
rect 38252 5956 38256 6012
rect 38192 5952 38256 5956
rect 34468 5748 34532 5812
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 39012 5468 39076 5472
rect 39012 5412 39016 5468
rect 39016 5412 39072 5468
rect 39072 5412 39076 5468
rect 39012 5408 39076 5412
rect 39092 5468 39156 5472
rect 39092 5412 39096 5468
rect 39096 5412 39152 5468
rect 39152 5412 39156 5468
rect 39092 5408 39156 5412
rect 39172 5468 39236 5472
rect 39172 5412 39176 5468
rect 39176 5412 39232 5468
rect 39232 5412 39236 5468
rect 39172 5408 39236 5412
rect 39252 5468 39316 5472
rect 39252 5412 39256 5468
rect 39256 5412 39312 5468
rect 39312 5412 39316 5468
rect 39252 5408 39316 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 37952 4924 38016 4928
rect 37952 4868 37956 4924
rect 37956 4868 38012 4924
rect 38012 4868 38016 4924
rect 37952 4864 38016 4868
rect 38032 4924 38096 4928
rect 38032 4868 38036 4924
rect 38036 4868 38092 4924
rect 38092 4868 38096 4924
rect 38032 4864 38096 4868
rect 38112 4924 38176 4928
rect 38112 4868 38116 4924
rect 38116 4868 38172 4924
rect 38172 4868 38176 4924
rect 38112 4864 38176 4868
rect 38192 4924 38256 4928
rect 38192 4868 38196 4924
rect 38196 4868 38252 4924
rect 38252 4868 38256 4924
rect 38192 4864 38256 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 39012 4380 39076 4384
rect 39012 4324 39016 4380
rect 39016 4324 39072 4380
rect 39072 4324 39076 4380
rect 39012 4320 39076 4324
rect 39092 4380 39156 4384
rect 39092 4324 39096 4380
rect 39096 4324 39152 4380
rect 39152 4324 39156 4380
rect 39092 4320 39156 4324
rect 39172 4380 39236 4384
rect 39172 4324 39176 4380
rect 39176 4324 39232 4380
rect 39232 4324 39236 4380
rect 39172 4320 39236 4324
rect 39252 4380 39316 4384
rect 39252 4324 39256 4380
rect 39256 4324 39312 4380
rect 39312 4324 39316 4380
rect 39252 4320 39316 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 37952 3836 38016 3840
rect 37952 3780 37956 3836
rect 37956 3780 38012 3836
rect 38012 3780 38016 3836
rect 37952 3776 38016 3780
rect 38032 3836 38096 3840
rect 38032 3780 38036 3836
rect 38036 3780 38092 3836
rect 38092 3780 38096 3836
rect 38032 3776 38096 3780
rect 38112 3836 38176 3840
rect 38112 3780 38116 3836
rect 38116 3780 38172 3836
rect 38172 3780 38176 3836
rect 38112 3776 38176 3780
rect 38192 3836 38256 3840
rect 38192 3780 38196 3836
rect 38196 3780 38252 3836
rect 38252 3780 38256 3836
rect 38192 3776 38256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 39012 3292 39076 3296
rect 39012 3236 39016 3292
rect 39016 3236 39072 3292
rect 39072 3236 39076 3292
rect 39012 3232 39076 3236
rect 39092 3292 39156 3296
rect 39092 3236 39096 3292
rect 39096 3236 39152 3292
rect 39152 3236 39156 3292
rect 39092 3232 39156 3236
rect 39172 3292 39236 3296
rect 39172 3236 39176 3292
rect 39176 3236 39232 3292
rect 39232 3236 39236 3292
rect 39172 3232 39236 3236
rect 39252 3292 39316 3296
rect 39252 3236 39256 3292
rect 39256 3236 39312 3292
rect 39312 3236 39316 3292
rect 39252 3232 39316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 37952 2748 38016 2752
rect 37952 2692 37956 2748
rect 37956 2692 38012 2748
rect 38012 2692 38016 2748
rect 37952 2688 38016 2692
rect 38032 2748 38096 2752
rect 38032 2692 38036 2748
rect 38036 2692 38092 2748
rect 38092 2692 38096 2748
rect 38032 2688 38096 2692
rect 38112 2748 38176 2752
rect 38112 2692 38116 2748
rect 38116 2692 38172 2748
rect 38172 2692 38176 2748
rect 38112 2688 38176 2692
rect 38192 2748 38256 2752
rect 38192 2692 38196 2748
rect 38196 2692 38252 2748
rect 38252 2692 38256 2748
rect 38192 2688 38256 2692
rect 34468 2484 34532 2548
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
rect 39012 2204 39076 2208
rect 39012 2148 39016 2204
rect 39016 2148 39072 2204
rect 39072 2148 39076 2204
rect 39012 2144 39076 2148
rect 39092 2204 39156 2208
rect 39092 2148 39096 2204
rect 39096 2148 39152 2204
rect 39152 2148 39156 2204
rect 39092 2144 39156 2148
rect 39172 2204 39236 2208
rect 39172 2148 39176 2204
rect 39176 2148 39232 2204
rect 39232 2148 39236 2204
rect 39172 2144 39236 2148
rect 39252 2204 39316 2208
rect 39252 2148 39256 2204
rect 39256 2148 39312 2204
rect 39312 2148 39316 2204
rect 39252 2144 39316 2148
<< metal4 >>
rect 1944 8192 2264 11250
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 8736 3324 11250
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11250
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 8736 9324 11250
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 8192 14264 11250
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13944 0 14264 2688
rect 15004 8736 15324 11250
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 8192 20264 11250
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19944 0 20264 2688
rect 21004 8736 21324 11250
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 21004 6560 21324 7584
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25944 8192 26264 11250
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25944 0 26264 2688
rect 27004 8736 27324 11250
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 31944 8192 32264 11250
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 0 32264 2688
rect 33004 8736 33324 11250
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 37944 8192 38264 11250
rect 37944 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38264 8192
rect 37944 7104 38264 8128
rect 37944 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38264 7104
rect 37944 6016 38264 7040
rect 37944 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38264 6016
rect 34467 5812 34533 5813
rect 34467 5748 34468 5812
rect 34532 5748 34533 5812
rect 34467 5747 34533 5748
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 34470 2549 34530 5747
rect 37944 4928 38264 5952
rect 37944 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38264 4928
rect 37944 3840 38264 4864
rect 37944 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38264 3840
rect 37944 2752 38264 3776
rect 37944 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38264 2752
rect 34467 2548 34533 2549
rect 34467 2484 34468 2548
rect 34532 2484 34533 2548
rect 34467 2483 34533 2484
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
rect 37944 0 38264 2688
rect 39004 8736 39324 11250
rect 39004 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39324 8736
rect 39004 7648 39324 8672
rect 39004 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39324 7648
rect 39004 6560 39324 7584
rect 39004 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39324 6560
rect 39004 5472 39324 6496
rect 39004 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39324 5472
rect 39004 4384 39324 5408
rect 39004 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39324 4384
rect 39004 3296 39324 4320
rect 39004 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39324 3296
rect 39004 2208 39324 3232
rect 39004 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39324 2208
rect 39004 0 39324 2144
use sky130_fd_sc_hd__buf_1  _000_
timestamp -3599
transform 1 0 21436 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _001_
timestamp -3599
transform 1 0 25668 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _002_
timestamp -3599
transform 1 0 26496 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _003_
timestamp -3599
transform 1 0 26772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _004_
timestamp -3599
transform 1 0 23368 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _005_
timestamp -3599
transform 1 0 21988 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _006_
timestamp -3599
transform 1 0 27048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _007_
timestamp -3599
transform 1 0 28428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _008_
timestamp -3599
transform 1 0 29992 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _009_
timestamp -3599
transform 1 0 27140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _010_
timestamp -3599
transform 1 0 28336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _011_
timestamp -3599
transform 1 0 27232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _012_
timestamp -3599
transform 1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _013_
timestamp -3599
transform 1 0 23552 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _014_
timestamp -3599
transform 1 0 19688 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _015_
timestamp -3599
transform 1 0 19964 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _016_
timestamp -3599
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _017_
timestamp -3599
transform 1 0 27508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _018_
timestamp -3599
transform 1 0 17664 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _019_
timestamp -3599
transform 1 0 25116 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _020_
timestamp -3599
transform 1 0 21344 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _021_
timestamp -3599
transform 1 0 17848 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _022_
timestamp -3599
transform 1 0 26036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _023_
timestamp -3599
transform 1 0 18952 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _024_
timestamp -3599
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _025_
timestamp -3599
transform 1 0 23552 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _026_
timestamp -3599
transform 1 0 26496 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _027_
timestamp -3599
transform 1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _028_
timestamp -3599
transform 1 0 21160 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _029_
timestamp -3599
transform 1 0 17664 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _030_
timestamp -3599
transform 1 0 19320 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _031_
timestamp -3599
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _032_
timestamp -3599
transform 1 0 9200 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _033_
timestamp -3599
transform 1 0 9752 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _034_
timestamp -3599
transform -1 0 17480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _035_
timestamp -3599
transform -1 0 22080 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _036_
timestamp -3599
transform -1 0 32476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _037_
timestamp -3599
transform -1 0 30360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _038_
timestamp -3599
transform -1 0 26312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _039_
timestamp -3599
transform 1 0 25484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp -3599
transform 1 0 28152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp -3599
transform 1 0 31004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp -3599
transform 1 0 31188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp -3599
transform 1 0 30728 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp -3599
transform 1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp -3599
transform 1 0 33672 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp -3599
transform 1 0 36892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp -3599
transform -1 0 35144 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp -3599
transform 1 0 37720 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp -3599
transform -1 0 38548 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp -3599
transform -1 0 39376 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp -3599
transform -1 0 41400 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _052_
timestamp -3599
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _053_
timestamp -3599
transform 1 0 2300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _054_
timestamp -3599
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _055_
timestamp -3599
transform 1 0 1840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _056_
timestamp -3599
transform 1 0 4048 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _057_
timestamp -3599
transform 1 0 4140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _058_
timestamp -3599
transform 1 0 3956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _059_
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _060_
timestamp -3599
transform 1 0 5888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _061_
timestamp -3599
transform 1 0 6624 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _062_
timestamp -3599
transform 1 0 7268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _063_
timestamp -3599
transform 1 0 7544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _064_
timestamp -3599
transform 1 0 12880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp -3599
transform -1 0 12696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _066_
timestamp -3599
transform 1 0 9384 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp -3599
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp -3599
transform -1 0 15272 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp -3599
transform -1 0 15732 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp -3599
transform -1 0 16192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp -3599
transform -1 0 17572 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp -3599
transform -1 0 16560 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _073_
timestamp -3599
transform 1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp -3599
transform -1 0 22448 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp -3599
transform 1 0 27324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp -3599
transform 1 0 27324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _077_
timestamp -3599
transform 1 0 13708 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp -3599
transform -1 0 18400 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp -3599
transform -1 0 18952 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _080_
timestamp -3599
transform 1 0 15272 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _081_
timestamp -3599
transform 1 0 16100 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _082_
timestamp -3599
transform 1 0 15824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _083_
timestamp -3599
transform 1 0 18492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp -3599
transform -1 0 20608 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp -3599
transform -1 0 23092 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _086_
timestamp -3599
transform 1 0 20332 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _087_
timestamp -3599
transform 1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp -3599
transform 1 0 38088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp -3599
transform 1 0 37260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp -3599
transform 1 0 35328 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp -3599
transform 1 0 34960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp -3599
transform 1 0 33396 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp -3599
transform 1 0 36800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp -3599
transform 1 0 35880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp -3599
transform 1 0 34500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp -3599
transform 1 0 34224 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp -3599
transform -1 0 33028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp -3599
transform -1 0 32752 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp -3599
transform -1 0 31832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp -3599
transform -1 0 30636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp -3599
transform -1 0 30360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp -3599
transform -1 0 27968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp -3599
transform -1 0 24472 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp -3599
transform -1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform -1 0 27232 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform 1 0 24656 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform 1 0 23368 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform 1 0 19504 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform -1 0 20424 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform -1 0 22264 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 27508 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform -1 0 17664 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform -1 0 25116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform -1 0 21344 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform -1 0 17848 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform -1 0 18952 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform -1 0 24840 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform 1 0 23368 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform 1 0 26312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform 1 0 20700 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp -3599
transform -1 0 21620 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp -3599
transform 1 0 17480 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp -3599
transform -1 0 26496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp -3599
transform -1 0 19780 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp -3599
transform -1 0 29992 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp -3599
transform -1 0 27232 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp -3599
transform 1 0 23184 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp -3599
transform -1 0 27048 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp -3599
transform -1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp -3599
transform -1 0 29992 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp -3599
transform -1 0 27140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp -3599
transform -1 0 9200 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp -3599
transform -1 0 9752 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp -3599
transform -1 0 17204 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp -3599
transform 1 0 33212 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp -3599
transform -1 0 35328 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp -3599
transform -1 0 37720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp -3599
transform 1 0 30176 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp -3599
transform 1 0 31372 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp -3599
transform 1 0 32292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp -3599
transform -1 0 33212 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp -3599
transform 1 0 34040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp -3599
transform -1 0 34960 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp -3599
transform 1 0 35696 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636964856
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636964856
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636964856
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636964856
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636964856
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636964856
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636964856
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636964856
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -3599
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636964856
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636964856
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -3599
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636964856
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636964856
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -3599
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636964856
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636964856
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp -3599
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_197
timestamp -3599
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -3599
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -3599
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -3599
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_325
timestamp -3599
transform 1 0 31004 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp -3599
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp -3599
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_373
timestamp 1636964856
transform 1 0 35420 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp -3599
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp -3599
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1636964856
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1636964856
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp -3599
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1636964856
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_433
timestamp -3599
transform 1 0 40940 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_441
timestamp -3599
transform 1 0 41676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_449
timestamp -3599
transform 1 0 42412 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7
timestamp -3599
transform 1 0 1748 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_11
timestamp 1636964856
transform 1 0 2116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_23
timestamp 1636964856
transform 1 0 3220 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_35
timestamp 1636964856
transform 1 0 4324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47
timestamp -3599
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -3599
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636964856
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_69
timestamp -3599
transform 1 0 7452 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_73
timestamp 1636964856
transform 1 0 7820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_85
timestamp 1636964856
transform 1 0 8924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_97
timestamp 1636964856
transform 1 0 10028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp -3599
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp -3599
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_121
timestamp -3599
transform 1 0 12236 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_126
timestamp 1636964856
transform 1 0 12696 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_138
timestamp -3599
transform 1 0 13800 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636964856
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_164
timestamp -3599
transform 1 0 16192 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636964856
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636964856
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636964856
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_205
timestamp -3599
transform 1 0 19964 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_210
timestamp -3599
transform 1 0 20424 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp -3599
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp -3599
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_231
timestamp 1636964856
transform 1 0 22356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_243
timestamp 1636964856
transform 1 0 23460 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_255
timestamp -3599
transform 1 0 24564 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_267
timestamp -3599
transform 1 0 25668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_273
timestamp -3599
transform 1 0 26220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp -3599
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_281
timestamp -3599
transform 1 0 26956 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_291
timestamp -3599
transform 1 0 27876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_295
timestamp -3599
transform 1 0 28244 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_304
timestamp -3599
transform 1 0 29072 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_310
timestamp -3599
transform 1 0 29624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_315
timestamp -3599
transform 1 0 30084 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_321
timestamp -3599
transform 1 0 30636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_327
timestamp -3599
transform 1 0 31188 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp -3599
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp -3599
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_357
timestamp -3599
transform 1 0 33948 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_371
timestamp -3599
transform 1 0 35236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_375
timestamp -3599
transform 1 0 35604 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_381
timestamp -3599
transform 1 0 36156 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_387
timestamp -3599
transform 1 0 36708 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp -3599
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp -3599
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_401
timestamp -3599
transform 1 0 37996 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1636964856
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1636964856
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1636964856
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp -3599
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp -3599
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_449
timestamp -3599
transform 1 0 42412 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636964856
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636964856
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636964856
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636964856
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636964856
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636964856
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636964856
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636964856
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636964856
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636964856
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp -3599
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp -3599
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636964856
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_153
timestamp -3599
transform 1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_159
timestamp 1636964856
transform 1 0 15732 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_171
timestamp 1636964856
transform 1 0 16836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_183
timestamp -3599
transform 1 0 17940 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp -3599
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_210
timestamp 1636964856
transform 1 0 20424 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_222
timestamp -3599
transform 1 0 21528 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_228
timestamp 1636964856
transform 1 0 22080 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_240
timestamp -3599
transform 1 0 23184 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp -3599
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp -3599
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp -3599
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_261
timestamp 1636964856
transform 1 0 25116 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_273
timestamp 1636964856
transform 1 0 26220 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_288
timestamp 1636964856
transform 1 0 27600 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_300
timestamp -3599
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_309
timestamp -3599
transform 1 0 29532 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_318
timestamp 1636964856
transform 1 0 30360 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_330
timestamp -3599
transform 1 0 31464 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_336
timestamp -3599
transform 1 0 32016 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_341
timestamp 1636964856
transform 1 0 32476 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_353
timestamp -3599
transform 1 0 33580 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_361
timestamp -3599
transform 1 0 34316 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636964856
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636964856
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636964856
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1636964856
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp -3599
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp -3599
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636964856
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636964856
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_445
timestamp -3599
transform 1 0 42044 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_453
timestamp -3599
transform 1 0 42780 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp -3599
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_13
timestamp 1636964856
transform 1 0 2300 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_25
timestamp -3599
transform 1 0 3404 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_31
timestamp -3599
transform 1 0 3956 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_35
timestamp 1636964856
transform 1 0 4324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp -3599
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -3599
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636964856
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636964856
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636964856
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636964856
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp -3599
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -3599
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636964856
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636964856
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636964856
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636964856
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp -3599
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -3599
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp -3599
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_178
timestamp 1636964856
transform 1 0 17480 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_190
timestamp 1636964856
transform 1 0 18584 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_202
timestamp 1636964856
transform 1 0 19688 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_214
timestamp -3599
transform 1 0 20792 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp -3599
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636964856
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636964856
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_249
timestamp -3599
transform 1 0 24012 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_254
timestamp 1636964856
transform 1 0 24472 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_266
timestamp 1636964856
transform 1 0 25576 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp -3599
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_281
timestamp -3599
transform 1 0 26956 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_292
timestamp 1636964856
transform 1 0 27968 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_304
timestamp 1636964856
transform 1 0 29072 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_316
timestamp 1636964856
transform 1 0 30176 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_328
timestamp -3599
transform 1 0 31280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_337
timestamp -3599
transform 1 0 32108 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_341
timestamp 1636964856
transform 1 0 32476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_353
timestamp 1636964856
transform 1 0 33580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_365
timestamp 1636964856
transform 1 0 34684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_377
timestamp 1636964856
transform 1 0 35788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_389
timestamp -3599
transform 1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636964856
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636964856
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1636964856
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1636964856
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp -3599
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp -3599
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_449
timestamp -3599
transform 1 0 42412 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_453
timestamp -3599
transform 1 0 42780 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636964856
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636964856
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636964856
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636964856
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636964856
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_65
timestamp -3599
transform 1 0 7084 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_70
timestamp 1636964856
transform 1 0 7544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp -3599
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636964856
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636964856
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636964856
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_121
timestamp -3599
transform 1 0 12236 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_129
timestamp -3599
transform 1 0 12972 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp -3599
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp -3599
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636964856
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636964856
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_165
timestamp -3599
transform 1 0 16284 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_173
timestamp -3599
transform 1 0 17020 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_179
timestamp 1636964856
transform 1 0 17572 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_191
timestamp -3599
transform 1 0 18676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp -3599
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636964856
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636964856
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_221
timestamp -3599
transform 1 0 21436 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_232
timestamp 1636964856
transform 1 0 22448 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_244
timestamp -3599
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636964856
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_265
timestamp -3599
transform 1 0 25484 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_273
timestamp -3599
transform 1 0 26220 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_284
timestamp -3599
transform 1 0 27232 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_292
timestamp -3599
transform 1 0 27968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_300
timestamp -3599
transform 1 0 28704 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_309
timestamp -3599
transform 1 0 29532 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_318
timestamp 1636964856
transform 1 0 30360 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_330
timestamp 1636964856
transform 1 0 31464 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_342
timestamp 1636964856
transform 1 0 32568 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_354
timestamp -3599
transform 1 0 33672 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp -3599
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636964856
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636964856
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1636964856
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1636964856
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp -3599
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp -3599
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636964856
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636964856
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_445
timestamp -3599
transform 1 0 42044 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_453
timestamp -3599
transform 1 0 42780 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_11
timestamp -3599
transform 1 0 2116 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_16
timestamp 1636964856
transform 1 0 2576 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_28
timestamp -3599
transform 1 0 3680 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_34
timestamp 1636964856
transform 1 0 4232 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_46
timestamp -3599
transform 1 0 5336 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp -3599
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636964856
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636964856
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_81
timestamp -3599
transform 1 0 8556 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_89
timestamp -3599
transform 1 0 9292 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_97
timestamp 1636964856
transform 1 0 10028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_109
timestamp -3599
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636964856
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636964856
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636964856
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636964856
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp -3599
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp -3599
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_177
timestamp -3599
transform 1 0 17388 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_183
timestamp -3599
transform 1 0 17940 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_188
timestamp 1636964856
transform 1 0 18400 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_200
timestamp 1636964856
transform 1 0 19504 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_212
timestamp 1636964856
transform 1 0 20608 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_230
timestamp -3599
transform 1 0 22264 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_238
timestamp -3599
transform 1 0 23000 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_245
timestamp 1636964856
transform 1 0 23644 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_257
timestamp -3599
transform 1 0 24748 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_265
timestamp -3599
transform 1 0 25484 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_270
timestamp -3599
transform 1 0 25944 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp -3599
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_281
timestamp -3599
transform 1 0 26956 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_290
timestamp 1636964856
transform 1 0 27784 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_302
timestamp 1636964856
transform 1 0 28888 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_314
timestamp 1636964856
transform 1 0 29992 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_326
timestamp -3599
transform 1 0 31096 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp -3599
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636964856
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_354
timestamp 1636964856
transform 1 0 33672 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_366
timestamp 1636964856
transform 1 0 34776 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_378
timestamp -3599
transform 1 0 35880 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_386
timestamp -3599
transform 1 0 36616 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_398
timestamp 1636964856
transform 1 0 37720 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_410
timestamp 1636964856
transform 1 0 38824 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_422
timestamp 1636964856
transform 1 0 39928 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_434
timestamp 1636964856
transform 1 0 41032 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_446
timestamp -3599
transform 1 0 42136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_449
timestamp -3599
transform 1 0 42412 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_453
timestamp -3599
transform 1 0 42780 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636964856
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636964856
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636964856
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636964856
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_53
timestamp -3599
transform 1 0 5980 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_59
timestamp -3599
transform 1 0 6532 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_63
timestamp 1636964856
transform 1 0 6900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp -3599
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp -3599
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636964856
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636964856
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636964856
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1636964856
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp -3599
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp -3599
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_141
timestamp -3599
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_149
timestamp -3599
transform 1 0 14812 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_157
timestamp 1636964856
transform 1 0 15548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_169
timestamp 1636964856
transform 1 0 16652 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_181
timestamp -3599
transform 1 0 17756 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp -3599
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636964856
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636964856
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_224
timestamp 1636964856
transform 1 0 21712 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_236
timestamp 1636964856
transform 1 0 22816 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp -3599
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636964856
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_265
timestamp -3599
transform 1 0 25484 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_274
timestamp 1636964856
transform 1 0 26312 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_286
timestamp -3599
transform 1 0 27416 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_294
timestamp -3599
transform 1 0 28152 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_299
timestamp -3599
transform 1 0 28612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp -3599
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636964856
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_321
timestamp -3599
transform 1 0 30636 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_325
timestamp 1636964856
transform 1 0 31004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_337
timestamp 1636964856
transform 1 0 32108 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_349
timestamp -3599
transform 1 0 33212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_353
timestamp -3599
transform 1 0 33580 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp -3599
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp -3599
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_365
timestamp -3599
transform 1 0 34684 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_369
timestamp -3599
transform 1 0 35052 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_375
timestamp 1636964856
transform 1 0 35604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_387
timestamp 1636964856
transform 1 0 36708 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_399
timestamp 1636964856
transform 1 0 37812 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_411
timestamp -3599
transform 1 0 38916 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp -3599
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1636964856
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1636964856
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_445
timestamp -3599
transform 1 0 42044 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_453
timestamp -3599
transform 1 0 42780 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636964856
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636964856
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636964856
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636964856
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_51
timestamp -3599
transform 1 0 5796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -3599
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636964856
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636964856
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_81
timestamp -3599
transform 1 0 8556 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_85
timestamp -3599
transform 1 0 8924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_91
timestamp 1636964856
transform 1 0 9476 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_103
timestamp -3599
transform 1 0 10580 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp -3599
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636964856
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636964856
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_140
timestamp 1636964856
transform 1 0 13984 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_152
timestamp 1636964856
transform 1 0 15088 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp -3599
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_169
timestamp -3599
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_177
timestamp -3599
transform 1 0 17388 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_185
timestamp 1636964856
transform 1 0 18124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_197
timestamp 1636964856
transform 1 0 19228 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_212
timestamp -3599
transform 1 0 20608 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp -3599
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636964856
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636964856
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636964856
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_261
timestamp -3599
transform 1 0 25116 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_268
timestamp 1636964856
transform 1 0 25760 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636964856
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1636964856
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1636964856
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_317
timestamp -3599
transform 1 0 30268 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_325
timestamp -3599
transform 1 0 31004 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_330
timestamp -3599
transform 1 0 31464 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1636964856
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1636964856
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1636964856
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1636964856
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp -3599
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp -3599
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_393
timestamp -3599
transform 1 0 37260 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_397
timestamp -3599
transform 1 0 37628 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_401
timestamp -3599
transform 1 0 37996 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_407
timestamp -3599
transform 1 0 38548 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_416
timestamp 1636964856
transform 1 0 39376 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_428
timestamp -3599
transform 1 0 40480 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_434
timestamp -3599
transform 1 0 41032 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_438
timestamp -3599
transform 1 0 41400 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_446
timestamp -3599
transform 1 0 42136 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_449
timestamp -3599
transform 1 0 42412 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_453
timestamp -3599
transform 1 0 42780 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_12
timestamp 1636964856
transform 1 0 2208 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp -3599
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636964856
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636964856
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636964856
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636964856
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp -3599
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp -3599
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_89
timestamp -3599
transform 1 0 9292 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_93
timestamp 1636964856
transform 1 0 9660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_105
timestamp 1636964856
transform 1 0 10764 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_117
timestamp -3599
transform 1 0 11868 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_125
timestamp -3599
transform 1 0 12604 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_131
timestamp -3599
transform 1 0 13156 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp -3599
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636964856
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_153
timestamp -3599
transform 1 0 15180 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_159
timestamp -3599
transform 1 0 15732 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_166
timestamp 1636964856
transform 1 0 16376 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_178
timestamp 1636964856
transform 1 0 17480 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_190
timestamp -3599
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636964856
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636964856
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1636964856
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_233
timestamp -3599
transform 1 0 22540 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_239
timestamp 1636964856
transform 1 0 23092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp -3599
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_253
timestamp -3599
transform 1 0 24380 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_264
timestamp 1636964856
transform 1 0 25392 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_276
timestamp -3599
transform 1 0 26496 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_280
timestamp -3599
transform 1 0 26864 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_286
timestamp 1636964856
transform 1 0 27416 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_298
timestamp -3599
transform 1 0 28520 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp -3599
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_309
timestamp -3599
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_317
timestamp 1636964856
transform 1 0 30268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_329
timestamp 1636964856
transform 1 0 31372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_341
timestamp 1636964856
transform 1 0 32476 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_353
timestamp -3599
transform 1 0 33580 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_361
timestamp -3599
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp -3599
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_370
timestamp 1636964856
transform 1 0 35144 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_382
timestamp 1636964856
transform 1 0 36248 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_394
timestamp 1636964856
transform 1 0 37352 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_406
timestamp 1636964856
transform 1 0 38456 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_418
timestamp -3599
transform 1 0 39560 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1636964856
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1636964856
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_445
timestamp -3599
transform 1 0 42044 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_453
timestamp -3599
transform 1 0 42780 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636964856
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636964856
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636964856
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1636964856
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp -3599
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -3599
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636964856
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636964856
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1636964856
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1636964856
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp -3599
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp -3599
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636964856
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1636964856
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1636964856
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1636964856
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp -3599
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp -3599
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636964856
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_181
timestamp -3599
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_189
timestamp -3599
transform 1 0 18492 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_197
timestamp 1636964856
transform 1 0 19228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_209
timestamp 1636964856
transform 1 0 20332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp -3599
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp -3599
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_230
timestamp 1636964856
transform 1 0 22264 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_242
timestamp 1636964856
transform 1 0 23368 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_254
timestamp 1636964856
transform 1 0 24472 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_266
timestamp 1636964856
transform 1 0 25576 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp -3599
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636964856
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1636964856
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1636964856
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_317
timestamp -3599
transform 1 0 30268 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_328
timestamp -3599
transform 1 0 31280 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1636964856
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1636964856
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1636964856
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1636964856
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp -3599
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp -3599
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1636964856
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1636964856
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1636964856
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1636964856
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp -3599
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp -3599
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_449
timestamp -3599
transform 1 0 42412 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_453
timestamp -3599
transform 1 0 42780 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636964856
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636964856
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -3599
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_32
timestamp -3599
transform 1 0 4048 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_36
timestamp 1636964856
transform 1 0 4416 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_48
timestamp 1636964856
transform 1 0 5520 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_60
timestamp 1636964856
transform 1 0 6624 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_72
timestamp 1636964856
transform 1 0 7728 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636964856
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1636964856
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1636964856
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1636964856
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp -3599
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp -3599
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1636964856
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_153
timestamp -3599
transform 1 0 15180 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_161
timestamp -3599
transform 1 0 15916 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1636964856
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_177
timestamp -3599
transform 1 0 17388 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_183
timestamp 1636964856
transform 1 0 17940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp -3599
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_197
timestamp -3599
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_203
timestamp -3599
transform 1 0 19780 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_212
timestamp -3599
transform 1 0 20608 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_223
timestamp 1636964856
transform 1 0 21620 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_235
timestamp -3599
transform 1 0 22724 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_241
timestamp -3599
transform 1 0 23276 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_247
timestamp -3599
transform 1 0 23828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp -3599
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_258
timestamp 1636964856
transform 1 0 24840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_270
timestamp -3599
transform 1 0 25944 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_279
timestamp -3599
transform 1 0 26772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_288
timestamp -3599
transform 1 0 27600 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_297
timestamp -3599
transform 1 0 28428 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_305
timestamp -3599
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_314
timestamp 1636964856
transform 1 0 29992 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_326
timestamp 1636964856
transform 1 0 31096 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_338
timestamp 1636964856
transform 1 0 32200 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_350
timestamp 1636964856
transform 1 0 33304 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp -3599
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1636964856
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1636964856
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1636964856
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1636964856
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp -3599
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp -3599
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1636964856
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_433
timestamp -3599
transform 1 0 40940 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_441
timestamp -3599
transform 1 0 41676 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_6
timestamp 1636964856
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_18
timestamp -3599
transform 1 0 2760 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_26
timestamp -3599
transform 1 0 3496 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_33
timestamp 1636964856
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_45
timestamp -3599
transform 1 0 5244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp -3599
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636964856
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_69
timestamp -3599
transform 1 0 7452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_76
timestamp -3599
transform 1 0 8096 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_85
timestamp -3599
transform 1 0 8924 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_93
timestamp -3599
transform 1 0 9660 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_99
timestamp 1636964856
transform 1 0 10212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp -3599
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_117
timestamp -3599
transform 1 0 11868 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_122
timestamp 1636964856
transform 1 0 12328 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_134
timestamp -3599
transform 1 0 13432 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_145
timestamp 1636964856
transform 1 0 14444 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_157
timestamp -3599
transform 1 0 15548 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_163
timestamp -3599
transform 1 0 16100 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1636964856
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_181
timestamp -3599
transform 1 0 17756 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_191
timestamp -3599
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_195
timestamp -3599
transform 1 0 19044 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_197
timestamp 1636964856
transform 1 0 19228 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_209
timestamp -3599
transform 1 0 20332 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_214
timestamp -3599
transform 1 0 20792 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp -3599
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp -3599
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1636964856
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_249
timestamp -3599
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_253
timestamp -3599
transform 1 0 24380 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_260
timestamp 1636964856
transform 1 0 25024 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_272
timestamp -3599
transform 1 0 26128 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_285
timestamp 1636964856
transform 1 0 27324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_297
timestamp -3599
transform 1 0 28428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_301
timestamp -3599
transform 1 0 28796 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_306
timestamp -3599
transform 1 0 29256 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_309
timestamp 1636964856
transform 1 0 29532 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_321
timestamp -3599
transform 1 0 30636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp -3599
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp -3599
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_337
timestamp -3599
transform 1 0 32108 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_345
timestamp -3599
transform 1 0 32844 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_352
timestamp 1636964856
transform 1 0 33488 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_365
timestamp -3599
transform 1 0 34684 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_375
timestamp 1636964856
transform 1 0 35604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_387
timestamp -3599
transform 1 0 36708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp -3599
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_393
timestamp -3599
transform 1 0 37260 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_398
timestamp 1636964856
transform 1 0 37720 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_410
timestamp -3599
transform 1 0 38824 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_418
timestamp -3599
transform 1 0 39560 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_425
timestamp -3599
transform 1 0 40204 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_433
timestamp -3599
transform 1 0 40940 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_449
timestamp -3599
transform 1 0 42412 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output1
timestamp -3599
transform 1 0 42504 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform 1 0 43240 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform 1 0 42872 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform 1 0 43240 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform 1 0 42872 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform 1 0 43240 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 42872 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform 1 0 43240 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 42872 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -3599
transform 1 0 43240 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -3599
transform 1 0 42872 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -3599
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp -3599
transform 1 0 43240 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp -3599
transform 1 0 43240 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp -3599
transform 1 0 42872 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp -3599
transform 1 0 43240 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp -3599
transform 1 0 43240 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -3599
transform 1 0 42872 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp -3599
transform 1 0 42504 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp -3599
transform 1 0 41952 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp -3599
transform 1 0 42504 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp -3599
transform 1 0 42872 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp -3599
transform 1 0 42504 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp -3599
transform 1 0 42136 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp -3599
transform 1 0 41768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp -3599
transform 1 0 42872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp -3599
transform 1 0 43240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp -3599
transform 1 0 42872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp -3599
transform 1 0 43240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp -3599
transform 1 0 42872 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp -3599
transform 1 0 43240 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp -3599
transform 1 0 42872 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp -3599
transform -1 0 4140 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp -3599
transform -1 0 25024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp -3599
transform -1 0 27324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp -3599
transform -1 0 29256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp -3599
transform -1 0 31372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp -3599
transform -1 0 33488 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp -3599
transform 1 0 35236 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp -3599
transform -1 0 37720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp -3599
transform 1 0 39836 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp -3599
transform 1 0 41584 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp -3599
transform 1 0 41216 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp -3599
transform -1 0 5980 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp -3599
transform -1 0 8096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp -3599
transform -1 0 10212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp -3599
transform -1 0 12328 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp -3599
transform -1 0 14444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp -3599
transform -1 0 16560 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp -3599
transform -1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp -3599
transform -1 0 20792 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp -3599
transform -1 0 22908 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp -3599
transform 1 0 19504 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp -3599
transform 1 0 20056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp -3599
transform 1 0 19872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp -3599
transform 1 0 20240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp -3599
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp -3599
transform 1 0 21160 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp -3599
transform 1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp -3599
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp -3599
transform 1 0 21988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp -3599
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp -3599
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp -3599
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp -3599
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp -3599
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp -3599
transform 1 0 23644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp -3599
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp -3599
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp -3599
transform 1 0 25116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp -3599
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp -3599
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp -3599
transform 1 0 25300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp -3599
transform 1 0 28796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp -3599
transform 1 0 28336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp -3599
transform 1 0 28704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform 1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform 1 0 30268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform 1 0 26220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform 1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform -1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform -1 0 26772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform 1 0 27692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform 1 0 27508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform -1 0 30084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform 1 0 33948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform 1 0 33212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform 1 0 33580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform 1 0 35052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform -1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform -1 0 31924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform -1 0 32476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform -1 0 31188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform -1 0 31556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform -1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform -1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform -1 0 32476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output105
timestamp -3599
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 43884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 43884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 43884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 43884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 43884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 43884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 43884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 43884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 43884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 43884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 43884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 43884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_38
timestamp -3599
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_39
timestamp -3599
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_45
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_46
timestamp -3599
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_47
timestamp -3599
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_48
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_49
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_50
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_52
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_53
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_54
timestamp -3599
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_55
timestamp -3599
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_56
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_57
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_58
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_59
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_60
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_61
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_62
timestamp -3599
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_63
timestamp -3599
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_65
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_66
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_67
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_68
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_69
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_70
timestamp -3599
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_71
timestamp -3599
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_73
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_74
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_75
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_76
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_77
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_78
timestamp -3599
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_79
timestamp -3599
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_80
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_81
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_82
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_83
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_84
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_85
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_86
timestamp -3599
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_87
timestamp -3599
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_88
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_89
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_90
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_91
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_92
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_93
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_94
timestamp -3599
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_95
timestamp -3599
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_96
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_97
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_98
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_99
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_100
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_101
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_102
timestamp -3599
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_103
timestamp -3599
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_104
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_105
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_106
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_107
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_108
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_109
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_110
timestamp -3599
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_111
timestamp -3599
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_112
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_113
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_114
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_115
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_116
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_117
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_118
timestamp -3599
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_119
timestamp -3599
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_121
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_122
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_123
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_124
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_125
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_126
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_127
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_128
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_129
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_130
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_131
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_132
timestamp -3599
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_133
timestamp -3599
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp -3599
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp -3599
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 9800 120 9920 0 FreeSans 480 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 44880 1368 45000 1488 0 FreeSans 480 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 44880 4088 45000 4208 0 FreeSans 480 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 44880 4360 45000 4480 0 FreeSans 480 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 44880 4632 45000 4752 0 FreeSans 480 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 44880 4904 45000 5024 0 FreeSans 480 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 44880 5176 45000 5296 0 FreeSans 480 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 44880 5448 45000 5568 0 FreeSans 480 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 44880 5720 45000 5840 0 FreeSans 480 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 44880 5992 45000 6112 0 FreeSans 480 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 44880 6264 45000 6384 0 FreeSans 480 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 44880 6536 45000 6656 0 FreeSans 480 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 44880 1640 45000 1760 0 FreeSans 480 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 44880 6808 45000 6928 0 FreeSans 480 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 44880 7080 45000 7200 0 FreeSans 480 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 44880 7352 45000 7472 0 FreeSans 480 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 44880 7624 45000 7744 0 FreeSans 480 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 44880 7896 45000 8016 0 FreeSans 480 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 44880 8168 45000 8288 0 FreeSans 480 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 44880 8440 45000 8560 0 FreeSans 480 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 44880 8712 45000 8832 0 FreeSans 480 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 44880 8984 45000 9104 0 FreeSans 480 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 44880 9256 45000 9376 0 FreeSans 480 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 44880 1912 45000 2032 0 FreeSans 480 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 44880 9528 45000 9648 0 FreeSans 480 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 44880 9800 45000 9920 0 FreeSans 480 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 44880 2184 45000 2304 0 FreeSans 480 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 44880 2456 45000 2576 0 FreeSans 480 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 44880 2728 45000 2848 0 FreeSans 480 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 44880 3000 45000 3120 0 FreeSans 480 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 44880 3272 45000 3392 0 FreeSans 480 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 44880 3544 45000 3664 0 FreeSans 480 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 44880 3816 45000 3936 0 FreeSans 480 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 34334 0 34390 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 37094 0 37150 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 37370 0 37426 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 37646 0 37702 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 37922 0 37978 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 38198 0 38254 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 38474 0 38530 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 38750 0 38806 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 39026 0 39082 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 39302 0 39358 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 39578 0 39634 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 34610 0 34666 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 34886 0 34942 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 35162 0 35218 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 35438 0 35494 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 35714 0 35770 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 35990 0 36046 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 36266 0 36322 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 36542 0 36598 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 36818 0 36874 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 3422 11194 3478 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 24582 11194 24638 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 26698 11194 26754 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 28814 11194 28870 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 30930 11194 30986 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 33046 11194 33102 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 35162 11194 35218 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 37278 11194 37334 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 39394 11194 39450 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 41510 11194 41566 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 43626 11194 43682 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 5538 11194 5594 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 7654 11194 7710 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 9770 11194 9826 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 11886 11194 11942 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 14002 11194 14058 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 16118 11194 16174 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 18234 11194 18290 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 20350 11194 20406 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 22466 11194 22522 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 5354 0 5410 56 0 FreeSans 224 0 0 0 N1END[0]
port 104 nsew signal input
flabel metal2 s 5630 0 5686 56 0 FreeSans 224 0 0 0 N1END[1]
port 105 nsew signal input
flabel metal2 s 5906 0 5962 56 0 FreeSans 224 0 0 0 N1END[2]
port 106 nsew signal input
flabel metal2 s 6182 0 6238 56 0 FreeSans 224 0 0 0 N1END[3]
port 107 nsew signal input
flabel metal2 s 8666 0 8722 56 0 FreeSans 224 0 0 0 N2END[0]
port 108 nsew signal input
flabel metal2 s 8942 0 8998 56 0 FreeSans 224 0 0 0 N2END[1]
port 109 nsew signal input
flabel metal2 s 9218 0 9274 56 0 FreeSans 224 0 0 0 N2END[2]
port 110 nsew signal input
flabel metal2 s 9494 0 9550 56 0 FreeSans 224 0 0 0 N2END[3]
port 111 nsew signal input
flabel metal2 s 9770 0 9826 56 0 FreeSans 224 0 0 0 N2END[4]
port 112 nsew signal input
flabel metal2 s 10046 0 10102 56 0 FreeSans 224 0 0 0 N2END[5]
port 113 nsew signal input
flabel metal2 s 10322 0 10378 56 0 FreeSans 224 0 0 0 N2END[6]
port 114 nsew signal input
flabel metal2 s 10598 0 10654 56 0 FreeSans 224 0 0 0 N2END[7]
port 115 nsew signal input
flabel metal2 s 6458 0 6514 56 0 FreeSans 224 0 0 0 N2MID[0]
port 116 nsew signal input
flabel metal2 s 6734 0 6790 56 0 FreeSans 224 0 0 0 N2MID[1]
port 117 nsew signal input
flabel metal2 s 7010 0 7066 56 0 FreeSans 224 0 0 0 N2MID[2]
port 118 nsew signal input
flabel metal2 s 7286 0 7342 56 0 FreeSans 224 0 0 0 N2MID[3]
port 119 nsew signal input
flabel metal2 s 7562 0 7618 56 0 FreeSans 224 0 0 0 N2MID[4]
port 120 nsew signal input
flabel metal2 s 7838 0 7894 56 0 FreeSans 224 0 0 0 N2MID[5]
port 121 nsew signal input
flabel metal2 s 8114 0 8170 56 0 FreeSans 224 0 0 0 N2MID[6]
port 122 nsew signal input
flabel metal2 s 8390 0 8446 56 0 FreeSans 224 0 0 0 N2MID[7]
port 123 nsew signal input
flabel metal2 s 10874 0 10930 56 0 FreeSans 224 0 0 0 N4END[0]
port 124 nsew signal input
flabel metal2 s 13634 0 13690 56 0 FreeSans 224 0 0 0 N4END[10]
port 125 nsew signal input
flabel metal2 s 13910 0 13966 56 0 FreeSans 224 0 0 0 N4END[11]
port 126 nsew signal input
flabel metal2 s 14186 0 14242 56 0 FreeSans 224 0 0 0 N4END[12]
port 127 nsew signal input
flabel metal2 s 14462 0 14518 56 0 FreeSans 224 0 0 0 N4END[13]
port 128 nsew signal input
flabel metal2 s 14738 0 14794 56 0 FreeSans 224 0 0 0 N4END[14]
port 129 nsew signal input
flabel metal2 s 15014 0 15070 56 0 FreeSans 224 0 0 0 N4END[15]
port 130 nsew signal input
flabel metal2 s 11150 0 11206 56 0 FreeSans 224 0 0 0 N4END[1]
port 131 nsew signal input
flabel metal2 s 11426 0 11482 56 0 FreeSans 224 0 0 0 N4END[2]
port 132 nsew signal input
flabel metal2 s 11702 0 11758 56 0 FreeSans 224 0 0 0 N4END[3]
port 133 nsew signal input
flabel metal2 s 11978 0 12034 56 0 FreeSans 224 0 0 0 N4END[4]
port 134 nsew signal input
flabel metal2 s 12254 0 12310 56 0 FreeSans 224 0 0 0 N4END[5]
port 135 nsew signal input
flabel metal2 s 12530 0 12586 56 0 FreeSans 224 0 0 0 N4END[6]
port 136 nsew signal input
flabel metal2 s 12806 0 12862 56 0 FreeSans 224 0 0 0 N4END[7]
port 137 nsew signal input
flabel metal2 s 13082 0 13138 56 0 FreeSans 224 0 0 0 N4END[8]
port 138 nsew signal input
flabel metal2 s 13358 0 13414 56 0 FreeSans 224 0 0 0 N4END[9]
port 139 nsew signal input
flabel metal2 s 15290 0 15346 56 0 FreeSans 224 0 0 0 NN4END[0]
port 140 nsew signal input
flabel metal2 s 18050 0 18106 56 0 FreeSans 224 0 0 0 NN4END[10]
port 141 nsew signal input
flabel metal2 s 18326 0 18382 56 0 FreeSans 224 0 0 0 NN4END[11]
port 142 nsew signal input
flabel metal2 s 18602 0 18658 56 0 FreeSans 224 0 0 0 NN4END[12]
port 143 nsew signal input
flabel metal2 s 18878 0 18934 56 0 FreeSans 224 0 0 0 NN4END[13]
port 144 nsew signal input
flabel metal2 s 19154 0 19210 56 0 FreeSans 224 0 0 0 NN4END[14]
port 145 nsew signal input
flabel metal2 s 19430 0 19486 56 0 FreeSans 224 0 0 0 NN4END[15]
port 146 nsew signal input
flabel metal2 s 15566 0 15622 56 0 FreeSans 224 0 0 0 NN4END[1]
port 147 nsew signal input
flabel metal2 s 15842 0 15898 56 0 FreeSans 224 0 0 0 NN4END[2]
port 148 nsew signal input
flabel metal2 s 16118 0 16174 56 0 FreeSans 224 0 0 0 NN4END[3]
port 149 nsew signal input
flabel metal2 s 16394 0 16450 56 0 FreeSans 224 0 0 0 NN4END[4]
port 150 nsew signal input
flabel metal2 s 16670 0 16726 56 0 FreeSans 224 0 0 0 NN4END[5]
port 151 nsew signal input
flabel metal2 s 16946 0 17002 56 0 FreeSans 224 0 0 0 NN4END[6]
port 152 nsew signal input
flabel metal2 s 17222 0 17278 56 0 FreeSans 224 0 0 0 NN4END[7]
port 153 nsew signal input
flabel metal2 s 17498 0 17554 56 0 FreeSans 224 0 0 0 NN4END[8]
port 154 nsew signal input
flabel metal2 s 17774 0 17830 56 0 FreeSans 224 0 0 0 NN4END[9]
port 155 nsew signal input
flabel metal2 s 19706 0 19762 56 0 FreeSans 224 0 0 0 S1BEG[0]
port 156 nsew signal output
flabel metal2 s 19982 0 20038 56 0 FreeSans 224 0 0 0 S1BEG[1]
port 157 nsew signal output
flabel metal2 s 20258 0 20314 56 0 FreeSans 224 0 0 0 S1BEG[2]
port 158 nsew signal output
flabel metal2 s 20534 0 20590 56 0 FreeSans 224 0 0 0 S1BEG[3]
port 159 nsew signal output
flabel metal2 s 20810 0 20866 56 0 FreeSans 224 0 0 0 S2BEG[0]
port 160 nsew signal output
flabel metal2 s 21086 0 21142 56 0 FreeSans 224 0 0 0 S2BEG[1]
port 161 nsew signal output
flabel metal2 s 21362 0 21418 56 0 FreeSans 224 0 0 0 S2BEG[2]
port 162 nsew signal output
flabel metal2 s 21638 0 21694 56 0 FreeSans 224 0 0 0 S2BEG[3]
port 163 nsew signal output
flabel metal2 s 21914 0 21970 56 0 FreeSans 224 0 0 0 S2BEG[4]
port 164 nsew signal output
flabel metal2 s 22190 0 22246 56 0 FreeSans 224 0 0 0 S2BEG[5]
port 165 nsew signal output
flabel metal2 s 22466 0 22522 56 0 FreeSans 224 0 0 0 S2BEG[6]
port 166 nsew signal output
flabel metal2 s 22742 0 22798 56 0 FreeSans 224 0 0 0 S2BEG[7]
port 167 nsew signal output
flabel metal2 s 23018 0 23074 56 0 FreeSans 224 0 0 0 S2BEGb[0]
port 168 nsew signal output
flabel metal2 s 23294 0 23350 56 0 FreeSans 224 0 0 0 S2BEGb[1]
port 169 nsew signal output
flabel metal2 s 23570 0 23626 56 0 FreeSans 224 0 0 0 S2BEGb[2]
port 170 nsew signal output
flabel metal2 s 23846 0 23902 56 0 FreeSans 224 0 0 0 S2BEGb[3]
port 171 nsew signal output
flabel metal2 s 24122 0 24178 56 0 FreeSans 224 0 0 0 S2BEGb[4]
port 172 nsew signal output
flabel metal2 s 24398 0 24454 56 0 FreeSans 224 0 0 0 S2BEGb[5]
port 173 nsew signal output
flabel metal2 s 24674 0 24730 56 0 FreeSans 224 0 0 0 S2BEGb[6]
port 174 nsew signal output
flabel metal2 s 24950 0 25006 56 0 FreeSans 224 0 0 0 S2BEGb[7]
port 175 nsew signal output
flabel metal2 s 25226 0 25282 56 0 FreeSans 224 0 0 0 S4BEG[0]
port 176 nsew signal output
flabel metal2 s 27986 0 28042 56 0 FreeSans 224 0 0 0 S4BEG[10]
port 177 nsew signal output
flabel metal2 s 28262 0 28318 56 0 FreeSans 224 0 0 0 S4BEG[11]
port 178 nsew signal output
flabel metal2 s 28538 0 28594 56 0 FreeSans 224 0 0 0 S4BEG[12]
port 179 nsew signal output
flabel metal2 s 28814 0 28870 56 0 FreeSans 224 0 0 0 S4BEG[13]
port 180 nsew signal output
flabel metal2 s 29090 0 29146 56 0 FreeSans 224 0 0 0 S4BEG[14]
port 181 nsew signal output
flabel metal2 s 29366 0 29422 56 0 FreeSans 224 0 0 0 S4BEG[15]
port 182 nsew signal output
flabel metal2 s 25502 0 25558 56 0 FreeSans 224 0 0 0 S4BEG[1]
port 183 nsew signal output
flabel metal2 s 25778 0 25834 56 0 FreeSans 224 0 0 0 S4BEG[2]
port 184 nsew signal output
flabel metal2 s 26054 0 26110 56 0 FreeSans 224 0 0 0 S4BEG[3]
port 185 nsew signal output
flabel metal2 s 26330 0 26386 56 0 FreeSans 224 0 0 0 S4BEG[4]
port 186 nsew signal output
flabel metal2 s 26606 0 26662 56 0 FreeSans 224 0 0 0 S4BEG[5]
port 187 nsew signal output
flabel metal2 s 26882 0 26938 56 0 FreeSans 224 0 0 0 S4BEG[6]
port 188 nsew signal output
flabel metal2 s 27158 0 27214 56 0 FreeSans 224 0 0 0 S4BEG[7]
port 189 nsew signal output
flabel metal2 s 27434 0 27490 56 0 FreeSans 224 0 0 0 S4BEG[8]
port 190 nsew signal output
flabel metal2 s 27710 0 27766 56 0 FreeSans 224 0 0 0 S4BEG[9]
port 191 nsew signal output
flabel metal2 s 29642 0 29698 56 0 FreeSans 224 0 0 0 SS4BEG[0]
port 192 nsew signal output
flabel metal2 s 32402 0 32458 56 0 FreeSans 224 0 0 0 SS4BEG[10]
port 193 nsew signal output
flabel metal2 s 32678 0 32734 56 0 FreeSans 224 0 0 0 SS4BEG[11]
port 194 nsew signal output
flabel metal2 s 32954 0 33010 56 0 FreeSans 224 0 0 0 SS4BEG[12]
port 195 nsew signal output
flabel metal2 s 33230 0 33286 56 0 FreeSans 224 0 0 0 SS4BEG[13]
port 196 nsew signal output
flabel metal2 s 33506 0 33562 56 0 FreeSans 224 0 0 0 SS4BEG[14]
port 197 nsew signal output
flabel metal2 s 33782 0 33838 56 0 FreeSans 224 0 0 0 SS4BEG[15]
port 198 nsew signal output
flabel metal2 s 29918 0 29974 56 0 FreeSans 224 0 0 0 SS4BEG[1]
port 199 nsew signal output
flabel metal2 s 30194 0 30250 56 0 FreeSans 224 0 0 0 SS4BEG[2]
port 200 nsew signal output
flabel metal2 s 30470 0 30526 56 0 FreeSans 224 0 0 0 SS4BEG[3]
port 201 nsew signal output
flabel metal2 s 30746 0 30802 56 0 FreeSans 224 0 0 0 SS4BEG[4]
port 202 nsew signal output
flabel metal2 s 31022 0 31078 56 0 FreeSans 224 0 0 0 SS4BEG[5]
port 203 nsew signal output
flabel metal2 s 31298 0 31354 56 0 FreeSans 224 0 0 0 SS4BEG[6]
port 204 nsew signal output
flabel metal2 s 31574 0 31630 56 0 FreeSans 224 0 0 0 SS4BEG[7]
port 205 nsew signal output
flabel metal2 s 31850 0 31906 56 0 FreeSans 224 0 0 0 SS4BEG[8]
port 206 nsew signal output
flabel metal2 s 32126 0 32182 56 0 FreeSans 224 0 0 0 SS4BEG[9]
port 207 nsew signal output
flabel metal2 s 34058 0 34114 56 0 FreeSans 224 0 0 0 UserCLK
port 208 nsew signal input
flabel metal2 s 1306 11194 1362 11250 0 FreeSans 224 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal4 s 3004 0 3324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 3004 11190 3324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 11190 9324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 11190 15324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 11190 21324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 11190 27324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 11190 33324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 0 39324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 0 39324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 11190 39324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 1944 11190 2264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 0 8264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 11190 8264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 0 14264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 11190 14264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 0 20264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 11190 20264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 0 26264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 11190 26264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 0 32264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 11190 32264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 0 38264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 0 38264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 11190 38264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
rlabel metal1 22494 8704 22494 8704 0 VGND
rlabel metal1 22494 8160 22494 8160 0 VPWR
rlabel metal3 528 1428 528 1428 0 FrameData[0]
rlabel metal3 666 4148 666 4148 0 FrameData[10]
rlabel metal3 712 4420 712 4420 0 FrameData[11]
rlabel metal3 3495 4692 3495 4692 0 FrameData[12]
rlabel metal3 942 4964 942 4964 0 FrameData[13]
rlabel metal2 19550 4369 19550 4369 0 FrameData[14]
rlabel metal3 1494 5508 1494 5508 0 FrameData[15]
rlabel metal1 18814 5236 18814 5236 0 FrameData[16]
rlabel metal3 919 6052 919 6052 0 FrameData[17]
rlabel metal1 13156 4998 13156 4998 0 FrameData[18]
rlabel metal3 1471 6596 1471 6596 0 FrameData[19]
rlabel metal2 7222 3417 7222 3417 0 FrameData[1]
rlabel metal1 21068 6426 21068 6426 0 FrameData[20]
rlabel metal3 919 7140 919 7140 0 FrameData[21]
rlabel metal3 712 7412 712 7412 0 FrameData[22]
rlabel metal3 1471 7684 1471 7684 0 FrameData[23]
rlabel metal1 24058 7854 24058 7854 0 FrameData[24]
rlabel metal3 942 8228 942 8228 0 FrameData[25]
rlabel metal2 26358 8279 26358 8279 0 FrameData[26]
rlabel metal3 1494 8772 1494 8772 0 FrameData[27]
rlabel metal1 21114 7854 21114 7854 0 FrameData[28]
rlabel metal1 16238 8058 16238 8058 0 FrameData[29]
rlabel metal3 2828 1972 2828 1972 0 FrameData[2]
rlabel metal2 19366 8721 19366 8721 0 FrameData[30]
rlabel metal3 666 9860 666 9860 0 FrameData[31]
rlabel metal3 1471 2244 1471 2244 0 FrameData[3]
rlabel metal2 7406 4063 7406 4063 0 FrameData[4]
rlabel metal3 919 2788 919 2788 0 FrameData[5]
rlabel metal2 13294 5168 13294 5168 0 FrameData[6]
rlabel metal3 1494 3332 1494 3332 0 FrameData[7]
rlabel metal2 14950 4624 14950 4624 0 FrameData[8]
rlabel metal3 942 3876 942 3876 0 FrameData[9]
rlabel metal3 43822 1428 43822 1428 0 FrameData_O[0]
rlabel metal3 44190 4148 44190 4148 0 FrameData_O[10]
rlabel metal3 44006 4420 44006 4420 0 FrameData_O[11]
rlabel metal3 44190 4692 44190 4692 0 FrameData_O[12]
rlabel metal3 44006 4964 44006 4964 0 FrameData_O[13]
rlabel metal3 44190 5236 44190 5236 0 FrameData_O[14]
rlabel metal3 44006 5508 44006 5508 0 FrameData_O[15]
rlabel metal3 44190 5780 44190 5780 0 FrameData_O[16]
rlabel metal3 44006 6052 44006 6052 0 FrameData_O[17]
rlabel metal3 44190 6324 44190 6324 0 FrameData_O[18]
rlabel metal3 44006 6596 44006 6596 0 FrameData_O[19]
rlabel metal3 43546 1700 43546 1700 0 FrameData_O[1]
rlabel metal3 44190 6868 44190 6868 0 FrameData_O[20]
rlabel metal3 44190 7140 44190 7140 0 FrameData_O[21]
rlabel metal3 44006 7412 44006 7412 0 FrameData_O[22]
rlabel metal3 44190 7684 44190 7684 0 FrameData_O[23]
rlabel metal3 44190 7956 44190 7956 0 FrameData_O[24]
rlabel metal3 44006 8228 44006 8228 0 FrameData_O[25]
rlabel metal3 43822 8500 43822 8500 0 FrameData_O[26]
rlabel metal2 42182 8687 42182 8687 0 FrameData_O[27]
rlabel metal1 42688 8058 42688 8058 0 FrameData_O[28]
rlabel metal1 43148 7514 43148 7514 0 FrameData_O[29]
rlabel metal3 43960 1972 43960 1972 0 FrameData_O[2]
rlabel metal2 42366 8823 42366 8823 0 FrameData_O[30]
rlabel metal2 41998 8959 41998 8959 0 FrameData_O[31]
rlabel metal3 44006 2244 44006 2244 0 FrameData_O[3]
rlabel metal3 44190 2516 44190 2516 0 FrameData_O[4]
rlabel metal3 44006 2788 44006 2788 0 FrameData_O[5]
rlabel metal3 44190 3060 44190 3060 0 FrameData_O[6]
rlabel metal3 44006 3332 44006 3332 0 FrameData_O[7]
rlabel metal3 44190 3604 44190 3604 0 FrameData_O[8]
rlabel metal3 44006 3876 44006 3876 0 FrameData_O[9]
rlabel metal2 9430 6239 9430 6239 0 FrameStrobe[0]
rlabel metal2 37122 735 37122 735 0 FrameStrobe[10]
rlabel metal2 33258 5950 33258 5950 0 FrameStrobe[11]
rlabel metal1 34822 6290 34822 6290 0 FrameStrobe[12]
rlabel metal2 37950 735 37950 735 0 FrameStrobe[13]
rlabel metal2 38226 735 38226 735 0 FrameStrobe[14]
rlabel metal1 36708 6766 36708 6766 0 FrameStrobe[15]
rlabel metal1 38364 6222 38364 6222 0 FrameStrobe[16]
rlabel metal2 39054 735 39054 735 0 FrameStrobe[17]
rlabel metal2 39330 735 39330 735 0 FrameStrobe[18]
rlabel metal1 40388 6290 40388 6290 0 FrameStrobe[19]
rlabel metal1 9982 5236 9982 5236 0 FrameStrobe[1]
rlabel via2 34914 55 34914 55 0 FrameStrobe[2]
rlabel metal1 22034 3604 22034 3604 0 FrameStrobe[3]
rlabel metal2 35466 650 35466 650 0 FrameStrobe[4]
rlabel metal2 35742 1401 35742 1401 0 FrameStrobe[5]
rlabel metal2 36018 1401 36018 1401 0 FrameStrobe[6]
rlabel metal1 33994 6392 33994 6392 0 FrameStrobe[7]
rlabel metal2 36570 1401 36570 1401 0 FrameStrobe[8]
rlabel metal2 36846 3744 36846 3744 0 FrameStrobe[9]
rlabel metal1 3680 8602 3680 8602 0 FrameStrobe_O[0]
rlabel metal1 24702 8602 24702 8602 0 FrameStrobe_O[10]
rlabel metal1 26910 8602 26910 8602 0 FrameStrobe_O[11]
rlabel metal1 28934 8602 28934 8602 0 FrameStrobe_O[12]
rlabel metal1 31050 8602 31050 8602 0 FrameStrobe_O[13]
rlabel metal1 33074 8602 33074 8602 0 FrameStrobe_O[14]
rlabel metal1 35328 8602 35328 8602 0 FrameStrobe_O[15]
rlabel metal1 37398 8602 37398 8602 0 FrameStrobe_O[16]
rlabel metal1 39744 8602 39744 8602 0 FrameStrobe_O[17]
rlabel metal1 41676 8602 41676 8602 0 FrameStrobe_O[18]
rlabel metal2 41446 8704 41446 8704 0 FrameStrobe_O[19]
rlabel metal1 5658 8602 5658 8602 0 FrameStrobe_O[1]
rlabel metal1 7774 8602 7774 8602 0 FrameStrobe_O[2]
rlabel metal1 9890 8602 9890 8602 0 FrameStrobe_O[3]
rlabel metal1 12006 8602 12006 8602 0 FrameStrobe_O[4]
rlabel metal1 14122 8602 14122 8602 0 FrameStrobe_O[5]
rlabel metal1 16238 8602 16238 8602 0 FrameStrobe_O[6]
rlabel metal1 18354 8602 18354 8602 0 FrameStrobe_O[7]
rlabel metal1 20470 8602 20470 8602 0 FrameStrobe_O[8]
rlabel metal1 22586 8602 22586 8602 0 FrameStrobe_O[9]
rlabel metal2 5382 1534 5382 1534 0 N1END[0]
rlabel metal2 5658 2044 5658 2044 0 N1END[1]
rlabel metal2 5934 2588 5934 2588 0 N1END[2]
rlabel metal2 6210 3404 6210 3404 0 N1END[3]
rlabel metal2 8694 2316 8694 2316 0 N2END[0]
rlabel metal2 8970 803 8970 803 0 N2END[1]
rlabel metal2 9246 55 9246 55 0 N2END[2]
rlabel metal2 9522 2860 9522 2860 0 N2END[3]
rlabel metal2 9798 1500 9798 1500 0 N2END[4]
rlabel metal2 10074 3404 10074 3404 0 N2END[5]
rlabel metal2 10350 1534 10350 1534 0 N2END[6]
rlabel metal2 10626 3404 10626 3404 0 N2END[7]
rlabel metal2 6486 1534 6486 1534 0 N2MID[0]
rlabel metal2 6762 2316 6762 2316 0 N2MID[1]
rlabel metal2 7038 2860 7038 2860 0 N2MID[2]
rlabel metal2 7314 3166 7314 3166 0 N2MID[3]
rlabel metal1 3818 7820 3818 7820 0 N2MID[4]
rlabel metal2 7866 55 7866 55 0 N2MID[5]
rlabel metal2 8142 55 8142 55 0 N2MID[6]
rlabel metal2 8418 2078 8418 2078 0 N2MID[7]
rlabel metal2 10902 3948 10902 3948 0 N4END[0]
rlabel metal1 13708 6290 13708 6290 0 N4END[10]
rlabel metal2 13938 242 13938 242 0 N4END[11]
rlabel metal2 14214 140 14214 140 0 N4END[12]
rlabel metal2 14490 718 14490 718 0 N4END[13]
rlabel metal1 10902 6256 10902 6256 0 N4END[14]
rlabel metal2 15042 735 15042 735 0 N4END[15]
rlabel metal2 11178 3642 11178 3642 0 N4END[1]
rlabel metal2 11454 1007 11454 1007 0 N4END[2]
rlabel metal2 11730 582 11730 582 0 N4END[3]
rlabel metal2 12006 2894 12006 2894 0 N4END[4]
rlabel metal2 12282 3370 12282 3370 0 N4END[5]
rlabel metal1 14352 6834 14352 6834 0 N4END[6]
rlabel metal2 12834 2792 12834 2792 0 N4END[7]
rlabel metal1 15916 3434 15916 3434 0 N4END[8]
rlabel metal2 13386 2248 13386 2248 0 N4END[9]
rlabel metal2 15318 242 15318 242 0 NN4END[0]
rlabel metal2 18078 55 18078 55 0 NN4END[10]
rlabel metal2 18354 327 18354 327 0 NN4END[11]
rlabel metal2 18630 191 18630 191 0 NN4END[12]
rlabel metal2 18906 1007 18906 1007 0 NN4END[13]
rlabel metal2 19182 55 19182 55 0 NN4END[14]
rlabel metal2 19458 1024 19458 1024 0 NN4END[15]
rlabel metal2 15594 174 15594 174 0 NN4END[1]
rlabel metal3 18170 3196 18170 3196 0 NN4END[2]
rlabel metal2 16146 208 16146 208 0 NN4END[3]
rlabel metal2 16422 259 16422 259 0 NN4END[4]
rlabel metal2 16698 1483 16698 1483 0 NN4END[5]
rlabel metal2 16974 990 16974 990 0 NN4END[6]
rlabel metal2 17250 106 17250 106 0 NN4END[7]
rlabel metal2 17526 123 17526 123 0 NN4END[8]
rlabel metal2 17802 735 17802 735 0 NN4END[9]
rlabel metal2 19734 1160 19734 1160 0 S1BEG[0]
rlabel metal2 20010 55 20010 55 0 S1BEG[1]
rlabel metal2 20286 1160 20286 1160 0 S1BEG[2]
rlabel metal2 20562 1160 20562 1160 0 S1BEG[3]
rlabel metal2 20838 1160 20838 1160 0 S2BEG[0]
rlabel metal2 21114 55 21114 55 0 S2BEG[1]
rlabel metal2 21390 1160 21390 1160 0 S2BEG[2]
rlabel metal2 21666 1160 21666 1160 0 S2BEG[3]
rlabel metal2 21942 1432 21942 1432 0 S2BEG[4]
rlabel metal2 22218 1160 22218 1160 0 S2BEG[5]
rlabel metal2 22494 1160 22494 1160 0 S2BEG[6]
rlabel metal2 22770 1160 22770 1160 0 S2BEG[7]
rlabel metal2 23046 1160 23046 1160 0 S2BEGb[0]
rlabel metal2 23322 1160 23322 1160 0 S2BEGb[1]
rlabel metal2 23598 1160 23598 1160 0 S2BEGb[2]
rlabel metal2 23874 1160 23874 1160 0 S2BEGb[3]
rlabel metal2 24150 1296 24150 1296 0 S2BEGb[4]
rlabel metal2 24426 718 24426 718 0 S2BEGb[5]
rlabel metal2 24702 1160 24702 1160 0 S2BEGb[6]
rlabel metal2 24978 1194 24978 1194 0 S2BEGb[7]
rlabel metal1 25392 2822 25392 2822 0 S4BEG[0]
rlabel metal2 28014 1194 28014 1194 0 S4BEG[10]
rlabel metal1 28428 2822 28428 2822 0 S4BEG[11]
rlabel metal2 28612 2822 28612 2822 0 S4BEG[12]
rlabel metal2 28842 1296 28842 1296 0 S4BEG[13]
rlabel metal2 29118 1160 29118 1160 0 S4BEG[14]
rlabel metal2 29394 1194 29394 1194 0 S4BEG[15]
rlabel metal2 25530 1296 25530 1296 0 S4BEG[1]
rlabel metal1 25944 2822 25944 2822 0 S4BEG[2]
rlabel metal2 26082 1160 26082 1160 0 S4BEG[3]
rlabel metal1 26450 2822 26450 2822 0 S4BEG[4]
rlabel metal2 26634 1296 26634 1296 0 S4BEG[5]
rlabel metal2 26910 1194 26910 1194 0 S4BEG[6]
rlabel metal2 27186 55 27186 55 0 S4BEG[7]
rlabel metal2 27508 2822 27508 2822 0 S4BEG[8]
rlabel metal2 27738 1296 27738 1296 0 S4BEG[9]
rlabel metal1 29762 2822 29762 2822 0 SS4BEG[0]
rlabel metal2 32430 1330 32430 1330 0 SS4BEG[10]
rlabel metal2 32706 735 32706 735 0 SS4BEG[11]
rlabel metal2 32982 735 32982 735 0 SS4BEG[12]
rlabel metal2 33258 684 33258 684 0 SS4BEG[13]
rlabel metal1 33672 2822 33672 2822 0 SS4BEG[14]
rlabel metal2 33810 599 33810 599 0 SS4BEG[15]
rlabel metal2 29946 1296 29946 1296 0 SS4BEG[1]
rlabel metal2 30222 1330 30222 1330 0 SS4BEG[2]
rlabel metal2 30498 599 30498 599 0 SS4BEG[3]
rlabel metal1 30866 2822 30866 2822 0 SS4BEG[4]
rlabel metal2 31050 1160 31050 1160 0 SS4BEG[5]
rlabel metal2 31326 1296 31326 1296 0 SS4BEG[6]
rlabel metal1 32982 2312 32982 2312 0 SS4BEG[7]
rlabel metal1 32062 3366 32062 3366 0 SS4BEG[8]
rlabel metal2 32154 1211 32154 1211 0 SS4BEG[9]
rlabel metal2 13478 4641 13478 4641 0 UserCLK
rlabel metal1 1380 8602 1380 8602 0 UserCLKo
rlabel metal2 42550 2465 42550 2465 0 net1
rlabel via2 43286 6307 43286 6307 0 net10
rlabel metal1 35650 3162 35650 3162 0 net100
rlabel metal1 33580 2074 33580 2074 0 net101
rlabel metal1 33810 2380 33810 2380 0 net102
rlabel metal2 34270 3332 34270 3332 0 net103
rlabel metal1 33120 2482 33120 2482 0 net104
rlabel metal1 3542 8398 3542 8398 0 net105
rlabel metal1 25346 6868 25346 6868 0 net11
rlabel metal2 33534 4998 33534 4998 0 net12
rlabel metal2 25438 5984 25438 5984 0 net13
rlabel metal2 18078 6936 18078 6936 0 net14
rlabel metal1 33258 5066 33258 5066 0 net15
rlabel metal2 20654 7106 20654 7106 0 net16
rlabel metal1 24748 8058 24748 8058 0 net17
rlabel metal2 23782 8296 23782 8296 0 net18
rlabel metal1 28060 8058 28060 8058 0 net19
rlabel metal2 36570 4488 36570 4488 0 net2
rlabel metal1 21390 7990 21390 7990 0 net20
rlabel metal2 21390 8160 21390 8160 0 net21
rlabel metal2 21298 7956 21298 7956 0 net22
rlabel metal2 40066 3638 40066 3638 0 net23
rlabel metal1 19550 7752 19550 7752 0 net24
rlabel metal2 29762 7616 29762 7616 0 net25
rlabel metal1 42918 2516 42918 2516 0 net26
rlabel metal1 43930 2176 43930 2176 0 net27
rlabel metal2 35650 6664 35650 6664 0 net28
rlabel metal1 31878 6120 31878 6120 0 net29
rlabel metal1 28106 2890 28106 2890 0 net3
rlabel metal1 31740 4488 31740 4488 0 net30
rlabel metal2 34454 5134 34454 5134 0 net31
rlabel metal2 29578 5338 29578 5338 0 net32
rlabel metal1 4968 8466 4968 8466 0 net33
rlabel metal1 29992 6086 29992 6086 0 net34
rlabel metal1 30774 5610 30774 5610 0 net35
rlabel metal1 30498 6426 30498 6426 0 net36
rlabel metal1 33580 5814 33580 5814 0 net37
rlabel metal1 35972 5338 35972 5338 0 net38
rlabel metal2 35098 7548 35098 7548 0 net39
rlabel metal1 31740 3604 31740 3604 0 net4
rlabel metal1 37720 6426 37720 6426 0 net40
rlabel metal1 39192 6426 39192 6426 0 net41
rlabel metal2 41630 7310 41630 7310 0 net42
rlabel metal1 41308 6426 41308 6426 0 net43
rlabel metal1 6394 8466 6394 8466 0 net44
rlabel metal1 12190 8466 12190 8466 0 net45
rlabel metal1 10166 8398 10166 8398 0 net46
rlabel metal2 12282 8704 12282 8704 0 net47
rlabel metal1 14398 8500 14398 8500 0 net48
rlabel metal2 16514 8772 16514 8772 0 net49
rlabel metal1 25070 3706 25070 3706 0 net5
rlabel metal2 18630 8738 18630 8738 0 net50
rlabel metal2 20746 8636 20746 8636 0 net51
rlabel metal2 31050 7990 31050 7990 0 net52
rlabel metal1 2162 6664 2162 6664 0 net53
rlabel metal2 2530 4896 2530 4896 0 net54
rlabel metal1 19826 2414 19826 2414 0 net55
rlabel metal2 7682 2652 7682 2652 0 net56
rlabel metal2 4278 3808 4278 3808 0 net57
rlabel metal2 4370 7616 4370 7616 0 net58
rlabel metal2 7498 3706 7498 3706 0 net59
rlabel metal2 19918 3417 19918 3417 0 net6
rlabel metal2 4002 7344 4002 7344 0 net60
rlabel metal2 9614 4828 9614 4828 0 net61
rlabel metal2 8510 5593 8510 5593 0 net62
rlabel metal2 10994 3536 10994 3536 0 net63
rlabel metal1 11040 2822 11040 2822 0 net64
rlabel metal1 13156 6630 13156 6630 0 net65
rlabel metal1 13754 3162 13754 3162 0 net66
rlabel metal2 9614 6766 9614 6766 0 net67
rlabel metal1 16054 2890 16054 2890 0 net68
rlabel metal2 15226 6120 15226 6120 0 net69
rlabel via2 20194 3621 20194 3621 0 net7
rlabel metal2 15686 3264 15686 3264 0 net70
rlabel metal2 16146 3468 16146 3468 0 net71
rlabel metal1 25806 2414 25806 2414 0 net72
rlabel metal1 25346 2958 25346 2958 0 net73
rlabel metal2 16054 4250 16054 4250 0 net74
rlabel metal1 21666 5712 21666 5712 0 net75
rlabel metal2 20562 5814 20562 5814 0 net76
rlabel metal2 29578 2587 29578 2587 0 net77
rlabel metal1 21758 7956 21758 7956 0 net78
rlabel metal3 19780 5304 19780 5304 0 net79
rlabel metal1 22034 5304 22034 5304 0 net8
rlabel metal2 11086 4301 11086 4301 0 net80
rlabel metal2 25898 3740 25898 3740 0 net81
rlabel metal2 27278 2587 27278 2587 0 net82
rlabel metal1 26726 3060 26726 3060 0 net83
rlabel metal1 14398 6086 14398 6086 0 net84
rlabel metal1 19504 4998 19504 4998 0 net85
rlabel metal2 18906 3230 18906 3230 0 net86
rlabel metal1 18492 5882 18492 5882 0 net87
rlabel metal1 18906 2074 18906 2074 0 net88
rlabel metal2 38134 3298 38134 3298 0 net89
rlabel via1 33166 5117 33166 5117 0 net9
rlabel metal1 33166 2890 33166 2890 0 net90
rlabel metal2 33212 2516 33212 2516 0 net91
rlabel metal1 33258 2992 33258 2992 0 net92
rlabel metal2 34730 3060 34730 3060 0 net93
rlabel metal2 33626 3502 33626 3502 0 net94
rlabel metal2 35098 2040 35098 2040 0 net95
rlabel metal2 37306 3400 37306 3400 0 net96
rlabel metal1 33856 1938 33856 1938 0 net97
rlabel metal1 33856 2006 33856 2006 0 net98
rlabel metal2 33442 4046 33442 4046 0 net99
<< properties >>
string FIXED_BBOX 0 0 45000 11250
<< end >>
