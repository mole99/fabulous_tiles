* NGSPICE file created from N_term_DSP.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

.subckt N_term_DSP FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1] N1END[2] N1END[3]
+ N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6] N2END[7] N2MID[0]
+ N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4END[0] NN4END[10] NN4END[11] NN4END[12]
+ NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3] NN4END[4] NN4END[5]
+ NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S2BEG[0]
+ S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1]
+ S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S4BEG[0] S4BEG[10] S4BEG[11]
+ S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5]
+ S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] SS4BEG[0] SS4BEG[10] SS4BEG[11] SS4BEG[12] SS4BEG[13]
+ SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4] SS4BEG[5] SS4BEG[6]
+ SS4BEG[7] SS4BEG[8] SS4BEG[9] UserCLK UserCLKo VGND VPWR
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_9_148 VPWR VGND sg13g2_fill_1
XFILLER_5_376 VPWR VGND sg13g2_fill_1
XFILLER_3_56 VPWR VGND sg13g2_decap_8
XFILLER_8_181 VPWR VGND sg13g2_decap_8
XFILLER_10_147 VPWR VGND sg13g2_decap_8
XFILLER_2_313 VPWR VGND sg13g2_decap_4
XFILLER_2_357 VPWR VGND sg13g2_decap_8
XFILLER_5_173 VPWR VGND sg13g2_decap_8
X_062_ N2MID[1] net63 VPWR VGND sg13g2_buf_1
XFILLER_9_88 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_2_187 VPWR VGND sg13g2_decap_8
XFILLER_11_231 VPWR VGND sg13g2_decap_8
XFILLER_11_220 VPWR VGND sg13g2_decap_8
XFILLER_7_213 VPWR VGND sg13g2_decap_8
X_045_ FrameStrobe[13] net37 VPWR VGND sg13g2_buf_1
XFILLER_4_238 VPWR VGND sg13g2_decap_8
X_028_ FrameData[28] net21 VPWR VGND sg13g2_buf_1
XFILLER_6_89 VPWR VGND sg13g2_decap_8
XFILLER_3_282 VPWR VGND sg13g2_fill_1
XFILLER_9_308 VPWR VGND sg13g2_decap_8
Xoutput20 net20 FrameData_O[27] VPWR VGND sg13g2_buf_1
Xoutput42 net42 FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
XFILLER_8_352 VPWR VGND sg13g2_decap_8
Xoutput7 net7 FrameData_O[15] VPWR VGND sg13g2_buf_1
Xoutput97 net97 SS4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput75 net75 S4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput86 net86 S4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput64 net64 S2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput53 net53 S1BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_0_285 VPWR VGND sg13g2_decap_8
Xoutput31 net31 FrameData_O[8] VPWR VGND sg13g2_buf_1
XFILLER_11_0 VPWR VGND sg13g2_decap_8
XFILLER_10_329 VPWR VGND sg13g2_decap_8
XFILLER_9_116 VPWR VGND sg13g2_decap_4
XFILLER_5_355 VPWR VGND sg13g2_decap_8
XFILLER_3_35 VPWR VGND sg13g2_decap_8
XFILLER_8_160 VPWR VGND sg13g2_decap_8
XFILLER_10_126 VPWR VGND sg13g2_decap_8
XFILLER_2_336 VPWR VGND sg13g2_decap_8
XFILLER_5_152 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_2_166 VPWR VGND sg13g2_decap_4
X_061_ N2MID[2] net62 VPWR VGND sg13g2_buf_1
XFILLER_7_269 VPWR VGND sg13g2_decap_8
X_044_ FrameStrobe[12] net36 VPWR VGND sg13g2_buf_1
X_027_ FrameData[27] net20 VPWR VGND sg13g2_buf_1
XFILLER_6_68 VPWR VGND sg13g2_decap_8
XFILLER_3_250 VPWR VGND sg13g2_decap_8
XFILLER_3_261 VPWR VGND sg13g2_decap_8
Xoutput43 net43 FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
Xoutput21 net21 FrameData_O[28] VPWR VGND sg13g2_buf_1
Xoutput10 net10 FrameData_O[18] VPWR VGND sg13g2_buf_1
Xoutput8 net8 FrameData_O[16] VPWR VGND sg13g2_buf_1
Xoutput98 net98 SS4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput76 net76 S4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput87 net87 S4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput65 net65 S2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput54 net54 S1BEG[1] VPWR VGND sg13g2_buf_1
Xoutput32 net32 FrameData_O[9] VPWR VGND sg13g2_buf_1
XFILLER_10_308 VPWR VGND sg13g2_decap_8
XFILLER_8_331 VPWR VGND sg13g2_decap_8
XFILLER_5_334 VPWR VGND sg13g2_decap_8
XFILLER_3_14 VPWR VGND sg13g2_decap_8
XFILLER_10_105 VPWR VGND sg13g2_decap_8
XFILLER_5_131 VPWR VGND sg13g2_decap_8
XFILLER_9_35 VPWR VGND sg13g2_decap_8
XFILLER_2_112 VPWR VGND sg13g2_decap_8
XFILLER_2_145 VPWR VGND sg13g2_decap_8
X_060_ N2MID[3] net61 VPWR VGND sg13g2_buf_1
XFILLER_9_46 VPWR VGND sg13g2_decap_8
XFILLER_7_248 VPWR VGND sg13g2_decap_8
X_043_ FrameStrobe[11] net35 VPWR VGND sg13g2_buf_1
XFILLER_6_292 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_1_91 VPWR VGND sg13g2_decap_8
XFILLER_4_207 VPWR VGND sg13g2_decap_8
X_026_ FrameData[26] net19 VPWR VGND sg13g2_buf_1
XFILLER_6_47 VPWR VGND sg13g2_decap_8
XFILLER_6_14 VPWR VGND sg13g2_fill_1
Xoutput44 net44 FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
Xoutput33 net33 FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
Xoutput22 net22 FrameData_O[29] VPWR VGND sg13g2_buf_1
Xoutput11 net11 FrameData_O[19] VPWR VGND sg13g2_buf_1
Xoutput9 net9 FrameData_O[17] VPWR VGND sg13g2_buf_1
Xoutput99 net99 SS4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput77 net77 S4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput88 net88 S4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput66 net66 S2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput55 net55 S1BEG[2] VPWR VGND sg13g2_buf_1
X_009_ FrameData[9] net32 VPWR VGND sg13g2_buf_1
XFILLER_8_310 VPWR VGND sg13g2_decap_8
XFILLER_9_129 VPWR VGND sg13g2_fill_2
XFILLER_8_195 VPWR VGND sg13g2_decap_8
XFILLER_5_313 VPWR VGND sg13g2_decap_8
XFILLER_5_7 VPWR VGND sg13g2_decap_8
XFILLER_5_187 VPWR VGND sg13g2_decap_8
XFILLER_5_110 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_9_69 VPWR VGND sg13g2_fill_1
XFILLER_9_58 VPWR VGND sg13g2_decap_8
XFILLER_9_14 VPWR VGND sg13g2_decap_8
XFILLER_11_267 VPWR VGND sg13g2_decap_8
XFILLER_11_256 VPWR VGND sg13g2_decap_8
X_042_ FrameStrobe[10] net34 VPWR VGND sg13g2_buf_1
XFILLER_7_227 VPWR VGND sg13g2_decap_8
XFILLER_6_271 VPWR VGND sg13g2_fill_2
XFILLER_1_70 VPWR VGND sg13g2_decap_8
X_025_ FrameData[25] net18 VPWR VGND sg13g2_buf_1
XFILLER_6_26 VPWR VGND sg13g2_decap_8
Xoutput34 net34 FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
Xoutput45 net45 FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
Xoutput89 net89 SS4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput78 net78 S4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput67 net67 S2BEGb[2] VPWR VGND sg13g2_buf_1
Xoutput56 net56 S1BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_0_299 VPWR VGND sg13g2_decap_8
Xoutput12 net12 FrameData_O[1] VPWR VGND sg13g2_buf_1
Xoutput23 net23 FrameData_O[2] VPWR VGND sg13g2_buf_1
XFILLER_8_366 VPWR VGND sg13g2_decap_8
X_008_ FrameData[8] net31 VPWR VGND sg13g2_buf_1
XFILLER_7_80 VPWR VGND sg13g2_decap_8
XFILLER_5_369 VPWR VGND sg13g2_decap_8
XFILLER_3_49 VPWR VGND sg13g2_decap_8
XFILLER_8_174 VPWR VGND sg13g2_decap_8
XFILLER_2_317 VPWR VGND sg13g2_fill_1
XFILLER_5_166 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_11_213 VPWR VGND sg13g2_decap_8
XFILLER_11_202 VPWR VGND sg13g2_decap_8
X_041_ FrameStrobe[9] net52 VPWR VGND sg13g2_buf_1
XFILLER_7_206 VPWR VGND sg13g2_decap_8
XFILLER_6_250 VPWR VGND sg13g2_decap_8
X_024_ FrameData[24] net17 VPWR VGND sg13g2_buf_1
XFILLER_10_91 VPWR VGND sg13g2_decap_8
XFILLER_3_275 VPWR VGND sg13g2_decap_8
Xoutput24 net24 FrameData_O[30] VPWR VGND sg13g2_buf_1
Xoutput35 net35 FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
Xoutput46 net46 FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
Xoutput13 net13 FrameData_O[20] VPWR VGND sg13g2_buf_1
Xoutput57 net57 S2BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_8_345 VPWR VGND sg13g2_decap_8
Xoutput79 net79 S4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput68 net68 S2BEGb[3] VPWR VGND sg13g2_buf_1
X_007_ FrameData[7] net30 VPWR VGND sg13g2_buf_1
XFILLER_9_109 VPWR VGND sg13g2_decap_8
XFILLER_5_348 VPWR VGND sg13g2_decap_8
XFILLER_3_28 VPWR VGND sg13g2_decap_8
XFILLER_8_153 VPWR VGND sg13g2_decap_8
XFILLER_10_119 VPWR VGND sg13g2_decap_8
XFILLER_2_307 VPWR VGND sg13g2_fill_2
XFILLER_2_329 VPWR VGND sg13g2_decap_8
XFILLER_5_145 VPWR VGND sg13g2_decap_8
XFILLER_4_71 VPWR VGND sg13g2_fill_1
XFILLER_2_159 VPWR VGND sg13g2_decap_8
X_040_ FrameStrobe[8] net51 VPWR VGND sg13g2_buf_1
XFILLER_10_280 VPWR VGND sg13g2_decap_8
XFILLER_6_273 VPWR VGND sg13g2_fill_1
XFILLER_10_70 VPWR VGND sg13g2_decap_8
X_023_ FrameData[23] net16 VPWR VGND sg13g2_buf_1
XFILLER_3_243 VPWR VGND sg13g2_decap_8
XFILLER_3_287 VPWR VGND sg13g2_decap_8
XFILLER_3_298 VPWR VGND sg13g2_decap_8
Xoutput36 net36 FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
Xoutput47 net47 FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
Xoutput25 net25 FrameData_O[31] VPWR VGND sg13g2_buf_1
Xoutput14 net14 FrameData_O[21] VPWR VGND sg13g2_buf_1
XFILLER_8_324 VPWR VGND sg13g2_decap_8
Xoutput69 net69 S2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput58 net58 S2BEG[1] VPWR VGND sg13g2_buf_1
X_006_ FrameData[6] net29 VPWR VGND sg13g2_buf_1
XFILLER_5_327 VPWR VGND sg13g2_decap_8
XFILLER_8_132 VPWR VGND sg13g2_decap_8
XFILLER_4_360 VPWR VGND sg13g2_decap_8
XFILLER_5_124 VPWR VGND sg13g2_decap_8
XFILLER_1_352 VPWR VGND sg13g2_decap_8
XFILLER_9_28 VPWR VGND sg13g2_decap_8
XFILLER_2_105 VPWR VGND sg13g2_decap_8
XFILLER_2_138 VPWR VGND sg13g2_decap_8
XFILLER_3_7 VPWR VGND sg13g2_decap_8
XFILLER_6_285 VPWR VGND sg13g2_decap_8
X_099_ NN4END[4] net91 VPWR VGND sg13g2_buf_1
XFILLER_1_84 VPWR VGND sg13g2_decap_8
X_022_ FrameData[22] net15 VPWR VGND sg13g2_buf_1
Xoutput37 net37 FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
Xoutput48 net48 FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
Xoutput15 net15 FrameData_O[22] VPWR VGND sg13g2_buf_1
XFILLER_8_303 VPWR VGND sg13g2_decap_8
Xoutput59 net59 S2BEG[2] VPWR VGND sg13g2_buf_1
Xoutput26 net26 FrameData_O[3] VPWR VGND sg13g2_buf_1
X_005_ FrameData[5] net28 VPWR VGND sg13g2_buf_1
XFILLER_7_94 VPWR VGND sg13g2_decap_8
XFILLER_5_306 VPWR VGND sg13g2_decap_8
XFILLER_8_188 VPWR VGND sg13g2_decap_8
XFILLER_8_111 VPWR VGND sg13g2_decap_8
XFILLER_8_100 VPWR VGND sg13g2_fill_2
XFILLER_1_331 VPWR VGND sg13g2_decap_8
XFILLER_5_103 VPWR VGND sg13g2_decap_8
XFILLER_1_172 VPWR VGND sg13g2_fill_1
XFILLER_1_161 VPWR VGND sg13g2_decap_8
XFILLER_11_249 VPWR VGND sg13g2_decap_8
XFILLER_11_238 VPWR VGND sg13g2_decap_8
XFILLER_9_294 VPWR VGND sg13g2_decap_8
XFILLER_9_283 VPWR VGND sg13g2_decap_8
XFILLER_6_264 VPWR VGND sg13g2_decap_8
X_098_ NN4END[5] net90 VPWR VGND sg13g2_buf_1
XFILLER_1_63 VPWR VGND sg13g2_decap_8
X_021_ FrameData[21] net14 VPWR VGND sg13g2_buf_1
XFILLER_6_19 VPWR VGND sg13g2_decap_8
Xoutput38 net38 FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
Xoutput49 net49 FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
Xoutput16 net16 FrameData_O[23] VPWR VGND sg13g2_buf_1
Xoutput27 net27 FrameData_O[4] VPWR VGND sg13g2_buf_1
XFILLER_11_7 VPWR VGND sg13g2_decap_4
XFILLER_8_359 VPWR VGND sg13g2_decap_8
X_004_ FrameData[4] net27 VPWR VGND sg13g2_buf_1
XFILLER_7_73 VPWR VGND sg13g2_decap_8
XFILLER_8_167 VPWR VGND sg13g2_decap_8
XFILLER_5_159 VPWR VGND sg13g2_decap_8
XFILLER_1_310 VPWR VGND sg13g2_decap_8
XFILLER_1_140 VPWR VGND sg13g2_decap_8
XFILLER_10_294 VPWR VGND sg13g2_decap_8
XFILLER_6_243 VPWR VGND sg13g2_decap_8
XFILLER_1_42 VPWR VGND sg13g2_decap_8
X_097_ NN4END[6] net104 VPWR VGND sg13g2_buf_1
X_020_ FrameData[20] net13 VPWR VGND sg13g2_buf_1
XFILLER_3_268 VPWR VGND sg13g2_fill_2
XFILLER_10_84 VPWR VGND sg13g2_decap_8
Xoutput39 net39 FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
Xoutput17 net17 FrameData_O[24] VPWR VGND sg13g2_buf_1
Xoutput28 net28 FrameData_O[5] VPWR VGND sg13g2_buf_1
XFILLER_8_338 VPWR VGND sg13g2_decap_8
X_003_ FrameData[3] net26 VPWR VGND sg13g2_buf_1
XFILLER_7_360 VPWR VGND sg13g2_decap_8
XFILLER_7_52 VPWR VGND sg13g2_decap_8
XFILLER_8_102 VPWR VGND sg13g2_fill_1
XFILLER_8_146 VPWR VGND sg13g2_decap_8
XFILLER_4_374 VPWR VGND sg13g2_fill_2
XFILLER_5_138 VPWR VGND sg13g2_decap_8
XFILLER_1_366 VPWR VGND sg13g2_decap_8
XFILLER_4_42 VPWR VGND sg13g2_decap_8
XFILLER_4_193 VPWR VGND sg13g2_decap_8
XFILLER_2_119 VPWR VGND sg13g2_decap_4
XFILLER_4_97 VPWR VGND sg13g2_decap_8
XFILLER_8_0 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_10_273 VPWR VGND sg13g2_decap_8
XFILLER_6_299 VPWR VGND sg13g2_decap_8
XFILLER_6_222 VPWR VGND sg13g2_decap_8
XFILLER_1_98 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
X_096_ NN4END[7] net103 VPWR VGND sg13g2_buf_1
XFILLER_10_63 VPWR VGND sg13g2_decap_8
Xoutput18 net18 FrameData_O[25] VPWR VGND sg13g2_buf_1
Xoutput29 net29 FrameData_O[6] VPWR VGND sg13g2_buf_1
X_079_ N4END[8] net86 VPWR VGND sg13g2_buf_1
XFILLER_8_317 VPWR VGND sg13g2_decap_8
X_002_ FrameData[2] net23 VPWR VGND sg13g2_buf_1
XFILLER_7_42 VPWR VGND sg13g2_decap_4
XFILLER_8_125 VPWR VGND sg13g2_decap_8
XFILLER_4_331 VPWR VGND sg13g2_decap_4
XFILLER_4_353 VPWR VGND sg13g2_decap_8
XFILLER_5_117 VPWR VGND sg13g2_decap_8
XFILLER_1_345 VPWR VGND sg13g2_decap_8
XFILLER_4_21 VPWR VGND sg13g2_decap_8
XFILLER_9_253 VPWR VGND sg13g2_fill_1
XFILLER_1_197 VPWR VGND sg13g2_decap_8
XFILLER_10_252 VPWR VGND sg13g2_decap_8
XFILLER_6_278 VPWR VGND sg13g2_decap_8
XFILLER_6_201 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
X_095_ NN4END[8] net102 VPWR VGND sg13g2_buf_1
XFILLER_10_42 VPWR VGND sg13g2_decap_8
XFILLER_3_204 VPWR VGND sg13g2_fill_2
X_078_ N4END[9] net85 VPWR VGND sg13g2_buf_1
Xoutput19 net19 FrameData_O[26] VPWR VGND sg13g2_buf_1
X_001_ FrameData[1] net12 VPWR VGND sg13g2_buf_1
XFILLER_7_87 VPWR VGND sg13g2_decap_8
XFILLER_7_21 VPWR VGND sg13g2_decap_8
XFILLER_4_310 VPWR VGND sg13g2_fill_2
XFILLER_4_376 VPWR VGND sg13g2_fill_1
XFILLER_7_192 VPWR VGND sg13g2_decap_8
XFILLER_1_324 VPWR VGND sg13g2_decap_8
XFILLER_4_88 VPWR VGND sg13g2_fill_1
XFILLER_9_265 VPWR VGND sg13g2_decap_4
XFILLER_1_154 VPWR VGND sg13g2_decap_8
XFILLER_10_231 VPWR VGND sg13g2_decap_8
XFILLER_6_257 VPWR VGND sg13g2_decap_8
X_094_ NN4END[9] net101 VPWR VGND sg13g2_buf_1
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_10_98 VPWR VGND sg13g2_decap_8
XFILLER_10_21 VPWR VGND sg13g2_decap_8
XFILLER_2_293 VPWR VGND sg13g2_decap_8
X_077_ N4END[10] net84 VPWR VGND sg13g2_buf_1
XFILLER_7_374 VPWR VGND sg13g2_fill_2
XFILLER_7_66 VPWR VGND sg13g2_decap_8
X_000_ FrameData[0] net1 VPWR VGND sg13g2_buf_1
XFILLER_7_171 VPWR VGND sg13g2_decap_8
XFILLER_1_303 VPWR VGND sg13g2_decap_8
XFILLER_4_56 VPWR VGND sg13g2_decap_8
XFILLER_9_222 VPWR VGND sg13g2_fill_2
XFILLER_9_200 VPWR VGND sg13g2_fill_1
XFILLER_1_133 VPWR VGND sg13g2_decap_8
XFILLER_10_287 VPWR VGND sg13g2_decap_8
XFILLER_10_210 VPWR VGND sg13g2_decap_8
XFILLER_6_236 VPWR VGND sg13g2_decap_8
XFILLER_6_0 VPWR VGND sg13g2_decap_8
X_093_ NN4END[10] net100 VPWR VGND sg13g2_buf_1
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_10_77 VPWR VGND sg13g2_decap_8
XFILLER_3_206 VPWR VGND sg13g2_fill_1
XFILLER_2_272 VPWR VGND sg13g2_fill_2
X_076_ N4END[11] net83 VPWR VGND sg13g2_buf_1
XFILLER_7_353 VPWR VGND sg13g2_decap_8
X_059_ N2MID[4] net60 VPWR VGND sg13g2_buf_1
XFILLER_8_139 VPWR VGND sg13g2_decap_8
XFILLER_4_312 VPWR VGND sg13g2_fill_1
XFILLER_7_150 VPWR VGND sg13g2_decap_8
XFILLER_4_367 VPWR VGND sg13g2_decap_8
XFILLER_1_359 VPWR VGND sg13g2_decap_8
XFILLER_4_35 VPWR VGND sg13g2_decap_8
XFILLER_4_142 VPWR VGND sg13g2_decap_8
XFILLER_4_153 VPWR VGND sg13g2_fill_1
XFILLER_4_186 VPWR VGND sg13g2_decap_8
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_9_245 VPWR VGND sg13g2_decap_4
XFILLER_10_266 VPWR VGND sg13g2_decap_8
XFILLER_6_215 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
X_092_ NN4END[11] net99 VPWR VGND sg13g2_buf_1
XFILLER_10_56 VPWR VGND sg13g2_decap_8
XFILLER_5_292 VPWR VGND sg13g2_decap_8
XFILLER_2_251 VPWR VGND sg13g2_decap_8
X_075_ N4END[12] net82 VPWR VGND sg13g2_buf_1
XFILLER_11_361 VPWR VGND sg13g2_fill_2
XFILLER_7_376 VPWR VGND sg13g2_fill_1
XFILLER_7_332 VPWR VGND sg13g2_decap_8
XFILLER_7_46 VPWR VGND sg13g2_fill_2
XFILLER_7_35 VPWR VGND sg13g2_decap_8
X_058_ N2MID[5] net59 VPWR VGND sg13g2_buf_1
XFILLER_8_118 VPWR VGND sg13g2_decap_8
XFILLER_4_324 VPWR VGND sg13g2_decap_8
XFILLER_4_346 VPWR VGND sg13g2_decap_8
XFILLER_1_338 VPWR VGND sg13g2_decap_8
XFILLER_4_14 VPWR VGND sg13g2_decap_8
XFILLER_1_168 VPWR VGND sg13g2_decap_4
XFILLER_9_235 VPWR VGND sg13g2_decap_4
XFILLER_9_213 VPWR VGND sg13g2_fill_1
XFILLER_8_290 VPWR VGND sg13g2_fill_2
XFILLER_10_245 VPWR VGND sg13g2_decap_8
X_091_ NN4END[12] net98 VPWR VGND sg13g2_buf_1
XFILLER_5_271 VPWR VGND sg13g2_decap_8
XFILLER_10_35 VPWR VGND sg13g2_decap_8
X_074_ N4END[13] net81 VPWR VGND sg13g2_buf_1
XFILLER_2_230 VPWR VGND sg13g2_decap_8
XFILLER_2_274 VPWR VGND sg13g2_fill_1
XFILLER_2_91 VPWR VGND sg13g2_decap_8
XFILLER_7_311 VPWR VGND sg13g2_decap_8
XFILLER_7_14 VPWR VGND sg13g2_decap_8
X_057_ N2MID[6] net58 VPWR VGND sg13g2_buf_1
XFILLER_4_303 VPWR VGND sg13g2_decap_8
XFILLER_7_185 VPWR VGND sg13g2_decap_8
XFILLER_1_317 VPWR VGND sg13g2_decap_8
XFILLER_4_111 VPWR VGND sg13g2_decap_8
XFILLER_4_122 VPWR VGND sg13g2_fill_2
XFILLER_1_147 VPWR VGND sg13g2_decap_8
XFILLER_9_269 VPWR VGND sg13g2_fill_2
XFILLER_9_258 VPWR VGND sg13g2_decap_8
XFILLER_10_224 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
X_090_ NN4END[13] net97 VPWR VGND sg13g2_buf_1
XFILLER_5_250 VPWR VGND sg13g2_decap_8
XFILLER_10_14 VPWR VGND sg13g2_decap_8
XFILLER_2_286 VPWR VGND sg13g2_fill_2
X_073_ N4END[14] net80 VPWR VGND sg13g2_buf_1
XFILLER_4_0 VPWR VGND sg13g2_decap_8
XFILLER_2_70 VPWR VGND sg13g2_decap_8
XFILLER_7_367 VPWR VGND sg13g2_decap_8
XFILLER_7_59 VPWR VGND sg13g2_decap_8
X_056_ N2MID[7] net57 VPWR VGND sg13g2_buf_1
X_039_ FrameStrobe[7] net50 VPWR VGND sg13g2_buf_1
XFILLER_7_164 VPWR VGND sg13g2_decap_8
XFILLER_3_370 VPWR VGND sg13g2_fill_2
XFILLER_8_91 VPWR VGND sg13g2_decap_4
XFILLER_0_362 VPWR VGND sg13g2_decap_8
XFILLER_4_49 VPWR VGND sg13g2_decap_8
XFILLER_8_7 VPWR VGND sg13g2_decap_8
XFILLER_1_126 VPWR VGND sg13g2_decap_8
XFILLER_10_203 VPWR VGND sg13g2_decap_8
XFILLER_6_229 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
X_072_ N4END[15] net73 VPWR VGND sg13g2_buf_1
XFILLER_2_265 VPWR VGND sg13g2_decap_8
XFILLER_11_375 VPWR VGND sg13g2_fill_2
XFILLER_7_346 VPWR VGND sg13g2_decap_8
X_055_ N1END[0] net56 VPWR VGND sg13g2_buf_1
X_038_ FrameStrobe[6] net49 VPWR VGND sg13g2_buf_1
XFILLER_7_143 VPWR VGND sg13g2_decap_8
XFILLER_8_70 VPWR VGND sg13g2_decap_8
XFILLER_0_341 VPWR VGND sg13g2_decap_8
XFILLER_4_28 VPWR VGND sg13g2_decap_8
XFILLER_4_135 VPWR VGND sg13g2_decap_8
XFILLER_4_179 VPWR VGND sg13g2_decap_8
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_10_259 VPWR VGND sg13g2_decap_8
XFILLER_6_208 VPWR VGND sg13g2_decap_8
XFILLER_5_82 VPWR VGND sg13g2_decap_8
XFILLER_5_285 VPWR VGND sg13g2_decap_8
XFILLER_10_49 VPWR VGND sg13g2_decap_8
X_071_ N2END[0] net72 VPWR VGND sg13g2_buf_1
XFILLER_2_244 VPWR VGND sg13g2_decap_8
XFILLER_2_288 VPWR VGND sg13g2_fill_1
XFILLER_11_321 VPWR VGND sg13g2_decap_8
XFILLER_11_310 VPWR VGND sg13g2_decap_8
XFILLER_7_325 VPWR VGND sg13g2_decap_8
XFILLER_7_28 VPWR VGND sg13g2_decap_8
X_054_ N1END[1] net55 VPWR VGND sg13g2_buf_1
XFILLER_4_317 VPWR VGND sg13g2_decap_8
XFILLER_4_339 VPWR VGND sg13g2_decap_8
XFILLER_11_195 VPWR VGND sg13g2_decap_8
XFILLER_11_184 VPWR VGND sg13g2_decap_8
X_037_ FrameStrobe[5] net48 VPWR VGND sg13g2_buf_1
XFILLER_7_199 VPWR VGND sg13g2_decap_8
XFILLER_7_122 VPWR VGND sg13g2_decap_8
XFILLER_3_372 VPWR VGND sg13g2_fill_1
XFILLER_0_320 VPWR VGND sg13g2_decap_8
XFILLER_4_158 VPWR VGND sg13g2_decap_8
XFILLER_4_169 VPWR VGND sg13g2_fill_2
XFILLER_3_191 VPWR VGND sg13g2_fill_2
XFILLER_9_239 VPWR VGND sg13g2_fill_2
XFILLER_9_228 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_4
XFILLER_10_238 VPWR VGND sg13g2_decap_8
XFILLER_8_272 VPWR VGND sg13g2_decap_8
XFILLER_5_61 VPWR VGND sg13g2_decap_8
XFILLER_5_264 VPWR VGND sg13g2_decap_8
XFILLER_10_28 VPWR VGND sg13g2_decap_8
XFILLER_2_201 VPWR VGND sg13g2_decap_8
XFILLER_2_223 VPWR VGND sg13g2_decap_8
X_070_ N2END[1] net71 VPWR VGND sg13g2_buf_1
XFILLER_2_84 VPWR VGND sg13g2_decap_8
XFILLER_7_304 VPWR VGND sg13g2_decap_8
XFILLER_2_0 VPWR VGND sg13g2_decap_8
X_053_ N1END[2] net54 VPWR VGND sg13g2_buf_1
XFILLER_11_141 VPWR VGND sg13g2_decap_8
XFILLER_11_130 VPWR VGND sg13g2_decap_8
XFILLER_7_101 VPWR VGND sg13g2_decap_8
X_036_ FrameStrobe[4] net47 VPWR VGND sg13g2_buf_1
XFILLER_7_178 VPWR VGND sg13g2_decap_8
XFILLER_4_104 VPWR VGND sg13g2_decap_8
X_019_ FrameData[19] net11 VPWR VGND sg13g2_buf_1
XFILLER_9_218 VPWR VGND sg13g2_decap_4
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_8_251 VPWR VGND sg13g2_decap_8
XFILLER_5_40 VPWR VGND sg13g2_decap_8
XFILLER_10_217 VPWR VGND sg13g2_decap_8
XFILLER_6_7 VPWR VGND sg13g2_decap_8
XFILLER_5_243 VPWR VGND sg13g2_decap_8
XFILLER_2_279 VPWR VGND sg13g2_decap_8
XFILLER_2_63 VPWR VGND sg13g2_decap_8
XFILLER_11_94 VPWR VGND sg13g2_decap_8
X_052_ N1END[3] net53 VPWR VGND sg13g2_buf_1
X_035_ FrameStrobe[3] net46 VPWR VGND sg13g2_buf_1
XFILLER_7_157 VPWR VGND sg13g2_decap_8
X_104_ UserCLK net105 VPWR VGND sg13g2_buf_1
XFILLER_3_363 VPWR VGND sg13g2_decap_8
XFILLER_8_95 VPWR VGND sg13g2_fill_1
XFILLER_8_84 VPWR VGND sg13g2_decap_8
X_018_ FrameData[18] net10 VPWR VGND sg13g2_buf_1
XFILLER_0_355 VPWR VGND sg13g2_decap_8
XFILLER_4_149 VPWR VGND sg13g2_decap_4
XFILLER_1_119 VPWR VGND sg13g2_decap_8
XFILLER_10_0 VPWR VGND sg13g2_decap_8
XFILLER_8_296 VPWR VGND sg13g2_decap_8
XFILLER_8_230 VPWR VGND sg13g2_decap_8
XFILLER_5_96 VPWR VGND sg13g2_decap_8
XFILLER_5_299 VPWR VGND sg13g2_decap_8
XFILLER_5_222 VPWR VGND sg13g2_decap_8
XFILLER_2_258 VPWR VGND sg13g2_decap_8
XFILLER_2_42 VPWR VGND sg13g2_decap_8
XFILLER_11_357 VPWR VGND sg13g2_decap_4
XFILLER_11_346 VPWR VGND sg13g2_decap_8
XFILLER_11_51 VPWR VGND sg13g2_decap_8
XFILLER_11_40 VPWR VGND sg13g2_decap_8
XFILLER_7_339 VPWR VGND sg13g2_decap_8
X_051_ FrameStrobe[19] net43 VPWR VGND sg13g2_buf_1
XFILLER_6_361 VPWR VGND sg13g2_decap_8
X_034_ FrameStrobe[2] net45 VPWR VGND sg13g2_buf_1
XFILLER_7_136 VPWR VGND sg13g2_decap_8
X_103_ NN4END[0] net95 VPWR VGND sg13g2_buf_1
XFILLER_3_320 VPWR VGND sg13g2_fill_2
XFILLER_3_342 VPWR VGND sg13g2_decap_8
XFILLER_8_63 VPWR VGND sg13g2_decap_8
XFILLER_6_180 VPWR VGND sg13g2_decap_8
XFILLER_0_334 VPWR VGND sg13g2_decap_8
XFILLER_4_128 VPWR VGND sg13g2_decap_8
X_017_ FrameData[17] net9 VPWR VGND sg13g2_buf_1
XFILLER_9_209 VPWR VGND sg13g2_decap_4
XFILLER_8_286 VPWR VGND sg13g2_decap_4
XFILLER_5_75 VPWR VGND sg13g2_decap_8
XFILLER_5_278 VPWR VGND sg13g2_decap_8
XFILLER_5_201 VPWR VGND sg13g2_decap_8
XFILLER_2_237 VPWR VGND sg13g2_decap_8
XFILLER_2_21 VPWR VGND sg13g2_decap_8
XFILLER_2_98 VPWR VGND sg13g2_decap_8
XFILLER_11_303 VPWR VGND sg13g2_decap_8
XFILLER_7_318 VPWR VGND sg13g2_decap_8
Xoutput100 net100 SS4BEG[5] VPWR VGND sg13g2_buf_1
X_050_ FrameStrobe[18] net42 VPWR VGND sg13g2_buf_1
XFILLER_6_340 VPWR VGND sg13g2_decap_8
XFILLER_11_177 VPWR VGND sg13g2_decap_8
XFILLER_11_166 VPWR VGND sg13g2_decap_8
XFILLER_7_115 VPWR VGND sg13g2_decap_8
X_033_ FrameStrobe[1] net44 VPWR VGND sg13g2_buf_1
XFILLER_0_0 VPWR VGND sg13g2_decap_8
X_102_ NN4END[1] net94 VPWR VGND sg13g2_buf_1
XFILLER_8_42 VPWR VGND sg13g2_decap_8
XFILLER_0_313 VPWR VGND sg13g2_decap_8
XFILLER_4_118 VPWR VGND sg13g2_decap_4
X_016_ FrameData[16] net8 VPWR VGND sg13g2_buf_1
XFILLER_8_265 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_5_54 VPWR VGND sg13g2_decap_8
XFILLER_5_257 VPWR VGND sg13g2_decap_8
XFILLER_4_7 VPWR VGND sg13g2_decap_8
XFILLER_1_282 VPWR VGND sg13g2_decap_8
XFILLER_2_77 VPWR VGND sg13g2_decap_8
XFILLER_9_371 VPWR VGND sg13g2_decap_4
Xoutput101 net101 SS4BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_11_123 VPWR VGND sg13g2_decap_8
XFILLER_11_112 VPWR VGND sg13g2_decap_8
X_101_ NN4END[2] net93 VPWR VGND sg13g2_buf_1
XFILLER_3_322 VPWR VGND sg13g2_fill_1
X_032_ FrameStrobe[0] net33 VPWR VGND sg13g2_buf_1
XFILLER_8_21 VPWR VGND sg13g2_decap_8
X_015_ FrameData[15] net7 VPWR VGND sg13g2_buf_1
XFILLER_3_141 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_8_244 VPWR VGND sg13g2_decap_8
XFILLER_5_33 VPWR VGND sg13g2_decap_8
XFILLER_5_236 VPWR VGND sg13g2_decap_8
XFILLER_2_56 VPWR VGND sg13g2_decap_8
XFILLER_9_350 VPWR VGND sg13g2_decap_8
Xoutput102 net102 SS4BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_11_87 VPWR VGND sg13g2_decap_8
XFILLER_11_76 VPWR VGND sg13g2_decap_8
XFILLER_6_375 VPWR VGND sg13g2_fill_2
X_031_ FrameData[31] net25 VPWR VGND sg13g2_buf_1
X_100_ NN4END[3] net92 VPWR VGND sg13g2_buf_1
XFILLER_8_77 VPWR VGND sg13g2_decap_8
XFILLER_6_194 VPWR VGND sg13g2_decap_8
XFILLER_3_312 VPWR VGND sg13g2_decap_4
XFILLER_3_356 VPWR VGND sg13g2_decap_8
X_014_ FrameData[14] net6 VPWR VGND sg13g2_buf_1
XFILLER_0_348 VPWR VGND sg13g2_decap_8
XFILLER_3_197 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_8_223 VPWR VGND sg13g2_decap_8
XFILLER_5_89 VPWR VGND sg13g2_decap_8
XFILLER_5_215 VPWR VGND sg13g2_decap_8
Xoutput103 net103 SS4BEG[8] VPWR VGND sg13g2_buf_1
XFILLER_2_35 VPWR VGND sg13g2_decap_8
XFILLER_11_339 VPWR VGND sg13g2_decap_8
XFILLER_11_328 VPWR VGND sg13g2_decap_8
XFILLER_11_33 VPWR VGND sg13g2_decap_8
XFILLER_11_22 VPWR VGND sg13g2_decap_8
XFILLER_10_350 VPWR VGND sg13g2_decap_8
XFILLER_6_354 VPWR VGND sg13g2_decap_8
XFILLER_9_170 VPWR VGND sg13g2_fill_1
X_030_ FrameData[30] net24 VPWR VGND sg13g2_buf_1
XFILLER_8_56 VPWR VGND sg13g2_decap_8
XFILLER_7_129 VPWR VGND sg13g2_decap_8
XFILLER_3_335 VPWR VGND sg13g2_decap_8
XFILLER_6_173 VPWR VGND sg13g2_decap_8
X_013_ FrameData[13] net5 VPWR VGND sg13g2_buf_1
XFILLER_0_327 VPWR VGND sg13g2_decap_8
XFILLER_3_110 VPWR VGND sg13g2_fill_1
XFILLER_8_279 VPWR VGND sg13g2_decap_8
XFILLER_8_202 VPWR VGND sg13g2_decap_8
XFILLER_5_68 VPWR VGND sg13g2_decap_8
XFILLER_7_290 VPWR VGND sg13g2_decap_8
XFILLER_4_271 VPWR VGND sg13g2_decap_8
XFILLER_4_282 VPWR VGND sg13g2_decap_8
XFILLER_2_208 VPWR VGND sg13g2_decap_8
XFILLER_9_0 VPWR VGND sg13g2_decap_8
Xoutput104 net104 SS4BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_1_296 VPWR VGND sg13g2_decap_8
XFILLER_2_14 VPWR VGND sg13g2_decap_8
XFILLER_2_7 VPWR VGND sg13g2_decap_8
XFILLER_6_333 VPWR VGND sg13g2_decap_8
XFILLER_3_90 VPWR VGND sg13g2_fill_1
XFILLER_11_159 VPWR VGND sg13g2_decap_8
XFILLER_11_148 VPWR VGND sg13g2_decap_8
XFILLER_7_108 VPWR VGND sg13g2_decap_8
XFILLER_8_35 VPWR VGND sg13g2_decap_8
XFILLER_6_152 VPWR VGND sg13g2_decap_8
X_089_ NN4END[14] net96 VPWR VGND sg13g2_buf_1
XFILLER_0_306 VPWR VGND sg13g2_decap_8
X_012_ FrameData[12] net4 VPWR VGND sg13g2_buf_1
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_8_258 VPWR VGND sg13g2_decap_8
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_5_14 VPWR VGND sg13g2_fill_1
XFILLER_5_47 VPWR VGND sg13g2_decap_8
XFILLER_9_375 VPWR VGND sg13g2_fill_2
XFILLER_9_364 VPWR VGND sg13g2_decap_8
XFILLER_1_275 VPWR VGND sg13g2_decap_8
Xoutput105 net105 UserCLKo VPWR VGND sg13g2_buf_1
XFILLER_11_105 VPWR VGND sg13g2_decap_8
XFILLER_10_182 VPWR VGND sg13g2_decap_8
XFILLER_8_14 VPWR VGND sg13g2_decap_8
XFILLER_6_131 VPWR VGND sg13g2_decap_8
X_088_ NN4END[15] net89 VPWR VGND sg13g2_buf_1
X_011_ FrameData[11] net3 VPWR VGND sg13g2_buf_1
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_8_237 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_5_26 VPWR VGND sg13g2_decap_8
XFILLER_10_7 VPWR VGND sg13g2_decap_8
XFILLER_5_229 VPWR VGND sg13g2_decap_8
XFILLER_2_49 VPWR VGND sg13g2_decap_8
XFILLER_9_343 VPWR VGND sg13g2_decap_8
XFILLER_11_69 VPWR VGND sg13g2_decap_8
XFILLER_11_58 VPWR VGND sg13g2_decap_8
XFILLER_10_364 VPWR VGND sg13g2_decap_4
XFILLER_6_313 VPWR VGND sg13g2_fill_2
XFILLER_9_184 VPWR VGND sg13g2_fill_1
XFILLER_6_368 VPWR VGND sg13g2_decap_8
XFILLER_3_70 VPWR VGND sg13g2_fill_2
XFILLER_3_81 VPWR VGND sg13g2_decap_8
XFILLER_3_305 VPWR VGND sg13g2_decap_8
XFILLER_3_349 VPWR VGND sg13g2_decap_8
XFILLER_10_161 VPWR VGND sg13g2_decap_8
XFILLER_6_187 VPWR VGND sg13g2_decap_8
XFILLER_6_110 VPWR VGND sg13g2_decap_8
XFILLER_2_371 VPWR VGND sg13g2_decap_4
X_087_ N4END[0] net79 VPWR VGND sg13g2_buf_1
X_010_ FrameData[10] net2 VPWR VGND sg13g2_buf_1
XFILLER_3_135 VPWR VGND sg13g2_fill_2
XFILLER_8_216 VPWR VGND sg13g2_decap_8
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_5_208 VPWR VGND sg13g2_decap_8
XFILLER_4_252 VPWR VGND sg13g2_fill_2
XFILLER_4_296 VPWR VGND sg13g2_decap_8
XFILLER_2_28 VPWR VGND sg13g2_decap_8
XFILLER_9_322 VPWR VGND sg13g2_decap_8
XFILLER_11_15 VPWR VGND sg13g2_decap_8
XFILLER_10_343 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_6_347 VPWR VGND sg13g2_decap_8
XFILLER_10_140 VPWR VGND sg13g2_decap_8
XFILLER_8_49 VPWR VGND sg13g2_decap_8
XFILLER_6_166 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
X_086_ N4END[1] net78 VPWR VGND sg13g2_buf_1
XFILLER_2_350 VPWR VGND sg13g2_decap_8
XFILLER_2_180 VPWR VGND sg13g2_decap_8
X_069_ N2END[2] net70 VPWR VGND sg13g2_buf_1
XFILLER_9_81 VPWR VGND sg13g2_decap_8
XFILLER_7_283 VPWR VGND sg13g2_decap_8
XFILLER_6_82 VPWR VGND sg13g2_decap_8
XFILLER_4_231 VPWR VGND sg13g2_decap_8
XFILLER_4_264 VPWR VGND sg13g2_decap_8
XFILLER_9_301 VPWR VGND sg13g2_decap_8
Xoutput90 net90 SS4BEG[10] VPWR VGND sg13g2_buf_1
XFILLER_1_289 VPWR VGND sg13g2_decap_8
XFILLER_10_322 VPWR VGND sg13g2_decap_8
XFILLER_6_326 VPWR VGND sg13g2_decap_8
XFILLER_9_175 VPWR VGND sg13g2_fill_1
XFILLER_9_153 VPWR VGND sg13g2_decap_8
XFILLER_9_131 VPWR VGND sg13g2_fill_1
XFILLER_9_120 VPWR VGND sg13g2_fill_1
XFILLER_3_72 VPWR VGND sg13g2_fill_1
XFILLER_8_28 VPWR VGND sg13g2_decap_8
XFILLER_10_196 VPWR VGND sg13g2_decap_8
XFILLER_6_145 VPWR VGND sg13g2_decap_8
X_085_ N4END[2] net77 VPWR VGND sg13g2_buf_1
XFILLER_3_148 VPWR VGND sg13g2_decap_8
XFILLER_2_170 VPWR VGND sg13g2_fill_2
X_068_ N2END[3] net69 VPWR VGND sg13g2_buf_1
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_7_262 VPWR VGND sg13g2_decap_8
XFILLER_4_254 VPWR VGND sg13g2_fill_1
XFILLER_6_61 VPWR VGND sg13g2_decap_8
XFILLER_9_357 VPWR VGND sg13g2_decap_8
Xoutput1 net1 FrameData_O[0] VPWR VGND sg13g2_buf_1
Xoutput80 net80 S4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput91 net91 SS4BEG[11] VPWR VGND sg13g2_buf_1
XFILLER_10_301 VPWR VGND sg13g2_decap_8
XFILLER_9_198 VPWR VGND sg13g2_fill_2
XFILLER_10_175 VPWR VGND sg13g2_decap_8
XFILLER_6_124 VPWR VGND sg13g2_decap_8
X_084_ N4END[3] net76 VPWR VGND sg13g2_buf_1
XFILLER_0_63 VPWR VGND sg13g2_decap_8
X_067_ N2END[4] net68 VPWR VGND sg13g2_buf_1
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_5_19 VPWR VGND sg13g2_decap_8
XFILLER_11_292 VPWR VGND sg13g2_decap_8
XFILLER_7_241 VPWR VGND sg13g2_decap_8
XFILLER_4_200 VPWR VGND sg13g2_decap_8
XFILLER_6_40 VPWR VGND sg13g2_decap_8
XFILLER_9_336 VPWR VGND sg13g2_decap_8
Xoutput81 net81 S4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput70 net70 S2BEGb[5] VPWR VGND sg13g2_buf_1
Xoutput92 net92 SS4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput2 net2 FrameData_O[10] VPWR VGND sg13g2_buf_1
XFILLER_10_368 VPWR VGND sg13g2_fill_1
XFILLER_10_357 VPWR VGND sg13g2_decap_8
XFILLER_6_306 VPWR VGND sg13g2_decap_8
XFILLER_3_63 VPWR VGND sg13g2_decap_8
XFILLER_10_154 VPWR VGND sg13g2_decap_8
XFILLER_6_103 VPWR VGND sg13g2_decap_8
XFILLER_2_364 VPWR VGND sg13g2_decap_8
XFILLER_2_375 VPWR VGND sg13g2_fill_2
X_083_ N4END[4] net75 VPWR VGND sg13g2_buf_1
XFILLER_5_0 VPWR VGND sg13g2_decap_8
XFILLER_5_180 VPWR VGND sg13g2_decap_8
XFILLER_3_106 VPWR VGND sg13g2_decap_4
XFILLER_9_95 VPWR VGND sg13g2_decap_8
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_2_194 VPWR VGND sg13g2_decap_8
X_066_ N2END[5] net67 VPWR VGND sg13g2_buf_1
XFILLER_8_209 VPWR VGND sg13g2_decap_8
XFILLER_7_297 VPWR VGND sg13g2_decap_8
XFILLER_7_220 VPWR VGND sg13g2_decap_8
X_049_ FrameStrobe[17] net41 VPWR VGND sg13g2_buf_1
XFILLER_4_245 VPWR VGND sg13g2_decap_8
XFILLER_4_289 VPWR VGND sg13g2_decap_8
XFILLER_6_96 VPWR VGND sg13g2_decap_8
XFILLER_9_7 VPWR VGND sg13g2_decap_8
XFILLER_1_204 VPWR VGND sg13g2_decap_8
XFILLER_9_315 VPWR VGND sg13g2_decap_8
Xoutput82 net82 S4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput71 net71 S2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput60 net60 S2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput93 net93 SS4BEG[13] VPWR VGND sg13g2_buf_1
XFILLER_0_292 VPWR VGND sg13g2_decap_8
Xoutput3 net3 FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_10_336 VPWR VGND sg13g2_decap_8
XFILLER_9_189 VPWR VGND sg13g2_fill_1
XFILLER_5_362 VPWR VGND sg13g2_decap_8
XFILLER_3_42 VPWR VGND sg13g2_decap_8
XFILLER_10_133 VPWR VGND sg13g2_decap_8
XFILLER_6_159 VPWR VGND sg13g2_decap_8
XFILLER_2_343 VPWR VGND sg13g2_decap_8
X_082_ N4END[5] net74 VPWR VGND sg13g2_buf_1
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
X_065_ N2END[6] net66 VPWR VGND sg13g2_buf_1
XFILLER_9_74 VPWR VGND sg13g2_decap_8
XFILLER_7_276 VPWR VGND sg13g2_decap_8
X_048_ FrameStrobe[16] net40 VPWR VGND sg13g2_buf_1
XFILLER_4_224 VPWR VGND sg13g2_decap_8
XFILLER_6_75 VPWR VGND sg13g2_decap_8
Xoutput50 net50 FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
Xoutput83 net83 S4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput72 net72 S2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput61 net61 S2BEG[4] VPWR VGND sg13g2_buf_1
Xoutput94 net94 SS4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput4 net4 FrameData_O[12] VPWR VGND sg13g2_buf_1
XFILLER_10_315 VPWR VGND sg13g2_decap_8
XFILLER_9_102 VPWR VGND sg13g2_decap_8
XFILLER_6_319 VPWR VGND sg13g2_decap_8
XFILLER_9_168 VPWR VGND sg13g2_fill_2
XFILLER_5_341 VPWR VGND sg13g2_decap_8
XFILLER_3_21 VPWR VGND sg13g2_decap_8
XFILLER_10_189 VPWR VGND sg13g2_decap_8
XFILLER_10_112 VPWR VGND sg13g2_decap_8
XFILLER_6_138 VPWR VGND sg13g2_decap_8
XFILLER_2_300 VPWR VGND sg13g2_decap_8
XFILLER_2_322 VPWR VGND sg13g2_decap_8
X_081_ N4END[6] net88 VPWR VGND sg13g2_buf_1
XFILLER_2_152 VPWR VGND sg13g2_decap_8
X_064_ N2END[7] net65 VPWR VGND sg13g2_buf_1
XFILLER_9_53 VPWR VGND sg13g2_fill_1
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_7_255 VPWR VGND sg13g2_decap_8
X_047_ FrameStrobe[15] net39 VPWR VGND sg13g2_buf_1
XFILLER_4_214 VPWR VGND sg13g2_fill_2
XFILLER_6_54 VPWR VGND sg13g2_decap_8
Xoutput40 net40 FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
Xoutput51 net51 FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
Xoutput84 net84 S4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput73 net73 S4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput62 net62 S2BEG[5] VPWR VGND sg13g2_buf_1
Xoutput95 net95 SS4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput5 net5 FrameData_O[13] VPWR VGND sg13g2_buf_1
XFILLER_9_136 VPWR VGND sg13g2_decap_4
XFILLER_5_320 VPWR VGND sg13g2_decap_8
XFILLER_3_88 VPWR VGND sg13g2_fill_2
XFILLER_3_99 VPWR VGND sg13g2_decap_8
XFILLER_10_168 VPWR VGND sg13g2_decap_8
XFILLER_6_117 VPWR VGND sg13g2_decap_8
X_080_ N4END[7] net87 VPWR VGND sg13g2_buf_1
XFILLER_5_194 VPWR VGND sg13g2_decap_8
XFILLER_2_131 VPWR VGND sg13g2_decap_8
XFILLER_3_0 VPWR VGND sg13g2_decap_8
X_063_ N2MID[0] net64 VPWR VGND sg13g2_buf_1
XFILLER_9_65 VPWR VGND sg13g2_decap_4
XFILLER_9_21 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_11_285 VPWR VGND sg13g2_decap_8
XFILLER_11_274 VPWR VGND sg13g2_decap_8
XFILLER_7_234 VPWR VGND sg13g2_decap_8
X_046_ FrameStrobe[14] net38 VPWR VGND sg13g2_buf_1
XFILLER_4_259 VPWR VGND sg13g2_fill_1
X_029_ FrameData[29] net22 VPWR VGND sg13g2_buf_1
XFILLER_6_33 VPWR VGND sg13g2_decap_8
XFILLER_3_270 VPWR VGND sg13g2_fill_1
Xoutput41 net41 FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
Xoutput52 net52 FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
XFILLER_9_329 VPWR VGND sg13g2_decap_8
Xoutput6 net6 FrameData_O[14] VPWR VGND sg13g2_buf_1
Xoutput30 net30 FrameData_O[7] VPWR VGND sg13g2_buf_1
XFILLER_8_373 VPWR VGND sg13g2_decap_4
Xoutput96 net96 SS4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput74 net74 S4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput85 net85 S4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput63 net63 S2BEG[6] VPWR VGND sg13g2_buf_1
.ends

