* NGSPICE file created from RegFile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

.subckt RegFile E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E1END[0] E1END[1] E1END[2] E1END[3]
+ E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3] E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7] E2BEGb[0]
+ E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4] E2BEGb[5] E2BEGb[6] E2BEGb[7] E2END[0] E2END[1]
+ E2END[2] E2END[3] E2END[4] E2END[5] E2END[6] E2END[7] E2MID[0] E2MID[1] E2MID[2]
+ E2MID[3] E2MID[4] E2MID[5] E2MID[6] E2MID[7] E6BEG[0] E6BEG[10] E6BEG[11] E6BEG[1]
+ E6BEG[2] E6BEG[3] E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8] E6BEG[9] E6END[0]
+ E6END[10] E6END[11] E6END[1] E6END[2] E6END[3] E6END[4] E6END[5] E6END[6] E6END[7]
+ E6END[8] E6END[9] EE4BEG[0] EE4BEG[10] EE4BEG[11] EE4BEG[12] EE4BEG[13] EE4BEG[14]
+ EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4] EE4BEG[5] EE4BEG[6] EE4BEG[7]
+ EE4BEG[8] EE4BEG[9] EE4END[0] EE4END[10] EE4END[11] EE4END[12] EE4END[13] EE4END[14]
+ EE4END[15] EE4END[1] EE4END[2] EE4END[3] EE4END[4] EE4END[5] EE4END[6] EE4END[7]
+ EE4END[8] EE4END[9] FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4]
+ N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5]
+ N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6]
+ N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7]
+ N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2]
+ N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12]
+ NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5]
+ NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] NN4END[0] NN4END[10] NN4END[11] NN4END[12]
+ NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3] NN4END[4] NN4END[5]
+ NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S1END[0]
+ S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5]
+ S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6]
+ S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7]
+ S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4BEG[0]
+ S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3]
+ S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] S4END[0] S4END[10] S4END[11]
+ S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5]
+ S4END[6] S4END[7] S4END[8] S4END[9] SS4BEG[0] SS4BEG[10] SS4BEG[11] SS4BEG[12] SS4BEG[13]
+ SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4] SS4BEG[5] SS4BEG[6]
+ SS4BEG[7] SS4BEG[8] SS4BEG[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13]
+ SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6]
+ SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR W1BEG[0] W1BEG[1] W1BEG[2]
+ W1BEG[3] W1END[0] W1END[1] W1END[2] W1END[3] W2BEG[0] W2BEG[1] W2BEG[2] W2BEG[3]
+ W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0] W2BEGb[1] W2BEGb[2] W2BEGb[3] W2BEGb[4]
+ W2BEGb[5] W2BEGb[6] W2BEGb[7] W2END[0] W2END[1] W2END[2] W2END[3] W2END[4] W2END[5]
+ W2END[6] W2END[7] W2MID[0] W2MID[1] W2MID[2] W2MID[3] W2MID[4] W2MID[5] W2MID[6]
+ W2MID[7] W6BEG[0] W6BEG[10] W6BEG[11] W6BEG[1] W6BEG[2] W6BEG[3] W6BEG[4] W6BEG[5]
+ W6BEG[6] W6BEG[7] W6BEG[8] W6BEG[9] W6END[0] W6END[10] W6END[11] W6END[1] W6END[2]
+ W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8] W6END[9] WW4BEG[0] WW4BEG[10]
+ WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15] WW4BEG[1] WW4BEG[2] WW4BEG[3]
+ WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8] WW4BEG[9] WW4END[0] WW4END[10]
+ WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15] WW4END[1] WW4END[2] WW4END[3]
+ WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8] WW4END[9]
XTAP_TAPCELL_ROW_65_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2037_ net621 net901 _0899_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__mux2_2
X_2106_ net600 net855 _0918_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__mux2_1
XFILLER_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2939_ Inst_RegFile_switch_matrix.JW2BEG4 VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_20_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold362 Inst_RegFile_32x4.mem\[23\]\[1\] VGND VGND VPWR VPWR net937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 Inst_RegFile_32x4.mem\[21\]\[2\] VGND VGND VPWR VPWR net926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold340 Inst_RegFile_32x4.mem\[7\]\[2\] VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_60_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_202 _1033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1270_ _0239_ _0240_ net675 VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1606_ net644 net634 net668 net640 Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q
+ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__mux4_1
X_2655_ net761 net738 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2724_ clknet_4_7_0_UserCLK_regs _0126_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1399_ net66 net8 net111 net122 Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q
+ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__mux4_2
X_2586_ net767 net719 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1537_ Inst_RegFile_32x4.mem\[18\]\[3\] Inst_RegFile_32x4.mem\[19\]\[3\] net609 VGND
+ VGND VPWR VPWR _0490_ sky130_fd_sc_hd__mux2_1
X_1468_ _0424_ _0425_ net413 VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__mux2_1
XFILLER_70_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout672 net673 VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__buf_2
XFILLER_37_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout694 net695 VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__clkbuf_2
Xfanout661 net662 VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__clkbuf_4
Xfanout650 _0163_ VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__clkbuf_2
Xfanout683 net684 VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__clkbuf_4
X_2440_ net750 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1253_ net73 net101 Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q VGND VGND VPWR VPWR
+ _0224_ sky130_fd_sc_hd__mux2_1
X_2371_ net757 net692 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1322_ net675 _0288_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__or2_1
X_1184_ net68 net10 net112 net124 Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q
+ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_47_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput286 net286 VGND VGND VPWR VPWR NN4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput264 net264 VGND VGND VPWR VPWR N4BEG[12] sky130_fd_sc_hd__buf_2
X_2569_ net749 net714 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput275 net275 VGND VGND VPWR VPWR N4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput253 net253 VGND VGND VPWR VPWR N2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput242 net242 VGND VGND VPWR VPWR N1BEG[1] sky130_fd_sc_hd__buf_4
Xoutput231 net231 VGND VGND VPWR VPWR FrameStrobe_O[19] sky130_fd_sc_hd__buf_2
Xoutput220 net220 VGND VGND VPWR VPWR FrameData_O[9] sky130_fd_sc_hd__buf_2
X_2638_ net747 net738 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2707_ clknet_4_2_0_UserCLK_regs _0109_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput297 net297 VGND VGND VPWR VPWR S2BEG[0] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_73_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1871_ net61 Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q
+ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_44_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1940_ _1018_ _0708_ _0824_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__a21oi_2
XFILLER_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2423_ net772 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1236_ _0961_ _0208_ Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q VGND VGND VPWR VPWR
+ _0209_ sky130_fd_sc_hd__o21a_1
X_2354_ net743 net691 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2285_ net748 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_29_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1305_ Inst_RegFile_32x4.mem\[22\]\[1\] Inst_RegFile_32x4.mem\[23\]\[1\] net628 VGND
+ VGND VPWR VPWR _0274_ sky130_fd_sc_hd__mux2_1
X_1167_ _0142_ _0143_ Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q VGND VGND VPWR VPWR
+ _0144_ sky130_fd_sc_hd__mux2_1
XFILLER_64_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1098_ Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__inv_1
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2070_ _0893_ _0909_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__nand2_2
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2972_ WW4END[13] VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__buf_1
X_1785_ net651 net644 Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q VGND VGND VPWR VPWR
+ _0713_ sky130_fd_sc_hd__mux2_1
X_1854_ Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q _0768_ Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q
+ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__a21bo_1
X_1923_ _0807_ _0806_ Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q VGND VGND VPWR VPWR
+ _0808_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2406_ net753 net695 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_72_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2337_ net759 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_44_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2268_ net765 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1219_ _0178_ Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q _0180_ _0191_ VGND VGND
+ VPWR VPWR _0192_ sky130_fd_sc_hd__a31o_4
X_2199_ clknet_4_10_0_UserCLK_regs _0023_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_60_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_5 E6END[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1570_ Inst_RegFile_32x4.mem\[0\]\[2\] Inst_RegFile_32x4.mem\[1\]\[2\] net606 VGND
+ VGND VPWR VPWR _0521_ sky130_fd_sc_hd__mux2_1
XFILLER_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2122_ net615 net928 _0921_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__mux2_4
X_2053_ net602 net847 _0905_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__mux2_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2955_ W6END[6] VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__buf_1
X_1837_ _0755_ _0754_ Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q VGND VGND VPWR VPWR
+ _0756_ sky130_fd_sc_hd__mux2_4
X_1906_ net635 net685 Inst_RegFile_switch_matrix.E2BEG1 net397 Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.S1BEG2
+ sky130_fd_sc_hd__mux4_2
X_1768_ net23 net777 net92 net120 Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q
+ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__mux4_1
X_2886_ Inst_RegFile_switch_matrix.JS2BEG4 VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__buf_6
X_1699_ Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q _0636_ VGND VGND VPWR VPWR _0637_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_68_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput131 W2MID[4] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
Xinput120 W2END[1] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_2
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1622_ Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q _0569_ VGND VGND VPWR VPWR _0570_
+ sky130_fd_sc_hd__nor2_1
X_2740_ net15 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_1
XFILLER_31_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2671_ clknet_4_12_0_UserCLK_regs Inst_RegFile_32x4.AD_comb\[1\] VGND VGND VPWR VPWR
+ Inst_RegFile_32x4.AD_reg\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1484_ Inst_RegFile_32x4.mem\[16\]\[0\] Inst_RegFile_32x4.mem\[17\]\[0\] net610 VGND
+ VGND VPWR VPWR _0441_ sky130_fd_sc_hd__mux2_1
X_1553_ Inst_RegFile_32x4.mem\[0\]\[3\] Inst_RegFile_32x4.mem\[1\]\[3\] net607 VGND
+ VGND VPWR VPWR _0506_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2036_ net617 net923 _0899_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__mux2_2
X_2105_ _0889_ _0909_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__nand2_4
XFILLER_50_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2938_ Inst_RegFile_switch_matrix.JW2BEG3 VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__buf_1
XFILLER_10_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold330 Inst_RegFile_32x4.mem\[28\]\[2\] VGND VGND VPWR VPWR net905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 Inst_RegFile_32x4.mem\[0\]\[2\] VGND VGND VPWR VPWR net916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 Inst_RegFile_32x4.mem\[25\]\[3\] VGND VGND VPWR VPWR net938 sky130_fd_sc_hd__dlygate4sd3_1
X_2869_ NN4END[11] VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__clkbuf_2
Xhold352 Inst_RegFile_32x4.mem\[22\]\[3\] VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 net679 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2723_ clknet_4_3_0_UserCLK_regs _0125_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1605_ net688 net670 net657 net653 Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q
+ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__mux4_2
X_2585_ net768 net718 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2654_ net762 net738 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1536_ Inst_RegFile_32x4.mem\[16\]\[3\] Inst_RegFile_32x4.mem\[17\]\[3\] net609 VGND
+ VGND VPWR VPWR _0489_ sky130_fd_sc_hd__mux2_1
XFILLER_8_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1398_ _0358_ _0357_ _0359_ _0945_ _0941_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__a221o_1
X_1467_ Inst_RegFile_32x4.mem\[14\]\[0\] Inst_RegFile_32x4.mem\[15\]\[0\] net410 VGND
+ VGND VPWR VPWR _0425_ sky130_fd_sc_hd__mux2_1
XFILLER_35_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2019_ net611 net815 _0892_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout640 net641 VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__clkbuf_4
Xfanout651 net652 VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__buf_2
XFILLER_73_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout684 _0363_ VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__buf_8
XFILLER_33_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout695 net58 VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__clkbuf_2
Xfanout673 AD0 VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__buf_2
Xfanout662 net663 VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1252_ Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q net129 Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q
+ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__o21a_1
X_2370_ net758 net692 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1321_ Inst_RegFile_32x4.mem\[2\]\[2\] Inst_RegFile_32x4.mem\[3\]\[2\] net627 VGND
+ VGND VPWR VPWR _0288_ sky130_fd_sc_hd__mux2_1
XFILLER_64_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1183_ net80 net123 net112 Inst_RegFile_switch_matrix.JS2BEG3 Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__mux4_2
XFILLER_24_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2706_ clknet_4_8_0_UserCLK_regs _0108_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput232 net232 VGND VGND VPWR VPWR FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput221 net221 VGND VGND VPWR VPWR FrameStrobe_O[0] sky130_fd_sc_hd__buf_2
Xoutput287 net287 VGND VGND VPWR VPWR NN4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput265 net265 VGND VGND VPWR VPWR N4BEG[13] sky130_fd_sc_hd__buf_2
X_2568_ net750 net714 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput276 net276 VGND VGND VPWR VPWR N4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput254 net254 VGND VGND VPWR VPWR N2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput210 net210 VGND VGND VPWR VPWR FrameData_O[29] sky130_fd_sc_hd__buf_2
Xoutput243 net243 VGND VGND VPWR VPWR N1BEG[2] sky130_fd_sc_hd__buf_4
X_2499_ net42 net709 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2637_ net49 net740 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1519_ Inst_RegFile_32x4.mem\[0\]\[1\] Inst_RegFile_32x4.mem\[1\]\[1\] net606 VGND
+ VGND VPWR VPWR _0474_ sky130_fd_sc_hd__mux2_1
Xoutput298 net298 VGND VGND VPWR VPWR S2BEG[1] sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1870_ net780 Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q VGND VGND VPWR VPWR _0784_
+ sky130_fd_sc_hd__nand2b_1
X_2353_ net744 net691 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2422_ net773 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1235_ net646 net679 net636 net640 Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q
+ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__mux4_1
X_1166_ net89 net97 net113 net115 Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q
+ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__mux4_1
XFILLER_49_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2284_ net751 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1304_ _0271_ _0272_ net662 VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__mux2_1
XFILLER_52_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1097_ Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__inv_1
X_1999_ Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q _0740_ VGND VGND VPWR VPWR _0881_
+ sky130_fd_sc_hd__or2_1
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_6_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_6_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1922_ _0740_ Inst_RegFile_switch_matrix.JN2BEG7 Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q
+ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__mux2_1
X_2971_ WW4END[12] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__buf_1
X_1784_ net84 net779 net112 net688 Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q
+ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__mux4_1
X_1853_ Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q _0146_ _0769_ Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q
+ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_12_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2336_ net39 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2405_ net755 net695 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2267_ net766 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_55_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1149_ net21 net95 net114 net123 Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q
+ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__mux4_1
XFILLER_52_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1218_ _0977_ _0188_ _0190_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__a21oi_1
X_2198_ clknet_4_8_0_UserCLK_regs _0022_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_6 E6END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2121_ net599 net852 _0921_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__mux2_1
X_2052_ _0889_ _0904_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__nand2_4
XFILLER_62_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1905_ net641 _0437_ Inst_RegFile_switch_matrix.E2BEG2 _0803_ Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.S1BEG3
+ sky130_fd_sc_hd__mux4_1
X_2885_ Inst_RegFile_switch_matrix.JS2BEG3 VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__buf_1
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2954_ W6END[5] VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__buf_1
X_1836_ net679 net636 net667 net640 Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q
+ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__mux4_1
X_1698_ net687 net669 net651 net644 Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q
+ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__mux4_1
X_1767_ net64 net80 net779 net6 Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q
+ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2319_ net746 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_68_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput110 S4END[3] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput132 W2MID[5] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
Xinput121 W2END[2] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_4
XFILLER_72_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1621_ net77 net19 net105 Inst_RegFile_switch_matrix.JN2BEG6 Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__mux4_1
X_1552_ Inst_RegFile_32x4.mem\[2\]\[3\] Inst_RegFile_32x4.mem\[3\]\[3\] net607 VGND
+ VGND VPWR VPWR _0505_ sky130_fd_sc_hd__mux2_1
X_2670_ clknet_4_7_0_UserCLK_regs Inst_RegFile_32x4.AD_comb\[0\] VGND VGND VPWR VPWR
+ Inst_RegFile_32x4.AD_reg\[0\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2104_ net612 net849 _0917_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__mux2_1
X_1483_ net619 _0427_ _0439_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_65_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2035_ net600 net841 _0899_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__mux2_1
X_2937_ Inst_RegFile_switch_matrix.JW2BEG2 VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__buf_4
XFILLER_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2868_ NN4END[10] VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__buf_2
X_2799_ net42 VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__buf_1
X_1819_ _0738_ _0739_ _0741_ Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q VGND VGND
+ VPWR VPWR _0742_ sky130_fd_sc_hd__a22o_1
Xhold331 Inst_RegFile_32x4.mem\[16\]\[2\] VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 Inst_RegFile_32x4.mem\[28\]\[1\] VGND VGND VPWR VPWR net917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 Inst_RegFile_32x4.mem\[31\]\[1\] VGND VGND VPWR VPWR net928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold320 Inst_RegFile_32x4.mem\[14\]\[3\] VGND VGND VPWR VPWR net895 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_204 net777 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2722_ clknet_4_7_0_UserCLK_regs _0124_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2584_ net770 net718 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2653_ net35 net741 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1604_ Inst_RegFile_32x4.BD_comb\[2\] Inst_RegFile_32x4.BD_reg\[2\] Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q
+ VGND VGND VPWR VPWR BD2 sky130_fd_sc_hd__mux2_4
X_1535_ Inst_RegFile_32x4.BD_comb\[1\] Inst_RegFile_32x4.BD_reg\[1\] Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q
+ VGND VGND VPWR VPWR BD1 sky130_fd_sc_hd__mux2_4
X_1397_ net81 net113 Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q VGND VGND VPWR VPWR
+ _0359_ sky130_fd_sc_hd__mux2_1
X_1466_ Inst_RegFile_32x4.mem\[12\]\[0\] Inst_RegFile_32x4.mem\[13\]\[0\] net410 VGND
+ VGND VPWR VPWR _0424_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2018_ net620 net813 _0892_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__mux2_1
Xfanout641 BD3 VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__buf_4
Xfanout685 _0348_ VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__clkbuf_4
Xfanout652 net655 VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__buf_8
Xfanout663 _0136_ VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__buf_4
Xfanout674 _0135_ VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__buf_6
Xfanout630 net632 VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__clkbuf_4
XFILLER_73_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout696 net697 VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__buf_2
XFILLER_33_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1320_ Inst_RegFile_32x4.mem\[0\]\[2\] Inst_RegFile_32x4.mem\[1\]\[2\] net627 VGND
+ VGND VPWR VPWR _0287_ sky130_fd_sc_hd__mux2_1
XFILLER_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1251_ _0216_ _0218_ _0221_ _0939_ _0937_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__a221o_1
X_1182_ _0154_ _0152_ _0157_ _0975_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JS2BEG3
+ sky130_fd_sc_hd__a22o_4
XTAP_TAPCELL_ROW_39_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput200 net200 VGND VGND VPWR VPWR FrameData_O[1] sky130_fd_sc_hd__buf_2
X_2636_ net46 net740 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_30_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2705_ clknet_4_11_0_UserCLK_regs _0107_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput222 net222 VGND VGND VPWR VPWR FrameStrobe_O[10] sky130_fd_sc_hd__buf_2
Xoutput233 net233 VGND VGND VPWR VPWR FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
Xoutput288 net288 VGND VGND VPWR VPWR NN4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput277 net277 VGND VGND VPWR VPWR NN4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput266 net266 VGND VGND VPWR VPWR N4BEG[14] sky130_fd_sc_hd__buf_2
X_2567_ net752 net714 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput244 net244 VGND VGND VPWR VPWR N1BEG[3] sky130_fd_sc_hd__buf_4
X_1449_ net88 net98 net90 net688 Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q
+ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__mux4_1
Xoutput255 net255 VGND VGND VPWR VPWR N2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput211 net211 VGND VGND VPWR VPWR FrameData_O[2] sky130_fd_sc_hd__buf_2
X_2498_ net41 net709 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1518_ Inst_RegFile_32x4.mem\[2\]\[1\] Inst_RegFile_32x4.mem\[3\]\[1\] net606 VGND
+ VGND VPWR VPWR _0473_ sky130_fd_sc_hd__mux2_1
Xoutput299 net299 VGND VGND VPWR VPWR S2BEG[2] sky130_fd_sc_hd__buf_6
XFILLER_67_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_14_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_14_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2352_ net745 net691 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2283_ net763 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2421_ net29 net700 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1303_ Inst_RegFile_32x4.mem\[18\]\[1\] Inst_RegFile_32x4.mem\[19\]\[1\] net631 VGND
+ VGND VPWR VPWR _0272_ sky130_fd_sc_hd__mux2_1
XFILLER_6_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1234_ Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q _0206_ VGND VGND VPWR VPWR _0207_
+ sky130_fd_sc_hd__or2_1
X_1165_ net61 net69 net780 net11 Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q
+ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__mux4_1
XFILLER_49_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1096_ Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__inv_1
XFILLER_52_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2619_ net766 net724 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1998_ Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q _0876_ _0879_ VGND VGND VPWR VPWR
+ _0880_ sky130_fd_sc_hd__a21o_1
XFILLER_68_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1852_ Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q net679 VGND VGND VPWR VPWR _0769_
+ sky130_fd_sc_hd__nor2_1
XFILLER_34_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1921_ Inst_RegFile_switch_matrix.JS2BEG7 Inst_RegFile_switch_matrix.JW2BEG7 Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q
+ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__mux2_1
X_2970_ WW4END[11] VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__buf_1
X_1783_ _0702_ _0711_ Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.W6BEG1 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2266_ net767 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2335_ net38 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2404_ net756 net695 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1148_ net61 net67 net79 net9 Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q
+ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__mux4_1
X_1079_ net75 VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__inv_1
XFILLER_25_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1217_ Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q _0189_ Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q
+ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__a21o_1
X_2197_ clknet_4_10_0_UserCLK_regs _0021_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_7 E6END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2120_ _0893_ _0895_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__nand2_4
XFILLER_66_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2051_ _0830_ _0901_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__nor2_8
X_1835_ _0707_ _0708_ _0147_ _0372_ Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q
+ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__mux4_2
X_2884_ Inst_RegFile_switch_matrix.JS2BEG2 VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_60_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1904_ net22 net108 net93 net673 Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.S4BEG0 sky130_fd_sc_hd__mux4_1
X_2953_ W6END[4] VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__clkbuf_1
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1697_ _0632_ _0630_ _0635_ _0993_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E2BEG1
+ sky130_fd_sc_hd__a22o_4
X_1766_ Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q _0695_ Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q
+ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_68_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ net50 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2249_ clknet_4_11_0_UserCLK_regs _0073_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[21\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput111 SS4END[0] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_4
Xinput100 S2MID[1] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__buf_2
Xinput133 W2MID[6] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
Xinput122 W2END[3] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__buf_2
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1620_ Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q _0567_ Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q
+ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__o21ai_1
X_1482_ _0438_ _0435_ Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q VGND VGND VPWR VPWR
+ _0439_ sky130_fd_sc_hd__mux2_4
X_1551_ net619 _0503_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__or2_1
X_2103_ net621 net897 _0917_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_65_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2034_ _0891_ _0898_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__nand2_4
X_2798_ net41 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__buf_1
X_1818_ _0372_ _0740_ Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q VGND VGND VPWR VPWR
+ _0741_ sky130_fd_sc_hd__mux2_1
X_2936_ Inst_RegFile_switch_matrix.JW2BEG1 VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_20_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold310 Inst_RegFile_32x4.mem\[2\]\[3\] VGND VGND VPWR VPWR net885 sky130_fd_sc_hd__dlygate4sd3_1
X_2867_ NN4END[9] VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__clkbuf_2
X_1749_ net676 net635 net666 net409 Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q
+ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__mux4_1
Xhold354 Inst_RegFile_32x4.mem\[18\]\[1\] VGND VGND VPWR VPWR net929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 Inst_RegFile_32x4.mem\[10\]\[2\] VGND VGND VPWR VPWR net918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 Inst_RegFile_32x4.mem\[8\]\[1\] VGND VGND VPWR VPWR net896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 Inst_RegFile_32x4.mem\[26\]\[1\] VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_205 net777 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_48_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2652_ net34 net741 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2721_ clknet_4_3_0_UserCLK_regs _0123_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2583_ net772 net719 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1603_ _0536_ _0553_ _0439_ VGND VGND VPWR VPWR Inst_RegFile_32x4.BD_comb\[2\] sky130_fd_sc_hd__mux2_4
X_1465_ _0421_ _0422_ net413 VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__mux2_1
X_1534_ _0464_ _0439_ _0472_ _0487_ _0488_ VGND VGND VPWR VPWR Inst_RegFile_32x4.BD_comb\[1\]
+ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_66_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1396_ Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q net121 Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q
+ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__o21a_1
X_2017_ net615 net907 _0892_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__mux2_4
X_2919_ SS4END[9] VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout664 net668 VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__buf_6
Xfanout653 net654 VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__buf_6
XFILLER_58_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout686 net136 VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__clkbuf_4
Xfanout697 net58 VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__clkbuf_2
Xfanout642 _0388_ VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__buf_4
Xfanout631 net632 VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__clkbuf_2
Xfanout675 _0135_ VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__buf_6
Xfanout620 net623 VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__clkbuf_2
XFILLER_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1250_ _0216_ _0218_ _0221_ _0939_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E2BEG6
+ sky130_fd_sc_hd__a22o_1
X_1181_ _0155_ _0156_ Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q VGND VGND VPWR VPWR
+ _0157_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput223 net223 VGND VGND VPWR VPWR FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
Xoutput234 net234 VGND VGND VPWR VPWR FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
Xoutput212 net212 VGND VGND VPWR VPWR FrameData_O[30] sky130_fd_sc_hd__buf_2
Xoutput201 net201 VGND VGND VPWR VPWR FrameData_O[20] sky130_fd_sc_hd__buf_2
X_2635_ net763 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_30_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2704_ clknet_4_14_0_UserCLK_regs _0106_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput278 net278 VGND VGND VPWR VPWR NN4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput289 net289 VGND VGND VPWR VPWR NN4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput267 net267 VGND VGND VPWR VPWR N4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput256 net256 VGND VGND VPWR VPWR N2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput245 net245 VGND VGND VPWR VPWR N2BEG[0] sky130_fd_sc_hd__buf_4
X_1448_ Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q _0406_ VGND VGND VPWR VPWR _0407_
+ sky130_fd_sc_hd__and2b_1
X_2566_ net753 net714 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2497_ net759 net706 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1517_ net619 _0471_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__or2_1
XFILLER_70_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1379_ _0331_ _0193_ _0335_ _0229_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__a31o_1
XFILLER_23_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2420_ net28 net700 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_24_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1233_ net117 net672 net659 net653 Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q
+ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__mux4_1
X_2282_ net27 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2351_ net746 net690 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1302_ Inst_RegFile_32x4.mem\[16\]\[1\] Inst_RegFile_32x4.mem\[17\]\[1\] net631 VGND
+ VGND VPWR VPWR _0271_ sky130_fd_sc_hd__mux2_1
X_1164_ _0972_ _0140_ Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q VGND VGND VPWR VPWR
+ _0141_ sky130_fd_sc_hd__o21a_1
X_1095_ Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__inv_2
X_1997_ Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q _0878_ Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q
+ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2618_ net767 net724 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2549_ net29 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_7_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1851_ _0372_ _0767_ Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q VGND VGND VPWR VPWR
+ _0768_ sky130_fd_sc_hd__mux2_1
X_1920_ net423 Inst_RegFile_switch_matrix.JW2BEG3 _0804_ _0805_ Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q
+ Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.N1BEG0
+ sky130_fd_sc_hd__mux4_1
X_1782_ _0710_ _0709_ Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q VGND VGND VPWR VPWR
+ _0711_ sky130_fd_sc_hd__mux2_1
X_2403_ net757 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_12_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2265_ net769 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2334_ net762 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1216_ net72 net14 net100 net128 Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q
+ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__mux4_1
X_2196_ clknet_4_8_0_UserCLK_regs _0020_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1147_ _0957_ _1037_ Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q VGND VGND VPWR VPWR
+ _1038_ sky130_fd_sc_hd__o21a_1
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1078_ Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__inv_1
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_8 E6END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_2_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_2_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
X_2050_ net614 net872 _0903_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__mux2_1
XFILLER_47_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2952_ W6END[3] VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__buf_1
XFILLER_15_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1834_ Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q _0752_ Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q
+ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_60_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1765_ net686 net423 net658 net645 Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q
+ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__mux4_1
X_1903_ net778 net94 net109 net660 Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.S4BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_30_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2883_ Inst_RegFile_switch_matrix.JS2BEG1 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__buf_4
X_1696_ _0633_ _0634_ _0992_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ net748 net734 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_38_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2179_ clknet_4_0_0_UserCLK_regs _0003_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[24\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2248_ clknet_4_9_0_UserCLK_regs _0072_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[21\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput112 SS4END[1] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_2
Xinput101 S2MID[2] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_2
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput134 W2MID[7] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
Xinput123 W2END[4] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_4
XFILLER_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1481_ net65 net93 _0436_ _0437_ Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q
+ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__mux4_2
X_1550_ _0499_ _0502_ net642 VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2102_ net616 net827 _0917_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__mux2_1
X_2033_ _0829_ _0897_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__nor2_8
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2935_ Inst_RegFile_switch_matrix.JW2BEG0 VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__clkbuf_2
X_2797_ net40 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_1
X_1748_ Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q _0679_ VGND VGND VPWR VPWR _0680_
+ sky130_fd_sc_hd__or2_1
X_1817_ net63 net91 net5 net140 Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q
+ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__mux4_2
Xhold311 Inst_RegFile_32x4.mem\[19\]\[1\] VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_20_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold333 Inst_RegFile_32x4.mem\[1\]\[2\] VGND VGND VPWR VPWR net908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 Inst_RegFile_32x4.mem\[22\]\[1\] VGND VGND VPWR VPWR net919 sky130_fd_sc_hd__dlygate4sd3_1
X_2866_ NN4END[8] VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__clkbuf_2
Xhold322 Inst_RegFile_32x4.mem\[20\]\[2\] VGND VGND VPWR VPWR net897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold300 Inst_RegFile_32x4.mem\[5\]\[1\] VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__dlygate4sd3_1
X_1679_ net93 net109 net112 net121 Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q
+ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__mux4_1
Xhold355 Inst_RegFile_32x4.mem\[12\]\[0\] VGND VGND VPWR VPWR net930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_41_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_206 net777 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2582_ net773 net719 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2651_ net33 net740 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2720_ clknet_4_2_0_UserCLK_regs _0122_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1602_ _0540_ _0545_ _0552_ net619 VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__o2bb2a_1
X_1395_ _0351_ _0353_ _0356_ _0944_ _0942_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__a221o_1
X_1464_ Inst_RegFile_32x4.mem\[10\]\[0\] Inst_RegFile_32x4.mem\[11\]\[0\] net608 VGND
+ VGND VPWR VPWR _0422_ sky130_fd_sc_hd__mux2_1
X_1533_ _0416_ _0479_ _0439_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__o21ba_1
XFILLER_67_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2016_ net599 net826 _0892_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__mux2_1
X_2918_ SS4END[8] VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__clkbuf_2
XFILLER_23_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2849_ N4END[7] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkbuf_2
Xfanout665 net668 VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout676 net678 VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__buf_2
Xfanout654 net655 VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__buf_2
Xfanout632 A_ADR0 VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__buf_6
Xfanout687 net135 VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__clkbuf_4
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout698 net699 VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__buf_2
Xfanout610 B_ADR0 VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__clkbuf_2
Xfanout643 _0388_ VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout621 net622 VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__clkbuf_2
XFILLER_73_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1180_ net778 net95 net107 net123 Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q
+ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_47_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput224 net224 VGND VGND VPWR VPWR FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
Xoutput235 net235 VGND VGND VPWR VPWR FrameStrobe_O[4] sky130_fd_sc_hd__buf_2
Xoutput213 net213 VGND VGND VPWR VPWR FrameData_O[31] sky130_fd_sc_hd__buf_2
Xoutput257 net257 VGND VGND VPWR VPWR N2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput246 net246 VGND VGND VPWR VPWR N2BEG[1] sky130_fd_sc_hd__buf_4
Xoutput268 net268 VGND VGND VPWR VPWR N4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput202 net202 VGND VGND VPWR VPWR FrameData_O[21] sky130_fd_sc_hd__buf_2
X_2565_ net44 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2634_ net776 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2703_ clknet_4_11_0_UserCLK_regs _0105_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1516_ _0467_ _0470_ net642 VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__mux2_4
Xoutput279 net279 VGND VGND VPWR VPWR NN4BEG[11] sky130_fd_sc_hd__buf_2
X_1447_ net62 net70 net779 net12 Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q
+ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_38_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2496_ net760 net706 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1378_ _0193_ _0342_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__nor2_1
XFILLER_63_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2281_ net48 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2350_ net747 net690 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1301_ _0265_ _0266_ net408 _0269_ net395 VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__a221o_1
X_1232_ _0164_ _0200_ _0204_ _0193_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__a211o_1
X_1094_ Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__inv_2
X_1163_ net647 net680 net636 net641 Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q
+ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__mux4_1
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1996_ _0877_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_15_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2617_ net768 net722 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2548_ net28 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_7_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2479_ net746 net707 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_43_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload0 clknet_4_0_0_UserCLK_regs VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinv_2
XFILLER_59_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_10_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_10_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_61_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1781_ net678 net634 net665 net638 Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q
+ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__mux4_1
X_1850_ net69 net11 net114 net125 Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q
+ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__mux4_1
X_2333_ net764 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2402_ net758 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2264_ net770 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1146_ net679 net636 net668 net640 Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q
+ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__mux4_2
X_1215_ net13 net127 net99 Inst_RegFile_switch_matrix.JW2BEG5 Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__mux4_1
X_2195_ clknet_4_5_0_UserCLK_regs _0019_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[28\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1077_ Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__inv_2
X_1979_ Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q _0863_ VGND VGND VPWR VPWR _0864_
+ sky130_fd_sc_hd__nor2_1
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 E6END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1902_ net91 net686 net110 net653 Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.S4BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_62_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2951_ W6END[2] VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__buf_1
XFILLER_15_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1833_ _0751_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__inv_2
X_1764_ _1009_ _0693_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__or2_1
X_2882_ Inst_RegFile_switch_matrix.JS2BEG0 VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__buf_1
X_1695_ net59 net65 net81 net84 Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q
+ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__mux4_1
X_2316_ net751 net734 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1129_ _0966_ _1020_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__or2_4
XFILLER_38_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2247_ clknet_4_11_0_UserCLK_regs _0071_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[20\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2178_ clknet_4_5_0_UserCLK_regs _0002_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[24\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_51_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput113 SS4END[2] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_2
Xinput102 S2MID[3] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput135 W6END[0] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput124 W2END[5] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1480_ net76 net18 net104 net132 Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q
+ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_65_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2032_ _0810_ _0820_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__or2_4
X_2101_ net600 net835 _0917_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__mux2_1
XFILLER_62_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2934_ Inst_RegFile_switch_matrix.W1BEG3 VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_20_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2865_ NN4END[7] VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkbuf_2
X_2796_ net39 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__buf_1
X_1816_ Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q _0146_ Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q
+ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1678_ net59 net7 net65 net778 Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q
+ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__mux4_1
X_1747_ net686 net423 net658 net645 Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q
+ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__mux4_1
Xhold312 Inst_RegFile_32x4.mem\[17\]\[3\] VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 Inst_RegFile_32x4.mem\[25\]\[1\] VGND VGND VPWR VPWR net931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 Inst_RegFile_32x4.mem\[0\]\[1\] VGND VGND VPWR VPWR net898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 Inst_RegFile_32x4.mem\[8\]\[3\] VGND VGND VPWR VPWR net920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold301 Inst_RegFile_32x4.mem\[29\]\[3\] VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 Inst_RegFile_32x4.mem\[24\]\[2\] VGND VGND VPWR VPWR net909 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_207 net777 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2581_ net774 net720 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2650_ net32 net740 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_12_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1532_ net619 _0486_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__or2_1
X_1601_ _0548_ _0551_ net642 VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__mux2_4
X_1394_ _0351_ _0353_ _0356_ _0944_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E2BEG4
+ sky130_fd_sc_hd__a22o_1
X_1463_ Inst_RegFile_32x4.mem\[8\]\[0\] Inst_RegFile_32x4.mem\[9\]\[0\] net608 VGND
+ VGND VPWR VPWR _0421_ sky130_fd_sc_hd__mux2_1
X_2015_ _0831_ _0891_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__nand2_4
X_2917_ SS4END[7] VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2848_ N4END[6] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_2
Xfanout633 net634 VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__buf_8
X_2779_ net51 VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_2
Xfanout622 net623 VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__clkbuf_2
Xfanout600 net601 VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__buf_4
Xfanout611 _0887_ VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__clkbuf_2
Xfanout677 net678 VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__buf_8
Xfanout644 net645 VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__buf_4
Xfanout688 net118 VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__clkbuf_4
Xfanout666 net668 VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__buf_2
Xfanout699 FrameStrobe[7] VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__clkbuf_2
Xfanout655 AD2 VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__buf_8
XFILLER_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2702_ clknet_4_11_0_UserCLK_regs _0104_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput236 net236 VGND VGND VPWR VPWR FrameStrobe_O[5] sky130_fd_sc_hd__buf_2
Xoutput225 net225 VGND VGND VPWR VPWR FrameStrobe_O[13] sky130_fd_sc_hd__buf_2
Xoutput258 net258 VGND VGND VPWR VPWR N2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput247 net247 VGND VGND VPWR VPWR N2BEG[2] sky130_fd_sc_hd__buf_6
Xoutput269 net269 VGND VGND VPWR VPWR N4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput203 net203 VGND VGND VPWR VPWR FrameData_O[22] sky130_fd_sc_hd__buf_2
X_2633_ net48 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput214 net214 VGND VGND VPWR VPWR FrameData_O[3] sky130_fd_sc_hd__buf_2
X_2564_ net43 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2495_ net761 net706 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1515_ _0468_ _0469_ net412 VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__mux2_1
X_1446_ Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q _0404_ Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q
+ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__a21boi_2
XTAP_TAPCELL_ROW_38_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1377_ _0338_ _0341_ net650 VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__mux2_1
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2280_ net47 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1162_ Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q _0138_ VGND VGND VPWR VPWR _0139_
+ sky130_fd_sc_hd__or2_1
X_1300_ _0267_ _0268_ net663 VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__mux2_1
X_1231_ net661 _0203_ _0202_ net650 VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__o211a_1
XFILLER_64_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1093_ Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__inv_1
XFILLER_60_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2616_ net770 net722 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1995_ net79 net778 Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q VGND VGND VPWR VPWR
+ _0877_ sky130_fd_sc_hd__mux2_1
XFILLER_9_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2547_ net742 net717 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2478_ net747 net707 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1429_ Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q _0385_ _0387_ _0374_ VGND VGND VPWR
+ VPWR _0389_ sky130_fd_sc_hd__a31o_1
XFILLER_43_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload1 clknet_4_1_0_UserCLK_regs VGND VGND VPWR VPWR clkload1/X sky130_fd_sc_hd__clkbuf_8
XFILLER_59_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1780_ _0707_ _0708_ _0147_ _0372_ Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q
+ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__mux4_2
XFILLER_6_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2332_ net765 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2401_ net759 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1214_ _0183_ _0976_ _0185_ _0187_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JW2BEG5
+ sky130_fd_sc_hd__o22a_4
XFILLER_65_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1145_ _1035_ Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q VGND VGND VPWR VPWR _1036_
+ sky130_fd_sc_hd__or2_4
XFILLER_37_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2263_ net772 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_25_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2194_ clknet_4_5_0_UserCLK_regs _0018_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[28\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1076_ Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__inv_2
X_1978_ net77 net105 Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q VGND VGND VPWR VPWR
+ _0863_ sky130_fd_sc_hd__mux2_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1832_ net672 net653 net659 net422 Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q
+ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__mux4_1
X_2881_ Inst_RegFile_switch_matrix.S1BEG3 VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__buf_4
X_1901_ net92 net687 net107 net421 Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.S4BEG3 sky130_fd_sc_hd__mux4_1
X_2950_ net134 VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_2
X_1694_ net7 net93 net21 net121 Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q
+ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__mux4_1
X_1763_ net676 net635 net666 net409 Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q
+ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__mux4_1
X_2315_ net763 net737 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2246_ clknet_4_9_0_UserCLK_regs _0070_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[20\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1128_ net647 net679 net636 net641 Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q
+ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__mux4_2
X_1059_ Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__inv_2
XFILLER_53_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2177_ clknet_4_1_0_UserCLK_regs _0001_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[24\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_51_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput114 SS4END[3] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
Xinput103 S2MID[4] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput136 W6END[1] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput125 W2END[6] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__buf_1
XFILLER_44_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2100_ _0859_ _0909_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_65_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2031_ net611 net900 _0896_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__mux2_4
X_2795_ net761 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__buf_1
X_1815_ Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q net680 VGND VGND VPWR VPWR _0738_
+ sky130_fd_sc_hd__or2_1
XFILLER_30_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2864_ NN4END[6] VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__buf_2
X_1746_ _0674_ _0675_ _0678_ _1004_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E2BEG7
+ sky130_fd_sc_hd__a22o_1
X_1677_ _0988_ _0617_ Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q VGND VGND VPWR VPWR
+ _0618_ sky130_fd_sc_hd__o21a_1
Xhold357 Inst_RegFile_32x4.mem\[25\]\[2\] VGND VGND VPWR VPWR net932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 Inst_RegFile_32x4.mem\[3\]\[3\] VGND VGND VPWR VPWR net921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 Inst_RegFile_32x4.mem\[12\]\[3\] VGND VGND VPWR VPWR net888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 Inst_RegFile_32x4.mem\[10\]\[1\] VGND VGND VPWR VPWR net899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold302 Inst_RegFile_32x4.mem\[27\]\[1\] VGND VGND VPWR VPWR net877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 Inst_RegFile_32x4.mem\[18\]\[3\] VGND VGND VPWR VPWR net910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2229_ clknet_4_6_0_UserCLK_regs _0053_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_36_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 net777 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2580_ net775 net720 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_26_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1531_ _0482_ _0485_ net642 VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__mux2_1
X_1462_ net643 _0419_ _0416_ _0392_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__a211o_1
X_1600_ _0550_ _0549_ net681 VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__mux2_1
XFILLER_67_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1393_ _0354_ _0355_ _0943_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__mux2_4
XFILLER_50_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2014_ _0853_ _0857_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__nor2_8
XFILLER_23_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2916_ SS4END[6] VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__clkbuf_2
X_2778_ net747 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__buf_2
X_2847_ N4END[5] VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_2
X_1729_ _0658_ _0660_ _0663_ _1001_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JS2BEG7
+ sky130_fd_sc_hd__a22o_1
Xfanout667 net668 VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__buf_8
Xfanout656 net658 VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__buf_2
Xfanout634 BD2 VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__buf_8
Xfanout645 AD3 VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__buf_6
Xfanout623 _0875_ VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__clkbuf_2
Xfanout612 net614 VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__clkbuf_2
Xfanout601 net602 VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__buf_2
XFILLER_73_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout689 net117 VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout678 BD0 VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__buf_8
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2632_ net47 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_30_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2701_ clknet_4_11_0_UserCLK_regs _0103_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput237 net237 VGND VGND VPWR VPWR FrameStrobe_O[6] sky130_fd_sc_hd__buf_2
Xoutput259 net259 VGND VGND VPWR VPWR N2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput226 net226 VGND VGND VPWR VPWR FrameStrobe_O[14] sky130_fd_sc_hd__buf_2
X_1445_ net645 net678 net665 BD3 Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q
+ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__mux4_2
Xoutput248 net248 VGND VGND VPWR VPWR N2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput204 net204 VGND VGND VPWR VPWR FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput215 net215 VGND VGND VPWR VPWR FrameData_O[4] sky130_fd_sc_hd__buf_2
X_2563_ net42 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2494_ net762 net706 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1514_ Inst_RegFile_32x4.mem\[30\]\[1\] Inst_RegFile_32x4.mem\[31\]\[1\] net603 VGND
+ VGND VPWR VPWR _0469_ sky130_fd_sc_hd__mux2_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1376_ _0339_ _0340_ net674 VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__mux2_1
XFILLER_58_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1161_ net689 net672 net660 net654 Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q
+ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__mux4_1
X_1092_ Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__inv_2
X_1230_ Inst_RegFile_32x4.mem\[20\]\[0\] Inst_RegFile_32x4.mem\[21\]\[0\] net627 VGND
+ VGND VPWR VPWR _0203_ sky130_fd_sc_hd__mux2_1
XFILLER_60_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1994_ net107 Inst_RegFile_switch_matrix.JW2BEG1 Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q
+ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2615_ net772 net722 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2546_ net743 net717 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2477_ net49 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1428_ Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q _0385_ _0387_ _0374_ VGND VGND VPWR
+ VPWR _0388_ sky130_fd_sc_hd__a31oi_1
XFILLER_51_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1359_ Inst_RegFile_32x4.mem\[6\]\[3\] Inst_RegFile_32x4.mem\[7\]\[3\] net630 VGND
+ VGND VPWR VPWR _0324_ sky130_fd_sc_hd__mux2_1
Xclkload2 clknet_4_2_0_UserCLK_regs VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_4
XFILLER_59_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2400_ net760 net695 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1213_ Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q _0186_ Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q
+ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__a21o_1
X_2331_ net766 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2262_ net773 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1144_ net687 net670 net657 net651 Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q
+ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__mux4_2
X_1075_ Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__inv_2
XFILLER_18_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2193_ clknet_4_0_0_UserCLK_regs _0017_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[28\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1977_ _0861_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__inv_1
X_2529_ net40 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_56_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1831_ Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q _0749_ VGND VGND VPWR VPWR _0750_
+ sky130_fd_sc_hd__or2_1
X_2880_ Inst_RegFile_switch_matrix.S1BEG2 VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__buf_6
X_1900_ net666 Inst_RegFile_switch_matrix.JS2BEG3 _0804_ _0805_ Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.W1BEG0
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_25_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1762_ _0687_ _0689_ _0692_ _1008_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JN2BEG7
+ sky130_fd_sc_hd__a22o_4
X_1693_ _0631_ Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q
+ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_68_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2314_ net776 net737 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2176_ clknet_4_0_0_UserCLK_regs _0000_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[24\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2245_ clknet_4_9_0_UserCLK_regs _0069_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[20\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1127_ Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__inv_2
XFILLER_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1058_ net131 VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__inv_2
XFILLER_21_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput104 S2MID[5] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput115 W1END[0] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_4
Xinput126 W2END[7] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput137 WW4END[0] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_4
XFILLER_72_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2030_ net620 net905 _0896_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__mux2_4
XFILLER_62_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2932_ Inst_RegFile_switch_matrix.W1BEG1 VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__clkbuf_2
X_1745_ _0676_ _0677_ _1003_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__mux2_1
X_2794_ net37 VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_1
X_1814_ net60 net2 net116 net673 Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q
+ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__mux4_1
X_2863_ NN4END[5] VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__clkbuf_2
X_1676_ net676 net635 net666 net639 Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q
+ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__mux4_1
Xhold336 Inst_RegFile_32x4.mem\[16\]\[1\] VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 Inst_RegFile_32x4.mem\[17\]\[2\] VGND VGND VPWR VPWR net889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 Inst_RegFile_32x4.mem\[10\]\[3\] VGND VGND VPWR VPWR net922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 Inst_RegFile_32x4.mem\[7\]\[0\] VGND VGND VPWR VPWR net933 sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 Inst_RegFile_32x4.mem\[28\]\[3\] VGND VGND VPWR VPWR net900 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold303 Inst_RegFile_32x4.mem\[29\]\[2\] VGND VGND VPWR VPWR net878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_209 net777 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2159_ net621 net916 _0929_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__mux2_2
X_2228_ clknet_4_6_0_UserCLK_regs _0052_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1392_ net60 net68 net2 net10 Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q
+ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__mux4_2
X_1530_ _0484_ _0483_ net412 VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__mux2_1
X_1461_ _0418_ _0417_ net683 VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__mux2_1
XFILLER_67_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2013_ net611 net938 _0890_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__mux2_4
X_2915_ SS4END[5] VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1728_ _0661_ _0662_ _1000_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__mux2_1
X_2777_ net49 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__buf_1
X_2846_ N4END[4] VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkbuf_2
Xfanout679 net680 VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__buf_6
Xfanout657 net658 VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__buf_6
X_1659_ net679 net636 net667 net640 Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q
+ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__mux4_1
Xfanout646 net647 VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__buf_8
Xfanout635 BD2 VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__buf_2
Xfanout602 _0869_ VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__buf_4
Xfanout668 BD1 VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__buf_8
Xfanout624 net626 VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__clkbuf_4
Xfanout613 net614 VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__buf_1
XFILLER_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput205 net205 VGND VGND VPWR VPWR FrameData_O[24] sky130_fd_sc_hd__buf_2
X_2631_ net752 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput216 net216 VGND VGND VPWR VPWR FrameData_O[5] sky130_fd_sc_hd__buf_2
X_2562_ net41 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_9_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2700_ clknet_4_11_0_UserCLK_regs _0102_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput238 net238 VGND VGND VPWR VPWR FrameStrobe_O[7] sky130_fd_sc_hd__buf_2
X_1444_ Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q _0402_ VGND VGND VPWR VPWR _0403_
+ sky130_fd_sc_hd__nand2b_1
Xoutput227 net227 VGND VGND VPWR VPWR FrameStrobe_O[15] sky130_fd_sc_hd__buf_2
Xoutput249 net249 VGND VGND VPWR VPWR N2BEG[4] sky130_fd_sc_hd__buf_2
X_2493_ net764 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1513_ Inst_RegFile_32x4.mem\[28\]\[1\] Inst_RegFile_32x4.mem\[29\]\[1\] net603 VGND
+ VGND VPWR VPWR _0468_ sky130_fd_sc_hd__mux2_1
X_1375_ Inst_RegFile_32x4.mem\[20\]\[3\] Inst_RegFile_32x4.mem\[21\]\[3\] net628 VGND
+ VGND VPWR VPWR _0340_ sky130_fd_sc_hd__mux2_1
XFILLER_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2829_ Inst_RegFile_switch_matrix.N1BEG3 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_2
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_63_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1091_ Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__inv_2
XFILLER_37_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1160_ Inst_RegFile_32x4.mem\[26\]\[0\] Inst_RegFile_32x4.mem\[27\]\[0\] net625 VGND
+ VGND VPWR VPWR _0137_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_72_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1993_ net620 net909 _0860_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_15_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2614_ net773 net722 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2545_ net53 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_9_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2476_ net46 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1427_ _0946_ _0386_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__nand2_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1358_ Inst_RegFile_32x4.mem\[4\]\[3\] Inst_RegFile_32x4.mem\[5\]\[3\] net630 VGND
+ VGND VPWR VPWR _0323_ sky130_fd_sc_hd__mux2_1
XFILLER_34_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1289_ Inst_RegFile_32x4.mem\[6\]\[1\] Inst_RegFile_32x4.mem\[7\]\[1\] net628 VGND
+ VGND VPWR VPWR _0258_ sky130_fd_sc_hd__mux2_1
XFILLER_50_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload3 clknet_4_3_0_UserCLK_regs VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_57_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1212_ net87 net97 net89 net689 Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q
+ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__mux4_1
XFILLER_69_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2261_ net774 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2330_ net32 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2192_ clknet_4_0_0_UserCLK_regs _0016_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[28\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1074_ Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__inv_2
X_1143_ _0968_ _1033_ Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q VGND VGND VPWR VPWR
+ _1034_ sky130_fd_sc_hd__o21ba_1
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1976_ net133 Inst_RegFile_switch_matrix.JN2BEG3 Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q
+ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__mux2_1
X_2528_ net39 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_56_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2459_ net766 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1761_ _0690_ _0691_ Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q VGND VGND VPWR VPWR
+ _0692_ sky130_fd_sc_hd__mux2_1
X_1830_ net86 net114 net780 net689 Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q
+ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__mux4_1
XFILLER_51_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1692_ net687 net673 net654 net647 Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q
+ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__mux4_1
X_2313_ net749 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1126_ Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__inv_2
X_2175_ net611 net888 _0932_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__mux2_1
X_2244_ clknet_4_9_0_UserCLK_regs _0068_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[20\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1057_ Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__inv_1
XFILLER_38_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1959_ Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q _0772_ Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q
+ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__o21ai_1
Xinput105 S2MID[6] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_2
Xinput116 W1END[1] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_4
Xinput127 W2MID[0] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
Xinput138 WW4END[1] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_4
XFILLER_56_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_6_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2931_ Inst_RegFile_switch_matrix.W1BEG0 VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__buf_2
X_1744_ net59 net1 net63 net5 Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q
+ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__mux4_1
X_1813_ _0736_ _0735_ Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.WW4BEG0 sky130_fd_sc_hd__mux2_1
X_2793_ net764 VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_1
X_2862_ NN4END[4] VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__clkbuf_2
Xhold326 Inst_RegFile_32x4.mem\[2\]\[2\] VGND VGND VPWR VPWR net901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 Inst_RegFile_32x4.mem\[0\]\[3\] VGND VGND VPWR VPWR net890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold304 Inst_RegFile_32x4.mem\[9\]\[0\] VGND VGND VPWR VPWR net879 sky130_fd_sc_hd__dlygate4sd3_1
X_1675_ Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q _0615_ VGND VGND VPWR VPWR _0616_
+ sky130_fd_sc_hd__or2_1
Xhold359 Inst_RegFile_32x4.mem\[16\]\[3\] VGND VGND VPWR VPWR net934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 Inst_RegFile_32x4.mem\[2\]\[1\] VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 Inst_RegFile_32x4.mem\[31\]\[3\] VGND VGND VPWR VPWR net912 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1109_ Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_64_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2089_ net613 net934 _0914_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2158_ net616 net898 _0929_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__mux2_4
X_2227_ clknet_4_6_0_UserCLK_regs _0051_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[14\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_36_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1391_ net26 net88 net90 net96 Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q
+ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__mux4_2
XFILLER_4_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1460_ Inst_RegFile_32x4.mem\[4\]\[0\] Inst_RegFile_32x4.mem\[5\]\[0\] net609 VGND
+ VGND VPWR VPWR _0418_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2012_ net620 net932 _0890_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__mux2_4
X_2914_ SS4END[4] VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_61_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2845_ net78 VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__clkbuf_2
X_1727_ net59 net1 net63 net5 Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q
+ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__mux4_1
X_1658_ net136 net673 net659 net646 Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q
+ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__mux4_1
X_2776_ net751 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__buf_4
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout669 net671 VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__buf_2
Xfanout636 net637 VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__clkbuf_4
Xfanout647 AD3 VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__buf_6
Xfanout658 AD1 VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__buf_8
X_1589_ _0389_ _0539_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__nand2_1
Xfanout625 net626 VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__clkbuf_2
Xfanout603 net604 VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__buf_6
Xfanout614 _0887_ VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__buf_2
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput239 net239 VGND VGND VPWR VPWR FrameStrobe_O[8] sky130_fd_sc_hd__buf_2
Xoutput228 net228 VGND VGND VPWR VPWR FrameStrobe_O[16] sky130_fd_sc_hd__buf_2
Xoutput206 net206 VGND VGND VPWR VPWR FrameData_O[25] sky130_fd_sc_hd__buf_2
X_2630_ net753 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput217 net217 VGND VGND VPWR VPWR FrameData_O[6] sky130_fd_sc_hd__buf_2
X_2492_ net765 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2561_ net759 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1512_ _0465_ _0466_ net412 VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__mux2_1
X_1443_ net138 net670 net657 net651 Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q
+ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__mux4_1
X_1374_ Inst_RegFile_32x4.mem\[22\]\[3\] Inst_RegFile_32x4.mem\[23\]\[3\] net628 VGND
+ VGND VPWR VPWR _0339_ sky130_fd_sc_hd__mux2_1
XFILLER_55_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2828_ Inst_RegFile_switch_matrix.N1BEG2 VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2759_ EE4END[5] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
XFILLER_73_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1090_ Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__inv_1
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1992_ _0707_ _0723_ _0437_ _0874_ Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q
+ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__mux4_1
Xclkload10 clknet_4_12_0_UserCLK_regs VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_15_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2613_ net774 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2475_ net36 net709 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2544_ net52 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1426_ net84 net10 net96 net124 Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q
+ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__mux4_2
XFILLER_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1357_ _0320_ _0321_ net661 VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__mux2_1
X_1288_ Inst_RegFile_32x4.mem\[4\]\[1\] Inst_RegFile_32x4.mem\[5\]\[1\] net630 VGND
+ VGND VPWR VPWR _0257_ sky130_fd_sc_hd__mux2_1
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload4 clknet_4_4_0_UserCLK_regs VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_57_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1211_ Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q _0184_ VGND VGND VPWR VPWR _0185_
+ sky130_fd_sc_hd__and2b_1
XFILLER_65_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2260_ net775 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_49_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1142_ net74 net16 net102 net130 Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q
+ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__mux4_2
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2191_ clknet_4_4_0_UserCLK_regs _0015_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[27\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_190 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1073_ Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__inv_2
XFILLER_25_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1975_ _0859_ _0831_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__nand2_4
X_1409_ _0369_ _0370_ Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q VGND VGND VPWR VPWR
+ _0371_ sky130_fd_sc_hd__mux2_1
X_2527_ net761 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2458_ net767 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2389_ net774 net696 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1760_ net5 net91 net87 net115 Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q
+ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__mux4_1
X_1691_ _0992_ _0629_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__or2_1
X_2312_ net750 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_53_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1125_ Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__inv_2
X_2243_ clknet_4_10_0_UserCLK_regs _0067_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2174_ net623 net823 _0932_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__mux2_1
X_1056_ Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_51_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1889_ _0719_ _0361_ Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q VGND VGND VPWR VPWR
+ _0799_ sky130_fd_sc_hd__mux2_1
X_1958_ _0839_ _0840_ _0842_ Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q
+ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__o221a_1
Xinput106 S2MID[7] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput128 W2MID[1] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__buf_2
Xclkbuf_4_9_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_9_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
Xinput117 W1END[2] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
Xinput139 WW4END[2] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_67_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_90 W6END[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2861_ Inst_RegFile_switch_matrix.N4BEG3 VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__buf_1
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2930_ clknet_1_0__leaf_UserCLK VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__buf_2
XFILLER_15_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1743_ net23 net89 net87 net91 Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q
+ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__mux4_1
X_2792_ net765 VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_2
X_1812_ net61 net89 net689 net656 Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q
+ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__mux4_1
X_1674_ net687 net671 net652 net645 Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q
+ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__mux4_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold305 Inst_RegFile_32x4.mem\[10\]\[0\] VGND VGND VPWR VPWR net880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 Inst_RegFile_32x4.mem\[3\]\[1\] VGND VGND VPWR VPWR net924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 Inst_RegFile_32x4.mem\[3\]\[2\] VGND VGND VPWR VPWR net913 sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 Inst_RegFile_32x4.mem\[28\]\[0\] VGND VGND VPWR VPWR net902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 Inst_RegFile_32x4.mem\[14\]\[0\] VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__dlygate4sd3_1
X_2226_ clknet_4_7_0_UserCLK_regs _0050_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[14\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1108_ Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2088_ net622 net906 _0914_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__mux2_4
X_2157_ net600 net812 _0929_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__mux2_1
XFILLER_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1390_ _0943_ _0352_ Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q VGND VGND VPWR VPWR
+ _0353_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_61_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2011_ net615 net931 _0890_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__mux2_4
XFILLER_50_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2913_ Inst_RegFile_switch_matrix.S4BEG3 VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__clkbuf_2
X_2844_ net77 VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_33_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1726_ net87 net91 net111 net115 Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q
+ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__mux4_1
X_1657_ _0600_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JS2BEG2 sky130_fd_sc_hd__inv_1
X_2775_ net36 VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__buf_1
X_1588_ _0537_ _0538_ net683 VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__mux2_1
Xfanout615 net618 VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__clkbuf_2
Xfanout604 net605 VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__buf_4
XFILLER_58_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout659 net660 VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__buf_2
Xfanout637 BD2 VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__clkbuf_2
X_2209_ clknet_4_3_0_UserCLK_regs _0033_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout648 _0164_ VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__buf_2
Xfanout626 net632 VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__buf_4
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput229 net229 VGND VGND VPWR VPWR FrameStrobe_O[17] sky130_fd_sc_hd__buf_2
Xoutput207 net207 VGND VGND VPWR VPWR FrameData_O[26] sky130_fd_sc_hd__buf_2
Xoutput218 net218 VGND VGND VPWR VPWR FrameData_O[7] sky130_fd_sc_hd__buf_2
X_2560_ net760 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2491_ net33 net709 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1442_ net64 net92 net26 net120 Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q
+ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__mux4_2
X_1511_ Inst_RegFile_32x4.mem\[26\]\[1\] Inst_RegFile_32x4.mem\[27\]\[1\] net604 VGND
+ VGND VPWR VPWR _0466_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1373_ _0336_ _0337_ net675 VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2827_ Inst_RegFile_switch_matrix.N1BEG1 VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__buf_4
X_2758_ EE4END[4] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_1
X_1709_ _0996_ _0645_ Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q VGND VGND VPWR VPWR
+ _0646_ sky130_fd_sc_hd__o21a_1
X_2689_ clknet_4_10_0_UserCLK_regs _0091_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_72_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2612_ net775 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1991_ net80 net686 net777 Inst_RegFile_switch_matrix.JS2BEG1 Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_15_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload11 clknet_4_13_0_UserCLK_regs VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__clkinvlp_4
X_2474_ net27 net709 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2543_ net51 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1425_ _0953_ _0382_ _0384_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__o21ai_1
XFILLER_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1287_ _0254_ _0255_ net661 VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__mux2_1
X_1356_ Inst_RegFile_32x4.mem\[2\]\[3\] Inst_RegFile_32x4.mem\[3\]\[3\] net627 VGND
+ VGND VPWR VPWR _0321_ sky130_fd_sc_hd__mux2_1
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload5 clknet_4_5_0_UserCLK_regs VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__clkinv_2
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1210_ net61 net69 net3 net11 Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q
+ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__mux4_1
X_1072_ Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__inv_1
X_1141_ _1027_ _1028_ _1030_ Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q VGND VGND
+ VPWR VPWR _1032_ sky130_fd_sc_hd__a211o_1
X_2190_ clknet_4_4_0_UserCLK_regs _0014_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[27\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_180 SS4END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_191 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1974_ _0853_ _0858_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__nor2_8
X_2526_ net762 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1408_ net90 net98 net112 net116 Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q
+ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__mux4_1
X_2388_ net775 net696 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2457_ net768 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_71_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1339_ Inst_RegFile_32x4.mem\[22\]\[2\] Inst_RegFile_32x4.mem\[23\]\[2\] net628 VGND
+ VGND VPWR VPWR _0306_ sky130_fd_sc_hd__mux2_1
XFILLER_51_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput390 net390 VGND VGND VPWR VPWR WW4BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1690_ net680 net637 net667 net641 Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q
+ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__mux4_1
X_2311_ net752 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2242_ clknet_4_8_0_UserCLK_regs _0066_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_69_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1124_ Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__inv_2
X_1055_ net103 VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__inv_1
X_2173_ net618 net851 _0932_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1957_ _0841_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__inv_1
X_1888_ _0794_ _0798_ Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.NN4BEG1 sky130_fd_sc_hd__mux2_4
X_2509_ net748 net711 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput107 S4END[0] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_67_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput118 W1END[3] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
Xinput129 W2MID[2] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_91 W6END[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_80 net347 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1811_ _0734_ _0733_ Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q VGND VGND VPWR VPWR
+ _0735_ sky130_fd_sc_hd__mux2_1
X_2860_ Inst_RegFile_switch_matrix.N4BEG2 VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_1
X_2791_ net766 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1742_ Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q _0672_ Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q
+ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__o21a_1
X_1673_ _0987_ _0614_ _0611_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JN2BEG2
+ sky130_fd_sc_hd__a21o_1
Xhold328 Inst_RegFile_32x4.mem\[16\]\[0\] VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 Inst_RegFile_32x4.mem\[8\]\[2\] VGND VGND VPWR VPWR net914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 Inst_RegFile_32x4.mem\[23\]\[3\] VGND VGND VPWR VPWR net892 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold306 Inst_RegFile_32x4.mem\[5\]\[3\] VGND VGND VPWR VPWR net881 sky130_fd_sc_hd__dlygate4sd3_1
X_2225_ clknet_4_6_0_UserCLK_regs _0049_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1107_ Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__inv_1
XFILLER_38_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2087_ net618 net911 _0914_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__mux2_4
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2156_ _0859_ _0898_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__nand2_4
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2010_ net599 net829 _0890_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__mux2_1
X_2912_ Inst_RegFile_switch_matrix.S4BEG2 VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_61_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1725_ Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q _0659_ Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q
+ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__o21a_1
X_2774_ net776 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_33_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2843_ net76 VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_2
X_1656_ Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q _0597_ _0599_ _0593_ _0595_ VGND
+ VGND VPWR VPWR _0600_ sky130_fd_sc_hd__o32a_1
Xfanout638 net639 VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__buf_8
X_1587_ Inst_RegFile_32x4.mem\[18\]\[2\] Inst_RegFile_32x4.mem\[19\]\[2\] net610 VGND
+ VGND VPWR VPWR _0538_ sky130_fd_sc_hd__mux2_1
Xfanout616 net617 VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__buf_4
Xfanout627 net628 VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__clkbuf_4
Xfanout605 B_ADR0 VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__buf_8
Xfanout649 _0163_ VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__buf_6
XFILLER_37_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2208_ clknet_4_7_0_UserCLK_regs _0032_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2139_ net622 net856 _0925_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__mux2_1
XFILLER_14_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer200 _0859_ VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__buf_6
XFILLER_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput208 net208 VGND VGND VPWR VPWR FrameData_O[27] sky130_fd_sc_hd__buf_2
Xoutput219 net219 VGND VGND VPWR VPWR FrameData_O[8] sky130_fd_sc_hd__buf_2
X_2490_ net32 net709 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1441_ net83 net778 net119 Inst_RegFile_switch_matrix.JW2BEG4 Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__mux4_2
XFILLER_4_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1510_ Inst_RegFile_32x4.mem\[24\]\[1\] Inst_RegFile_32x4.mem\[25\]\[1\] net603 VGND
+ VGND VPWR VPWR _0465_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1372_ Inst_RegFile_32x4.mem\[16\]\[3\] Inst_RegFile_32x4.mem\[17\]\[3\] net631 VGND
+ VGND VPWR VPWR _0337_ sky130_fd_sc_hd__mux2_1
XFILLER_63_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1708_ net644 net411 net664 net415 Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q
+ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__mux4_1
X_2826_ Inst_RegFile_switch_matrix.N1BEG0 VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_2
X_2688_ clknet_4_8_0_UserCLK_regs _0090_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1639_ _0581_ _0582_ _0584_ _0583_ Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q
+ VGND VGND VPWR VPWR A_ADR0 sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_72_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_32_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1990_ net615 net833 _0860_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__mux2_1
X_2611_ net742 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2542_ net747 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_41_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload12 clknet_4_14_0_UserCLK_regs VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__clkinv_2
XPHY_EDGE_ROW_50_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1424_ Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q _0383_ Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q
+ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__o21a_1
X_2473_ net749 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1355_ Inst_RegFile_32x4.mem\[0\]\[3\] Inst_RegFile_32x4.mem\[1\]\[3\] net627 VGND
+ VGND VPWR VPWR _0320_ sky130_fd_sc_hd__mux2_1
XFILLER_68_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1286_ Inst_RegFile_32x4.mem\[2\]\[1\] Inst_RegFile_32x4.mem\[3\]\[1\] net627 VGND
+ VGND VPWR VPWR _0255_ sky130_fd_sc_hd__mux2_1
XFILLER_51_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload6 clknet_4_6_0_UserCLK_regs VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__clkinvlp_4
X_2809_ net715 VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__buf_1
XFILLER_3_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1071_ Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__inv_1
X_1140_ _1028_ _1027_ _1030_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__a21o_1
XFILLER_18_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_170 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_192 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1973_ Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q _0854_ _0856_ VGND VGND VPWR VPWR
+ _0858_ sky130_fd_sc_hd__o21a_2
XANTENNA_181 WW4END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2525_ net764 net712 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1407_ net62 net70 net4 net12 Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q
+ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__mux4_1
XFILLER_68_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2387_ net742 net696 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2456_ net770 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1338_ _0303_ _0304_ net662 VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1269_ Inst_RegFile_32x4.mem\[8\]\[0\] Inst_RegFile_32x4.mem\[9\]\[0\] net629 VGND
+ VGND VPWR VPWR _0240_ sky130_fd_sc_hd__mux2_1
Xoutput380 net380 VGND VGND VPWR VPWR WW4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput391 net391 VGND VGND VPWR VPWR WW4BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_59_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2310_ net753 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2241_ clknet_4_10_0_UserCLK_regs _0065_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2172_ net602 net930 _0932_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__mux2_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1123_ Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__inv_2
X_1054_ Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__inv_2
X_1887_ Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q _0797_ _0796_ VGND VGND VPWR VPWR
+ _0798_ sky130_fd_sc_hd__a21bo_1
X_1956_ net8 net114 Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q VGND VGND VPWR VPWR
+ _0841_ sky130_fd_sc_hd__mux2_1
XFILLER_33_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput108 S4END[1] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__buf_2
X_2508_ net751 net711 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_71_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2439_ net45 net700 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput119 W2END[0] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_2
XFILLER_72_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_70 S4END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_92 W6END[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_81 net349 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1741_ _1003_ _0673_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__or2_1
X_2790_ net767 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_2
X_1810_ net664 _0718_ Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q VGND VGND VPWR VPWR
+ _0734_ sky130_fd_sc_hd__mux2_1
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1672_ _0612_ _0613_ _0986_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__mux2_1
Xhold318 Inst_RegFile_32x4.mem\[11\]\[0\] VGND VGND VPWR VPWR net893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold307 Inst_RegFile_32x4.mem\[21\]\[1\] VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 Inst_RegFile_32x4.mem\[14\]\[1\] VGND VGND VPWR VPWR net904 sky130_fd_sc_hd__dlygate4sd3_1
X_1106_ Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__inv_1
XFILLER_38_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2155_ net614 net920 _0928_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__mux2_2
X_2224_ clknet_4_6_0_UserCLK_regs _0048_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2086_ net602 net903 _0914_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__mux2_4
Xinput90 S1END[3] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_6
X_1939_ Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q _0823_ Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q
+ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__a21o_1
XFILLER_44_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_5_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_5_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2911_ Inst_RegFile_switch_matrix.S4BEG1 VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_33_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1724_ net689 net669 net656 net651 Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q
+ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__mux4_1
X_2773_ Inst_RegFile_switch_matrix.EE4BEG3 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__buf_1
X_2842_ net75 VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__buf_2
X_1655_ _0983_ _0598_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__nor2_1
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout639 BD3 VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__buf_8
Xfanout617 net618 VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__buf_4
X_1586_ Inst_RegFile_32x4.mem\[16\]\[2\] Inst_RegFile_32x4.mem\[17\]\[2\] net610 VGND
+ VGND VPWR VPWR _0537_ sky130_fd_sc_hd__mux2_1
Xfanout606 net607 VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__clkbuf_4
Xfanout628 net629 VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__clkbuf_4
X_2069_ net612 net927 _0910_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__mux2_4
X_2207_ clknet_4_2_0_UserCLK_regs _0031_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2138_ net617 net875 _0925_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__mux2_1
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput209 net209 VGND VGND VPWR VPWR FrameData_O[28] sky130_fd_sc_hd__buf_2
XFILLER_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1440_ _0396_ _0394_ _0399_ _0956_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JW2BEG4
+ sky130_fd_sc_hd__a22o_4
X_1371_ Inst_RegFile_32x4.mem\[18\]\[3\] Inst_RegFile_32x4.mem\[19\]\[3\] net630 VGND
+ VGND VPWR VPWR _0336_ sky130_fd_sc_hd__mux2_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2825_ FrameStrobe[19] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_46_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1707_ Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q _0643_ VGND VGND VPWR VPWR _0644_
+ sky130_fd_sc_hd__or2_1
X_2756_ Inst_RegFile_switch_matrix.E6BEG0 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_1
X_1638_ net70 net98 net25 net126 Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q
+ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__mux4_1
X_2687_ clknet_4_10_0_UserCLK_regs _0089_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1569_ Inst_RegFile_32x4.BD_comb\[3\] Inst_RegFile_32x4.BD_reg\[3\] Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q
+ VGND VGND VPWR VPWR BD3 sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_72_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2610_ net743 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2541_ net748 net714 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2472_ net750 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1423_ net22 net108 Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q VGND VGND VPWR VPWR
+ _0383_ sky130_fd_sc_hd__mux2_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1285_ Inst_RegFile_32x4.mem\[0\]\[1\] Inst_RegFile_32x4.mem\[1\]\[1\] net627 VGND
+ VGND VPWR VPWR _0254_ sky130_fd_sc_hd__mux2_1
X_1354_ net648 _0314_ _0318_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__a21oi_1
XFILLER_55_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2808_ net721 VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_1
Xclkload7 clknet_4_7_0_UserCLK_regs VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__clkinv_2
X_2739_ net14 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1070_ Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__inv_1
XANTENNA_160 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_193 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_171 FrameStrobe[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1972_ Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q _0854_ _0856_ VGND VGND VPWR VPWR
+ _0857_ sky130_fd_sc_hd__o21ai_4
XPHY_EDGE_ROW_23_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_182 WW4END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2524_ net765 net712 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2455_ net772 net705 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1406_ _0948_ _0367_ Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q VGND VGND VPWR VPWR
+ _0368_ sky130_fd_sc_hd__o21a_1
XFILLER_68_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2386_ net54 net696 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1337_ Inst_RegFile_32x4.mem\[18\]\[2\] Inst_RegFile_32x4.mem\[19\]\[2\] net630 VGND
+ VGND VPWR VPWR _0304_ sky130_fd_sc_hd__mux2_1
X_1268_ Inst_RegFile_32x4.mem\[10\]\[0\] Inst_RegFile_32x4.mem\[11\]\[0\] net629 VGND
+ VGND VPWR VPWR _0239_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1199_ _0172_ _0173_ Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q VGND VGND VPWR VPWR
+ _0174_ sky130_fd_sc_hd__mux2_1
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput370 net370 VGND VGND VPWR VPWR W6BEG[2] sky130_fd_sc_hd__buf_2
Xoutput381 net381 VGND VGND VPWR VPWR WW4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput392 net392 VGND VGND VPWR VPWR WW4BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_59_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1122_ Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__inv_1
X_2171_ _0859_ _0904_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__nand2_4
X_2240_ clknet_4_8_0_UserCLK_regs _0064_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1053_ Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__inv_2
XFILLER_21_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1886_ _0708_ _0133_ Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q VGND VGND VPWR VPWR
+ _0797_ sky130_fd_sc_hd__mux2_4
X_1955_ net139 Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q
+ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__o21ai_1
Xinput109 S4END[2] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_4
X_2507_ net763 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2438_ net753 net700 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_67_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2369_ net759 net693 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
Xclkbuf_4_13_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_13_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_12_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_71 S4END[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 W6END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 net352 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_60 N4END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1740_ net644 net411 net665 net415 Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q
+ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__mux4_1
X_1671_ net66 net2 net82 net8 Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q
+ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__mux4_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold308 Inst_RegFile_32x4.mem\[27\]\[3\] VGND VGND VPWR VPWR net883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 Inst_RegFile_32x4.mem\[18\]\[2\] VGND VGND VPWR VPWR net894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1105_ Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_64_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2085_ _0859_ _0907_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__nand2_8
X_2154_ net621 net914 _0928_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__mux2_2
X_2223_ clknet_4_11_0_UserCLK_regs _0047_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[23\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput91 S2END[0] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_2
X_1869_ net667 _0718_ _0719_ _0567_ Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q
+ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__mux4_1
X_1938_ net76 net18 net104 net132 Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q
+ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__mux4_1
Xinput80 N4END[1] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2841_ net74 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__buf_1
XFILLER_31_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2910_ Inst_RegFile_switch_matrix.S4BEG0 VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__buf_1
X_1723_ _1000_ _0657_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__or2_1
X_1654_ net777 net94 net110 net122 Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q
+ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__mux4_1
X_2772_ Inst_RegFile_switch_matrix.EE4BEG2 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
Xfanout618 _0873_ VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__buf_4
X_2206_ clknet_4_9_0_UserCLK_regs _0030_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout629 net632 VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__buf_2
Xfanout607 net608 VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__clkbuf_4
X_1585_ _0524_ _0528_ net619 _0535_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__o22a_1
X_2068_ net622 net935 _0910_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__mux2_4
X_2137_ net601 net837 _0925_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__mux2_1
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1370_ net649 _0334_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_46_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2824_ FrameStrobe[18] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_1
XFILLER_31_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2755_ E6END[11] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__buf_1
X_1706_ net137 net669 net656 net651 Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q
+ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__mux4_1
X_1637_ net82 net8 net122 Inst_RegFile_switch_matrix.JN2BEG3 Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__mux4_2
X_2686_ clknet_4_8_0_UserCLK_regs _0088_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1499_ _0455_ _0415_ _0439_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__o21a_1
X_1568_ _0439_ _0496_ _0504_ _0520_ _0519_ VGND VGND VPWR VPWR Inst_RegFile_32x4.BD_comb\[3\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_72_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2540_ net751 net714 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1422_ net140 Inst_RegFile_switch_matrix.JS2BEG4 Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q
+ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__mux2_1
X_2471_ net45 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1284_ _0249_ _0252_ net649 VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__mux2_1
X_1353_ net649 _0317_ _0192_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__a21o_1
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2807_ net726 VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_1
X_2738_ net13 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
Xclkload8 clknet_4_9_0_UserCLK_regs VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_14_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2669_ clknet_4_12_0_UserCLK_regs Inst_RegFile_32x4.BD_comb\[3\] VGND VGND VPWR VPWR
+ Inst_RegFile_32x4.BD_reg\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_150 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_161 net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_172 FrameStrobe[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_194 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_183 _0264_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1971_ Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q _0805_ _0855_ VGND VGND VPWR VPWR
+ _0856_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_11_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1405_ net646 net679 net668 net640 Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q
+ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__mux4_2
XFILLER_68_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2523_ net766 net712 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2385_ net53 net696 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2454_ net773 net705 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1198_ net778 net95 net107 net123 Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q
+ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__mux4_1
XFILLER_36_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 E1END[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_4
X_1336_ Inst_RegFile_32x4.mem\[16\]\[2\] Inst_RegFile_32x4.mem\[17\]\[2\] net630 VGND
+ VGND VPWR VPWR _0303_ sky130_fd_sc_hd__mux2_1
X_1267_ net650 _0237_ _0234_ _0193_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__a211o_1
XFILLER_51_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput371 net371 VGND VGND VPWR VPWR W6BEG[3] sky130_fd_sc_hd__buf_2
Xoutput382 net382 VGND VGND VPWR VPWR WW4BEG[13] sky130_fd_sc_hd__buf_8
Xoutput393 net393 VGND VGND VPWR VPWR WW4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput360 net360 VGND VGND VPWR VPWR W2BEGb[2] sky130_fd_sc_hd__buf_2
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1121_ Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__inv_1
X_1052_ Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__inv_2
XFILLER_38_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2170_ net614 net839 _0931_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__mux2_1
X_1954_ _0987_ _0614_ _0611_ _1016_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__a211oi_1
XPHY_EDGE_ROW_38_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1885_ Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q _0706_ _0795_ Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q
+ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_47_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2506_ net776 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2437_ net755 net701 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2368_ net760 net693 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_67_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2299_ net766 net730 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1319_ net648 _0281_ _0284_ _0285_ _0192_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__a221o_1
XANTENNA_72 S4END[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_50 net242 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_83 net356 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_94 W6END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput190 net190 VGND VGND VPWR VPWR FrameData_O[10] sky130_fd_sc_hd__buf_2
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_UserCLK clknet_0_UserCLK VGND VGND VPWR VPWR clknet_1_0__leaf_UserCLK
+ sky130_fd_sc_hd__clkbuf_16
X_1670_ net777 net94 net122 net139 Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q
+ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__mux4_1
Xhold309 Inst_RegFile_32x4.mem\[14\]\[2\] VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__dlygate4sd3_1
X_2222_ clknet_4_9_0_UserCLK_regs _0046_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[23\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1104_ Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_64_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2153_ net616 net896 _0928_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__mux2_2
X_2084_ _0887_ net817 _0913_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__mux2_1
XFILLER_34_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1937_ _0810_ _0820_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__nand2_1
Xinput92 S2END[1] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_2
X_1799_ _0725_ _0724_ Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.WW4BEG3 sky130_fd_sc_hd__mux2_4
X_1868_ Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q _0778_ _0782_ VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.EE4BEG1 sky130_fd_sc_hd__o21a_1
Xinput81 N4END[2] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_2
Xinput70 N2END[7] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_4
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2840_ net73 VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__buf_4
X_1722_ net644 net677 net664 net633 Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q
+ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__mux4_1
X_1653_ Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q _0596_ VGND VGND VPWR VPWR _0597_
+ sky130_fd_sc_hd__nor2_1
XFILLER_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1584_ _0531_ _0534_ net642 VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__mux2_4
X_2205_ clknet_4_2_0_UserCLK_regs _0029_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout608 B_ADR0 VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__buf_6
Xfanout619 _0415_ VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__buf_2
XFILLER_53_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2136_ _0889_ _0923_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__nand2_2
X_2067_ net617 net919 _0910_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_32_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2969_ WW4END[10] VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__buf_1
XFILLER_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_1_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_1_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_63_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2823_ FrameStrobe[17] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_1
X_2754_ E6END[10] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_1
X_1705_ _0637_ _0639_ _0642_ _0995_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JN2BEG1
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1636_ net78 net20 net106 net134 Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q
+ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__mux4_2
X_2685_ clknet_4_4_0_UserCLK_regs _0087_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[31\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1567_ _0416_ _0511_ _0439_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__o21ba_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ _0451_ _0454_ net642 VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__mux2_1
X_2119_ net611 net876 _0920_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__mux2_1
XFILLER_10_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1421_ _0378_ _0376_ _0381_ _0952_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JS2BEG4
+ sky130_fd_sc_hd__a22o_4
X_2470_ net753 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1283_ _0250_ _0251_ net396 VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__mux2_1
X_1352_ _0315_ _0316_ net663 VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__mux2_1
XFILLER_36_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2737_ Inst_RegFile_switch_matrix.E2BEG7 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__buf_4
X_2806_ net740 VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__buf_1
X_2668_ clknet_4_12_0_UserCLK_regs Inst_RegFile_32x4.BD_comb\[2\] VGND VGND VPWR VPWR
+ Inst_RegFile_32x4.BD_reg\[2\] sky130_fd_sc_hd__dfxtp_1
Xclkload9 clknet_4_10_0_UserCLK_regs VGND VGND VPWR VPWR clkload9/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_14_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2599_ net752 net720 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1619_ net70 net12 net98 net137 Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q
+ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_6_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout780 net3 VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__clkbuf_4
XANTENNA_173 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_162 net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_151 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_184 net636 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_140 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_195 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1970_ _1017_ _0791_ Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q VGND VGND VPWR VPWR
+ _0855_ sky130_fd_sc_hd__a21bo_1
X_2522_ net767 net712 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1404_ Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q _0365_ VGND VGND VPWR VPWR _0366_
+ sky130_fd_sc_hd__or2_1
X_2453_ net774 net704 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2384_ net745 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1335_ net408 _0301_ net395 VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__a21oi_2
XFILLER_68_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1197_ net61 net67 net86 net9 Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q
+ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__mux4_1
XFILLER_36_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 E1END[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_6
XFILLER_24_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1266_ _0235_ _0236_ net662 VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__mux2_1
Xoutput350 net350 VGND VGND VPWR VPWR W2BEG[0] sky130_fd_sc_hd__buf_4
Xoutput361 net361 VGND VGND VPWR VPWR W2BEGb[3] sky130_fd_sc_hd__buf_2
XFILLER_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput372 net372 VGND VGND VPWR VPWR W6BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput383 net383 VGND VGND VPWR VPWR WW4BEG[14] sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_53_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1051_ Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__inv_2
X_1120_ Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__inv_1
XFILLER_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1884_ Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q net636 VGND VGND VPWR VPWR _0795_
+ sky130_fd_sc_hd__nor2_1
X_1953_ _0837_ _0835_ Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q VGND VGND VPWR VPWR
+ _0838_ sky130_fd_sc_hd__mux2_4
X_2505_ net749 net706 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_56_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2298_ net767 net730 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2367_ net38 net693 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2436_ net756 net701 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1318_ net663 _0282_ net408 VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__o21a_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1249_ _0219_ _0220_ Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q VGND VGND VPWR VPWR
+ _0221_ sky130_fd_sc_hd__mux2_1
XFILLER_24_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_62 net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_40 FrameStrobe[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 net249 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_73 S4END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_95 W6END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 net360 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput191 net191 VGND VGND VPWR VPWR FrameData_O[11] sky130_fd_sc_hd__buf_2
Xoutput180 net180 VGND VGND VPWR VPWR EE4BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_47_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2152_ net600 net811 _0928_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__mux2_1
X_2221_ clknet_4_10_0_UserCLK_regs _0045_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[23\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1103_ Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__inv_1
XFILLER_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2083_ net620 net859 _0913_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__mux2_1
X_1867_ _0779_ Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q _0780_ _0781_ _1012_ VGND
+ VGND VPWR VPWR _0782_ sky130_fd_sc_hd__a221o_1
X_1936_ _0812_ _0813_ _0819_ Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q VGND VGND
+ VPWR VPWR _0821_ sky130_fd_sc_hd__a2bb2o_1
Xinput93 S2END[2] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_4
X_1798_ net60 net88 net116 net670 Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q
+ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__mux4_1
Xinput60 N1END[1] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_12
Xinput71 N2MID[0] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput82 N4END[3] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_2
XFILLER_72_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2419_ net742 net700 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2770_ Inst_RegFile_switch_matrix.EE4BEG0 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
X_1721_ _0651_ _0653_ _0656_ _0999_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JW2BEG0
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1652_ net66 net8 net2 net25 Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q
+ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__mux4_1
X_1583_ _0532_ _0533_ net684 VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__mux2_1
Xfanout609 B_ADR0 VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__clkbuf_4
XFILLER_66_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2204_ clknet_4_2_0_UserCLK_regs _0028_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2135_ net613 net820 _0924_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__mux2_1
XFILLER_22_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2066_ net601 net862 _0910_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__mux2_1
X_2899_ S4END[5] VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__buf_4
X_1919_ net645 _0582_ Inst_RegFile_switch_matrix.JW2BEG0 _0158_ Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q
+ Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.N1BEG1
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_32_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2968_ WW4END[9] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__buf_1
XFILLER_27_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclone30 net655 VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__clkbuf_1
XFILLER_25_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2753_ E6END[9] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_1
X_2822_ FrameStrobe[16] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_1
X_1704_ _0640_ _0641_ Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q VGND VGND VPWR VPWR
+ _0642_ sky130_fd_sc_hd__mux2_1
X_2684_ clknet_4_5_0_UserCLK_regs _0086_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[31\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1635_ net77 net19 net133 Inst_RegFile_switch_matrix.JN2BEG5 Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__mux4_1
X_1497_ _0453_ _0452_ net412 VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__mux2_1
X_1566_ net619 _0518_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__or2_4
XFILLER_54_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2049_ net621 net864 _0903_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__mux2_1
X_2118_ net620 net878 _0920_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__mux2_1
XFILLER_22_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1420_ _0379_ _0380_ _0951_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__mux2_1
X_1351_ Inst_RegFile_32x4.mem\[14\]\[3\] Inst_RegFile_32x4.mem\[15\]\[3\] net626 VGND
+ VGND VPWR VPWR _0316_ sky130_fd_sc_hd__mux2_1
XFILLER_63_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1282_ Inst_RegFile_32x4.mem\[12\]\[1\] Inst_RegFile_32x4.mem\[13\]\[1\] net626 VGND
+ VGND VPWR VPWR _0251_ sky130_fd_sc_hd__mux2_1
X_2805_ net749 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2736_ Inst_RegFile_switch_matrix.E2BEG6 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__buf_1
X_1618_ _0563_ _0562_ _0565_ Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q
+ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__o221a_4
X_2667_ clknet_4_12_0_UserCLK_regs Inst_RegFile_32x4.BD_comb\[1\] VGND VGND VPWR VPWR
+ Inst_RegFile_32x4.BD_reg\[1\] sky130_fd_sc_hd__dfxtp_1
X_2598_ net754 net720 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_6_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1549_ _0500_ _0501_ net681 VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__mux2_1
XFILLER_67_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold290 Inst_RegFile_32x4.mem\[21\]\[3\] VGND VGND VPWR VPWR net865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout770 net771 VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__clkbuf_4
XFILLER_18_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_regs_0_UserCLK UserCLK VGND VGND VPWR VPWR UserCLK_regs sky130_fd_sc_hd__clkbuf_16
XFILLER_73_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_130 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_174 net260 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_185 net754 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_196 net195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_152 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_163 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_141 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2521_ net768 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_11_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1403_ net688 net672 net659 net653 Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q
+ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__mux4_1
X_2452_ net775 net704 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2383_ net746 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1265_ Inst_RegFile_32x4.mem\[6\]\[0\] Inst_RegFile_32x4.mem\[7\]\[0\] net630 VGND
+ VGND VPWR VPWR _0236_ sky130_fd_sc_hd__mux2_1
X_1334_ _0299_ _0300_ net663 VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__mux2_1
X_1196_ _0170_ _0978_ Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q VGND VGND VPWR VPWR
+ _0171_ sky130_fd_sc_hd__o21a_1
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput3 E1END[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput373 net373 VGND VGND VPWR VPWR W6BEG[5] sky130_fd_sc_hd__buf_2
Xoutput384 net384 VGND VGND VPWR VPWR WW4BEG[15] sky130_fd_sc_hd__buf_8
Xoutput351 net351 VGND VGND VPWR VPWR W2BEG[1] sky130_fd_sc_hd__buf_4
X_2719_ clknet_4_2_0_UserCLK_regs _0121_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput340 net340 VGND VGND VPWR VPWR SS4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput362 net362 VGND VGND VPWR VPWR W2BEGb[4] sky130_fd_sc_hd__buf_2
XFILLER_19_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1050_ Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__inv_1
X_1883_ net62 net779 net688 net653 Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q
+ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__mux4_1
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1952_ net66 net94 _0836_ _0823_ Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q
+ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2435_ net757 net699 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2504_ net750 net706 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_67_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1248_ net24 net88 net90 net98 Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q
+ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__mux4_1
X_2297_ net769 net730 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2366_ net37 net693 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1317_ net396 _0283_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__or2_1
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1179_ net67 net9 net780 net26 Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q
+ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__mux4_1
XFILLER_24_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_52 net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 FrameStrobe[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_30 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_63 net298 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 W6END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_74 S4END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 net364 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput192 net192 VGND VGND VPWR VPWR FrameData_O[12] sky130_fd_sc_hd__buf_2
Xoutput170 net170 VGND VGND VPWR VPWR E6BEG[7] sky130_fd_sc_hd__buf_2
Xoutput181 net181 VGND VGND VPWR VPWR EE4BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1102_ Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__inv_1
X_2151_ _0859_ _0902_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__nand2_4
X_2220_ clknet_4_9_0_UserCLK_regs _0044_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[23\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2082_ net615 net857 _0913_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1797_ net411 _0147_ _0372_ _0723_ Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q
+ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__mux4_2
Xinput50 FrameData[4] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_2
X_1866_ Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q _0706_ Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q
+ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1935_ Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q _0819_ _0813_ _0812_ VGND VGND
+ VPWR VPWR _0820_ sky130_fd_sc_hd__o2bb2a_1
Xinput61 N1END[2] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_4
Xinput72 N2MID[1] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput94 S2END[3] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_2
XFILLER_69_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2418_ net743 net699 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput83 NN4END[0] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_4
X_2349_ net748 net690 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_29_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1651_ _0983_ _0594_ Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q VGND VGND VPWR VPWR
+ _0595_ sky130_fd_sc_hd__o21ai_1
X_1720_ _0654_ _0655_ Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q VGND VGND VPWR VPWR
+ _0656_ sky130_fd_sc_hd__mux2_1
X_1582_ Inst_RegFile_32x4.mem\[14\]\[2\] Inst_RegFile_32x4.mem\[15\]\[2\] net605 VGND
+ VGND VPWR VPWR _0533_ sky130_fd_sc_hd__mux2_1
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2065_ _0891_ _0909_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__nand2_4
X_2203_ clknet_4_4_0_UserCLK_regs _0027_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[30\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2134_ net622 net825 _0924_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2967_ WW4END[8] VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_14_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1849_ net60 net2 net88 net673 Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q
+ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__mux4_1
X_1918_ net676 net685 Inst_RegFile_switch_matrix.JW2BEG1 net394 Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q
+ Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.N1BEG2
+ sky130_fd_sc_hd__mux4_1
X_2898_ S4END[4] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclone20 _0363_ VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__buf_6
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2821_ FrameStrobe[15] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_46_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2752_ E6END[8] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_1
X_1634_ _0577_ _0576_ _0580_ _0964_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JN2BEG3
+ sky130_fd_sc_hd__a22o_4
X_1703_ net24 net778 net93 net121 Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q
+ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__mux4_1
X_2683_ clknet_4_1_0_UserCLK_regs _0085_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[31\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1496_ Inst_RegFile_32x4.mem\[28\]\[0\] Inst_RegFile_32x4.mem\[29\]\[0\] net603 VGND
+ VGND VPWR VPWR _0453_ sky130_fd_sc_hd__mux2_1
X_1565_ _0514_ _0517_ net642 VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__mux2_4
XFILLER_66_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2117_ net615 net860 _0920_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__mux2_1
X_2048_ net616 net853 _0903_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__mux2_1
XFILLER_13_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1350_ Inst_RegFile_32x4.mem\[12\]\[3\] Inst_RegFile_32x4.mem\[13\]\[3\] net626 VGND
+ VGND VPWR VPWR _0315_ sky130_fd_sc_hd__mux2_1
X_1281_ Inst_RegFile_32x4.mem\[14\]\[1\] Inst_RegFile_32x4.mem\[15\]\[1\] net626 VGND
+ VGND VPWR VPWR _0250_ sky130_fd_sc_hd__mux2_1
XFILLER_63_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2804_ net750 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_2
X_2597_ net755 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2735_ Inst_RegFile_switch_matrix.E2BEG5 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
X_1617_ _0564_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__inv_1
X_2666_ clknet_4_12_0_UserCLK_regs Inst_RegFile_32x4.BD_comb\[0\] VGND VGND VPWR VPWR
+ Inst_RegFile_32x4.BD_reg\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1479_ net15 net129 net101 Inst_RegFile_switch_matrix.E2BEG3 Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__mux4_2
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1548_ Inst_RegFile_32x4.mem\[30\]\[3\] Inst_RegFile_32x4.mem\[31\]\[3\] net603 VGND
+ VGND VPWR VPWR _0501_ sky130_fd_sc_hd__mux2_1
XFILLER_54_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_UserCLK_regs UserCLK_regs VGND VGND VPWR VPWR clknet_0_UserCLK_regs sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_17_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout760 net39 VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__buf_4
XFILLER_49_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold291 Inst_RegFile_32x4.mem\[24\]\[3\] VGND VGND VPWR VPWR net866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold280 Inst_RegFile_32x4.mem\[21\]\[0\] VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_131 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout771 FrameData[14] VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_56_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_142 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_120 net755 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_197 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_153 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_164 net141 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_186 net760 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_175 N4END[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2520_ net770 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2451_ net742 net705 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1402_ Inst_RegFile_32x4.mem\[0\]\[0\] Inst_RegFile_32x4.mem\[1\]\[0\] net606 VGND
+ VGND VPWR VPWR _0364_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 E1END[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
X_2382_ net50 net697 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1264_ Inst_RegFile_32x4.mem\[4\]\[0\] Inst_RegFile_32x4.mem\[5\]\[0\] net630 VGND
+ VGND VPWR VPWR _0235_ sky130_fd_sc_hd__mux2_1
X_1333_ Inst_RegFile_32x4.mem\[30\]\[2\] Inst_RegFile_32x4.mem\[31\]\[2\] net624 VGND
+ VGND VPWR VPWR _0300_ sky130_fd_sc_hd__mux2_1
XFILLER_64_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1195_ net676 net633 net664 net638 Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q
+ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__mux4_2
XFILLER_51_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2718_ clknet_4_2_0_UserCLK_regs _0120_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2649_ net768 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput374 net374 VGND VGND VPWR VPWR W6BEG[6] sky130_fd_sc_hd__buf_2
Xoutput330 net330 VGND VGND VPWR VPWR SS4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput341 net341 VGND VGND VPWR VPWR SS4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput352 net352 VGND VGND VPWR VPWR W2BEG[2] sky130_fd_sc_hd__buf_4
Xoutput385 net385 VGND VGND VPWR VPWR WW4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput363 net363 VGND VGND VPWR VPWR W2BEGb[5] sky130_fd_sc_hd__buf_2
XFILLER_70_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1882_ _0793_ _0792_ Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.NN4BEG2 sky130_fd_sc_hd__mux2_1
X_1951_ net73 net129 net15 Inst_RegFile_switch_matrix.E2BEG4 Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__mux4_2
X_2365_ net764 net692 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2503_ net752 net707 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2434_ net758 net699 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_67_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1247_ net62 net70 net779 net12 Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q
+ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__mux4_1
X_2296_ net771 net730 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1178_ _0974_ _0153_ Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q VGND VGND VPWR VPWR
+ _0154_ sky130_fd_sc_hd__o21a_1
XFILLER_37_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1316_ Inst_RegFile_32x4.mem\[14\]\[2\] Inst_RegFile_32x4.mem\[15\]\[2\] net626 VGND
+ VGND VPWR VPWR _0283_ sky130_fd_sc_hd__mux2_1
XANTENNA_31 FrameStrobe[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_20 EE4END[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_75 S4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 net257 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_86 net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 FrameStrobe[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_97 W6END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 net317 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput193 net193 VGND VGND VPWR VPWR FrameData_O[13] sky130_fd_sc_hd__buf_2
Xoutput171 net171 VGND VGND VPWR VPWR E6BEG[8] sky130_fd_sc_hd__buf_2
Xoutput182 net182 VGND VGND VPWR VPWR EE4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput160 net160 VGND VGND VPWR VPWR E2BEGb[7] sky130_fd_sc_hd__buf_2
XFILLER_70_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1101_ Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__inv_1
X_2150_ net612 net936 _0927_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__mux2_2
X_2081_ net599 net831 _0913_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1934_ Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q _0816_ _0818_ _0814_ VGND VGND
+ VPWR VPWR _0819_ sky130_fd_sc_hd__a31o_1
XFILLER_34_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput95 S2END[4] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_2
Xinput40 FrameData[23] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
Xinput51 FrameData[5] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_2
X_1796_ net67 net95 net23 net123 Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q
+ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__mux4_2
X_1865_ Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q net637 VGND VGND VPWR VPWR _0780_
+ sky130_fd_sc_hd__or2_1
Xinput84 NN4END[1] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_2
Xinput73 N2MID[2] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_2
Xinput62 N1END[3] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_4
X_2348_ net751 net691 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2417_ net744 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2279_ net45 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_27_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1650_ net677 net633 net664 net638 Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q
+ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__mux4_1
XFILLER_7_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1581_ Inst_RegFile_32x4.mem\[12\]\[2\] Inst_RegFile_32x4.mem\[13\]\[2\] net605 VGND
+ VGND VPWR VPWR _0532_ sky130_fd_sc_hd__mux2_1
X_2202_ clknet_4_5_0_UserCLK_regs _0026_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[30\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2064_ _0830_ _0906_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__nor2_2
X_2133_ net617 net828 _0924_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__mux2_1
X_1917_ net664 _0437_ Inst_RegFile_switch_matrix.JW2BEG2 _0803_ Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q
+ Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.N1BEG3
+ sky130_fd_sc_hd__mux4_1
XFILLER_34_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2897_ net106 VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__buf_1
XFILLER_22_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2966_ WW4END[7] VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__buf_1
X_1848_ _0762_ _0765_ Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.E6BEG0 sky130_fd_sc_hd__mux2_1
X_1779_ net75 net103 net17 Inst_RegFile_switch_matrix.JS2BEG4 Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__mux4_2
XFILLER_69_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2751_ E6END[7] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_1
X_2820_ FrameStrobe[14] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_46_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1633_ _0578_ _0579_ Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q VGND VGND VPWR VPWR
+ _0580_ sky130_fd_sc_hd__mux2_1
X_1702_ net65 net1 net81 net7 Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q
+ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__mux4_1
X_2682_ clknet_4_1_0_UserCLK_regs _0084_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[31\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1564_ _0516_ _0515_ net684 VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__mux2_4
X_1495_ Inst_RegFile_32x4.mem\[30\]\[0\] Inst_RegFile_32x4.mem\[31\]\[0\] net604 VGND
+ VGND VPWR VPWR _0452_ sky130_fd_sc_hd__mux2_1
X_2116_ net599 net838 _0920_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__mux2_1
X_2047_ net600 net879 _0903_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__mux2_1
X_2949_ net133 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1280_ _0247_ _0248_ net675 VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2803_ net752 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_2
X_2734_ Inst_RegFile_switch_matrix.E2BEG4 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_14_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2596_ net756 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1616_ net82 net23 Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q VGND VGND VPWR VPWR
+ _0564_ sky130_fd_sc_hd__mux2_1
X_2665_ net749 net738 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_6_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1547_ Inst_RegFile_32x4.mem\[28\]\[3\] Inst_RegFile_32x4.mem\[29\]\[3\] net603 VGND
+ VGND VPWR VPWR _0500_ sky130_fd_sc_hd__mux2_1
XFILLER_67_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1478_ _0179_ Inst_RegFile_switch_matrix.JS2BEG6 Inst_RegFile_switch_matrix.JN2BEG6
+ Inst_RegFile_switch_matrix.JW2BEG6 Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q
+ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_40_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout750 net47 VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__clkbuf_4
Xfanout761 net38 VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__buf_4
Xfanout772 net31 VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__clkbuf_4
Xhold270 Inst_RegFile_32x4.mem\[19\]\[3\] VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 Inst_RegFile_32x4.mem\[13\]\[3\] VGND VGND VPWR VPWR net867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 Inst_RegFile_32x4.mem\[5\]\[2\] VGND VGND VPWR VPWR net856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_154 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_143 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_110 _0133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_165 E6END[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_121 net755 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_176 N4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_187 net762 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_198 net326 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1401_ _0360_ Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q _0362_ _0347_ _0349_ VGND
+ VGND VPWR VPWR _0363_ sky130_fd_sc_hd__a32o_2
X_2450_ net743 net705 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2381_ net748 net697 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1194_ Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q _0168_ VGND VGND VPWR VPWR _0169_
+ sky130_fd_sc_hd__or2_1
Xinput5 E2END[0] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_19_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1263_ net661 _0231_ _0233_ _0164_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__o211a_1
X_1332_ Inst_RegFile_32x4.mem\[28\]\[2\] Inst_RegFile_32x4.mem\[29\]\[2\] net624 VGND
+ VGND VPWR VPWR _0299_ sky130_fd_sc_hd__mux2_1
XFILLER_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2717_ clknet_4_3_0_UserCLK_regs _0119_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2579_ net742 net720 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2648_ net770 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput375 net375 VGND VGND VPWR VPWR W6BEG[7] sky130_fd_sc_hd__buf_2
Xoutput353 net353 VGND VGND VPWR VPWR W2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput331 net331 VGND VGND VPWR VPWR SS4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput320 net320 VGND VGND VPWR VPWR S4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput342 net342 VGND VGND VPWR VPWR SS4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput364 net364 VGND VGND VPWR VPWR W2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput386 net386 VGND VGND VPWR VPWR WW4BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_70_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1950_ _0832_ _0833_ _0834_ Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q VGND VGND
+ VPWR VPWR _0835_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_16_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1881_ net59 net1 net115 net422 Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q
+ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__mux4_1
X_2502_ net753 net707 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2364_ net765 net690 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2433_ net759 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1315_ Inst_RegFile_32x4.mem\[12\]\[2\] Inst_RegFile_32x4.mem\[13\]\[2\] net626 VGND
+ VGND VPWR VPWR _0282_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1246_ _0938_ _0217_ Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q VGND VGND VPWR VPWR
+ _0218_ sky130_fd_sc_hd__o21a_1
X_1177_ net676 net635 net666 net409 Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q
+ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__mux4_1
X_2295_ net31 net732 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_24_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_54 net259 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 E6END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 FrameStrobe[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_43 FrameStrobe[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 EE4END[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_65 net320 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput161 net161 VGND VGND VPWR VPWR E6BEG[0] sky130_fd_sc_hd__buf_2
Xoutput150 net150 VGND VGND VPWR VPWR E2BEG[5] sky130_fd_sc_hd__buf_6
XANTENNA_87 net375 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 net336 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 W6END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput194 net194 VGND VGND VPWR VPWR FrameData_O[14] sky130_fd_sc_hd__buf_2
Xoutput172 net172 VGND VGND VPWR VPWR E6BEG[9] sky130_fd_sc_hd__buf_2
Xoutput183 net183 VGND VGND VPWR VPWR EE4BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1100_ Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__inv_2
XFILLER_19_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2080_ _0893_ _0904_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__nand2_4
X_1933_ net111 _1019_ _0817_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__o21ai_1
Xinput96 S2END[5] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_6
Xinput41 FrameData[24] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
X_1795_ _0717_ _0722_ Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.W6BEG0 sky130_fd_sc_hd__mux2_1
Xinput30 FrameData[12] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_2
Xinput52 FrameData[6] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_2
X_1864_ _0708_ _0584_ Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q VGND VGND VPWR VPWR
+ _0779_ sky130_fd_sc_hd__mux2_4
Xinput74 N2MID[3] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
Xinput85 NN4END[2] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_4
Xinput63 N2END[0] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_2
X_2278_ net754 net729 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2347_ net763 net691 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2416_ net745 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_52_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1229_ net675 _0201_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__or2_1
XFILLER_40_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_35_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_44_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1580_ _0529_ _0530_ net413 VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__mux2_4
XFILLER_66_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2201_ clknet_4_1_0_UserCLK_regs _0025_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[30\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2132_ net601 net819 _0924_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_53_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2063_ net613 net887 _0908_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_62_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1847_ _0764_ _0763_ Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q VGND VGND VPWR VPWR
+ _0765_ sky130_fd_sc_hd__mux2_1
X_2896_ net105 VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__buf_1
X_1916_ net65 net80 net777 net676 Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.N4BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_30_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2965_ WW4END[6] VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__buf_1
X_1778_ _0706_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__clkinv_2
XFILLER_1_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_71_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclone22 net634 VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2750_ E6END[6] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_1
X_1701_ _0994_ _0638_ Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q VGND VGND VPWR VPWR
+ _0639_ sky130_fd_sc_hd__o21a_1
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2681_ clknet_4_5_0_UserCLK_regs _0083_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[29\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1632_ net778 net95 net123 net140 Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q
+ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__mux4_1
X_1563_ Inst_RegFile_32x4.mem\[12\]\[3\] Inst_RegFile_32x4.mem\[13\]\[3\] net605 VGND
+ VGND VPWR VPWR _0516_ sky130_fd_sc_hd__mux2_2
X_1494_ _0449_ _0450_ net412 VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__mux2_1
XFILLER_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2115_ _0889_ _0895_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__nand2_4
X_2046_ _0889_ _0902_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__nand2_4
X_2879_ Inst_RegFile_switch_matrix.S1BEG1 VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__clkbuf_2
X_2948_ net132 VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__buf_1
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2802_ net754 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_2
X_2733_ Inst_RegFile_switch_matrix.E2BEG3 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_1
X_2664_ net750 net738 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_14_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1477_ _0431_ _0429_ _0434_ _0934_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JN2BEG6
+ sky130_fd_sc_hd__a22o_4
X_2595_ net757 net720 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1615_ Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q net110 Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q
+ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_6_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1546_ _0497_ _0498_ net681 VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__mux2_1
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2029_ net615 net917 _0896_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__mux2_4
XFILLER_40_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold271 Inst_RegFile_32x4.mem\[13\]\[1\] VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold260 Inst_RegFile_32x4.mem\[20\]\[0\] VGND VGND VPWR VPWR net835 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout762 net37 VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__buf_4
XFILLER_58_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout773 net30 VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__clkbuf_4
Xfanout751 net46 VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__buf_4
Xfanout740 FrameStrobe[0] VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__buf_2
Xhold293 Inst_RegFile_32x4.mem\[27\]\[0\] VGND VGND VPWR VPWR net868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 Inst_RegFile_32x4.mem\[15\]\[1\] VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_177 net284 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_199 _0718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_155 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_111 _0213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_188 net777 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_144 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_166 E6END[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_122 net755 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_100 WW4END[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1400_ Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q _0361_ VGND VGND VPWR VPWR _0362_
+ sky130_fd_sc_hd__or2_1
X_2380_ net46 net697 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1331_ net648 _0297_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__nand2_1
X_1193_ net687 net669 net656 net651 Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q
+ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__mux4_1
Xinput6 E2END[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_19_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1262_ net675 _0232_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__or2_1
X_2647_ net772 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput332 net332 VGND VGND VPWR VPWR SS4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput321 net321 VGND VGND VPWR VPWR S4BEG[2] sky130_fd_sc_hd__buf_2
X_2716_ clknet_4_2_0_UserCLK_regs _0118_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput343 net343 VGND VGND VPWR VPWR SS4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput310 net310 VGND VGND VPWR VPWR S2BEGb[5] sky130_fd_sc_hd__buf_2
X_2578_ net743 net720 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput376 net376 VGND VGND VPWR VPWR W6BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1529_ Inst_RegFile_32x4.mem\[12\]\[1\] Inst_RegFile_32x4.mem\[13\]\[1\] net410 VGND
+ VGND VPWR VPWR _0484_ sky130_fd_sc_hd__mux2_1
Xoutput365 net365 VGND VGND VPWR VPWR W2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput354 net354 VGND VGND VPWR VPWR W2BEG[4] sky130_fd_sc_hd__buf_4
Xoutput387 net387 VGND VGND VPWR VPWR WW4BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_70_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_443 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1880_ net641 _1033_ net685 _0791_ Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q
+ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2501_ net755 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2363_ net766 net690 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2294_ net30 net732 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2432_ net760 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1314_ _0279_ _0280_ net675 VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__mux2_1
X_1245_ net422 net680 net667 net641 Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q
+ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1176_ Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q _0151_ VGND VGND VPWR VPWR _0152_
+ sky130_fd_sc_hd__or2_4
XANTENNA_11 E6END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 net263 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 FrameStrobe[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_22 EE4END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 net377 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_99 WW4END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_66 net321 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 net343 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput195 net195 VGND VGND VPWR VPWR FrameData_O[15] sky130_fd_sc_hd__buf_2
Xoutput162 net162 VGND VGND VPWR VPWR E6BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput184 net184 VGND VGND VPWR VPWR EE4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput173 net173 VGND VGND VPWR VPWR EE4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput151 net151 VGND VGND VPWR VPWR E2BEG[6] sky130_fd_sc_hd__buf_4
XFILLER_28_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput31 FrameData[13] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
X_1863_ net62 net779 net90 net654 Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q
+ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__mux4_1
X_1932_ net79 Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q
+ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__o21ba_1
Xinput20 E2MID[7] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
Xinput97 S2END[6] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
Xinput42 FrameData[25] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
X_1794_ _0721_ _0720_ Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q VGND VGND VPWR VPWR
+ _0722_ sky130_fd_sc_hd__mux2_1
Xinput53 FrameData[7] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_2
X_2415_ net51 net699 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput75 N2MID[4] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_2
Xinput64 N2END[1] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_2
Xinput86 NN4END[3] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_2
X_2277_ net44 net729 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2346_ net776 net691 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_27_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1228_ Inst_RegFile_32x4.mem\[22\]\[0\] Inst_RegFile_32x4.mem\[23\]\[0\] net627 VGND
+ VGND VPWR VPWR _0201_ sky130_fd_sc_hd__mux2_1
XFILLER_52_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1159_ Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q _0132_ _0134_ _1032_ _1034_ VGND
+ VGND VPWR VPWR _0136_ sky130_fd_sc_hd__a32o_1
XFILLER_25_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2062_ net623 net889 _0908_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__mux2_1
X_2200_ clknet_4_1_0_UserCLK_regs _0024_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[30\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2131_ _0859_ _0923_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_49_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2964_ WW4END[5] VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__buf_1
X_1846_ net679 net636 net667 net640 Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q
+ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__mux4_1
X_1915_ net66 net81 net778 net665 Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.N4BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_30_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1777_ Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q _0703_ _0704_ _0705_ VGND VGND VPWR
+ VPWR _0706_ sky130_fd_sc_hd__a2bb2o_2
X_2895_ net104 VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__buf_1
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2329_ net769 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1700_ net677 net633 net664 net638 Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q
+ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__mux4_1
X_1631_ net67 net79 net780 net9 Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q
+ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__mux4_1
X_2680_ clknet_4_5_0_UserCLK_regs _0082_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[29\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1493_ Inst_RegFile_32x4.mem\[26\]\[0\] Inst_RegFile_32x4.mem\[27\]\[0\] net604 VGND
+ VGND VPWR VPWR _0450_ sky130_fd_sc_hd__mux2_1
X_1562_ Inst_RegFile_32x4.mem\[14\]\[3\] Inst_RegFile_32x4.mem\[15\]\[3\] net605 VGND
+ VGND VPWR VPWR _0515_ sky130_fd_sc_hd__mux2_2
XFILLER_39_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2114_ net613 net845 _0919_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__mux2_1
X_2045_ _0901_ _0829_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__nor2_8
XFILLER_62_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2947_ net131 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkbuf_2
X_1829_ _0748_ _0747_ Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.SS4BEG0 sky130_fd_sc_hd__mux2_1
X_2878_ Inst_RegFile_switch_matrix.S1BEG0 VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_9_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_8_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_8_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_71_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2801_ net755 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2594_ net758 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1614_ Inst_RegFile_switch_matrix.JN2BEG4 _0935_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__nor2_2
X_2732_ Inst_RegFile_switch_matrix.E2BEG2 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
X_2663_ net752 net740 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_14_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1476_ _0432_ _0433_ Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q VGND VGND VPWR VPWR
+ _0434_ sky130_fd_sc_hd__mux2_1
XFILLER_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1545_ Inst_RegFile_32x4.mem\[26\]\[3\] Inst_RegFile_32x4.mem\[27\]\[3\] net604 VGND
+ VGND VPWR VPWR _0498_ sky130_fd_sc_hd__mux2_1
XFILLER_35_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2028_ net599 net902 _0896_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__mux2_4
XFILLER_50_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold283 Inst_RegFile_32x4.mem\[31\]\[2\] VGND VGND VPWR VPWR net858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 Inst_RegFile_32x4.mem\[13\]\[2\] VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 Inst_RegFile_32x4.mem\[23\]\[0\] VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 Inst_RegFile_32x4.mem\[13\]\[0\] VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold250 Inst_RegFile_32x4.mem\[4\]\[2\] VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout730 net731 VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__clkbuf_2
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout774 net29 VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__buf_4
Xfanout763 net36 VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__clkbuf_4
Xfanout741 FrameStrobe[0] VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__clkbuf_2
Xfanout752 net45 VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_56_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_189 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_112 _0213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_156 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_145 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_123 net755 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_167 EE4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_101 WW4END[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_178 NN4END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1261_ Inst_RegFile_32x4.mem\[2\]\[0\] Inst_RegFile_32x4.mem\[3\]\[0\] net627 VGND
+ VGND VPWR VPWR _0232_ sky130_fd_sc_hd__mux2_1
X_1330_ _0295_ _0296_ net674 VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__mux2_1
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 E2END[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_19_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1192_ net648 _0166_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__nand2_1
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2646_ net773 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2577_ net744 net718 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput377 net377 VGND VGND VPWR VPWR W6BEG[9] sky130_fd_sc_hd__buf_2
Xoutput366 net366 VGND VGND VPWR VPWR W6BEG[0] sky130_fd_sc_hd__buf_2
Xoutput333 Inst_RegFile_switch_matrix.SS4BEG1 VGND VGND VPWR VPWR SS4BEG[13] sky130_fd_sc_hd__buf_8
Xoutput322 net322 VGND VGND VPWR VPWR S4BEG[3] sky130_fd_sc_hd__buf_2
X_2715_ clknet_4_2_0_UserCLK_regs _0117_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput300 net300 VGND VGND VPWR VPWR S2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput311 net311 VGND VGND VPWR VPWR S2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput344 net344 VGND VGND VPWR VPWR SS4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput355 Inst_RegFile_switch_matrix.JW2BEG5 VGND VGND VPWR VPWR W2BEG[5] sky130_fd_sc_hd__buf_8
XFILLER_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1528_ Inst_RegFile_32x4.mem\[14\]\[1\] Inst_RegFile_32x4.mem\[15\]\[1\] net410 VGND
+ VGND VPWR VPWR _0483_ sky130_fd_sc_hd__mux2_1
X_1459_ Inst_RegFile_32x4.mem\[6\]\[0\] Inst_RegFile_32x4.mem\[7\]\[0\] net609 VGND
+ VGND VPWR VPWR _0417_ sky130_fd_sc_hd__mux2_1
Xoutput388 net388 VGND VGND VPWR VPWR WW4BEG[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_53_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2500_ net43 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2431_ net761 net701 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2362_ net767 net690 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1244_ Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q _0215_ VGND VGND VPWR VPWR _0216_
+ sky130_fd_sc_hd__or2_1
X_2293_ net29 net732 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1313_ Inst_RegFile_32x4.mem\[8\]\[2\] Inst_RegFile_32x4.mem\[9\]\[2\] net629 VGND
+ VGND VPWR VPWR _0280_ sky130_fd_sc_hd__mux2_1
XFILLER_64_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1175_ net687 net671 net658 net652 Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q
+ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__mux4_2
XFILLER_37_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_45 net224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 W6END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_12 E6END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 net270 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 FrameStrobe[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 EE4END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 SS4END[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 net323 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2629_ net755 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput196 net196 VGND VGND VPWR VPWR FrameData_O[16] sky130_fd_sc_hd__buf_2
Xoutput163 Inst_RegFile_switch_matrix.E6BEG1 VGND VGND VPWR VPWR E6BEG[11] sky130_fd_sc_hd__buf_6
Xoutput174 net174 VGND VGND VPWR VPWR EE4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput185 net185 VGND VGND VPWR VPWR EE4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput152 net152 VGND VGND VPWR VPWR E2BEG[7] sky130_fd_sc_hd__buf_4
Xoutput141 net141 VGND VGND VPWR VPWR E1BEG[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput43 FrameData[26] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
Xinput32 FrameData[16] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
X_1793_ net411 net415 net664 net638 Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q
+ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__mux4_1
Xinput54 FrameData[8] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_4
X_1862_ _1011_ _0773_ _0777_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.EE4BEG2
+ sky130_fd_sc_hd__o21a_1
Xinput21 E6END[0] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlymetal6s2s_1
X_1931_ _1019_ Inst_RegFile_switch_matrix.JW2BEG2 _0815_ VGND VGND VPWR VPWR _0816_
+ sky130_fd_sc_hd__o21ai_1
Xinput10 E2END[5] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_6
Xinput98 S2END[7] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_2
Xinput87 S1END[0] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_2
XFILLER_69_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2414_ net50 net699 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput76 N2MID[5] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_2
Xinput65 N2END[2] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_4
X_2276_ net756 net729 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2345_ net749 net734 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1158_ _0132_ Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q _0134_ _1032_ _1034_ VGND
+ VGND VPWR VPWR _0135_ sky130_fd_sc_hd__a32oi_4
X_1227_ _0198_ _0199_ net662 VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__mux2_1
X_1089_ Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__inv_1
XFILLER_52_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2061_ net617 net840 _0908_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__mux2_1
XFILLER_19_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2130_ _0830_ _0897_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__nor2_8
X_1914_ net63 net686 net82 net415 Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.N4BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_34_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2963_ WW4END[4] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__buf_1
X_1845_ _0718_ _0719_ _1033_ net685 Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q
+ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__mux4_1
X_1776_ _0950_ Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q
+ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__o21a_1
X_2894_ net103 VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__buf_1
X_2328_ net771 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_72_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2259_ net742 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_25_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1630_ Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q _0574_ Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q
+ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__o21a_1
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1492_ Inst_RegFile_32x4.mem\[24\]\[0\] Inst_RegFile_32x4.mem\[25\]\[0\] net603 VGND
+ VGND VPWR VPWR _0449_ sky130_fd_sc_hd__mux2_1
X_1561_ _0512_ _0513_ net681 VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__mux2_4
XFILLER_47_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2113_ net622 net842 _0919_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__mux2_1
X_2044_ _0821_ _0810_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_45_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2946_ net130 VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__buf_1
XFILLER_22_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1759_ net59 net63 net83 net1 Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q
+ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__mux4_1
X_1828_ net61 net780 net689 net660 Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q
+ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__mux4_1
XFILLER_1_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2800_ net43 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__buf_1
XFILLER_44_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2731_ Inst_RegFile_switch_matrix.E2BEG1 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_14_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2593_ net40 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1613_ Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q _0559_ _0561_ _0557_ VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix.JN2BEG4 sky130_fd_sc_hd__o31ai_4
X_2662_ net753 net740 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1544_ Inst_RegFile_32x4.mem\[24\]\[3\] Inst_RegFile_32x4.mem\[25\]\[3\] net604 VGND
+ VGND VPWR VPWR _0497_ sky130_fd_sc_hd__mux2_1
XFILLER_12_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1475_ net12 net90 net98 net116 Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q
+ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__mux4_1
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_59_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2027_ net593 _0895_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__nand2_8
X_2929_ Inst_RegFile_switch_matrix.SS4BEG3 VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__clkbuf_2
Xfanout720 net721 VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_68_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout742 net55 VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__clkbuf_4
Xfanout731 net732 VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__buf_2
Xhold284 Inst_RegFile_32x4.mem\[15\]\[2\] VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 Inst_RegFile_32x4.mem\[3\]\[0\] VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 Inst_RegFile_32x4.mem\[11\]\[1\] VGND VGND VPWR VPWR net870 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold251 Inst_RegFile_32x4.mem\[26\]\[0\] VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 Inst_RegFile_32x4.mem\[26\]\[3\] VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 Inst_RegFile_32x4.mem\[5\]\[0\] VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout753 net754 VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__buf_4
XFILLER_65_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout764 net35 VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__buf_4
Xfanout775 net28 VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__buf_4
XANTENNA_113 _0213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_124 net755 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_102 WW4END[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_135 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_146 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_157 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_168 EE4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_179 net326 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput8 E2END[3] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
X_1260_ Inst_RegFile_32x4.mem\[0\]\[0\] Inst_RegFile_32x4.mem\[1\]\[0\] net627 VGND
+ VGND VPWR VPWR _0231_ sky130_fd_sc_hd__mux2_1
X_1191_ _0137_ _0165_ net396 VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__mux2_1
XFILLER_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2714_ clknet_4_2_0_UserCLK_regs _0116_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput345 net345 VGND VGND VPWR VPWR UserCLKo sky130_fd_sc_hd__buf_1
X_2645_ net774 net740 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2576_ net745 net718 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput367 net367 VGND VGND VPWR VPWR W6BEG[10] sky130_fd_sc_hd__buf_4
Xoutput312 net312 VGND VGND VPWR VPWR S2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput334 net334 VGND VGND VPWR VPWR SS4BEG[14] sky130_fd_sc_hd__buf_8
Xoutput301 net301 VGND VGND VPWR VPWR S2BEG[4] sky130_fd_sc_hd__buf_8
Xoutput323 net323 VGND VGND VPWR VPWR S4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput356 net356 VGND VGND VPWR VPWR W2BEG[6] sky130_fd_sc_hd__buf_4
X_1527_ _0480_ _0481_ net413 VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__mux2_1
Xoutput378 net378 VGND VGND VPWR VPWR WW4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput389 net389 VGND VGND VPWR VPWR WW4BEG[5] sky130_fd_sc_hd__buf_2
X_1389_ net421 net637 net667 net641 Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q
+ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__mux4_2
XFILLER_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1458_ net619 VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_53_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2361_ net768 net691 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2430_ net762 net701 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1243_ net688 net672 net659 net653 Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q
+ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__mux4_1
X_2292_ net28 net730 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1174_ Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q _0146_ _0149_ VGND VGND VPWR VPWR
+ _0150_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_22_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1312_ Inst_RegFile_32x4.mem\[10\]\[2\] Inst_RegFile_32x4.mem\[11\]\[2\] net629 VGND
+ VGND VPWR VPWR _0279_ sky130_fd_sc_hd__mux2_1
XANTENNA_13 E6END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_46 net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 FrameStrobe[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 EE4END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_79 net346 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 net324 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 N4END[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2628_ net756 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput197 net197 VGND VGND VPWR VPWR FrameData_O[17] sky130_fd_sc_hd__buf_2
X_2559_ net761 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput164 net164 VGND VGND VPWR VPWR E6BEG[1] sky130_fd_sc_hd__buf_2
Xoutput175 net175 VGND VGND VPWR VPWR EE4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput186 net186 VGND VGND VPWR VPWR EE4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput153 net153 VGND VGND VPWR VPWR E2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput142 net142 VGND VGND VPWR VPWR E1BEG[1] sky130_fd_sc_hd__buf_4
XFILLER_28_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1930_ net135 Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q
+ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__o21a_1
Xinput88 S1END[1] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_6
Xinput44 FrameData[27] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
Xinput33 FrameData[17] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_2
X_1792_ _0718_ _0719_ _1033_ net685 Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q
+ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__mux4_1
Xinput55 FrameData[9] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_2
X_1861_ _0774_ _0775_ _0776_ Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q
+ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__a221o_1
Xinput22 E6END[1] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
Xinput11 E2END[6] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_4
Xinput77 N2MID[6] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_2
Xinput66 N2END[3] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_4
Xinput99 S2MID[0] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2344_ net750 net734 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2413_ net49 net700 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2275_ net757 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_63_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1157_ Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q _0133_ VGND VGND VPWR VPWR _0134_
+ sky130_fd_sc_hd__or2_1
XFILLER_25_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1226_ Inst_RegFile_32x4.mem\[18\]\[0\] Inst_RegFile_32x4.mem\[19\]\[0\] net631 VGND
+ VGND VPWR VPWR _0199_ sky130_fd_sc_hd__mux2_1
XFILLER_52_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1088_ Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__inv_1
XFILLER_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2060_ net601 net844 _0908_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__mux2_1
X_2962_ Inst_RegFile_switch_matrix.W6BEG1 VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_60_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1913_ net64 net79 net687 net409 Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.N4BEG3 sky130_fd_sc_hd__mux4_1
X_2893_ net102 VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_32_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1844_ Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q _0757_ _0760_ _0761_ VGND VGND
+ VPWR VPWR _0762_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_31_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1775_ Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q Inst_RegFile_switch_matrix.JS2BEG3
+ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__nand2_1
XFILLER_57_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2327_ net31 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2258_ net743 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1209_ _0181_ _0182_ Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q VGND VGND VPWR VPWR
+ _0183_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_48_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2189_ clknet_4_1_0_UserCLK_regs _0013_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[27\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1560_ Inst_RegFile_32x4.mem\[10\]\[3\] Inst_RegFile_32x4.mem\[11\]\[3\] net410 VGND
+ VGND VPWR VPWR _0513_ sky130_fd_sc_hd__mux2_2
X_2112_ net617 net886 _0919_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__mux2_1
X_1491_ _0389_ _0443_ _0447_ _0416_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__a211o_1
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2043_ net611 net821 _0900_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__mux2_1
X_2876_ Inst_RegFile_switch_matrix.NN4BEG2 VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__clkbuf_2
X_1827_ net667 _0718_ _0719_ _0401_ Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q
+ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__mux4_1
X_2945_ net129 VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__buf_4
XFILLER_30_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1758_ Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q _0688_ Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q
+ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__o21a_1
X_1689_ _0623_ _0625_ _0628_ _0991_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JS2BEG1
+ sky130_fd_sc_hd__a22o_1
XFILLER_57_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2661_ net44 net741 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2730_ Inst_RegFile_switch_matrix.E2BEG0 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
XFILLER_8_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1474_ net62 net70 net84 net779 Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q
+ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__mux4_1
X_2592_ net760 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1612_ _0936_ _0560_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__nor2_1
X_1543_ net643 _0495_ _0492_ _0416_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__a211o_1
XFILLER_50_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2026_ _0822_ _0830_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__nor2_2
X_2859_ Inst_RegFile_switch_matrix.N4BEG1 VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_1
X_2928_ Inst_RegFile_switch_matrix.SS4BEG2 VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__buf_6
XFILLER_40_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout754 FrameData[28] VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__buf_2
Xfanout721 net57 VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__clkbuf_2
Xfanout710 net711 VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__clkbuf_2
Xfanout765 net34 VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__buf_4
Xfanout732 FrameStrobe[11] VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__clkbuf_2
Xfanout776 net27 VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__buf_4
Xfanout743 net54 VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__buf_4
Xhold241 Inst_RegFile_32x4.mem\[18\]\[0\] VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 Inst_RegFile_32x4.mem\[29\]\[1\] VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 Inst_RegFile_32x4.mem\[1\]\[3\] VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 Inst_RegFile_32x4.mem\[29\]\[0\] VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 Inst_RegFile_32x4.mem\[20\]\[1\] VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 Inst_RegFile_32x4.mem\[20\]\[3\] VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_114 _0707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 net762 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_136 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_147 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_158 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_103 WW4END[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_169 net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_4_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_4_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_5_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 E2END[4] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1190_ Inst_RegFile_32x4.mem\[24\]\[0\] Inst_RegFile_32x4.mem\[25\]\[0\] net624 VGND
+ VGND VPWR VPWR _0165_ sky130_fd_sc_hd__mux2_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2644_ net775 net740 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2713_ clknet_4_10_0_UserCLK_regs _0115_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2575_ net746 net718 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput368 net368 VGND VGND VPWR VPWR W6BEG[11] sky130_fd_sc_hd__buf_4
X_1457_ _0412_ Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q _0414_ VGND VGND VPWR VPWR
+ _0415_ sky130_fd_sc_hd__a21oi_2
Xoutput379 net379 VGND VGND VPWR VPWR WW4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput346 net346 VGND VGND VPWR VPWR W1BEG[0] sky130_fd_sc_hd__buf_4
Xoutput313 net313 VGND VGND VPWR VPWR S4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput335 net335 VGND VGND VPWR VPWR SS4BEG[15] sky130_fd_sc_hd__buf_4
Xoutput302 Inst_RegFile_switch_matrix.JS2BEG5 VGND VGND VPWR VPWR S2BEG[5] sky130_fd_sc_hd__buf_6
X_1526_ Inst_RegFile_32x4.mem\[10\]\[1\] Inst_RegFile_32x4.mem\[11\]\[1\] net608 VGND
+ VGND VPWR VPWR _0481_ sky130_fd_sc_hd__mux2_1
Xoutput324 net324 VGND VGND VPWR VPWR S4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput357 net357 VGND VGND VPWR VPWR W2BEG[7] sky130_fd_sc_hd__buf_4
X_1388_ Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q _0350_ VGND VGND VPWR VPWR _0351_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_53_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2009_ _0831_ _0889_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__nand2_8
XFILLER_2_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2360_ net771 net691 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2291_ net55 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1311_ Inst_RegFile_32x4.AD_comb\[1\] Inst_RegFile_32x4.AD_reg\[1\] Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q
+ VGND VGND VPWR VPWR AD1 sky130_fd_sc_hd__mux2_4
XFILLER_37_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1242_ _0213_ Inst_RegFile_switch_matrix.JN2BEG5 Inst_RegFile_switch_matrix.JS2BEG5
+ Inst_RegFile_switch_matrix.JW2BEG5 Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q
+ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__mux4_1
X_1173_ Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q _0148_ Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q
+ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_14 E6END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 FrameStrobe[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_25 EE4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 Inst_RegFile_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2627_ net757 net724 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput143 net143 VGND VGND VPWR VPWR E1BEG[2] sky130_fd_sc_hd__buf_4
XFILLER_21_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_69 net327 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_58 N4END[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput198 net198 VGND VGND VPWR VPWR FrameData_O[18] sky130_fd_sc_hd__buf_2
X_2558_ net762 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput165 net165 VGND VGND VPWR VPWR E6BEG[2] sky130_fd_sc_hd__buf_2
Xoutput176 net176 VGND VGND VPWR VPWR EE4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput187 net187 VGND VGND VPWR VPWR EE4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput154 net154 VGND VGND VPWR VPWR E2BEGb[1] sky130_fd_sc_hd__buf_2
X_2489_ net768 net706 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1509_ net643 _0463_ _0460_ _0416_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__a211o_1
XFILLER_43_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1860_ net87 net422 Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q VGND VGND VPWR VPWR
+ _0776_ sky130_fd_sc_hd__mux2_1
XFILLER_36_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput89 S1END[2] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
Xinput45 FrameData[29] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
Xinput34 FrameData[18] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_4
Xinput12 E2END[7] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
X_1791_ net74 net16 net102 net130 Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q
+ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__mux4_2
Xinput23 EE4END[0] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
Xinput67 N2END[4] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_2
Xinput78 N2MID[7] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_2
Xinput56 FrameStrobe[12] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2274_ net758 net729 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2343_ net752 net734 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2412_ net46 net700 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_63_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1156_ net66 net8 net94 net138 Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q
+ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__mux4_2
X_1087_ Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__inv_1
XFILLER_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1225_ Inst_RegFile_32x4.mem\[16\]\[0\] Inst_RegFile_32x4.mem\[17\]\[0\] net631 VGND
+ VGND VPWR VPWR _0198_ sky130_fd_sc_hd__mux2_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1989_ _0870_ _0872_ Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q VGND VGND VPWR VPWR
+ _0873_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2961_ Inst_RegFile_switch_matrix.W6BEG0 VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__buf_1
X_1843_ Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q _0758_ Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q
+ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_60_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1912_ net421 Inst_RegFile_switch_matrix.JN2BEG3 _0804_ _0805_ Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E1BEG0
+ sky130_fd_sc_hd__mux4_1
X_2892_ net101 VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_32_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1774_ net75 net17 Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q VGND VGND VPWR VPWR
+ _0703_ sky130_fd_sc_hd__mux2_1
X_1208_ net646 net679 net636 net640 Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q
+ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__mux4_2
X_2326_ net30 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2257_ net744 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_27_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1139_ net15 _0965_ _1029_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__o21a_1
XFILLER_25_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2188_ clknet_4_1_0_UserCLK_regs _0012_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[27\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclone15 _0163_ VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__buf_6
XFILLER_44_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1490_ net682 _0446_ _0445_ net643 VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__o211a_1
XFILLER_39_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2111_ net601 net861 _0919_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__mux2_1
X_2042_ net620 net850 _0900_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__mux2_1
XFILLER_62_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1826_ _0745_ _0746_ Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.SS4BEG1 sky130_fd_sc_hd__mux2_4
X_2944_ net128 VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__clkbuf_1
X_1757_ net689 net669 net656 net651 Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q
+ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1688_ _0626_ _0627_ Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q VGND VGND VPWR VPWR
+ _0628_ sky130_fd_sc_hd__mux2_1
X_2309_ net44 net730 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_12_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_12_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_5_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1611_ net10 net88 net96 net116 Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q
+ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__mux4_1
X_2660_ net756 net741 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_42_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1473_ Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q _0430_ Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q
+ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__o21a_1
X_2591_ net38 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1542_ _0494_ _0493_ net682 VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__mux2_1
XFILLER_39_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2025_ net611 net883 _0894_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__mux2_1
XFILLER_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1809_ _0719_ _0386_ Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q VGND VGND VPWR VPWR
+ _0733_ sky130_fd_sc_hd__mux2_1
X_2789_ net769 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
X_2858_ Inst_RegFile_switch_matrix.N4BEG0 VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__buf_1
Xhold253 Inst_RegFile_32x4.mem\[4\]\[1\] VGND VGND VPWR VPWR net828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 Inst_RegFile_32x4.mem\[15\]\[3\] VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout711 net712 VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__clkbuf_2
Xfanout755 net44 VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__buf_4
Xfanout722 net725 VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__buf_2
XFILLER_49_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout733 FrameStrobe[11] VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__buf_2
Xfanout766 net33 VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__buf_4
Xfanout744 net53 VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__buf_4
Xfanout700 FrameStrobe[7] VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__buf_2
Xfanout777 net22 VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__clkbuf_4
Xhold286 Inst_RegFile_32x4.mem\[19\]\[0\] VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 Inst_RegFile_32x4.mem\[30\]\[2\] VGND VGND VPWR VPWR net850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 Inst_RegFile_32x4.mem\[11\]\[3\] VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 Inst_RegFile_32x4.mem\[9\]\[3\] VGND VGND VPWR VPWR net872 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_148 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_115 _0788_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_137 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_126 net766 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_159 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_104 WW4END[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2643_ net55 net740 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2574_ net747 net718 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2712_ clknet_4_8_0_UserCLK_regs _0114_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput303 net303 VGND VGND VPWR VPWR S2BEG[6] sky130_fd_sc_hd__buf_6
Xoutput314 net314 VGND VGND VPWR VPWR S4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput325 net325 VGND VGND VPWR VPWR S4BEG[6] sky130_fd_sc_hd__buf_2
X_1387_ net116 net673 net660 net654 Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q
+ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__mux4_1
Xoutput369 net369 VGND VGND VPWR VPWR W6BEG[1] sky130_fd_sc_hd__buf_2
X_1456_ _0410_ Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q _0413_ VGND VGND VPWR VPWR
+ _0414_ sky130_fd_sc_hd__o21a_1
Xoutput336 net336 VGND VGND VPWR VPWR SS4BEG[1] sky130_fd_sc_hd__buf_2
X_1525_ Inst_RegFile_32x4.mem\[8\]\[1\] Inst_RegFile_32x4.mem\[9\]\[1\] net608 VGND
+ VGND VPWR VPWR _0480_ sky130_fd_sc_hd__mux2_1
Xoutput347 net347 VGND VGND VPWR VPWR W1BEG[1] sky130_fd_sc_hd__buf_4
Xoutput358 net358 VGND VGND VPWR VPWR W2BEGb[0] sky130_fd_sc_hd__buf_2
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2008_ _0858_ _0888_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__nor2_8
XFILLER_51_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2290_ net743 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_49_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1241_ net63 net91 net24 net119 Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q
+ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__mux4_2
X_1310_ _0228_ _0278_ _0270_ _0261_ _0262_ VGND VGND VPWR VPWR Inst_RegFile_32x4.AD_comb\[1\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_52_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1172_ net76 net18 net104 net132 Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q
+ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__mux4_2
XANTENNA_37 FrameStrobe[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 Inst_RegFile_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_26 FrameData[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_15 EE4END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_59 N4END[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2626_ net758 net724 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput166 net166 VGND VGND VPWR VPWR E6BEG[3] sky130_fd_sc_hd__buf_2
Xoutput177 Inst_RegFile_switch_matrix.EE4BEG1 VGND VGND VPWR VPWR EE4BEG[13] sky130_fd_sc_hd__buf_6
X_2557_ net35 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput155 net155 VGND VGND VPWR VPWR E2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput144 net144 VGND VGND VPWR VPWR E1BEG[3] sky130_fd_sc_hd__buf_4
Xoutput199 net199 VGND VGND VPWR VPWR FrameData_O[19] sky130_fd_sc_hd__buf_2
X_1439_ _0397_ _0398_ Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q VGND VGND VPWR VPWR
+ _0399_ sky130_fd_sc_hd__mux2_1
Xoutput188 net188 VGND VGND VPWR VPWR EE4BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2488_ net770 net706 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1508_ _0462_ _0461_ net682 VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1790_ net74 net16 net102 net130 Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q
+ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__mux4_2
Xinput13 E2MID[0] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput35 FrameData[19] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_4
Xinput46 FrameData[2] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
X_2411_ net763 net701 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput24 EE4END[1] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_2
Xinput79 N4END[0] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_2
Xinput68 N2END[5] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_6
Xinput57 FrameStrobe[2] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_2
X_2273_ net759 net729 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2342_ net753 net734 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1224_ net408 _0196_ net395 VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_63_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1086_ Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_35_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1155_ _0130_ _0129_ _0131_ _0970_ _0968_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__a221o_1
XFILLER_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1988_ _0788_ _0871_ Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q VGND VGND VPWR VPWR
+ _0872_ sky130_fd_sc_hd__mux2_1
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2609_ net744 net722 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2960_ W6END[11] VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_60_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1773_ _0700_ _0701_ Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q VGND VGND VPWR VPWR
+ _0702_ sky130_fd_sc_hd__mux2_1
XFILLER_63_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1842_ Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q _0759_ VGND VGND VPWR VPWR _0760_
+ sky130_fd_sc_hd__and2b_1
X_1911_ net676 _0582_ Inst_RegFile_switch_matrix.JN2BEG0 _0158_ Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E1BEG1
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_32_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2891_ net100 VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1207_ net139 net672 net659 net653 Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q
+ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__mux4_1
X_2325_ net29 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2256_ net745 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_27_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2187_ clknet_4_4_0_UserCLK_regs _0011_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[26\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1069_ Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone16 BD3 VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__clkbuf_1
X_1138_ net73 Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q
+ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__o21ba_1
XFILLER_25_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2110_ _0893_ _0907_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__nand2_2
X_2041_ net615 net832 _0900_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__mux2_1
XFILLER_50_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2943_ net127 VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__buf_1
X_1756_ _1007_ _0686_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__or2_1
X_2874_ Inst_RegFile_switch_matrix.NN4BEG0 VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__clkbuf_2
X_1825_ net637 _0707_ _0708_ _0179_ Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q
+ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__mux4_2
X_2308_ net43 net730 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1687_ net93 net109 net121 net138 Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q
+ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__mux4_1
XFILLER_53_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2239_ clknet_4_15_0_UserCLK_regs _0063_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[18\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2590_ net37 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1610_ Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q _0558_ VGND VGND VPWR VPWR _0559_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_14_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1472_ net688 net670 net657 net655 Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q
+ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__mux4_1
XFILLER_39_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1541_ Inst_RegFile_32x4.mem\[20\]\[3\] Inst_RegFile_32x4.mem\[21\]\[3\] net607 VGND
+ VGND VPWR VPWR _0494_ sky130_fd_sc_hd__mux2_1
XFILLER_67_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2024_ net620 net834 _0894_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__mux2_1
XFILLER_50_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2926_ Inst_RegFile_switch_matrix.SS4BEG0 VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_28_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2857_ N4END[15] VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__clkbuf_2
X_1739_ net115 net669 net656 net651 Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q
+ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__mux4_1
X_2788_ net771 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_2
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1808_ _0732_ _0731_ Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.WW4BEG1 sky130_fd_sc_hd__mux2_4
Xhold265 Inst_RegFile_32x4.mem\[17\]\[1\] VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 Inst_RegFile_32x4.mem\[25\]\[0\] VGND VGND VPWR VPWR net829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 Inst_RegFile_32x4.mem\[12\]\[1\] VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 Inst_RegFile_32x4.mem\[6\]\[1\] VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 Inst_RegFile_32x4.mem\[22\]\[0\] VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout712 net713 VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__buf_2
Xfanout723 net725 VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__buf_2
XFILLER_58_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout756 net43 VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__buf_4
Xfanout778 net21 VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__buf_2
Xfanout734 net737 VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__buf_2
Xfanout745 net52 VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_37_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout767 net32 VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__buf_4
Xfanout701 FrameStrobe[7] VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold298 Inst_RegFile_32x4.mem\[1\]\[1\] VGND VGND VPWR VPWR net873 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_116 net623 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_127 net772 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_105 WW4END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2711_ clknet_4_8_0_UserCLK_regs _0113_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2642_ net54 net741 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2573_ net748 net718 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput304 net304 VGND VGND VPWR VPWR S2BEG[7] sky130_fd_sc_hd__buf_4
Xoutput337 net337 VGND VGND VPWR VPWR SS4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput315 net315 VGND VGND VPWR VPWR S4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput326 net326 VGND VGND VPWR VPWR S4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput348 Inst_RegFile_switch_matrix.W1BEG2 VGND VGND VPWR VPWR W1BEG[2] sky130_fd_sc_hd__buf_6
Xoutput359 net359 VGND VGND VPWR VPWR W2BEGb[1] sky130_fd_sc_hd__buf_2
X_1524_ _0475_ _0478_ net643 VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__mux2_1
XFILLER_55_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1386_ _0941_ _0348_ Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q VGND VGND VPWR VPWR
+ _0349_ sky130_fd_sc_hd__o21ba_1
X_1455_ _0954_ _0411_ Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q VGND VGND VPWR VPWR
+ _0413_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_53_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2007_ _0852_ _0838_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__nand2b_4
X_2909_ S4END[15] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1240_ _0209_ _0207_ _0212_ _0962_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JN2BEG5
+ sky130_fd_sc_hd__a22o_4
X_1171_ _0146_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__inv_2
XFILLER_49_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_0_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_0_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_49 net241 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 FrameStrobe[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_27 net195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_16 EE4END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2625_ net40 net726 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput189 net189 VGND VGND VPWR VPWR FrameData_O[0] sky130_fd_sc_hd__buf_2
X_2487_ net772 net707 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput167 net167 VGND VGND VPWR VPWR E6BEG[4] sky130_fd_sc_hd__buf_2
Xoutput178 net178 VGND VGND VPWR VPWR EE4BEG[14] sky130_fd_sc_hd__clkbuf_4
X_2556_ net765 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput156 net156 VGND VGND VPWR VPWR E2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput145 net145 VGND VGND VPWR VPWR E2BEG[0] sky130_fd_sc_hd__buf_4
X_1507_ Inst_RegFile_32x4.mem\[20\]\[1\] Inst_RegFile_32x4.mem\[21\]\[1\] net607 VGND
+ VGND VPWR VPWR _0462_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1438_ net88 net96 net90 net116 Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q
+ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__mux4_1
XFILLER_55_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1369_ _0332_ _0333_ net663 VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__mux2_1
XFILLER_36_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput36 FrameData[1] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_2
XFILLER_42_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput25 EE4END[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_2
Xinput14 E2MID[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput47 FrameData[30] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
X_2410_ net27 net701 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2341_ net755 net734 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput69 N2END[6] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_4
Xinput58 FrameStrobe[8] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_2
X_2272_ net760 net729 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1154_ net85 net7 Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q VGND VGND VPWR VPWR
+ _0131_ sky130_fd_sc_hd__mux2_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1223_ _0194_ _0195_ net663 VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1085_ Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__inv_2
XFILLER_20_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1987_ net25 net126 net109 Inst_RegFile_switch_matrix.E2BEG1 Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__mux4_1
X_2608_ net745 net722 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2539_ net763 net714 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1910_ net666 net685 Inst_RegFile_switch_matrix.JN2BEG1 net394 Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E1BEG2
+ sky130_fd_sc_hd__mux4_2
XFILLER_30_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2890_ net99 VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__buf_1
X_1772_ net670 net655 net657 net645 Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q
+ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__mux4_1
X_1841_ net672 net659 Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q VGND VGND VPWR VPWR
+ _0759_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2324_ net775 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2255_ net746 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1137_ net101 Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q
+ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__o21a_1
X_1206_ _0977_ _0179_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__nand2_1
X_2186_ clknet_4_4_0_UserCLK_regs _0010_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[26\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xclone28 AD3 VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__buf_6
Xclone17 B_ADR0 VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__buf_6
X_1068_ Inst_RegFile_32x4.mem\[22\]\[2\] VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__inv_1
XFILLER_68_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2040_ net599 net843 _0900_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2942_ Inst_RegFile_switch_matrix.JW2BEG7 VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__buf_1
X_2873_ NN4END[15] VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__buf_2
X_1755_ net644 net411 net664 net415 Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q
+ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__mux4_1
X_1824_ net62 net779 net688 net654 Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q
+ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__mux4_1
X_1686_ net65 net7 net1 net778 Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q
+ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__mux4_1
X_2307_ net42 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2238_ clknet_4_13_0_UserCLK_regs _0062_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[18\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_13_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2169_ net621 net874 _0931_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1540_ Inst_RegFile_32x4.mem\[22\]\[3\] Inst_RegFile_32x4.mem\[23\]\[3\] net607 VGND
+ VGND VPWR VPWR _0493_ sky130_fd_sc_hd__mux2_1
XFILLER_8_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1471_ _0933_ _0428_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__or2_4
XFILLER_39_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2023_ net615 net877 _0894_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__mux2_1
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1807_ net62 net90 net688 net423 Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q
+ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__mux4_1
X_2925_ SS4END[15] VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__buf_1
X_2856_ N4END[14] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkbuf_2
Xfanout713 FrameStrobe[4] VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__clkbuf_2
Xfanout724 net725 VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__dlymetal6s2s_1
X_1669_ _0986_ _0610_ _0609_ Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q VGND VGND
+ VPWR VPWR _0611_ sky130_fd_sc_hd__o211a_1
X_2787_ net31 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_1
X_1738_ _0667_ _0671_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JS2BEG0 sky130_fd_sc_hd__or2_1
Xfanout702 net704 VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__clkbuf_2
Xhold299 Inst_RegFile_32x4.mem\[11\]\[2\] VGND VGND VPWR VPWR net874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 Inst_RegFile_32x4.mem\[1\]\[0\] VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 Inst_RegFile_32x4.mem\[2\]\[0\] VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold277 Inst_RegFile_32x4.mem\[31\]\[0\] VGND VGND VPWR VPWR net852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 Inst_RegFile_32x4.mem\[23\]\[2\] VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 Inst_RegFile_32x4.mem\[4\]\[0\] VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout779 net4 VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout757 net42 VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__clkbuf_4
Xfanout768 net769 VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__clkbuf_4
Xfanout735 net736 VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__buf_2
Xfanout746 net51 VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__clkbuf_4
XANTENNA_106 WW4END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 net687 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_139 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2710_ clknet_4_8_0_UserCLK_regs _0112_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2572_ net751 net718 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2641_ net744 net738 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1454_ _0400_ _0401_ _0954_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__mux2_2
Xoutput305 net305 VGND VGND VPWR VPWR S2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput338 net338 VGND VGND VPWR VPWR SS4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput349 net349 VGND VGND VPWR VPWR W1BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput327 net327 VGND VGND VPWR VPWR S4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput316 net316 VGND VGND VPWR VPWR S4BEG[12] sky130_fd_sc_hd__buf_2
X_1523_ _0477_ _0476_ net682 VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__mux2_1
XFILLER_67_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1385_ net74 net16 net102 net130 Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q
+ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__mux4_2
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2006_ net611 net866 _0860_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__mux2_1
X_2908_ S4END[14] VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2839_ net72 VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__clkbuf_2
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1170_ _0971_ _0950_ _0947_ _0145_ Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q
+ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_50_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2624_ net39 net726 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_39 FrameStrobe[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_28 net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 EE4END[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1437_ net60 net68 net2 net10 Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q
+ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__mux4_1
X_2486_ net773 net707 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput168 net168 VGND VGND VPWR VPWR E6BEG[5] sky130_fd_sc_hd__buf_2
Xoutput179 net179 VGND VGND VPWR VPWR EE4BEG[15] sky130_fd_sc_hd__clkbuf_4
X_2555_ net33 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput157 net157 VGND VGND VPWR VPWR E2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput146 net146 VGND VGND VPWR VPWR E2BEG[1] sky130_fd_sc_hd__buf_6
X_1506_ Inst_RegFile_32x4.mem\[22\]\[1\] Inst_RegFile_32x4.mem\[23\]\[1\] net606 VGND
+ VGND VPWR VPWR _0461_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1299_ Inst_RegFile_32x4.mem\[30\]\[1\] Inst_RegFile_32x4.mem\[31\]\[1\] net624 VGND
+ VGND VPWR VPWR _0268_ sky130_fd_sc_hd__mux2_1
X_1368_ Inst_RegFile_32x4.mem\[30\]\[3\] Inst_RegFile_32x4.mem\[31\]\[3\] net624 VGND
+ VGND VPWR VPWR _0333_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput48 FrameData[31] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_2
Xinput37 FrameData[20] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
Xinput26 EE4END[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_6
Xinput15 E2MID[2] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
Xinput59 N1END[0] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_4
X_2271_ net761 net729 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2340_ net756 net734 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1084_ Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__inv_1
XFILLER_37_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1153_ Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q net109 Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q
+ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__o21a_1
X_1222_ Inst_RegFile_32x4.mem\[30\]\[0\] Inst_RegFile_32x4.mem\[31\]\[0\] net624 VGND
+ VGND VPWR VPWR _0195_ sky130_fd_sc_hd__mux2_1
XFILLER_60_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1986_ net420 _0718_ Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q VGND VGND VPWR VPWR
+ _0870_ sky130_fd_sc_hd__mux2_1
XFILLER_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2607_ net746 net722 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2538_ net776 net714 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2469_ net755 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1840_ net653 net422 Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q VGND VGND VPWR VPWR
+ _0758_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1771_ net85 net780 net113 net689 Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q
+ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__mux4_1
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2323_ net55 net737 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2254_ net747 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1136_ _1021_ _1023_ _1026_ _0967_ _0965_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_48_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1205_ net85 net6 net92 net120 Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q
+ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__mux4_2
X_1067_ Inst_RegFile_32x4.mem\[22\]\[0\] VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__inv_1
X_2185_ clknet_4_1_0_UserCLK_regs _0009_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[26\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclone18 net678 VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__clkbuf_1
Xclone29 net647 VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__clkbuf_1
X_1969_ _0719_ _0836_ _1017_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__mux2_1
XFILLER_21_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2941_ Inst_RegFile_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__buf_2
X_1823_ _0744_ _0743_ Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.SS4BEG2 sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_45_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2872_ NN4END[14] VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__clkbuf_2
X_1685_ _0990_ _0624_ Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q VGND VGND VPWR VPWR
+ _0625_ sky130_fd_sc_hd__o21a_1
X_1754_ _0680_ _0682_ _0685_ _1006_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E2BEG0
+ sky130_fd_sc_hd__a22o_1
X_2306_ net41 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2237_ clknet_4_15_0_UserCLK_regs _0061_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[18\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1119_ Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__inv_1
X_2099_ net612 net871 _0916_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2168_ net616 net870 _0931_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1470_ net398 net678 net665 net638 Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q
+ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__mux4_2
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2022_ net599 net868 _0894_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__mux2_1
X_2924_ SS4END[14] VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkbuf_2
X_2786_ net30 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_1
X_1806_ net635 _0707_ _0708_ _0159_ Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q
+ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_13_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2855_ N4END[13] VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__clkbuf_2
Xfanout725 net726 VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__clkbuf_2
X_1668_ net680 net636 net668 net640 Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q
+ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout758 net41 VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__clkbuf_4
Xfanout714 net717 VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__buf_2
Xfanout736 net737 VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__clkbuf_2
X_1737_ Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q _0670_ VGND VGND VPWR VPWR _0671_
+ sky130_fd_sc_hd__and2b_1
Xfanout703 net704 VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout747 net50 VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__clkbuf_4
Xhold267 Inst_RegFile_32x4.mem\[19\]\[2\] VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold278 Inst_RegFile_32x4.mem\[9\]\[1\] VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__dlygate4sd3_1
Xhold289 Inst_RegFile_32x4.mem\[9\]\[2\] VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 Inst_RegFile_32x4.mem\[15\]\[0\] VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__dlygate4sd3_1
X_1599_ Inst_RegFile_32x4.mem\[28\]\[2\] Inst_RegFile_32x4.mem\[29\]\[2\] net603 VGND
+ VGND VPWR VPWR _0550_ sky130_fd_sc_hd__mux2_1
Xhold245 Inst_RegFile_32x4.mem\[4\]\[3\] VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_129 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_118 net689 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout769 FrameData[15] VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__buf_2
XFILLER_26_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_107 WW4END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2640_ net745 net738 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_10_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2571_ net763 net718 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1453_ net72 net14 net100 net128 Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q
+ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__mux4_1
Xoutput306 net306 VGND VGND VPWR VPWR S2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput328 net328 VGND VGND VPWR VPWR S4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput339 net339 VGND VGND VPWR VPWR SS4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput317 net317 VGND VGND VPWR VPWR S4BEG[13] sky130_fd_sc_hd__buf_2
X_1522_ Inst_RegFile_32x4.mem\[4\]\[1\] Inst_RegFile_32x4.mem\[5\]\[1\] net609 VGND
+ VGND VPWR VPWR _0477_ sky130_fd_sc_hd__mux2_1
XFILLER_67_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1384_ _0222_ _0223_ _0224_ _0940_ Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q VGND
+ VGND VPWR VPWR _0347_ sky130_fd_sc_hd__a221o_1
X_2005_ Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q _0880_ _0881_ _0886_ VGND VGND
+ VPWR VPWR _0887_ sky130_fd_sc_hd__a31o_1
X_2907_ S4END[13] VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkbuf_2
XFILLER_63_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2769_ EE4END[15] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
X_2838_ net71 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_2
Xfanout599 net602 VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__clkbuf_2
XFILLER_73_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_29 net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_18 EE4END[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2623_ net761 net726 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2554_ net32 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1436_ Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q _0395_ Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q
+ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__o21a_1
Xoutput169 net169 VGND VGND VPWR VPWR E6BEG[6] sky130_fd_sc_hd__buf_2
X_2485_ net774 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput158 net158 VGND VGND VPWR VPWR E2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput147 net147 VGND VGND VPWR VPWR E2BEG[2] sky130_fd_sc_hd__buf_6
X_1367_ Inst_RegFile_32x4.mem\[28\]\[3\] Inst_RegFile_32x4.mem\[29\]\[3\] net624 VGND
+ VGND VPWR VPWR _0332_ sky130_fd_sc_hd__mux2_1
X_1505_ _0389_ _0459_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_66_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1298_ Inst_RegFile_32x4.mem\[28\]\[1\] Inst_RegFile_32x4.mem\[29\]\[1\] net624 VGND
+ VGND VPWR VPWR _0267_ sky130_fd_sc_hd__mux2_1
XFILLER_11_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput38 FrameData[21] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
Xinput49 FrameData[3] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_2
Xinput27 FrameData[0] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_2
Xinput16 E2MID[3] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
XFILLER_6_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2270_ net762 net729 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1221_ Inst_RegFile_32x4.mem\[28\]\[0\] Inst_RegFile_32x4.mem\[29\]\[0\] net624 VGND
+ VGND VPWR VPWR _0194_ sky130_fd_sc_hd__mux2_1
XFILLER_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1152_ _1038_ _1036_ _0128_ _0958_ _0969_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__a221o_2
X_1083_ Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__inv_1
XFILLER_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1985_ net599 net814 _0860_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__mux2_1
X_2537_ net48 net711 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2606_ net747 net722 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1419_ net60 net68 net2 net10 Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q
+ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__mux4_1
X_2468_ net756 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2399_ net761 net697 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_36_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1770_ _0694_ _0696_ _0699_ _1010_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JN2BEG0
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2322_ net54 net737 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1204_ _0980_ _0175_ _0177_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__o21ai_4
X_2253_ net748 net56 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2184_ clknet_4_1_0_UserCLK_regs _0008_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[26\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1135_ _1021_ _1023_ _1026_ _0967_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E2BEG5
+ sky130_fd_sc_hd__a22o_1
X_1066_ Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1899_ net81 net126 net7 Inst_RegFile_switch_matrix.E2BEG2 Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_31_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1968_ _0838_ _0852_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__nand2_8
Xclone19 net684 VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_3_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1822_ net59 net1 net115 net421 Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q
+ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__mux4_2
X_1753_ _0683_ _0684_ _1005_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__mux2_1
XFILLER_30_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2871_ NN4END[13] VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__clkbuf_2
X_1684_ net676 net635 net666 net639 Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q
+ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__mux4_1
XFILLER_65_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2305_ net759 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2236_ clknet_4_13_0_UserCLK_regs _0060_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[18\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2167_ net600 net893 _0931_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__mux2_1
XFILLER_53_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1118_ Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__inv_1
X_1049_ Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__inv_2
XFILLER_21_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2098_ net621 net908 _0916_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_0_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2021_ _0831_ _0893_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__nand2_2
X_2923_ SS4END[13] VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__clkbuf_2
X_2785_ net774 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__buf_2
X_1805_ _0730_ _0729_ Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.WW4BEG2 sky130_fd_sc_hd__mux2_1
X_1736_ _0668_ _0669_ Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q VGND VGND VPWR VPWR
+ _0670_ sky130_fd_sc_hd__mux2_1
XFILLER_7_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2854_ N4END[12] VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__clkbuf_2
Xfanout726 FrameStrobe[1] VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__clkbuf_2
Xfanout737 FrameStrobe[10] VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__clkbuf_2
Xfanout759 net40 VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__buf_4
X_1667_ Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q _0608_ VGND VGND VPWR VPWR _0609_
+ sky130_fd_sc_hd__or2_1
Xfanout715 net716 VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__clkbuf_2
Xfanout748 net49 VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__buf_4
Xfanout704 net705 VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold268 Inst_RegFile_32x4.mem\[30\]\[0\] VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 Inst_RegFile_32x4.mem\[30\]\[1\] VGND VGND VPWR VPWR net832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 Inst_RegFile_32x4.mem\[6\]\[3\] VGND VGND VPWR VPWR net854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 Inst_RegFile_32x4.mem\[30\]\[3\] VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__dlygate4sd3_1
X_1598_ Inst_RegFile_32x4.mem\[30\]\[2\] Inst_RegFile_32x4.mem\[31\]\[2\] net603 VGND
+ VGND VPWR VPWR _0549_ sky130_fd_sc_hd__mux2_1
XANTENNA_119 net689 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2219_ clknet_4_10_0_UserCLK_regs _0043_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[22\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_108 WW4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2570_ net776 net718 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput307 net307 VGND VGND VPWR VPWR S2BEGb[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_10_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1452_ net71 net13 net127 Inst_RegFile_switch_matrix.JW2BEG6 Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__mux4_2
X_1383_ _0345_ Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q _0346_ VGND VGND VPWR VPWR
+ AD3 sky130_fd_sc_hd__o21ai_4
Xoutput318 net318 VGND VGND VPWR VPWR S4BEG[14] sky130_fd_sc_hd__buf_6
Xoutput329 net329 VGND VGND VPWR VPWR SS4BEG[0] sky130_fd_sc_hd__buf_2
X_1521_ Inst_RegFile_32x4.mem\[6\]\[1\] Inst_RegFile_32x4.mem\[7\]\[1\] net607 VGND
+ VGND VPWR VPWR _0476_ sky130_fd_sc_hd__mux2_1
XFILLER_67_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2004_ Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q _0882_ _0885_ VGND VGND VPWR VPWR
+ _0886_ sky130_fd_sc_hd__o21a_1
X_2906_ S4END[12] VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__buf_2
XFILLER_23_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2837_ Inst_RegFile_switch_matrix.JN2BEG7 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__clkbuf_1
X_1719_ net92 net108 net111 net120 Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q
+ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__mux4_1
X_2768_ EE4END[14] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_1
X_2699_ clknet_4_11_0_UserCLK_regs _0101_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_19 EE4END[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2622_ net762 net726 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2553_ net768 net714 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput159 net159 VGND VGND VPWR VPWR E2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput148 net148 VGND VGND VPWR VPWR E2BEG[3] sky130_fd_sc_hd__buf_6
X_1504_ _0457_ _0458_ net683 VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__mux2_1
X_1435_ net140 net670 net657 net655 Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q
+ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__mux4_1
X_2484_ net775 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1366_ net648 _0330_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_66_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1297_ net663 _0263_ net648 VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__o21a_1
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput39 FrameData[22] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
Xinput28 FrameData[10] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_4
Xinput17 E2MID[4] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1151_ net414 _1038_ _0128_ _0958_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E2BEG3
+ sky130_fd_sc_hd__a22o_4
X_1220_ _0192_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_63_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1082_ Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__inv_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1984_ _0865_ _0867_ _0868_ _1014_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_33_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2536_ net47 net711 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2605_ net748 net725 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2467_ net757 net704 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1418_ net88 net96 net114 net116 Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q
+ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__mux4_1
X_2398_ net762 net697 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1349_ _0312_ _0313_ net674 VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__mux2_1
XFILLER_51_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2321_ net53 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1134_ _1024_ _1025_ _0966_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__mux2_1
X_1203_ Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q _0176_ Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q
+ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__o21a_1
X_2252_ net751 net56 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2183_ clknet_4_0_0_UserCLK_regs _0007_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[25\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1065_ Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_48_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1967_ Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q _0849_ _0851_ _0843_ _0844_ VGND
+ VGND VPWR VPWR _0852_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_31_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1898_ net72 net14 net100 net128 Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q
+ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__mux4_2
X_2519_ net772 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_71_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone2 _0178_ Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q _0180_ _0191_ VGND VGND
+ VPWR VPWR net395 sky130_fd_sc_hd__a31o_4
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2870_ NN4END[12] VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__clkbuf_2
X_1821_ net641 _1033_ net685 _0213_ Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q
+ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__mux4_1
X_1752_ net62 net64 net80 net83 Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q
+ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__mux4_1
X_1683_ Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q _0622_ VGND VGND VPWR VPWR _0623_
+ sky130_fd_sc_hd__or2_1
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2304_ net760 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_65_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1117_ Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__inv_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2235_ clknet_4_15_0_UserCLK_regs _0059_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[16\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2166_ _0893_ _0902_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__nand2_4
X_2097_ net617 net873 _0916_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1048_ Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__inv_2
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2020_ _0857_ _0888_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__nor2_8
X_2922_ SS4END[12] VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkbuf_2
X_2853_ N4END[11] VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkbuf_2
X_1666_ net686 net672 net659 net646 Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q
+ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__mux4_1
X_1804_ net59 net87 net115 net644 Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q
+ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__mux4_1
X_2784_ net28 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__buf_1
X_1735_ net92 net120 net108 net137 Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q
+ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__mux4_1
Xhold269 Inst_RegFile_32x4.mem\[17\]\[0\] VGND VGND VPWR VPWR net844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 Inst_RegFile_32x4.mem\[8\]\[0\] VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 Inst_RegFile_32x4.mem\[24\]\[1\] VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 Inst_RegFile_32x4.mem\[6\]\[0\] VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_13_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout749 net48 VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__clkbuf_4
Xfanout727 net729 VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__buf_2
Xfanout716 net717 VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__buf_2
Xfanout738 net739 VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__clkbuf_2
Xfanout705 FrameStrobe[6] VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1597_ _0546_ _0547_ net681 VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__mux2_1
XFILLER_66_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_109 _0129_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2218_ clknet_4_13_0_UserCLK_regs _0042_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[22\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2149_ net622 net915 _0927_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__mux2_2
XFILLER_49_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1520_ _0474_ _0473_ net682 VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__mux2_1
Xoutput319 net319 VGND VGND VPWR VPWR S4BEG[15] sky130_fd_sc_hd__buf_4
Xoutput308 net308 VGND VGND VPWR VPWR S2BEGb[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_10_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1451_ _0403_ _0405_ _0407_ _0409_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JW2BEG6
+ sky130_fd_sc_hd__o2bb2a_4
X_1382_ Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q Inst_RegFile_32x4.AD_reg\[3\] VGND
+ VGND VPWR VPWR _0346_ sky130_fd_sc_hd__nand2_1
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2003_ Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q _0884_ Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q
+ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__a21oi_1
X_2905_ S4END[11] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__buf_2
X_2836_ Inst_RegFile_switch_matrix.JN2BEG6 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__buf_4
XFILLER_50_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1649_ Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q _0592_ VGND VGND VPWR VPWR _0593_
+ sky130_fd_sc_hd__nor2_1
X_1718_ net62 net64 net6 net777 Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q
+ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__mux4_1
X_2767_ EE4END[13] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_1
X_2698_ clknet_4_14_0_UserCLK_regs _0100_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2621_ net764 net724 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2552_ net770 net714 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2483_ net55 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_34_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput149 net149 VGND VGND VPWR VPWR E2BEG[4] sky130_fd_sc_hd__buf_6
X_1503_ Inst_RegFile_32x4.mem\[18\]\[1\] Inst_RegFile_32x4.mem\[19\]\[1\] net609 VGND
+ VGND VPWR VPWR _0458_ sky130_fd_sc_hd__mux2_1
X_1434_ _0955_ _0393_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__or2_4
XFILLER_55_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1365_ _0328_ _0329_ net674 VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__mux2_4
X_1296_ net396 _0264_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_66_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2819_ FrameStrobe[13] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_52_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 E2MID[5] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_70_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput29 FrameData[11] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_4
X_1150_ _1039_ _1040_ Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q VGND VGND VPWR VPWR
+ _0128_ sky130_fd_sc_hd__mux2_1
X_1081_ Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2604_ net751 net725 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1983_ _0767_ _0803_ Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q VGND VGND VPWR VPWR
+ _0868_ sky130_fd_sc_hd__mux2_1
X_2535_ net752 net711 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1417_ _0377_ _0951_ Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q VGND VGND VPWR VPWR
+ _0378_ sky130_fd_sc_hd__o21a_1
X_2466_ net758 net704 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2397_ net35 net696 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_36_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1348_ Inst_RegFile_32x4.mem\[8\]\[3\] Inst_RegFile_32x4.mem\[9\]\[3\] net629 VGND
+ VGND VPWR VPWR _0313_ sky130_fd_sc_hd__mux2_1
X_1279_ Inst_RegFile_32x4.mem\[8\]\[1\] Inst_RegFile_32x4.mem\[9\]\[1\] net629 VGND
+ VGND VPWR VPWR _0248_ sky130_fd_sc_hd__mux2_1
XFILLER_22_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_5_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2320_ net52 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2251_ clknet_4_11_0_UserCLK_regs _0075_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[21\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1064_ Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__inv_1
X_1133_ net61 net69 net780 net11 Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q
+ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__mux4_1
X_1202_ net26 net107 Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q VGND VGND VPWR VPWR
+ _0176_ sky130_fd_sc_hd__mux2_1
X_2182_ clknet_4_5_0_UserCLK_regs _0006_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[25\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_48_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1966_ _1015_ _0850_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_31_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1897_ net635 _0582_ Inst_RegFile_switch_matrix.JS2BEG0 _0158_ Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.W1BEG1
+ sky130_fd_sc_hd__mux4_1
XFILLER_68_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2518_ net773 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2449_ net744 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_56_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone3 _0135_ VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1820_ _0737_ _0742_ Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.SS4BEG3 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1751_ net6 net92 net777 net120 Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q
+ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__mux4_1
X_1682_ net687 net671 net423 net645 Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q
+ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__mux4_1
X_2303_ net38 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2234_ clknet_4_15_0_UserCLK_regs _0058_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[16\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1116_ Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__inv_1
XFILLER_65_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1047_ Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__inv_2
X_2096_ net600 net830 _0916_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2165_ net614 net922 _0930_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__mux2_2
X_1949_ _0401_ Inst_RegFile_switch_matrix.JN2BEG0 Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q
+ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__mux2_1
XFILLER_21_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2921_ SS4END[11] VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__clkbuf_2
X_2783_ net742 VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__buf_1
X_1803_ _0728_ _0727_ Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q VGND VGND VPWR VPWR
+ _0729_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2852_ N4END[10] VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__clkbuf_2
X_1665_ _0603_ _0604_ _0607_ _0985_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E2BEG2
+ sky130_fd_sc_hd__a22o_1
Xfanout706 FrameStrobe[5] VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__buf_2
X_1734_ net64 net6 net779 net777 Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q
+ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__mux4_1
Xhold237 Inst_RegFile_32x4.mem\[0\]\[0\] VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__dlygate4sd3_1
X_1596_ Inst_RegFile_32x4.mem\[26\]\[2\] Inst_RegFile_32x4.mem\[27\]\[2\] net604 VGND
+ VGND VPWR VPWR _0547_ sky130_fd_sc_hd__mux2_1
Xhold259 Inst_RegFile_32x4.mem\[27\]\[2\] VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 Inst_RegFile_32x4.mem\[12\]\[2\] VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_439 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout717 FrameStrobe[3] VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout728 net729 VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout739 FrameStrobe[0] VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2217_ clknet_4_10_0_UserCLK_regs _0041_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[22\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2148_ net616 net925 _0927_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__mux2_2
X_2079_ _0887_ net895 _0912_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1450_ Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q _0408_ Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q
+ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__a21o_1
XFILLER_4_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput309 net309 VGND VGND VPWR VPWR S2BEGb[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_10_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1381_ _0345_ VGND VGND VPWR VPWR Inst_RegFile_32x4.AD_comb\[3\] sky130_fd_sc_hd__inv_1
XFILLER_35_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2002_ _0883_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_18_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2904_ S4END[10] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__buf_2
XFILLER_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2766_ EE4END[12] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_1
X_1648_ net686 net669 net656 net644 Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q
+ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__mux4_1
X_1717_ _0998_ _0652_ Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q VGND VGND VPWR VPWR
+ _0653_ sky130_fd_sc_hd__o21a_1
X_1579_ Inst_RegFile_32x4.mem\[10\]\[2\] Inst_RegFile_32x4.mem\[11\]\[2\] net608 VGND
+ VGND VPWR VPWR _0530_ sky130_fd_sc_hd__mux2_1
X_2697_ clknet_4_14_0_UserCLK_regs _0099_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_52_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2620_ net765 net724 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_32_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1433_ AD3 net634 net665 net638 Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q
+ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__mux4_1
X_2551_ net772 net717 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2482_ net54 net709 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1502_ Inst_RegFile_32x4.mem\[16\]\[1\] Inst_RegFile_32x4.mem\[17\]\[1\] net610 VGND
+ VGND VPWR VPWR _0457_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1295_ Inst_RegFile_32x4.mem\[26\]\[1\] Inst_RegFile_32x4.mem\[27\]\[1\] net625 VGND
+ VGND VPWR VPWR _0264_ sky130_fd_sc_hd__mux2_1
X_1364_ Inst_RegFile_32x4.mem\[24\]\[3\] Inst_RegFile_32x4.mem\[25\]\[3\] net625 VGND
+ VGND VPWR VPWR _0329_ sky130_fd_sc_hd__mux2_1
XFILLER_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2749_ E6END[5] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_1
X_2818_ net56 VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_21_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_7_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_52_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput19 E2MID[6] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
XFILLER_35_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1080_ Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__inv_1
XFILLER_18_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1982_ Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q _0866_ Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q
+ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__a21oi_1
XFILLER_33_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2534_ net753 net711 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2603_ net763 net722 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_21_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1416_ net647 net637 net667 net641 Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q
+ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__mux4_2
X_2396_ net34 net696 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2465_ net759 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1347_ Inst_RegFile_32x4.mem\[10\]\[3\] Inst_RegFile_32x4.mem\[11\]\[3\] net626 VGND
+ VGND VPWR VPWR _0312_ sky130_fd_sc_hd__mux2_1
X_1278_ Inst_RegFile_32x4.mem\[10\]\[1\] Inst_RegFile_32x4.mem\[11\]\[1\] net629 VGND
+ VGND VPWR VPWR _0247_ sky130_fd_sc_hd__mux2_1
XFILLER_24_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1201_ net138 Inst_RegFile_switch_matrix.JW2BEG3 Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q
+ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__mux2_4
X_2250_ clknet_4_9_0_UserCLK_regs _0074_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[21\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1132_ net25 net87 net89 net97 Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q
+ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__mux4_1
X_1063_ Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__inv_1
XFILLER_18_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2181_ clknet_4_0_0_UserCLK_regs _0005_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[25\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1965_ net78 net20 net106 net134 Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q
+ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_31_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2517_ net774 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1896_ net409 net685 Inst_RegFile_switch_matrix.JS2BEG1 net394 Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.W1BEG2
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_39_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2379_ net36 net697 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2448_ net745 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_33_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1750_ _1005_ _0681_ Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q VGND VGND VPWR VPWR
+ _0682_ sky130_fd_sc_hd__o21a_1
X_1681_ _0616_ _0618_ _0621_ _0989_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JW2BEG1
+ sky130_fd_sc_hd__a22o_1
X_2302_ net37 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2233_ clknet_4_15_0_UserCLK_regs _0057_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[16\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2164_ net621 net918 _0930_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__mux2_2
X_1115_ Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__inv_1
XFILLER_65_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1046_ Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_0_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2095_ _0898_ _0889_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__nand2_4
X_1879_ net65 net93 net7 net139 Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q
+ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__mux4_2
X_1948_ Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q Inst_RegFile_switch_matrix.JW2BEG0
+ Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__a21bo_1
XFILLER_21_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2920_ SS4END[10] VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__clkbuf_2
XFILLER_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2782_ net743 VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_2
X_1802_ net638 _1033_ Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q VGND VGND VPWR VPWR
+ _0728_ sky130_fd_sc_hd__mux2_1
XFILLER_43_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1733_ _1002_ _0664_ _0666_ Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q VGND VGND VPWR
+ VPWR _0667_ sky130_fd_sc_hd__o211a_1
X_2851_ N4END[9] VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__clkbuf_2
X_1664_ _0605_ _0606_ _0984_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__mux2_1
Xfanout707 FrameStrobe[5] VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout718 net719 VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__clkbuf_2
Xfanout729 net56 VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold238 Inst_RegFile_32x4.mem\[26\]\[2\] VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 Inst_RegFile_32x4.mem\[6\]\[2\] VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__dlygate4sd3_1
X_1595_ Inst_RegFile_32x4.mem\[24\]\[2\] Inst_RegFile_32x4.mem\[25\]\[2\] net603 VGND
+ VGND VPWR VPWR _0546_ sky130_fd_sc_hd__mux2_1
XFILLER_66_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2216_ clknet_4_11_0_UserCLK_regs _0040_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[22\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2147_ net601 net933 _0927_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__mux2_2
XFILLER_53_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2078_ net620 net884 _0912_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__mux2_2
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1380_ _0228_ _0319_ _0327_ _0344_ _0343_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__o32a_4
XFILLER_48_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2001_ net72 net14 net100 net128 Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q
+ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__mux4_1
X_2903_ S4END[9] VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_18_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2834_ Inst_RegFile_switch_matrix.JN2BEG4 VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__buf_1
X_1716_ net678 net635 net666 net639 Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q
+ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__mux4_1
X_2765_ EE4END[11] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_1
X_2696_ clknet_4_14_0_UserCLK_regs _0098_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[5\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1647_ _0586_ _0588_ _0591_ _0982_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JW2BEG2
+ sky130_fd_sc_hd__a22o_1
X_1578_ Inst_RegFile_32x4.mem\[8\]\[2\] Inst_RegFile_32x4.mem\[9\]\[2\] net608 VGND
+ VGND VPWR VPWR _0529_ sky130_fd_sc_hd__mux2_1
XFILLER_54_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_15_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_15_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_52_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2550_ net773 net717 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2481_ net744 net706 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1501_ Inst_RegFile_32x4.BD_comb\[0\] Inst_RegFile_32x4.BD_reg\[0\] Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q
+ VGND VGND VPWR VPWR BD0 sky130_fd_sc_hd__mux2_4
X_1363_ Inst_RegFile_32x4.mem\[26\]\[3\] Inst_RegFile_32x4.mem\[27\]\[3\] net625 VGND
+ VGND VPWR VPWR _0328_ sky130_fd_sc_hd__mux2_1
X_1432_ _0389_ _0391_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_66_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1294_ Inst_RegFile_32x4.mem\[24\]\[1\] Inst_RegFile_32x4.mem\[25\]\[1\] net624 VGND
+ VGND VPWR VPWR _0263_ sky130_fd_sc_hd__mux2_1
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2817_ net730 VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__buf_1
X_2748_ E6END[4] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_1
X_2679_ clknet_4_0_0_UserCLK_regs _0081_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[29\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1981_ net78 net20 net106 net134 Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q
+ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__mux4_1
X_2533_ net755 net712 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2602_ net776 net722 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1415_ Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q _0375_ VGND VGND VPWR VPWR _0376_
+ sky130_fd_sc_hd__or2_1
X_2395_ net766 net695 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2464_ net760 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1346_ Inst_RegFile_32x4.AD_comb\[2\] Inst_RegFile_32x4.AD_reg\[2\] Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q
+ VGND VGND VPWR VPWR AD2 sky130_fd_sc_hd__mux2_4
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1277_ Inst_RegFile_32x4.AD_comb\[0\] Inst_RegFile_32x4.AD_reg\[0\] Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q
+ VGND VGND VPWR VPWR AD0 sky130_fd_sc_hd__mux2_4
XFILLER_51_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1200_ _0171_ _0169_ _0174_ _0979_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JW2BEG3
+ sky130_fd_sc_hd__a22o_4
X_2180_ clknet_4_0_0_UserCLK_regs _0004_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[25\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1131_ Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q _1022_ Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q
+ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__o21a_1
X_1062_ Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__inv_2
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1895_ net671 _0437_ Inst_RegFile_switch_matrix.JS2BEG2 _0803_ Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.W1BEG3
+ sky130_fd_sc_hd__mux4_1
X_1964_ _0845_ _0846_ _0848_ Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q _1015_ VGND
+ VGND VPWR VPWR _0849_ sky130_fd_sc_hd__o221a_1
XFILLER_33_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2516_ net775 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2447_ net51 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2378_ net776 net58 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1329_ Inst_RegFile_32x4.mem\[24\]\[2\] Inst_RegFile_32x4.mem\[25\]\[2\] net625 VGND
+ VGND VPWR VPWR _0296_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_49_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput290 net290 VGND VGND VPWR VPWR NN4BEG[7] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_58_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2301_ net764 net730 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1680_ _0619_ _0620_ Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q VGND VGND VPWR VPWR
+ _0621_ sky130_fd_sc_hd__mux2_1
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1114_ Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__inv_1
X_2232_ clknet_4_12_0_UserCLK_regs _0056_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[16\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2163_ net616 net899 _0930_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__mux2_2
XFILLER_46_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1045_ Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__inv_1
X_2094_ net613 net910 _0915_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__mux2_4
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1878_ _0790_ _0789_ Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.NN4BEG3 sky130_fd_sc_hd__mux2_4
X_1947_ _0667_ _0671_ Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q VGND VGND VPWR VPWR
+ _0832_ sky130_fd_sc_hd__o21ba_1
XFILLER_56_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2850_ N4END[8] VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkbuf_2
X_1801_ net685 _0726_ Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q VGND VGND VPWR VPWR
+ _0727_ sky130_fd_sc_hd__mux2_1
X_1663_ net60 net66 net82 net8 Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q
+ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__mux4_1
X_1732_ Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q _0665_ VGND VGND VPWR VPWR _0666_
+ sky130_fd_sc_hd__or2_1
X_2781_ net744 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__buf_4
XFILLER_7_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout719 net720 VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout708 FrameStrobe[5] VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__buf_2
Xhold239 Inst_RegFile_32x4.mem\[24\]\[0\] VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1594_ _0389_ _0542_ _0544_ net619 VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__o31a_1
XFILLER_66_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2215_ clknet_4_15_0_UserCLK_regs _0039_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[17\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2146_ _0893_ _0923_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__nand2_4
X_2077_ net615 net904 _0912_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__mux2_2
XFILLER_61_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2000_ net71 net13 net99 Inst_RegFile_switch_matrix.JW2BEG3 Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_18_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2902_ S4END[8] VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__buf_2
X_2833_ Inst_RegFile_switch_matrix.JN2BEG3 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__buf_1
XFILLER_43_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1646_ _0589_ _0590_ Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q VGND VGND VPWR VPWR
+ _0591_ sky130_fd_sc_hd__mux2_1
X_1715_ Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q _0650_ VGND VGND VPWR VPWR _0651_
+ sky130_fd_sc_hd__or2_1
X_2764_ EE4END[10] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2695_ clknet_4_14_0_UserCLK_regs _0097_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1577_ net642 _0527_ net619 VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__a21bo_1
XFILLER_66_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer21 _1036_ VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__buf_6
XFILLER_39_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2129_ net612 net921 _0922_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__mux2_2
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2480_ net745 net706 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1500_ _0420_ _0440_ _0456_ _0448_ VGND VGND VPWR VPWR Inst_RegFile_32x4.BD_comb\[0\]
+ sky130_fd_sc_hd__a22o_1
X_1431_ _0364_ _0390_ net682 VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__mux2_1
X_1293_ _0192_ _0253_ _0229_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__o21a_1
X_1362_ net648 _0322_ _0326_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_66_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2816_ net737 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__buf_1
X_1629_ _0575_ _0963_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__or2_4
X_2747_ E6END[3] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_1
X_2678_ clknet_4_3_0_UserCLK_regs _0080_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[29\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1980_ Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q _0862_ _0864_ Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q
+ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__a211o_1
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2532_ net756 net712 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2601_ net48 net720 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer1 _0400_ VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__buf_6
X_2463_ net761 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_9_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1414_ net118 net673 net660 net654 Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q
+ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__mux4_1
X_2394_ net767 net695 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1276_ _0246_ _0238_ _0229_ _0230_ _0205_ VGND VGND VPWR VPWR Inst_RegFile_32x4.AD_comb\[0\]
+ sky130_fd_sc_hd__a32o_1
X_1345_ _0229_ _0286_ _0294_ _0310_ _0311_ VGND VGND VPWR VPWR Inst_RegFile_32x4.AD_comb\[2\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_34_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_3_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_3_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
X_1130_ net689 net672 net660 net653 Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q
+ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_48_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1061_ Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__inv_1
X_1894_ net86 net110 net137 Inst_RegFile_switch_matrix.JN2BEG1 Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__mux4_2
X_1963_ _0847_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__inv_1
XFILLER_21_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2515_ net742 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2446_ net50 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2377_ net749 net690 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_39_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1328_ Inst_RegFile_32x4.mem\[26\]\[2\] Inst_RegFile_32x4.mem\[27\]\[2\] net625 VGND
+ VGND VPWR VPWR _0295_ sky130_fd_sc_hd__mux2_1
X_1259_ _0167_ _0197_ _0229_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__a21oi_1
XFILLER_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput280 net280 VGND VGND VPWR VPWR NN4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput291 net291 VGND VGND VPWR VPWR NN4BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_58_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2300_ net34 net730 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2231_ clknet_4_6_0_UserCLK_regs _0055_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[15\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1044_ Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__inv_2
X_1113_ Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__inv_2
X_2093_ net622 net894 _0915_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__mux2_4
X_2162_ net600 net880 _0930_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__mux2_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1877_ net60 net2 net116 net672 Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q
+ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__mux4_1
X_1946_ _0822_ _0829_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__nor2_2
X_2429_ net35 net701 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_29_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1800_ net67 net9 net113 net123 Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q
+ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__mux4_2
XFILLER_50_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1662_ net777 net94 net113 net122 Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q
+ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__mux4_1
X_2780_ net52 VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_2
X_1731_ net686 net652 net658 net645 Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q
+ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_13_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout709 FrameStrobe[5] VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__clkbuf_2
X_2214_ clknet_4_15_0_UserCLK_regs _0038_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[17\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1593_ net682 _0543_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__nor2_1
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2145_ net612 net854 _0926_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__mux2_1
X_2076_ net599 net891 _0912_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__mux2_2
X_2978_ Inst_RegFile_switch_matrix.WW4BEG3 VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__buf_8
X_1929_ Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q _0213_ VGND VGND VPWR VPWR _0814_
+ sky130_fd_sc_hd__nor2_1
XFILLER_39_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2901_ S4END[7] VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__buf_4
X_2832_ Inst_RegFile_switch_matrix.JN2BEG2 VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2763_ EE4END[9] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1645_ net777 net94 net110 net122 Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q
+ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__mux4_1
X_1714_ net686 net652 net658 net645 Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q
+ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__mux4_1
X_1576_ _0526_ _0525_ net683 VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__mux2_1
X_2694_ clknet_4_13_0_UserCLK_regs _0096_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2059_ _0889_ _0907_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__nand2_4
XFILLER_22_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2128_ net621 net913 _0922_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__mux2_2
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1430_ Inst_RegFile_32x4.mem\[2\]\[0\] Inst_RegFile_32x4.mem\[3\]\[0\] net606 VGND
+ VGND VPWR VPWR _0390_ sky130_fd_sc_hd__mux2_1
XFILLER_68_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1361_ net649 _0325_ _0192_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__a21bo_1
X_1292_ _0193_ _0260_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__or2_1
XFILLER_23_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2746_ E6END[2] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_1
X_2815_ net693 VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_1
X_1628_ net677 net633 net664 net638 Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q
+ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__mux4_2
X_2677_ clknet_4_15_0_UserCLK_regs _0079_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[19\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1559_ Inst_RegFile_32x4.mem\[8\]\[3\] Inst_RegFile_32x4.mem\[9\]\[3\] net608 VGND
+ VGND VPWR VPWR _0512_ sky130_fd_sc_hd__mux2_4
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_11_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_11_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_33_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2600_ net47 net720 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_71_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2531_ net757 net712 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2462_ net762 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2393_ net768 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1413_ _0946_ _0372_ _0373_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1275_ net648 _0241_ _0245_ _0244_ net395 VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__a221o_1
X_1344_ _0302_ _0298_ _0229_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__a21oi_1
XFILLER_36_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2729_ Inst_RegFile_switch_matrix.E1BEG3 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1060_ Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__inv_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1962_ net19 net105 Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q VGND VGND VPWR VPWR
+ _0847_ sky130_fd_sc_hd__mux2_1
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1893_ _0802_ _0801_ Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.NN4BEG0 sky130_fd_sc_hd__mux2_1
X_2514_ net743 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2445_ net748 net704 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2376_ net750 net693 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1258_ _0228_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__inv_2
X_1327_ net408 _0293_ _0290_ _0193_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__a211o_1
X_1189_ _0150_ _0162_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__nand2_1
XFILLER_33_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput270 net270 VGND VGND VPWR VPWR N4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput281 Inst_RegFile_switch_matrix.NN4BEG1 VGND VGND VPWR VPWR NN4BEG[13] sky130_fd_sc_hd__buf_8
Xoutput292 net292 VGND VGND VPWR VPWR NN4BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_58_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2230_ clknet_4_7_0_UserCLK_regs _0054_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[15\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1112_ Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__inv_1
XFILLER_65_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1043_ Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__inv_1
X_2092_ net617 net929 _0915_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__mux2_4
X_2161_ _0891_ _0902_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_44_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1945_ Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q _0828_ _0825_ VGND VGND VPWR VPWR
+ _0830_ sky130_fd_sc_hd__a21o_2
X_1876_ net679 _0147_ _0372_ _0788_ Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q
+ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__mux4_2
XFILLER_69_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2359_ net772 net691 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2428_ net34 net700 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1661_ Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q _0601_ Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q
+ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__o21a_1
X_1730_ net676 net635 net666 net639 Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q
+ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__mux4_1
X_1592_ Inst_RegFile_32x4.mem\[20\]\[2\] Inst_RegFile_32x4.mem\[21\]\[2\] net607 VGND
+ VGND VPWR VPWR _0543_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2213_ clknet_4_15_0_UserCLK_regs _0037_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[17\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2144_ net622 net824 _0926_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__mux2_1
XFILLER_34_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2075_ _0891_ _0904_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__nand2_4
X_2977_ Inst_RegFile_switch_matrix.WW4BEG2 VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__clkbuf_2
X_1859_ net59 Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q
+ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__o21ba_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1928_ Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q _0804_ Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q
+ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_12_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2900_ S4END[6] VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_18_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1713_ _0644_ _0646_ _0649_ _0997_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JW2BEG7
+ sky130_fd_sc_hd__a22o_1
X_2831_ Inst_RegFile_switch_matrix.JN2BEG1 VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__buf_1
XFILLER_31_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2762_ EE4END[8] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_1
X_1644_ net60 net66 net85 net8 Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q
+ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__mux4_1
X_1575_ Inst_RegFile_32x4.mem\[4\]\[2\] Inst_RegFile_32x4.mem\[5\]\[2\] net609 VGND
+ VGND VPWR VPWR _0526_ sky130_fd_sc_hd__mux2_1
X_2693_ clknet_4_14_0_UserCLK_regs _0095_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2127_ net616 net924 _0922_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_52_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2058_ _0829_ _0906_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__nor2_2
XFILLER_22_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1360_ _0323_ _0324_ net661 VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__mux2_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1291_ _0256_ _0259_ net650 VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__mux2_1
XFILLER_63_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2814_ net696 VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__buf_1
X_2745_ net20 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__buf_1
X_2676_ clknet_4_13_0_UserCLK_regs _0078_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[19\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1627_ net687 net669 net656 net651 Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q
+ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__mux4_1
X_1489_ Inst_RegFile_32x4.mem\[20\]\[0\] Inst_RegFile_32x4.mem\[21\]\[0\] net606 VGND
+ VGND VPWR VPWR _0446_ sky130_fd_sc_hd__mux2_1
X_1558_ _0507_ _0510_ net642 VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2530_ net758 net712 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_71_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2461_ net764 net704 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2392_ net770 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1412_ Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q _0226_ Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q
+ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__a21o_1
X_1343_ net648 _0305_ _0309_ _0193_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__a211o_1
X_1274_ net663 _0242_ net649 VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_62_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2659_ net757 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2728_ Inst_RegFile_switch_matrix.E1BEG2 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__buf_6
XFILLER_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout690 net692 VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1892_ net61 net780 net689 net659 Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q
+ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__mux4_1
X_1961_ net133 Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q
+ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_31_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2513_ net744 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_39_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2444_ net751 net704 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2375_ net752 net693 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1326_ _0291_ _0292_ net661 VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__mux2_1
XFILLER_49_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1257_ _0227_ _0214_ Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q VGND VGND VPWR VPWR
+ _0228_ sky130_fd_sc_hd__mux2_2
X_1188_ _0150_ _0162_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__and2_4
Xoutput282 net282 VGND VGND VPWR VPWR NN4BEG[14] sky130_fd_sc_hd__buf_4
Xoutput271 net271 VGND VGND VPWR VPWR N4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput260 net260 VGND VGND VPWR VPWR N2BEGb[7] sky130_fd_sc_hd__buf_2
XFILLER_59_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput293 net293 VGND VGND VPWR VPWR S1BEG[0] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_73_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2160_ net612 net890 _0929_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__mux2_2
X_1042_ Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__inv_1
X_1111_ Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__inv_2
XFILLER_61_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2091_ net601 net816 _0915_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1875_ net83 net93 net7 net121 Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q
+ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__mux4_2
X_1944_ Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q _0828_ _0825_ VGND VGND VPWR VPWR
+ _0829_ sky130_fd_sc_hd__a21oi_4
X_2427_ net33 net700 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2358_ net773 net691 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_56_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2289_ net53 net732 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_29_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1309_ _0164_ _0273_ _0277_ _0193_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__a211o_1
XFILLER_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1660_ _0984_ _0602_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__or2_1
XFILLER_3_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1591_ _0960_ net607 net683 _0541_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__o211a_1
XFILLER_66_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2212_ clknet_4_12_0_UserCLK_regs _0036_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[17\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2143_ net616 net818 _0926_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__mux2_1
X_2074_ net612 net892 _0911_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__mux2_1
X_1858_ net1 Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q VGND VGND VPWR VPWR _0774_
+ sky130_fd_sc_hd__nand2b_1
X_2976_ Inst_RegFile_switch_matrix.WW4BEG1 VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__buf_6
X_1927_ Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q _0811_ VGND VGND VPWR VPWR _0812_
+ sky130_fd_sc_hd__and2b_1
X_1789_ Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q _0712_ _0715_ _0716_ VGND VGND
+ VPWR VPWR _0717_ sky130_fd_sc_hd__o22a_1
XFILLER_39_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2830_ Inst_RegFile_switch_matrix.JN2BEG0 VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_26_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1712_ _0647_ _0648_ Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q VGND VGND VPWR VPWR
+ _0649_ sky130_fd_sc_hd__mux2_1
X_1643_ _0981_ _0587_ Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q VGND VGND VPWR VPWR
+ _0588_ sky130_fd_sc_hd__o21a_1
XANTENNA_1 net142 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2761_ EE4END[7] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
X_2692_ clknet_4_15_0_UserCLK_regs _0094_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1574_ Inst_RegFile_32x4.mem\[6\]\[2\] Inst_RegFile_32x4.mem\[7\]\[2\] net609 VGND
+ VGND VPWR VPWR _0525_ sky130_fd_sc_hd__mux2_1
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2057_ _0810_ _0821_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__nand2_1
X_2126_ net600 net848 _0922_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2959_ W6END[10] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_68_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1290_ _0257_ _0258_ net661 VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__mux2_1
XFILLER_63_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2813_ net701 VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__buf_1
X_1626_ _0568_ _0566_ _0573_ VGND VGND VPWR VPWR B_ADR0 sky130_fd_sc_hd__o21ai_4
X_2744_ net19 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__buf_1
X_2675_ clknet_4_15_0_UserCLK_regs _0077_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[19\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1488_ _0959_ net606 net682 _0444_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__o211ai_1
X_1557_ _0509_ _0508_ net683 VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2109_ net612 net865 _0918_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__mux2_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_210 net777 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2460_ net765 net704 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer4 _0400_ VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__dlymetal6s2s_1
X_2391_ net31 net696 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1411_ net17 net103 net131 Inst_RegFile_switch_matrix.JS2BEG6 Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__mux4_2
X_1273_ net396 _0243_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__or2_1
X_1342_ net661 _0308_ _0307_ net650 VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_62_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2589_ net764 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1609_ net60 net68 net86 net2 Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q
+ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__mux4_1
X_2658_ net758 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2727_ Inst_RegFile_switch_matrix.E1BEG1 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
XFILLER_67_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout691 net692 VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__clkbuf_2
Xfanout680 BD0 VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__buf_6
X_1891_ _0800_ _0799_ Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q VGND VGND VPWR VPWR
+ _0801_ sky130_fd_sc_hd__mux2_1
X_1960_ Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q _0559_ _0561_ Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q
+ _0557_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_31_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2512_ net745 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2443_ net763 net705 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_39_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2374_ net754 net693 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1256_ net64 net92 _0225_ _0226_ Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q
+ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__mux4_1
X_1325_ Inst_RegFile_32x4.mem\[6\]\[2\] Inst_RegFile_32x4.mem\[7\]\[2\] net630 VGND
+ VGND VPWR VPWR _0292_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1187_ _0158_ Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q _0161_ VGND VGND VPWR VPWR
+ _0162_ sky130_fd_sc_hd__a21o_1
XFILLER_20_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput272 net272 VGND VGND VPWR VPWR N4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput250 Inst_RegFile_switch_matrix.JN2BEG5 VGND VGND VPWR VPWR N2BEG[5] sky130_fd_sc_hd__buf_8
Xoutput283 Inst_RegFile_switch_matrix.NN4BEG3 VGND VGND VPWR VPWR NN4BEG[15] sky130_fd_sc_hd__buf_8
Xoutput261 net261 VGND VGND VPWR VPWR N4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput294 net294 VGND VGND VPWR VPWR S1BEG[1] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_73_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1110_ Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__inv_1
X_2090_ _0907_ _0891_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__nand2_8
XFILLER_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1041_ Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__inv_1
XFILLER_61_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1874_ _1013_ _0783_ _0787_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.EE4BEG0
+ sky130_fd_sc_hd__o21a_1
X_1943_ _1018_ _0826_ _0827_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__o21ai_2
X_2426_ net767 net700 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_UserCLK UserCLK VGND VGND VPWR VPWR clknet_0_UserCLK sky130_fd_sc_hd__clkbuf_16
X_1239_ _0210_ _0211_ _0961_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__mux2_1
X_2357_ net774 net690 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2288_ net52 net732 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1308_ net661 _0276_ _0275_ net650 VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__o211a_1
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1590_ Inst_RegFile_32x4.mem\[23\]\[2\] net607 VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__nand2_1
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2211_ clknet_4_3_0_UserCLK_regs _0035_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2073_ net622 net863 _0911_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__mux2_1
X_2142_ net601 net822 _0926_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__mux2_1
X_2975_ Inst_RegFile_switch_matrix.WW4BEG0 VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__buf_1
XFILLER_22_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1788_ Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q _0713_ Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q
+ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__a21bo_1
X_1857_ net640 _1033_ net685 _0772_ Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q
+ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__mux4_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1926_ net71 net127 net99 Inst_RegFile_switch_matrix.JW2BEG4 Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_55_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2409_ net749 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_64_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_73_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1711_ net87 net91 net89 net115 Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q
+ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__mux4_1
X_1642_ net677 net634 net665 net638 Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q
+ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__mux4_1
X_2760_ EE4END[6] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_1
XFILLER_31_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_2 net143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2691_ clknet_4_14_0_UserCLK_regs _0093_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1573_ _0389_ _0523_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__and2_1
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2056_ net611 net867 _0905_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__mux2_1
X_2125_ _0893_ _0898_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_52_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1909_ net637 _0437_ Inst_RegFile_switch_matrix.JN2BEG2 _0803_ Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E1BEG3
+ sky130_fd_sc_hd__mux4_1
X_2958_ W6END[9] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__buf_4
X_2889_ Inst_RegFile_switch_matrix.JS2BEG7 VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_68_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2812_ net705 VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_2
X_2743_ net18 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__buf_1
X_1625_ Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q _0572_ _0570_ Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q
+ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__a211o_1
X_2674_ clknet_4_13_0_UserCLK_regs _0076_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[19\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1556_ Inst_RegFile_32x4.mem\[4\]\[3\] Inst_RegFile_32x4.mem\[5\]\[3\] net609 VGND
+ VGND VPWR VPWR _0509_ sky130_fd_sc_hd__mux2_1
XFILLER_39_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1487_ Inst_RegFile_32x4.mem\[23\]\[0\] net606 VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_37_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2108_ net621 net926 _0918_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__mux2_4
X_2039_ _0891_ _0895_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__nand2_4
XFILLER_50_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold360 Inst_RegFile_32x4.mem\[22\]\[2\] VGND VGND VPWR VPWR net935 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_200 _0718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_211 net777 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1410_ _0366_ _0368_ _0371_ _0949_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JS2BEG6
+ sky130_fd_sc_hd__a22o_4
Xrebuffer5 AD3 VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2390_ net30 net696 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1272_ Inst_RegFile_32x4.mem\[14\]\[0\] Inst_RegFile_32x4.mem\[15\]\[0\] net626 VGND
+ VGND VPWR VPWR _0243_ sky130_fd_sc_hd__mux2_1
X_1341_ Inst_RegFile_32x4.mem\[20\]\[2\] Inst_RegFile_32x4.mem\[21\]\[2\] net628 VGND
+ VGND VPWR VPWR _0308_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2726_ Inst_RegFile_switch_matrix.E1BEG0 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_34_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2588_ net765 net57 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1608_ Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q _0554_ _0556_ VGND VGND VPWR VPWR
+ _0557_ sky130_fd_sc_hd__o21ai_4
X_2657_ net759 net738 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1539_ _0389_ _0491_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__and2_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout670 net671 VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__buf_8
Xfanout692 net693 VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__buf_2
Xfanout681 net684 VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__buf_8
XFILLER_33_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1890_ net667 _0718_ Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q VGND VGND VPWR VPWR
+ _0800_ sky130_fd_sc_hd__mux2_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2511_ net746 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2442_ net776 net705 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2373_ net755 net692 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1186_ Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q _0160_ Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q
+ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__o21ai_1
X_1255_ net76 net18 net104 net132 Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q
+ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__mux4_1
X_1324_ Inst_RegFile_32x4.mem\[4\]\[2\] Inst_RegFile_32x4.mem\[5\]\[2\] net630 VGND
+ VGND VPWR VPWR _0291_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2709_ clknet_4_3_0_UserCLK_regs _0111_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput240 net240 VGND VGND VPWR VPWR FrameStrobe_O[9] sky130_fd_sc_hd__buf_2
Xoutput262 net262 VGND VGND VPWR VPWR N4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput273 net273 VGND VGND VPWR VPWR N4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput251 net251 VGND VGND VPWR VPWR N2BEG[6] sky130_fd_sc_hd__buf_6
Xoutput284 net284 VGND VGND VPWR VPWR NN4BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_58_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput295 net295 VGND VGND VPWR VPWR S1BEG[2] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_73_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1942_ Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q _0726_ VGND VGND VPWR VPWR _0827_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1873_ _0784_ _0785_ _0786_ Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q
+ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__a221o_1
X_2356_ net775 net690 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2425_ net768 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1238_ net61 net85 net69 net780 Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q
+ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__mux4_1
X_2287_ net746 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1169_ _0145_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JS2BEG5 sky130_fd_sc_hd__inv_4
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1307_ Inst_RegFile_32x4.mem\[20\]\[1\] Inst_RegFile_32x4.mem\[21\]\[1\] net628 VGND
+ VGND VPWR VPWR _0276_ sky130_fd_sc_hd__mux2_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ clknet_4_7_0_UserCLK_regs _0034_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2072_ net617 net937 _0911_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__mux2_1
X_2141_ _0891_ _0923_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__nand2_4
X_1925_ _0809_ _0808_ Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q VGND VGND VPWR VPWR
+ _0810_ sky130_fd_sc_hd__mux2_4
X_2974_ WW4END[15] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__buf_1
X_1787_ Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q _0714_ VGND VGND VPWR VPWR _0715_
+ sky130_fd_sc_hd__and2b_1
X_1856_ net86 net11 net97 net125 Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q
+ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__mux4_1
X_2339_ net757 net734 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2408_ net750 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_3 E6END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1710_ net59 net1 net63 net5 Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q
+ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__mux4_1
X_1641_ Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q _0585_ VGND VGND VPWR VPWR _0586_
+ sky130_fd_sc_hd__or2_1
X_1572_ _0521_ _0522_ net682 VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__mux2_1
X_2690_ clknet_4_14_0_UserCLK_regs _0092_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2124_ net611 net912 _0921_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__mux2_2
XFILLER_62_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2055_ net623 net836 _0905_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__mux2_1
X_1839_ net83 net111 net779 net688 Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q
+ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__mux4_1
X_1908_ net680 Inst_RegFile_switch_matrix.E2BEG3 _0804_ _0805_ Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.S1BEG0
+ sky130_fd_sc_hd__mux4_1
X_2888_ Inst_RegFile_switch_matrix.JS2BEG6 VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__buf_1
X_2957_ W6END[8] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__buf_1
XFILLER_1_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput140 WW4END[3] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_4
XFILLER_51_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2811_ net708 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__buf_1
X_2742_ net17 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__buf_1
X_1624_ _0571_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__inv_2
X_2673_ clknet_4_7_0_UserCLK_regs Inst_RegFile_32x4.AD_comb\[3\] VGND VGND VPWR VPWR
+ Inst_RegFile_32x4.AD_reg\[3\] sky130_fd_sc_hd__dfxtp_1
X_1555_ Inst_RegFile_32x4.mem\[6\]\[3\] Inst_RegFile_32x4.mem\[7\]\[3\] net609 VGND
+ VGND VPWR VPWR _0508_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1486_ _0441_ _0442_ net683 VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__mux2_1
X_2107_ net616 net882 _0918_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__mux2_1
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2038_ net612 net885 _0899_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_20_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold361 Inst_RegFile_32x4.mem\[7\]\[3\] VGND VGND VPWR VPWR net936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold350 Inst_RegFile_32x4.mem\[7\]\[1\] VGND VGND VPWR VPWR net925 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_201 _1033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1340_ net674 _0306_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__or2_1
XFILLER_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1271_ Inst_RegFile_32x4.mem\[12\]\[0\] Inst_RegFile_32x4.mem\[13\]\[0\] net632 VGND
+ VGND VPWR VPWR _0242_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_62_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2656_ net760 net738 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2725_ clknet_4_3_0_UserCLK_regs _0127_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1607_ _0936_ _0555_ Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q VGND VGND VPWR VPWR
+ _0556_ sky130_fd_sc_hd__o21a_1
X_2587_ net766 net719 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1538_ _0489_ _0490_ net683 VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__mux2_1
X_1469_ _0423_ _0426_ net642 VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__mux2_1
XFILLER_67_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout693 FrameStrobe[9] VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__buf_2
Xfanout660 AD1 VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__buf_2
Xfanout671 AD0 VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__buf_8
Xfanout682 net683 VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__clkbuf_4
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2510_ net747 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_31_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2372_ net756 net692 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2441_ net749 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1323_ net661 _0287_ _0289_ net648 VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__o211a_1
XFILLER_68_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1254_ _0222_ _0223_ _0224_ _0940_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__a22o_1
X_1185_ _0159_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__inv_1
XFILLER_32_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput252 net252 VGND VGND VPWR VPWR N2BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput241 net241 VGND VGND VPWR VPWR N1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput230 net230 VGND VGND VPWR VPWR FrameStrobe_O[18] sky130_fd_sc_hd__buf_2
X_2639_ net746 net738 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2708_ clknet_4_8_0_UserCLK_regs _0110_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput285 net285 VGND VGND VPWR VPWR NN4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput263 net263 VGND VGND VPWR VPWR N4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput274 net274 VGND VGND VPWR VPWR N4BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput296 net296 VGND VGND VPWR VPWR S1BEG[3] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_73_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1872_ net89 net659 Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q VGND VGND VPWR VPWR
+ _0786_ sky130_fd_sc_hd__mux2_1
X_1941_ net84 net24 net108 Inst_RegFile_switch_matrix.JS2BEG2 Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_44_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2355_ net742 net690 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2286_ net747 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2424_ net770 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1306_ net675 _0274_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__or2_1
X_1237_ net11 net89 net97 net115 Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q
+ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__mux4_1
X_1168_ _0141_ _0139_ _0144_ _0973_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__a22oi_4
XFILLER_64_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1099_ Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_7_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ net613 net881 _0925_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__mux2_1
XFILLER_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2071_ net601 net869 _0911_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__mux2_1
X_1855_ Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q _0766_ _0770_ _0771_ VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix.EE4BEG3 sky130_fd_sc_hd__o22a_1
X_1924_ net63 net91 _1031_ _0148_ Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q
+ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__mux4_2
X_2973_ WW4END[14] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__buf_1
X_1786_ net669 net656 Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q VGND VGND VPWR VPWR
+ _0714_ sky130_fd_sc_hd__mux2_1
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2338_ net758 net734 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2269_ net764 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2407_ net45 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_55_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_4 E6END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1640_ net686 net669 net656 net644 Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q
+ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__mux4_1
X_1571_ Inst_RegFile_32x4.mem\[2\]\[2\] Inst_RegFile_32x4.mem\[3\]\[2\] net606 VGND
+ VGND VPWR VPWR _0522_ sky130_fd_sc_hd__mux2_1
XFILLER_66_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer27 _0436_ VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__dlygate4sd1_1
X_2123_ net620 net858 _0921_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2054_ net618 net846 _0905_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__mux2_1
X_1838_ _0750_ _0753_ Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q _0756_ VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix.E6BEG1 sky130_fd_sc_hd__a22o_1
X_1907_ net666 _0582_ Inst_RegFile_switch_matrix.E2BEG0 _0158_ Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.S1BEG1
+ sky130_fd_sc_hd__mux4_1
X_2956_ W6END[7] VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__buf_1
X_1769_ _0697_ _0698_ Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q VGND VGND VPWR VPWR
+ _0699_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput130 W2MID[3] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_2
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2810_ net713 VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_1
X_2741_ net16 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
X_2672_ clknet_4_12_0_UserCLK_regs Inst_RegFile_32x4.AD_comb\[2\] VGND VGND VPWR VPWR
+ Inst_RegFile_32x4.AD_reg\[2\] sky130_fd_sc_hd__dfxtp_1
X_1623_ net78 net20 net106 net134 Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q
+ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__mux4_1
X_1485_ Inst_RegFile_32x4.mem\[18\]\[0\] Inst_RegFile_32x4.mem\[19\]\[0\] net610 VGND
+ VGND VPWR VPWR _0442_ sky130_fd_sc_hd__mux2_1
X_1554_ _0506_ _0505_ net682 VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__mux2_1
.ends

