magic
tech ihp-sg13g2
magscale 1 2
timestamp 1743691610
<< metal1 >>
rect 1152 10604 45216 10628
rect 1152 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 45216 10604
rect 1152 10540 45216 10564
rect 1467 10436 1509 10445
rect 1467 10396 1468 10436
rect 1508 10396 1509 10436
rect 1467 10387 1509 10396
rect 3003 10436 3045 10445
rect 3003 10396 3004 10436
rect 3044 10396 3045 10436
rect 3003 10387 3045 10396
rect 3867 10436 3909 10445
rect 3867 10396 3868 10436
rect 3908 10396 3909 10436
rect 3867 10387 3909 10396
rect 5307 10436 5349 10445
rect 5307 10396 5308 10436
rect 5348 10396 5349 10436
rect 5307 10387 5349 10396
rect 5883 10436 5925 10445
rect 5883 10396 5884 10436
rect 5924 10396 5925 10436
rect 5883 10387 5925 10396
rect 7803 10436 7845 10445
rect 7803 10396 7804 10436
rect 7844 10396 7845 10436
rect 7803 10387 7845 10396
rect 8091 10436 8133 10445
rect 8091 10396 8092 10436
rect 8132 10396 8133 10436
rect 8091 10387 8133 10396
rect 9147 10436 9189 10445
rect 9147 10396 9148 10436
rect 9188 10396 9189 10436
rect 9147 10387 9189 10396
rect 11355 10436 11397 10445
rect 11355 10396 11356 10436
rect 11396 10396 11397 10436
rect 11355 10387 11397 10396
rect 11739 10436 11781 10445
rect 11739 10396 11740 10436
rect 11780 10396 11781 10436
rect 11739 10387 11781 10396
rect 16731 10436 16773 10445
rect 16731 10396 16732 10436
rect 16772 10396 16773 10436
rect 16731 10387 16773 10396
rect 17403 10436 17445 10445
rect 17403 10396 17404 10436
rect 17444 10396 17445 10436
rect 17403 10387 17445 10396
rect 19707 10436 19749 10445
rect 19707 10396 19708 10436
rect 19748 10396 19749 10436
rect 19707 10387 19749 10396
rect 24027 10436 24069 10445
rect 24027 10396 24028 10436
rect 24068 10396 24069 10436
rect 24027 10387 24069 10396
rect 27387 10436 27429 10445
rect 27387 10396 27388 10436
rect 27428 10396 27429 10436
rect 27387 10387 27429 10396
rect 27771 10436 27813 10445
rect 27771 10396 27772 10436
rect 27812 10396 27813 10436
rect 27771 10387 27813 10396
rect 29883 10436 29925 10445
rect 29883 10396 29884 10436
rect 29924 10396 29925 10436
rect 29883 10387 29925 10396
rect 32283 10436 32325 10445
rect 32283 10396 32284 10436
rect 32324 10396 32325 10436
rect 32283 10387 32325 10396
rect 34683 10436 34725 10445
rect 34683 10396 34684 10436
rect 34724 10396 34725 10436
rect 34683 10387 34725 10396
rect 36795 10436 36837 10445
rect 36795 10396 36796 10436
rect 36836 10396 36837 10436
rect 36795 10387 36837 10396
rect 37563 10436 37605 10445
rect 37563 10396 37564 10436
rect 37604 10396 37605 10436
rect 37563 10387 37605 10396
rect 38139 10436 38181 10445
rect 38139 10396 38140 10436
rect 38180 10396 38181 10436
rect 38139 10387 38181 10396
rect 38811 10436 38853 10445
rect 38811 10396 38812 10436
rect 38852 10396 38853 10436
rect 38811 10387 38853 10396
rect 40587 10436 40629 10445
rect 40587 10396 40588 10436
rect 40628 10396 40629 10436
rect 40587 10387 40629 10396
rect 42555 10436 42597 10445
rect 42555 10396 42556 10436
rect 42596 10396 42597 10436
rect 42555 10387 42597 10396
rect 42939 10436 42981 10445
rect 42939 10396 42940 10436
rect 42980 10396 42981 10436
rect 42939 10387 42981 10396
rect 44091 10436 44133 10445
rect 44091 10396 44092 10436
rect 44132 10396 44133 10436
rect 44091 10387 44133 10396
rect 44475 10436 44517 10445
rect 44475 10396 44476 10436
rect 44516 10396 44517 10436
rect 44475 10387 44517 10396
rect 8763 10352 8805 10361
rect 8763 10312 8764 10352
rect 8804 10312 8805 10352
rect 8763 10303 8805 10312
rect 32667 10352 32709 10361
rect 32667 10312 32668 10352
rect 32708 10312 32709 10352
rect 32667 10303 32709 10312
rect 38955 10352 38997 10361
rect 38955 10312 38956 10352
rect 38996 10312 38997 10352
rect 38955 10303 38997 10312
rect 42171 10352 42213 10361
rect 42171 10312 42172 10352
rect 42212 10312 42213 10352
rect 42171 10303 42213 10312
rect 44859 10352 44901 10361
rect 44859 10312 44860 10352
rect 44900 10312 44901 10352
rect 44859 10303 44901 10312
rect 6795 10268 6837 10277
rect 6795 10228 6796 10268
rect 6836 10228 6837 10268
rect 6795 10219 6837 10228
rect 6939 10268 6981 10277
rect 6939 10228 6940 10268
rect 6980 10228 6981 10268
rect 6939 10219 6981 10228
rect 7083 10268 7125 10277
rect 7083 10228 7084 10268
rect 7124 10228 7125 10268
rect 7083 10219 7125 10228
rect 7197 10268 7255 10269
rect 7197 10228 7206 10268
rect 7246 10228 7255 10268
rect 7197 10227 7255 10228
rect 7324 10268 7382 10269
rect 7324 10228 7333 10268
rect 7373 10228 7382 10268
rect 7324 10227 7382 10228
rect 9291 10268 9333 10277
rect 11883 10268 11925 10277
rect 13515 10268 13557 10277
rect 15147 10268 15189 10277
rect 17547 10268 17589 10277
rect 21483 10268 21525 10277
rect 9291 10228 9292 10268
rect 9332 10228 9333 10268
rect 9291 10219 9333 10228
rect 10539 10259 10581 10268
rect 10539 10219 10540 10259
rect 10580 10219 10581 10259
rect 11883 10228 11884 10268
rect 11924 10228 11925 10268
rect 11883 10219 11925 10228
rect 13131 10259 13173 10268
rect 13131 10219 13132 10259
rect 13172 10219 13173 10259
rect 13515 10228 13516 10268
rect 13556 10228 13557 10268
rect 13515 10219 13557 10228
rect 14763 10259 14805 10268
rect 14763 10219 14764 10259
rect 14804 10219 14805 10259
rect 15147 10228 15148 10268
rect 15188 10228 15189 10268
rect 15147 10219 15189 10228
rect 16395 10259 16437 10268
rect 16395 10219 16396 10259
rect 16436 10219 16437 10259
rect 17547 10228 17548 10268
rect 17588 10228 17589 10268
rect 17547 10219 17589 10228
rect 18795 10259 18837 10268
rect 18795 10219 18796 10259
rect 18836 10219 18837 10259
rect 10539 10210 10581 10219
rect 13131 10210 13173 10219
rect 14763 10210 14805 10219
rect 16395 10210 16437 10219
rect 18795 10210 18837 10219
rect 20235 10259 20277 10268
rect 20235 10219 20236 10259
rect 20276 10219 20277 10259
rect 21483 10228 21484 10268
rect 21524 10228 21525 10268
rect 21483 10219 21525 10228
rect 21867 10268 21909 10277
rect 24171 10268 24213 10277
rect 25803 10268 25845 10277
rect 28299 10268 28341 10277
rect 30315 10268 30357 10277
rect 21867 10228 21868 10268
rect 21908 10228 21909 10268
rect 21867 10219 21909 10228
rect 23115 10259 23157 10268
rect 23115 10219 23116 10259
rect 23156 10219 23157 10259
rect 24171 10228 24172 10268
rect 24212 10228 24213 10268
rect 24171 10219 24213 10228
rect 25419 10259 25461 10268
rect 25419 10219 25420 10259
rect 25460 10219 25461 10259
rect 25803 10228 25804 10268
rect 25844 10228 25845 10268
rect 25803 10219 25845 10228
rect 27051 10259 27093 10268
rect 27051 10219 27052 10259
rect 27092 10219 27093 10259
rect 28299 10228 28300 10268
rect 28340 10228 28341 10268
rect 28299 10219 28341 10228
rect 29547 10259 29589 10268
rect 29547 10219 29548 10259
rect 29588 10219 29589 10259
rect 30315 10228 30316 10268
rect 30356 10228 30357 10268
rect 30315 10219 30357 10228
rect 31563 10268 31621 10269
rect 31563 10228 31572 10268
rect 31612 10228 31621 10268
rect 31563 10227 31621 10228
rect 33099 10268 33141 10277
rect 35211 10268 35253 10277
rect 40395 10268 40437 10277
rect 42027 10268 42069 10277
rect 33099 10228 33100 10268
rect 33140 10228 33141 10268
rect 33099 10219 33141 10228
rect 34347 10259 34389 10268
rect 34347 10219 34348 10259
rect 34388 10219 34389 10259
rect 35211 10228 35212 10268
rect 35252 10228 35253 10268
rect 35211 10219 35253 10228
rect 36459 10259 36501 10268
rect 36459 10219 36460 10259
rect 36500 10219 36501 10259
rect 20235 10210 20277 10219
rect 23115 10210 23157 10219
rect 25419 10210 25461 10219
rect 27051 10210 27093 10219
rect 29547 10210 29589 10219
rect 34347 10210 34389 10219
rect 36459 10210 36501 10219
rect 39147 10259 39189 10268
rect 39147 10219 39148 10259
rect 39188 10219 39189 10259
rect 40395 10228 40396 10268
rect 40436 10228 40437 10268
rect 40395 10219 40437 10228
rect 40779 10259 40821 10268
rect 40779 10219 40780 10259
rect 40820 10219 40821 10259
rect 42027 10228 42028 10268
rect 42068 10228 42069 10268
rect 42027 10219 42069 10228
rect 39147 10210 39189 10219
rect 40779 10210 40821 10219
rect 1227 10184 1269 10193
rect 1227 10144 1228 10184
rect 1268 10144 1269 10184
rect 1227 10135 1269 10144
rect 1611 10184 1653 10193
rect 1611 10144 1612 10184
rect 1652 10144 1653 10184
rect 1611 10135 1653 10144
rect 1995 10184 2037 10193
rect 1995 10144 1996 10184
rect 2036 10144 2037 10184
rect 1995 10135 2037 10144
rect 2379 10184 2421 10193
rect 2379 10144 2380 10184
rect 2420 10144 2421 10184
rect 2379 10135 2421 10144
rect 2763 10184 2805 10193
rect 2763 10144 2764 10184
rect 2804 10144 2805 10184
rect 2763 10135 2805 10144
rect 3627 10184 3669 10193
rect 3627 10144 3628 10184
rect 3668 10144 3669 10184
rect 3627 10135 3669 10144
rect 4971 10184 5013 10193
rect 4971 10144 4972 10184
rect 5012 10144 5013 10184
rect 4971 10135 5013 10144
rect 5547 10184 5589 10193
rect 5547 10144 5548 10184
rect 5588 10144 5589 10184
rect 5547 10135 5589 10144
rect 6123 10184 6165 10193
rect 6123 10144 6124 10184
rect 6164 10144 6165 10184
rect 6123 10135 6165 10144
rect 7563 10184 7605 10193
rect 7563 10144 7564 10184
rect 7604 10144 7605 10184
rect 7563 10135 7605 10144
rect 8331 10184 8373 10193
rect 8331 10144 8332 10184
rect 8372 10144 8373 10184
rect 8331 10135 8373 10144
rect 8523 10184 8565 10193
rect 8523 10144 8524 10184
rect 8564 10144 8565 10184
rect 8523 10135 8565 10144
rect 8907 10184 8949 10193
rect 8907 10144 8908 10184
rect 8948 10144 8949 10184
rect 8907 10135 8949 10144
rect 11115 10184 11157 10193
rect 11115 10144 11116 10184
rect 11156 10144 11157 10184
rect 11115 10135 11157 10144
rect 11499 10184 11541 10193
rect 11499 10144 11500 10184
rect 11540 10144 11541 10184
rect 11499 10135 11541 10144
rect 16971 10184 17013 10193
rect 16971 10144 16972 10184
rect 17012 10144 17013 10184
rect 16971 10135 17013 10144
rect 17163 10184 17205 10193
rect 17163 10144 17164 10184
rect 17204 10144 17205 10184
rect 17163 10135 17205 10144
rect 19467 10184 19509 10193
rect 19467 10144 19468 10184
rect 19508 10144 19509 10184
rect 19467 10135 19509 10144
rect 23787 10184 23829 10193
rect 23787 10144 23788 10184
rect 23828 10144 23829 10184
rect 23787 10135 23829 10144
rect 27627 10184 27669 10193
rect 27627 10144 27628 10184
rect 27668 10144 27669 10184
rect 27627 10135 27669 10144
rect 28011 10184 28053 10193
rect 28011 10144 28012 10184
rect 28052 10144 28053 10184
rect 28011 10135 28053 10144
rect 30123 10184 30165 10193
rect 30123 10144 30124 10184
rect 30164 10144 30165 10184
rect 30123 10135 30165 10144
rect 31947 10184 31989 10193
rect 31947 10144 31948 10184
rect 31988 10144 31989 10184
rect 31947 10135 31989 10144
rect 32187 10184 32229 10193
rect 32187 10144 32188 10184
rect 32228 10144 32229 10184
rect 32187 10135 32229 10144
rect 32523 10184 32565 10193
rect 32523 10144 32524 10184
rect 32564 10144 32565 10184
rect 32523 10135 32565 10144
rect 32907 10184 32949 10193
rect 32907 10144 32908 10184
rect 32948 10144 32949 10184
rect 32907 10135 32949 10144
rect 34923 10184 34965 10193
rect 34923 10144 34924 10184
rect 34964 10144 34965 10184
rect 34923 10135 34965 10144
rect 37035 10184 37077 10193
rect 37035 10144 37036 10184
rect 37076 10144 37077 10184
rect 37035 10135 37077 10144
rect 37227 10184 37269 10193
rect 37227 10144 37228 10184
rect 37268 10144 37269 10184
rect 37227 10135 37269 10144
rect 37803 10184 37845 10193
rect 37803 10144 37804 10184
rect 37844 10144 37845 10184
rect 37803 10135 37845 10144
rect 38379 10184 38421 10193
rect 38379 10144 38380 10184
rect 38420 10144 38421 10184
rect 38379 10135 38421 10144
rect 38571 10184 38613 10193
rect 38571 10144 38572 10184
rect 38612 10144 38613 10184
rect 38571 10135 38613 10144
rect 42411 10184 42453 10193
rect 42411 10144 42412 10184
rect 42452 10144 42453 10184
rect 42411 10135 42453 10144
rect 42795 10184 42837 10193
rect 42795 10144 42796 10184
rect 42836 10144 42837 10184
rect 42795 10135 42837 10144
rect 43179 10184 43221 10193
rect 43179 10144 43180 10184
rect 43220 10144 43221 10184
rect 43179 10135 43221 10144
rect 43563 10184 43605 10193
rect 43563 10144 43564 10184
rect 43604 10144 43605 10184
rect 43563 10135 43605 10144
rect 43707 10184 43749 10193
rect 43707 10144 43708 10184
rect 43748 10144 43749 10184
rect 43707 10135 43749 10144
rect 43947 10184 43989 10193
rect 43947 10144 43948 10184
rect 43988 10144 43989 10184
rect 43947 10135 43989 10144
rect 44331 10184 44373 10193
rect 44331 10144 44332 10184
rect 44372 10144 44373 10184
rect 44331 10135 44373 10144
rect 44715 10184 44757 10193
rect 44715 10144 44716 10184
rect 44756 10144 44757 10184
rect 44715 10135 44757 10144
rect 45099 10184 45141 10193
rect 45099 10144 45100 10184
rect 45140 10144 45141 10184
rect 45099 10135 45141 10144
rect 2235 10100 2277 10109
rect 2235 10060 2236 10100
rect 2276 10060 2277 10100
rect 2235 10051 2277 10060
rect 5211 10100 5253 10109
rect 5211 10060 5212 10100
rect 5252 10060 5253 10100
rect 5211 10051 5253 10060
rect 7179 10100 7221 10109
rect 7179 10060 7180 10100
rect 7220 10060 7221 10100
rect 7179 10051 7221 10060
rect 16587 10100 16629 10109
rect 16587 10060 16588 10100
rect 16628 10060 16629 10100
rect 16587 10051 16629 10060
rect 25611 10100 25653 10109
rect 25611 10060 25612 10100
rect 25652 10060 25653 10100
rect 25611 10051 25653 10060
rect 27243 10100 27285 10109
rect 27243 10060 27244 10100
rect 27284 10060 27285 10100
rect 27243 10051 27285 10060
rect 37467 10100 37509 10109
rect 37467 10060 37468 10100
rect 37508 10060 37509 10100
rect 37467 10051 37509 10060
rect 43323 10100 43365 10109
rect 43323 10060 43324 10100
rect 43364 10060 43365 10100
rect 43323 10051 43365 10060
rect 1851 10016 1893 10025
rect 1851 9976 1852 10016
rect 1892 9976 1893 10016
rect 1851 9967 1893 9976
rect 2619 10016 2661 10025
rect 2619 9976 2620 10016
rect 2660 9976 2661 10016
rect 2619 9967 2661 9976
rect 10731 10016 10773 10025
rect 10731 9976 10732 10016
rect 10772 9976 10773 10016
rect 10731 9967 10773 9976
rect 13323 10016 13365 10025
rect 13323 9976 13324 10016
rect 13364 9976 13365 10016
rect 13323 9967 13365 9976
rect 14955 10016 14997 10025
rect 14955 9976 14956 10016
rect 14996 9976 14997 10016
rect 14955 9967 14997 9976
rect 18987 10016 19029 10025
rect 18987 9976 18988 10016
rect 19028 9976 19029 10016
rect 18987 9967 19029 9976
rect 20043 10016 20085 10025
rect 20043 9976 20044 10016
rect 20084 9976 20085 10016
rect 20043 9967 20085 9976
rect 23307 10016 23349 10025
rect 23307 9976 23308 10016
rect 23348 9976 23349 10016
rect 23307 9967 23349 9976
rect 29739 10016 29781 10025
rect 29739 9976 29740 10016
rect 29780 9976 29781 10016
rect 29739 9967 29781 9976
rect 31755 10016 31797 10025
rect 31755 9976 31756 10016
rect 31796 9976 31797 10016
rect 31755 9967 31797 9976
rect 34539 10016 34581 10025
rect 34539 9976 34540 10016
rect 34580 9976 34581 10016
rect 34539 9967 34581 9976
rect 36651 10016 36693 10025
rect 36651 9976 36652 10016
rect 36692 9976 36693 10016
rect 36651 9967 36693 9976
rect 1152 9848 45216 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 45216 9848
rect 1152 9784 45216 9808
rect 5739 9680 5781 9689
rect 5739 9640 5740 9680
rect 5780 9640 5781 9680
rect 5739 9631 5781 9640
rect 7371 9680 7413 9689
rect 7371 9640 7372 9680
rect 7412 9640 7413 9680
rect 7371 9631 7413 9640
rect 13947 9680 13989 9689
rect 13947 9640 13948 9680
rect 13988 9640 13989 9680
rect 13947 9631 13989 9640
rect 14811 9680 14853 9689
rect 14811 9640 14812 9680
rect 14852 9640 14853 9680
rect 14811 9631 14853 9640
rect 18171 9680 18213 9689
rect 18171 9640 18172 9680
rect 18212 9640 18213 9680
rect 18171 9631 18213 9640
rect 20763 9680 20805 9689
rect 20763 9640 20764 9680
rect 20804 9640 20805 9680
rect 20763 9631 20805 9640
rect 26235 9680 26277 9689
rect 26235 9640 26236 9680
rect 26276 9640 26277 9680
rect 26235 9631 26277 9640
rect 33147 9680 33189 9689
rect 33147 9640 33148 9680
rect 33188 9640 33189 9680
rect 33147 9631 33189 9640
rect 33915 9680 33957 9689
rect 33915 9640 33916 9680
rect 33956 9640 33957 9680
rect 33915 9631 33957 9640
rect 44187 9680 44229 9689
rect 44187 9640 44188 9680
rect 44228 9640 44229 9680
rect 44187 9631 44229 9640
rect 44571 9680 44613 9689
rect 44571 9640 44572 9680
rect 44612 9640 44613 9680
rect 44571 9631 44613 9640
rect 21435 9596 21477 9605
rect 21435 9556 21436 9596
rect 21476 9556 21477 9596
rect 21435 9547 21477 9556
rect 43035 9596 43077 9605
rect 43035 9556 43036 9596
rect 43076 9556 43077 9596
rect 43035 9547 43077 9556
rect 1227 9512 1269 9521
rect 1227 9472 1228 9512
rect 1268 9472 1269 9512
rect 1227 9463 1269 9472
rect 1611 9512 1653 9521
rect 1611 9472 1612 9512
rect 1652 9472 1653 9512
rect 1611 9463 1653 9472
rect 1995 9512 2037 9521
rect 1995 9472 1996 9512
rect 2036 9472 2037 9512
rect 1995 9463 2037 9472
rect 2235 9512 2277 9521
rect 2235 9472 2236 9512
rect 2276 9472 2277 9512
rect 2235 9463 2277 9472
rect 8139 9512 8181 9521
rect 8139 9472 8140 9512
rect 8180 9472 8181 9512
rect 8139 9463 8181 9472
rect 8523 9512 8565 9521
rect 8523 9472 8524 9512
rect 8564 9472 8565 9512
rect 8523 9463 8565 9472
rect 9003 9512 9045 9521
rect 9003 9472 9004 9512
rect 9044 9472 9045 9512
rect 9003 9463 9045 9472
rect 11979 9512 12021 9521
rect 11979 9472 11980 9512
rect 12020 9472 12021 9512
rect 11979 9463 12021 9472
rect 13258 9512 13316 9513
rect 13258 9472 13267 9512
rect 13307 9472 13316 9512
rect 13258 9471 13316 9472
rect 13419 9512 13461 9521
rect 13419 9472 13420 9512
rect 13460 9472 13461 9512
rect 13419 9463 13461 9472
rect 14187 9512 14229 9521
rect 14187 9472 14188 9512
rect 14228 9472 14229 9512
rect 14187 9463 14229 9472
rect 14571 9512 14613 9521
rect 14571 9472 14572 9512
rect 14612 9472 14613 9512
rect 14571 9463 14613 9472
rect 15531 9512 15573 9521
rect 15531 9472 15532 9512
rect 15572 9472 15573 9512
rect 15531 9463 15573 9472
rect 16971 9512 17013 9521
rect 16971 9472 16972 9512
rect 17012 9472 17013 9512
rect 16971 9463 17013 9472
rect 17931 9512 17973 9521
rect 17931 9472 17932 9512
rect 17972 9472 17973 9512
rect 17931 9463 17973 9472
rect 18891 9512 18933 9521
rect 18891 9472 18892 9512
rect 18932 9472 18933 9512
rect 18891 9463 18933 9472
rect 20170 9512 20228 9513
rect 20170 9472 20179 9512
rect 20219 9472 20228 9512
rect 20170 9471 20228 9472
rect 20331 9512 20373 9521
rect 20331 9472 20332 9512
rect 20372 9472 20373 9512
rect 20331 9463 20373 9472
rect 21003 9512 21045 9521
rect 21003 9472 21004 9512
rect 21044 9472 21045 9512
rect 21003 9463 21045 9472
rect 21226 9512 21284 9513
rect 21226 9472 21235 9512
rect 21275 9472 21284 9512
rect 21226 9471 21284 9472
rect 22155 9512 22197 9521
rect 22155 9472 22156 9512
rect 22196 9472 22197 9512
rect 22155 9463 22197 9472
rect 23434 9512 23492 9513
rect 23434 9472 23443 9512
rect 23483 9472 23492 9512
rect 23434 9471 23492 9472
rect 23595 9512 23637 9521
rect 23595 9472 23596 9512
rect 23636 9472 23637 9512
rect 23595 9463 23637 9472
rect 24843 9512 24885 9521
rect 24843 9472 24844 9512
rect 24884 9472 24885 9512
rect 24843 9463 24885 9472
rect 26475 9512 26517 9521
rect 26475 9472 26476 9512
rect 26516 9472 26517 9512
rect 26475 9463 26517 9472
rect 26698 9512 26756 9513
rect 26698 9472 26707 9512
rect 26747 9472 26756 9512
rect 26698 9471 26756 9472
rect 26907 9512 26949 9521
rect 26907 9472 26908 9512
rect 26948 9472 26949 9512
rect 26907 9463 26949 9472
rect 27819 9512 27861 9521
rect 27819 9472 27820 9512
rect 27860 9472 27861 9512
rect 27819 9463 27861 9472
rect 29242 9512 29300 9513
rect 29242 9472 29251 9512
rect 29291 9472 29300 9512
rect 29242 9471 29300 9472
rect 31755 9512 31797 9521
rect 31755 9472 31756 9512
rect 31796 9472 31797 9512
rect 31755 9463 31797 9472
rect 33387 9512 33429 9521
rect 33387 9472 33388 9512
rect 33428 9472 33429 9512
rect 33387 9463 33429 9472
rect 33771 9512 33813 9521
rect 33771 9472 33772 9512
rect 33812 9472 33813 9512
rect 33771 9463 33813 9472
rect 34155 9512 34197 9521
rect 34155 9472 34156 9512
rect 34196 9472 34197 9512
rect 34155 9463 34197 9472
rect 35019 9512 35061 9521
rect 35019 9472 35020 9512
rect 35060 9472 35061 9512
rect 35019 9463 35061 9472
rect 36555 9512 36597 9521
rect 36555 9472 36556 9512
rect 36596 9472 36597 9512
rect 36555 9463 36597 9472
rect 42027 9512 42069 9521
rect 42027 9472 42028 9512
rect 42068 9472 42069 9512
rect 42027 9463 42069 9472
rect 42651 9512 42693 9521
rect 42651 9472 42652 9512
rect 42692 9472 42693 9512
rect 42651 9463 42693 9472
rect 42891 9512 42933 9521
rect 42891 9472 42892 9512
rect 42932 9472 42933 9512
rect 42891 9463 42933 9472
rect 43275 9512 43317 9521
rect 43275 9472 43276 9512
rect 43316 9472 43317 9512
rect 43275 9463 43317 9472
rect 43659 9512 43701 9521
rect 43659 9472 43660 9512
rect 43700 9472 43701 9512
rect 43659 9463 43701 9472
rect 44043 9512 44085 9521
rect 44043 9472 44044 9512
rect 44084 9472 44085 9512
rect 44043 9463 44085 9472
rect 44427 9512 44469 9521
rect 44427 9472 44428 9512
rect 44468 9472 44469 9512
rect 44427 9463 44469 9472
rect 44811 9512 44853 9521
rect 44811 9472 44812 9512
rect 44852 9472 44853 9512
rect 44811 9463 44853 9472
rect 4299 9428 4341 9437
rect 4299 9388 4300 9428
rect 4340 9388 4341 9428
rect 4299 9379 4341 9388
rect 5539 9428 5597 9429
rect 5539 9388 5548 9428
rect 5588 9388 5597 9428
rect 5539 9387 5597 9388
rect 5931 9428 5973 9437
rect 5931 9388 5932 9428
rect 5972 9388 5973 9428
rect 5931 9379 5973 9388
rect 7171 9428 7229 9429
rect 7171 9388 7180 9428
rect 7220 9388 7229 9428
rect 7171 9387 7229 9388
rect 7659 9428 7701 9437
rect 7659 9388 7660 9428
rect 7700 9388 7701 9428
rect 7659 9379 7701 9388
rect 7778 9428 7820 9437
rect 7778 9388 7779 9428
rect 7819 9388 7820 9428
rect 7778 9379 7820 9388
rect 7890 9428 7932 9437
rect 7890 9388 7891 9428
rect 7931 9388 7932 9428
rect 7890 9379 7932 9388
rect 9675 9428 9717 9437
rect 9675 9388 9676 9428
rect 9716 9388 9717 9428
rect 9675 9379 9717 9388
rect 10915 9428 10973 9429
rect 10915 9388 10924 9428
rect 10964 9388 10973 9428
rect 10915 9387 10973 9388
rect 11469 9428 11511 9437
rect 11469 9388 11470 9428
rect 11510 9388 11511 9428
rect 12075 9428 12117 9437
rect 11469 9379 11511 9388
rect 11578 9400 11636 9401
rect 11578 9360 11587 9400
rect 11627 9360 11636 9400
rect 12075 9388 12076 9428
rect 12116 9388 12117 9428
rect 12075 9379 12117 9388
rect 12547 9428 12605 9429
rect 12547 9388 12556 9428
rect 12596 9388 12605 9428
rect 12547 9387 12605 9388
rect 13066 9428 13124 9429
rect 13066 9388 13075 9428
rect 13115 9388 13124 9428
rect 13066 9387 13124 9388
rect 15021 9428 15063 9437
rect 15021 9388 15022 9428
rect 15062 9388 15063 9428
rect 15021 9379 15063 9388
rect 15147 9428 15189 9437
rect 15147 9388 15148 9428
rect 15188 9388 15189 9428
rect 15147 9379 15189 9388
rect 15627 9428 15669 9437
rect 15627 9388 15628 9428
rect 15668 9388 15669 9428
rect 15627 9379 15669 9388
rect 16099 9428 16157 9429
rect 16099 9388 16108 9428
rect 16148 9388 16157 9428
rect 16099 9387 16157 9388
rect 16587 9428 16645 9429
rect 16587 9388 16596 9428
rect 16636 9388 16645 9428
rect 16587 9387 16645 9388
rect 18394 9428 18452 9429
rect 18394 9388 18403 9428
rect 18443 9388 18452 9428
rect 18394 9387 18452 9388
rect 18507 9428 18549 9437
rect 18507 9388 18508 9428
rect 18548 9388 18549 9428
rect 18507 9379 18549 9388
rect 18987 9428 19029 9437
rect 18987 9388 18988 9428
rect 19028 9388 19029 9428
rect 18987 9379 19029 9388
rect 19459 9428 19517 9429
rect 19459 9388 19468 9428
rect 19508 9388 19517 9428
rect 19459 9387 19517 9388
rect 19978 9428 20036 9429
rect 19978 9388 19987 9428
rect 20027 9388 20036 9428
rect 19978 9387 20036 9388
rect 21658 9428 21716 9429
rect 21658 9388 21667 9428
rect 21707 9388 21716 9428
rect 21658 9387 21716 9388
rect 21771 9428 21813 9437
rect 21771 9388 21772 9428
rect 21812 9388 21813 9428
rect 21771 9379 21813 9388
rect 22251 9428 22293 9437
rect 22251 9388 22252 9428
rect 22292 9388 22293 9428
rect 22251 9379 22293 9388
rect 22723 9428 22781 9429
rect 22723 9388 22732 9428
rect 22772 9388 22781 9428
rect 22723 9387 22781 9388
rect 23242 9428 23300 9429
rect 23242 9388 23251 9428
rect 23291 9388 23300 9428
rect 23242 9387 23300 9388
rect 24346 9428 24404 9429
rect 24346 9388 24355 9428
rect 24395 9388 24404 9428
rect 24346 9387 24404 9388
rect 24459 9428 24501 9437
rect 24459 9388 24460 9428
rect 24500 9388 24501 9428
rect 24459 9379 24501 9388
rect 24939 9428 24981 9437
rect 24939 9388 24940 9428
rect 24980 9388 24981 9428
rect 24939 9379 24981 9388
rect 25411 9428 25469 9429
rect 25411 9388 25420 9428
rect 25460 9388 25469 9428
rect 25411 9387 25469 9388
rect 25899 9428 25957 9429
rect 25899 9388 25908 9428
rect 25948 9388 25957 9428
rect 25899 9387 25957 9388
rect 27322 9428 27380 9429
rect 27322 9388 27331 9428
rect 27371 9388 27380 9428
rect 27322 9387 27380 9388
rect 27435 9428 27477 9437
rect 27435 9388 27436 9428
rect 27476 9388 27477 9428
rect 27435 9379 27477 9388
rect 27915 9428 27957 9437
rect 27915 9388 27916 9428
rect 27956 9388 27957 9428
rect 27915 9379 27957 9388
rect 28387 9428 28445 9429
rect 28387 9388 28396 9428
rect 28436 9388 28445 9428
rect 28387 9387 28445 9388
rect 28906 9428 28964 9429
rect 28906 9388 28915 9428
rect 28955 9388 28964 9428
rect 28906 9387 28964 9388
rect 29443 9428 29501 9429
rect 29443 9388 29452 9428
rect 29492 9388 29501 9428
rect 29443 9387 29501 9388
rect 30699 9428 30741 9437
rect 30699 9388 30700 9428
rect 30740 9388 30741 9428
rect 30699 9379 30741 9388
rect 31258 9428 31316 9429
rect 31258 9388 31267 9428
rect 31307 9388 31316 9428
rect 31258 9387 31316 9388
rect 31371 9428 31413 9437
rect 31371 9388 31372 9428
rect 31412 9388 31413 9428
rect 31371 9379 31413 9388
rect 31851 9428 31893 9437
rect 31851 9388 31852 9428
rect 31892 9388 31893 9428
rect 31851 9379 31893 9388
rect 32323 9428 32381 9429
rect 32323 9388 32332 9428
rect 32372 9388 32381 9428
rect 32323 9387 32381 9388
rect 32811 9428 32869 9429
rect 32811 9388 32820 9428
rect 32860 9388 32869 9428
rect 32811 9387 32869 9388
rect 34518 9428 34576 9429
rect 34518 9388 34527 9428
rect 34567 9388 34576 9428
rect 34518 9387 34576 9388
rect 34635 9428 34677 9437
rect 34635 9388 34636 9428
rect 34676 9388 34677 9428
rect 34635 9379 34677 9388
rect 35115 9428 35157 9437
rect 35115 9388 35116 9428
rect 35156 9388 35157 9428
rect 35115 9379 35157 9388
rect 35587 9428 35645 9429
rect 35587 9388 35596 9428
rect 35636 9388 35645 9428
rect 35587 9387 35645 9388
rect 36106 9428 36164 9429
rect 36106 9388 36115 9428
rect 36155 9388 36164 9428
rect 36106 9387 36164 9388
rect 37123 9428 37181 9429
rect 37123 9388 37132 9428
rect 37172 9388 37181 9428
rect 37123 9387 37181 9388
rect 38379 9428 38421 9437
rect 38379 9388 38380 9428
rect 38420 9388 38421 9428
rect 38379 9379 38421 9388
rect 38763 9428 38805 9437
rect 38763 9388 38764 9428
rect 38804 9388 38805 9428
rect 38763 9379 38805 9388
rect 40003 9428 40061 9429
rect 40003 9388 40012 9428
rect 40052 9388 40061 9428
rect 40003 9387 40061 9388
rect 40400 9428 40442 9437
rect 40400 9388 40401 9428
rect 40441 9388 40442 9428
rect 40400 9379 40442 9388
rect 41635 9428 41693 9429
rect 41635 9388 41644 9428
rect 41684 9388 41693 9428
rect 41635 9387 41693 9388
rect 11578 9359 11636 9360
rect 7563 9344 7605 9353
rect 7563 9304 7564 9344
rect 7604 9304 7605 9344
rect 7563 9295 7605 9304
rect 20571 9344 20613 9353
rect 20571 9304 20572 9344
rect 20612 9304 20613 9344
rect 20571 9295 20613 9304
rect 36939 9344 36981 9353
rect 36939 9304 36940 9344
rect 36980 9304 36981 9344
rect 36939 9295 36981 9304
rect 43803 9344 43845 9353
rect 43803 9304 43804 9344
rect 43844 9304 43845 9344
rect 43803 9295 43845 9304
rect 1467 9260 1509 9269
rect 1467 9220 1468 9260
rect 1508 9220 1509 9260
rect 1467 9211 1509 9220
rect 1851 9260 1893 9269
rect 1851 9220 1852 9260
rect 1892 9220 1893 9260
rect 1851 9211 1893 9220
rect 7371 9260 7413 9269
rect 7371 9220 7372 9260
rect 7412 9220 7413 9260
rect 7371 9211 7413 9220
rect 8379 9260 8421 9269
rect 8379 9220 8380 9260
rect 8420 9220 8421 9260
rect 8379 9211 8421 9220
rect 8763 9260 8805 9269
rect 8763 9220 8764 9260
rect 8804 9220 8805 9260
rect 8763 9211 8805 9220
rect 9243 9260 9285 9269
rect 9243 9220 9244 9260
rect 9284 9220 9285 9260
rect 9243 9211 9285 9220
rect 11115 9260 11157 9269
rect 11115 9220 11116 9260
rect 11156 9220 11157 9260
rect 11115 9211 11157 9220
rect 13659 9260 13701 9269
rect 13659 9220 13660 9260
rect 13700 9220 13701 9260
rect 13659 9211 13701 9220
rect 16779 9260 16821 9269
rect 16779 9220 16780 9260
rect 16820 9220 16821 9260
rect 16779 9211 16821 9220
rect 17211 9260 17253 9269
rect 17211 9220 17212 9260
rect 17252 9220 17253 9260
rect 17211 9211 17253 9220
rect 23835 9260 23877 9269
rect 23835 9220 23836 9260
rect 23876 9220 23877 9260
rect 23835 9211 23877 9220
rect 26091 9260 26133 9269
rect 26091 9220 26092 9260
rect 26132 9220 26133 9260
rect 26091 9211 26133 9220
rect 29067 9260 29109 9269
rect 29067 9220 29068 9260
rect 29108 9220 29109 9260
rect 29067 9211 29109 9220
rect 33003 9260 33045 9269
rect 33003 9220 33004 9260
rect 33044 9220 33045 9260
rect 33003 9211 33045 9220
rect 33531 9260 33573 9269
rect 33531 9220 33532 9260
rect 33572 9220 33573 9260
rect 33531 9211 33573 9220
rect 36267 9260 36309 9269
rect 36267 9220 36268 9260
rect 36308 9220 36309 9260
rect 36267 9211 36309 9220
rect 36795 9260 36837 9269
rect 36795 9220 36796 9260
rect 36836 9220 36837 9260
rect 36795 9211 36837 9220
rect 40203 9260 40245 9269
rect 40203 9220 40204 9260
rect 40244 9220 40245 9260
rect 40203 9211 40245 9220
rect 41835 9260 41877 9269
rect 41835 9220 41836 9260
rect 41876 9220 41877 9260
rect 41835 9211 41877 9220
rect 42267 9260 42309 9269
rect 42267 9220 42268 9260
rect 42308 9220 42309 9260
rect 42267 9211 42309 9220
rect 43419 9260 43461 9269
rect 43419 9220 43420 9260
rect 43460 9220 43461 9260
rect 43419 9211 43461 9220
rect 1152 9092 45216 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 45216 9092
rect 1152 9028 45216 9052
rect 1851 8924 1893 8933
rect 1851 8884 1852 8924
rect 1892 8884 1893 8924
rect 1851 8875 1893 8884
rect 12459 8924 12501 8933
rect 12459 8884 12460 8924
rect 12500 8884 12501 8924
rect 12459 8875 12501 8884
rect 12651 8924 12693 8933
rect 12651 8884 12652 8924
rect 12692 8884 12693 8924
rect 12651 8875 12693 8884
rect 15723 8924 15765 8933
rect 15723 8884 15724 8924
rect 15764 8884 15765 8924
rect 15723 8875 15765 8884
rect 17355 8924 17397 8933
rect 17355 8884 17356 8924
rect 17396 8884 17397 8924
rect 17355 8875 17397 8884
rect 19371 8924 19413 8933
rect 19371 8884 19372 8924
rect 19412 8884 19413 8924
rect 19371 8875 19413 8884
rect 19707 8924 19749 8933
rect 19707 8884 19708 8924
rect 19748 8884 19749 8924
rect 19707 8875 19749 8884
rect 21675 8924 21717 8933
rect 21675 8884 21676 8924
rect 21716 8884 21717 8924
rect 21675 8875 21717 8884
rect 22107 8924 22149 8933
rect 22107 8884 22108 8924
rect 22148 8884 22149 8924
rect 22107 8875 22149 8884
rect 24267 8924 24309 8933
rect 24267 8884 24268 8924
rect 24308 8884 24309 8924
rect 24267 8875 24309 8884
rect 31755 8924 31797 8933
rect 31755 8884 31756 8924
rect 31796 8884 31797 8924
rect 31755 8875 31797 8884
rect 33387 8924 33429 8933
rect 33387 8884 33388 8924
rect 33428 8884 33429 8924
rect 33387 8875 33429 8884
rect 44475 8924 44517 8933
rect 44475 8884 44476 8924
rect 44516 8884 44517 8924
rect 44475 8875 44517 8884
rect 9675 8840 9717 8849
rect 9675 8800 9676 8840
rect 9716 8800 9717 8840
rect 9675 8791 9717 8800
rect 10491 8840 10533 8849
rect 10491 8800 10492 8840
rect 10532 8800 10533 8840
rect 10491 8791 10533 8800
rect 29403 8840 29445 8849
rect 29403 8800 29404 8840
rect 29444 8800 29445 8840
rect 29403 8791 29445 8800
rect 36219 8840 36261 8849
rect 36219 8800 36220 8840
rect 36260 8800 36261 8840
rect 36219 8791 36261 8800
rect 42171 8840 42213 8849
rect 42171 8800 42172 8840
rect 42212 8800 42213 8840
rect 42171 8791 42213 8800
rect 43035 8840 43077 8849
rect 43035 8800 43036 8840
rect 43076 8800 43077 8840
rect 43035 8791 43077 8800
rect 4299 8756 4341 8765
rect 5931 8756 5973 8765
rect 7710 8756 7768 8757
rect 4299 8716 4300 8756
rect 4340 8716 4341 8756
rect 4299 8707 4341 8716
rect 5547 8747 5589 8756
rect 5547 8707 5548 8747
rect 5588 8707 5589 8747
rect 5931 8716 5932 8756
rect 5972 8716 5973 8756
rect 5931 8707 5973 8716
rect 7179 8747 7221 8756
rect 7179 8707 7180 8747
rect 7220 8707 7221 8747
rect 7710 8716 7719 8756
rect 7759 8716 7768 8756
rect 7930 8756 7988 8757
rect 7710 8715 7768 8716
rect 7836 8736 7878 8745
rect 5547 8698 5589 8707
rect 7179 8698 7221 8707
rect 7836 8696 7837 8736
rect 7877 8696 7878 8736
rect 7930 8716 7939 8756
rect 7979 8716 7988 8756
rect 7930 8715 7988 8716
rect 8235 8756 8277 8765
rect 10714 8756 10772 8757
rect 8235 8716 8236 8756
rect 8276 8716 8277 8756
rect 8235 8707 8277 8716
rect 9483 8747 9525 8756
rect 9483 8707 9484 8747
rect 9524 8707 9525 8747
rect 10714 8716 10723 8756
rect 10763 8716 10772 8756
rect 10714 8715 10772 8716
rect 10827 8756 10869 8765
rect 10827 8716 10828 8756
rect 10868 8716 10869 8756
rect 10827 8707 10869 8716
rect 11211 8756 11253 8765
rect 12827 8756 12885 8757
rect 11211 8716 11212 8756
rect 11252 8716 11253 8756
rect 11211 8707 11253 8716
rect 11787 8747 11829 8756
rect 11787 8707 11788 8747
rect 11828 8707 11829 8747
rect 9483 8698 9525 8707
rect 11787 8698 11829 8707
rect 12267 8747 12309 8756
rect 12267 8707 12268 8747
rect 12308 8707 12309 8747
rect 12827 8716 12836 8756
rect 12876 8716 12885 8756
rect 12827 8715 12885 8716
rect 14091 8756 14133 8765
rect 14091 8716 14092 8756
rect 14132 8716 14133 8756
rect 14091 8707 14133 8716
rect 14283 8756 14325 8765
rect 15915 8756 15957 8765
rect 17626 8756 17684 8757
rect 14283 8716 14284 8756
rect 14324 8716 14325 8756
rect 14283 8707 14325 8716
rect 15531 8747 15573 8756
rect 15531 8707 15532 8747
rect 15572 8707 15573 8747
rect 15915 8716 15916 8756
rect 15956 8716 15957 8756
rect 15915 8707 15957 8716
rect 17163 8747 17205 8756
rect 17163 8707 17164 8747
rect 17204 8707 17205 8747
rect 17626 8716 17635 8756
rect 17675 8716 17684 8756
rect 17626 8715 17684 8716
rect 17739 8756 17781 8765
rect 17739 8716 17740 8756
rect 17780 8716 17781 8756
rect 17739 8707 17781 8716
rect 18123 8756 18165 8765
rect 20235 8756 20277 8765
rect 22827 8756 22869 8765
rect 25227 8756 25269 8765
rect 27051 8756 27093 8765
rect 30010 8756 30068 8757
rect 18123 8716 18124 8756
rect 18164 8716 18165 8756
rect 18123 8707 18165 8716
rect 18699 8747 18741 8756
rect 18699 8707 18700 8747
rect 18740 8707 18741 8747
rect 12267 8698 12309 8707
rect 15531 8698 15573 8707
rect 17163 8698 17205 8707
rect 18699 8698 18741 8707
rect 19179 8747 19221 8756
rect 19179 8707 19180 8747
rect 19220 8707 19221 8747
rect 20235 8716 20236 8756
rect 20276 8716 20277 8756
rect 20235 8707 20277 8716
rect 21483 8747 21525 8756
rect 21483 8707 21484 8747
rect 21524 8707 21525 8747
rect 22827 8716 22828 8756
rect 22868 8716 22869 8756
rect 22827 8707 22869 8716
rect 24075 8747 24117 8756
rect 24075 8707 24076 8747
rect 24116 8707 24117 8747
rect 25227 8716 25228 8756
rect 25268 8716 25269 8756
rect 25227 8707 25269 8716
rect 26475 8747 26517 8756
rect 26475 8707 26476 8747
rect 26516 8707 26517 8747
rect 27051 8716 27052 8756
rect 27092 8716 27093 8756
rect 27051 8707 27093 8716
rect 28299 8747 28341 8756
rect 28299 8707 28300 8747
rect 28340 8707 28341 8747
rect 30010 8716 30019 8756
rect 30059 8716 30068 8756
rect 30010 8715 30068 8716
rect 30123 8756 30165 8765
rect 30123 8716 30124 8756
rect 30164 8716 30165 8756
rect 30123 8707 30165 8716
rect 30507 8756 30549 8765
rect 31947 8756 31989 8765
rect 34330 8756 34388 8757
rect 30507 8716 30508 8756
rect 30548 8716 30549 8756
rect 30507 8707 30549 8716
rect 31083 8747 31125 8756
rect 31083 8707 31084 8747
rect 31124 8707 31125 8747
rect 19179 8698 19221 8707
rect 21483 8698 21525 8707
rect 24075 8698 24117 8707
rect 26475 8698 26517 8707
rect 28299 8698 28341 8707
rect 31083 8698 31125 8707
rect 31563 8747 31605 8756
rect 31563 8707 31564 8747
rect 31604 8707 31605 8747
rect 31947 8716 31948 8756
rect 31988 8716 31989 8756
rect 31947 8707 31989 8716
rect 33195 8747 33237 8756
rect 33195 8707 33196 8747
rect 33236 8707 33237 8747
rect 34330 8716 34339 8756
rect 34379 8716 34388 8756
rect 34330 8715 34388 8716
rect 34443 8756 34485 8765
rect 34443 8716 34444 8756
rect 34484 8716 34485 8756
rect 34443 8707 34485 8716
rect 34827 8756 34869 8765
rect 36747 8756 36789 8765
rect 38379 8756 38421 8765
rect 40282 8756 40340 8757
rect 34827 8716 34828 8756
rect 34868 8716 34869 8756
rect 34827 8707 34869 8716
rect 35403 8747 35445 8756
rect 35403 8707 35404 8747
rect 35444 8707 35445 8747
rect 31563 8698 31605 8707
rect 33195 8698 33237 8707
rect 35403 8698 35445 8707
rect 35883 8747 35925 8756
rect 35883 8707 35884 8747
rect 35924 8707 35925 8747
rect 36747 8716 36748 8756
rect 36788 8716 36789 8756
rect 36747 8707 36789 8716
rect 37995 8747 38037 8756
rect 37995 8707 37996 8747
rect 38036 8707 38037 8747
rect 38379 8716 38380 8756
rect 38420 8716 38421 8756
rect 38379 8707 38421 8716
rect 39627 8747 39669 8756
rect 39627 8707 39628 8747
rect 39668 8707 39669 8747
rect 40282 8716 40291 8756
rect 40331 8716 40340 8756
rect 40282 8715 40340 8716
rect 40384 8756 40442 8757
rect 40384 8716 40393 8756
rect 40433 8716 40442 8756
rect 40384 8715 40442 8716
rect 40779 8756 40821 8765
rect 40779 8716 40780 8756
rect 40820 8716 40821 8756
rect 40779 8707 40821 8716
rect 41355 8747 41397 8756
rect 41355 8707 41356 8747
rect 41396 8707 41397 8747
rect 35883 8698 35925 8707
rect 37995 8698 38037 8707
rect 39627 8698 39669 8707
rect 41355 8698 41397 8707
rect 41835 8747 41877 8756
rect 41835 8707 41836 8747
rect 41876 8707 41877 8747
rect 41835 8698 41877 8707
rect 7836 8687 7878 8696
rect 1227 8672 1269 8681
rect 1227 8632 1228 8672
rect 1268 8632 1269 8672
rect 1227 8623 1269 8632
rect 1611 8672 1653 8681
rect 1611 8632 1612 8672
rect 1652 8632 1653 8672
rect 1611 8623 1653 8632
rect 2571 8672 2613 8681
rect 2571 8632 2572 8672
rect 2612 8632 2613 8672
rect 2571 8623 2613 8632
rect 2811 8672 2853 8681
rect 2811 8632 2812 8672
rect 2852 8632 2853 8672
rect 2811 8623 2853 8632
rect 3915 8672 3957 8681
rect 3915 8632 3916 8672
rect 3956 8632 3957 8672
rect 3915 8623 3957 8632
rect 4155 8672 4197 8681
rect 4155 8632 4156 8672
rect 4196 8632 4197 8672
rect 4155 8623 4197 8632
rect 10251 8672 10293 8681
rect 10251 8632 10252 8672
rect 10292 8632 10293 8672
rect 10251 8623 10293 8632
rect 11307 8672 11349 8681
rect 11307 8632 11308 8672
rect 11348 8632 11349 8672
rect 11307 8623 11349 8632
rect 18219 8672 18261 8681
rect 18219 8632 18220 8672
rect 18260 8632 18261 8672
rect 18219 8623 18261 8632
rect 19947 8672 19989 8681
rect 19947 8632 19948 8672
rect 19988 8632 19989 8672
rect 19947 8623 19989 8632
rect 21867 8672 21909 8681
rect 21867 8632 21868 8672
rect 21908 8632 21909 8672
rect 21867 8623 21909 8632
rect 29115 8672 29157 8681
rect 29115 8632 29116 8672
rect 29156 8632 29157 8672
rect 29115 8623 29157 8632
rect 29547 8672 29589 8681
rect 29547 8632 29548 8672
rect 29588 8632 29589 8672
rect 29547 8623 29589 8632
rect 30603 8672 30645 8681
rect 30603 8632 30604 8672
rect 30644 8632 30645 8672
rect 30603 8623 30645 8632
rect 34923 8672 34965 8681
rect 34923 8632 34924 8672
rect 34964 8632 34965 8672
rect 34923 8623 34965 8632
rect 36106 8672 36164 8673
rect 36106 8632 36115 8672
rect 36155 8632 36164 8672
rect 36106 8631 36164 8632
rect 36459 8672 36501 8681
rect 36459 8632 36460 8672
rect 36500 8632 36501 8672
rect 36459 8623 36501 8632
rect 40875 8672 40917 8681
rect 40875 8632 40876 8672
rect 40916 8632 40917 8672
rect 40875 8623 40917 8632
rect 42058 8672 42116 8673
rect 42058 8632 42067 8672
rect 42107 8632 42116 8672
rect 42058 8631 42116 8632
rect 42411 8672 42453 8681
rect 42411 8632 42412 8672
rect 42452 8632 42453 8672
rect 42411 8623 42453 8632
rect 42795 8672 42837 8681
rect 42795 8632 42796 8672
rect 42836 8632 42837 8672
rect 42795 8623 42837 8632
rect 43371 8672 43413 8681
rect 43371 8632 43372 8672
rect 43412 8632 43413 8672
rect 43371 8623 43413 8632
rect 43755 8672 43797 8681
rect 43755 8632 43756 8672
rect 43796 8632 43797 8672
rect 43755 8623 43797 8632
rect 44091 8672 44133 8681
rect 44091 8632 44092 8672
rect 44132 8632 44133 8672
rect 44091 8623 44133 8632
rect 44331 8672 44373 8681
rect 44331 8632 44332 8672
rect 44372 8632 44373 8672
rect 44331 8623 44373 8632
rect 44715 8672 44757 8681
rect 44715 8632 44716 8672
rect 44756 8632 44757 8672
rect 44715 8623 44757 8632
rect 44907 8672 44949 8681
rect 44907 8632 44908 8672
rect 44948 8632 44949 8672
rect 44907 8623 44949 8632
rect 45147 8672 45189 8681
rect 45147 8632 45148 8672
rect 45188 8632 45189 8672
rect 45147 8623 45189 8632
rect 7371 8588 7413 8597
rect 7371 8548 7372 8588
rect 7412 8548 7413 8588
rect 7371 8539 7413 8548
rect 43995 8588 44037 8597
rect 43995 8548 43996 8588
rect 44036 8548 44037 8588
rect 43995 8539 44037 8548
rect 1467 8504 1509 8513
rect 1467 8464 1468 8504
rect 1508 8464 1509 8504
rect 1467 8455 1509 8464
rect 5739 8504 5781 8513
rect 5739 8464 5740 8504
rect 5780 8464 5781 8504
rect 5739 8455 5781 8464
rect 7563 8504 7605 8513
rect 7563 8464 7564 8504
rect 7604 8464 7605 8504
rect 7563 8455 7605 8464
rect 26667 8504 26709 8513
rect 26667 8464 26668 8504
rect 26708 8464 26709 8504
rect 26667 8455 26709 8464
rect 28491 8504 28533 8513
rect 28491 8464 28492 8504
rect 28532 8464 28533 8504
rect 28491 8455 28533 8464
rect 29787 8504 29829 8513
rect 29787 8464 29788 8504
rect 29828 8464 29829 8504
rect 29787 8455 29829 8464
rect 38187 8504 38229 8513
rect 38187 8464 38188 8504
rect 38228 8464 38229 8504
rect 38187 8455 38229 8464
rect 39819 8504 39861 8513
rect 39819 8464 39820 8504
rect 39860 8464 39861 8504
rect 39819 8455 39861 8464
rect 43131 8504 43173 8513
rect 43131 8464 43132 8504
rect 43172 8464 43173 8504
rect 43131 8455 43173 8464
rect 1152 8336 45216 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 45216 8336
rect 1152 8272 45216 8296
rect 11643 8168 11685 8177
rect 11643 8128 11644 8168
rect 11684 8128 11685 8168
rect 11643 8119 11685 8128
rect 12027 8168 12069 8177
rect 12027 8128 12028 8168
rect 12068 8128 12069 8168
rect 12027 8119 12069 8128
rect 13755 8168 13797 8177
rect 13755 8128 13756 8168
rect 13796 8128 13797 8168
rect 13755 8119 13797 8128
rect 15387 8168 15429 8177
rect 15387 8128 15388 8168
rect 15428 8128 15429 8168
rect 15387 8119 15429 8128
rect 23163 8168 23205 8177
rect 23163 8128 23164 8168
rect 23204 8128 23205 8168
rect 23163 8119 23205 8128
rect 34443 8168 34485 8177
rect 34443 8128 34444 8168
rect 34484 8128 34485 8168
rect 34443 8119 34485 8128
rect 36267 8168 36309 8177
rect 36267 8128 36268 8168
rect 36308 8128 36309 8168
rect 36267 8119 36309 8128
rect 37083 8168 37125 8177
rect 37083 8128 37084 8168
rect 37124 8128 37125 8168
rect 37083 8119 37125 8128
rect 41691 8168 41733 8177
rect 41691 8128 41692 8168
rect 41732 8128 41733 8168
rect 41691 8119 41733 8128
rect 42555 8168 42597 8177
rect 42555 8128 42556 8168
rect 42596 8128 42597 8168
rect 42555 8119 42597 8128
rect 42939 8168 42981 8177
rect 42939 8128 42940 8168
rect 42980 8128 42981 8168
rect 42939 8119 42981 8128
rect 43323 8168 43365 8177
rect 43323 8128 43324 8168
rect 43364 8128 43365 8168
rect 43323 8119 43365 8128
rect 4203 8084 4245 8093
rect 15003 8084 15045 8093
rect 4203 8044 4204 8084
rect 4244 8044 4245 8084
rect 4203 8035 4245 8044
rect 10299 8075 10341 8084
rect 10299 8035 10300 8075
rect 10340 8035 10341 8075
rect 15003 8044 15004 8084
rect 15044 8044 15045 8084
rect 15003 8035 15045 8044
rect 26571 8084 26613 8093
rect 26571 8044 26572 8084
rect 26612 8044 26613 8084
rect 26571 8035 26613 8044
rect 44091 8084 44133 8093
rect 44091 8044 44092 8084
rect 44132 8044 44133 8084
rect 44091 8035 44133 8044
rect 10299 8026 10341 8035
rect 1227 8000 1269 8009
rect 1227 7960 1228 8000
rect 1268 7960 1269 8000
rect 1227 7951 1269 7960
rect 1611 8000 1653 8009
rect 1611 7960 1612 8000
rect 1652 7960 1653 8000
rect 1611 7951 1653 7960
rect 6123 8000 6165 8009
rect 6123 7960 6124 8000
rect 6164 7960 6165 8000
rect 6123 7951 6165 7960
rect 7778 8000 7820 8009
rect 7778 7960 7779 8000
rect 7819 7960 7820 8000
rect 7224 7949 7266 7958
rect 7778 7951 7820 7960
rect 8122 8000 8180 8001
rect 8122 7960 8131 8000
rect 8171 7960 8180 8000
rect 8122 7959 8180 7960
rect 8523 8000 8565 8009
rect 8523 7960 8524 8000
rect 8564 7960 8565 8000
rect 8523 7951 8565 7960
rect 11499 8000 11541 8009
rect 11499 7960 11500 8000
rect 11540 7960 11541 8000
rect 11499 7951 11541 7960
rect 11883 8000 11925 8009
rect 11883 7960 11884 8000
rect 11924 7960 11925 8000
rect 11883 7951 11925 7960
rect 12267 8000 12309 8009
rect 12267 7960 12268 8000
rect 12308 7960 12309 8000
rect 12267 7951 12309 7960
rect 12459 8000 12501 8009
rect 12459 7960 12460 8000
rect 12500 7960 12501 8000
rect 12459 7951 12501 7960
rect 13035 8000 13077 8009
rect 13035 7960 13036 8000
rect 13076 7960 13077 8000
rect 13035 7951 13077 7960
rect 13515 8000 13557 8009
rect 13515 7960 13516 8000
rect 13556 7960 13557 8000
rect 13515 7951 13557 7960
rect 13995 8000 14037 8009
rect 13995 7960 13996 8000
rect 14036 7960 14037 8000
rect 13995 7951 14037 7960
rect 14235 8000 14277 8009
rect 14235 7960 14236 8000
rect 14276 7960 14277 8000
rect 14235 7951 14277 7960
rect 14379 8000 14421 8009
rect 14379 7960 14380 8000
rect 14420 7960 14421 8000
rect 14379 7951 14421 7960
rect 14763 8000 14805 8009
rect 14763 7960 14764 8000
rect 14804 7960 14805 8000
rect 14763 7951 14805 7960
rect 15147 8000 15189 8009
rect 15147 7960 15148 8000
rect 15188 7960 15189 8000
rect 15147 7951 15189 7960
rect 15723 8000 15765 8009
rect 15723 7960 15724 8000
rect 15764 7960 15765 8000
rect 15723 7951 15765 7960
rect 15915 8000 15957 8009
rect 15915 7960 15916 8000
rect 15956 7960 15957 8000
rect 15915 7951 15957 7960
rect 16299 8000 16341 8009
rect 16299 7960 16300 8000
rect 16340 7960 16341 8000
rect 16299 7951 16341 7960
rect 18315 8000 18357 8009
rect 18315 7960 18316 8000
rect 18356 7960 18357 8000
rect 18315 7951 18357 7960
rect 18699 8000 18741 8009
rect 18699 7960 18700 8000
rect 18740 7960 18741 8000
rect 18699 7951 18741 7960
rect 19083 8000 19125 8009
rect 19083 7960 19084 8000
rect 19124 7960 19125 8000
rect 19083 7951 19125 7960
rect 19755 8000 19797 8009
rect 19755 7960 19756 8000
rect 19796 7960 19797 8000
rect 19755 7951 19797 7960
rect 20331 8000 20373 8009
rect 20331 7960 20332 8000
rect 20372 7960 20373 8000
rect 20331 7951 20373 7960
rect 23403 8000 23445 8009
rect 23403 7960 23404 8000
rect 23444 7960 23445 8000
rect 23403 7951 23445 7960
rect 23787 8000 23829 8009
rect 23787 7960 23788 8000
rect 23828 7960 23829 8000
rect 23787 7951 23829 7960
rect 27435 8000 27477 8009
rect 27435 7960 27436 8000
rect 27476 7960 27477 8000
rect 27435 7951 27477 7960
rect 28714 8000 28772 8001
rect 28714 7960 28723 8000
rect 28763 7960 28772 8000
rect 28714 7959 28772 7960
rect 29067 8000 29109 8009
rect 29067 7960 29068 8000
rect 29108 7960 29109 8000
rect 29067 7951 29109 7960
rect 29451 8000 29493 8009
rect 29451 7960 29452 8000
rect 29492 7960 29493 8000
rect 29451 7951 29493 7960
rect 29835 8000 29877 8009
rect 29835 7960 29836 8000
rect 29876 7960 29877 8000
rect 29835 7951 29877 7960
rect 30795 8000 30837 8009
rect 30795 7960 30796 8000
rect 30836 7960 30837 8000
rect 30795 7951 30837 7960
rect 32074 8000 32132 8001
rect 32074 7960 32083 8000
rect 32123 7960 32132 8000
rect 32074 7959 32132 7960
rect 32235 8000 32277 8009
rect 32235 7960 32236 8000
rect 32276 7960 32277 8000
rect 32235 7951 32277 7960
rect 32811 8000 32853 8009
rect 32811 7960 32812 8000
rect 32852 7960 32853 8000
rect 32811 7951 32853 7960
rect 36651 8000 36693 8009
rect 36651 7960 36652 8000
rect 36692 7960 36693 8000
rect 36651 7951 36693 7960
rect 36843 8000 36885 8009
rect 36843 7960 36844 8000
rect 36884 7960 36885 8000
rect 36843 7951 36885 7960
rect 38571 8000 38613 8009
rect 38571 7960 38572 8000
rect 38612 7960 38613 8000
rect 38571 7951 38613 7960
rect 41931 8000 41973 8009
rect 41931 7960 41932 8000
rect 41972 7960 41973 8000
rect 41931 7951 41973 7960
rect 42315 8000 42357 8009
rect 42315 7960 42316 8000
rect 42356 7960 42357 8000
rect 42315 7951 42357 7960
rect 42699 8000 42741 8009
rect 42699 7960 42700 8000
rect 42740 7960 42741 8000
rect 42699 7951 42741 7960
rect 43083 8000 43125 8009
rect 43083 7960 43084 8000
rect 43124 7960 43125 8000
rect 43083 7951 43125 7960
rect 43659 8000 43701 8009
rect 43659 7960 43660 8000
rect 43700 7960 43701 8000
rect 43659 7951 43701 7960
rect 44331 8000 44373 8009
rect 44331 7960 44332 8000
rect 44372 7960 44373 8000
rect 44331 7951 44373 7960
rect 44523 8000 44565 8009
rect 44523 7960 44524 8000
rect 44564 7960 44565 8000
rect 44523 7951 44565 7960
rect 44907 8000 44949 8009
rect 44907 7960 44908 8000
rect 44948 7960 44949 8000
rect 44907 7951 44949 7960
rect 2763 7916 2805 7925
rect 2763 7876 2764 7916
rect 2804 7876 2805 7916
rect 2763 7867 2805 7876
rect 4003 7916 4061 7917
rect 4003 7876 4012 7916
rect 4052 7876 4061 7916
rect 4003 7875 4061 7876
rect 5146 7916 5204 7917
rect 5146 7876 5155 7916
rect 5195 7876 5204 7916
rect 5146 7875 5204 7876
rect 5635 7916 5693 7917
rect 5635 7876 5644 7916
rect 5684 7876 5693 7916
rect 5635 7875 5693 7876
rect 6219 7916 6261 7925
rect 6219 7876 6220 7916
rect 6260 7876 6261 7916
rect 6219 7867 6261 7876
rect 6603 7916 6645 7925
rect 6603 7876 6604 7916
rect 6644 7876 6645 7916
rect 6984 7916 7042 7917
rect 6603 7867 6645 7876
rect 6716 7896 6758 7905
rect 6716 7856 6717 7896
rect 6757 7856 6758 7896
rect 6984 7876 6993 7916
rect 7033 7876 7042 7916
rect 6984 7875 7042 7876
rect 7101 7916 7159 7917
rect 7101 7876 7110 7916
rect 7150 7876 7159 7916
rect 7224 7909 7225 7949
rect 7265 7909 7266 7949
rect 7224 7900 7266 7909
rect 7323 7916 7365 7925
rect 7101 7875 7159 7876
rect 7323 7876 7324 7916
rect 7364 7876 7365 7916
rect 7323 7867 7365 7876
rect 7659 7916 7701 7925
rect 7659 7876 7660 7916
rect 7700 7876 7701 7916
rect 7659 7867 7701 7876
rect 7890 7916 7932 7925
rect 7890 7876 7891 7916
rect 7931 7876 7932 7916
rect 7890 7867 7932 7876
rect 7995 7916 8037 7925
rect 7995 7876 7996 7916
rect 8036 7876 8037 7916
rect 7995 7867 8037 7876
rect 8235 7916 8277 7925
rect 8235 7876 8236 7916
rect 8276 7876 8277 7916
rect 8235 7867 8277 7876
rect 9003 7916 9045 7925
rect 9003 7876 9004 7916
rect 9044 7876 9045 7916
rect 9003 7867 9045 7876
rect 9291 7916 9333 7925
rect 9291 7876 9292 7916
rect 9332 7876 9333 7916
rect 9291 7867 9333 7876
rect 9579 7916 9621 7925
rect 9579 7876 9580 7916
rect 9620 7876 9621 7916
rect 9579 7867 9621 7876
rect 10051 7916 10109 7917
rect 10051 7876 10060 7916
rect 10100 7876 10109 7916
rect 10051 7875 10109 7876
rect 10330 7916 10388 7917
rect 10330 7876 10339 7916
rect 10379 7876 10388 7916
rect 10330 7875 10388 7876
rect 10731 7916 10773 7925
rect 10731 7876 10732 7916
rect 10772 7876 10773 7916
rect 10731 7867 10773 7876
rect 10923 7916 10965 7925
rect 10923 7876 10924 7916
rect 10964 7876 10965 7916
rect 10923 7867 10965 7876
rect 16683 7916 16725 7925
rect 16683 7876 16684 7916
rect 16724 7876 16725 7916
rect 16683 7867 16725 7876
rect 17923 7916 17981 7917
rect 17923 7876 17932 7916
rect 17972 7876 17981 7916
rect 17923 7875 17981 7876
rect 20715 7916 20757 7925
rect 20715 7876 20716 7916
rect 20756 7876 20757 7916
rect 20715 7867 20757 7876
rect 21955 7916 22013 7917
rect 21955 7876 21964 7916
rect 22004 7876 22013 7916
rect 21955 7875 22013 7876
rect 24171 7916 24213 7925
rect 24171 7876 24172 7916
rect 24212 7876 24213 7916
rect 24171 7867 24213 7876
rect 25411 7916 25469 7917
rect 25411 7876 25420 7916
rect 25460 7876 25469 7916
rect 25411 7875 25469 7876
rect 25899 7916 25941 7925
rect 25899 7876 25900 7916
rect 25940 7876 25941 7916
rect 25899 7867 25941 7876
rect 26146 7916 26204 7917
rect 26146 7876 26155 7916
rect 26195 7876 26204 7916
rect 26146 7875 26204 7876
rect 26266 7916 26324 7917
rect 26266 7876 26275 7916
rect 26315 7876 26324 7916
rect 26266 7875 26324 7876
rect 26938 7916 26996 7917
rect 26938 7876 26947 7916
rect 26987 7876 26996 7916
rect 26938 7875 26996 7876
rect 27051 7916 27093 7925
rect 27051 7876 27052 7916
rect 27092 7876 27093 7916
rect 27051 7867 27093 7876
rect 27531 7916 27573 7925
rect 27531 7876 27532 7916
rect 27572 7876 27573 7916
rect 27531 7867 27573 7876
rect 28003 7916 28061 7917
rect 28003 7876 28012 7916
rect 28052 7876 28061 7916
rect 28003 7875 28061 7876
rect 28491 7916 28549 7917
rect 28491 7876 28500 7916
rect 28540 7876 28549 7916
rect 28491 7875 28549 7876
rect 30298 7916 30356 7917
rect 30298 7876 30307 7916
rect 30347 7876 30356 7916
rect 30298 7875 30356 7876
rect 30411 7916 30453 7925
rect 30411 7876 30412 7916
rect 30452 7876 30453 7916
rect 30411 7867 30453 7876
rect 30891 7916 30933 7925
rect 30891 7876 30892 7916
rect 30932 7876 30933 7916
rect 30891 7867 30933 7876
rect 31363 7916 31421 7917
rect 31363 7876 31372 7916
rect 31412 7876 31421 7916
rect 31363 7875 31421 7876
rect 31882 7916 31940 7917
rect 31882 7876 31891 7916
rect 31931 7876 31940 7916
rect 31882 7875 31940 7876
rect 33003 7916 33045 7925
rect 33003 7876 33004 7916
rect 33044 7876 33045 7916
rect 33003 7867 33045 7876
rect 34243 7916 34301 7917
rect 34243 7876 34252 7916
rect 34292 7876 34301 7916
rect 34243 7875 34301 7876
rect 34827 7916 34869 7925
rect 34827 7876 34828 7916
rect 34868 7876 34869 7916
rect 34827 7867 34869 7876
rect 36067 7916 36125 7917
rect 36067 7876 36076 7916
rect 36116 7876 36125 7916
rect 36067 7875 36125 7876
rect 37978 7916 38036 7917
rect 37978 7876 37987 7916
rect 38027 7876 38036 7916
rect 37978 7875 38036 7876
rect 38091 7916 38133 7925
rect 38091 7876 38092 7916
rect 38132 7876 38133 7916
rect 38091 7867 38133 7876
rect 38468 7916 38510 7925
rect 38468 7876 38469 7916
rect 38509 7876 38510 7916
rect 38468 7867 38510 7876
rect 39043 7916 39101 7917
rect 39043 7876 39052 7916
rect 39092 7876 39101 7916
rect 39043 7875 39101 7876
rect 39562 7916 39620 7917
rect 39562 7876 39571 7916
rect 39611 7876 39620 7916
rect 39562 7875 39620 7876
rect 40107 7916 40149 7925
rect 40107 7876 40108 7916
rect 40148 7876 40149 7916
rect 40107 7867 40149 7876
rect 41347 7916 41405 7917
rect 41347 7876 41356 7916
rect 41396 7876 41405 7916
rect 41347 7875 41405 7876
rect 6716 7847 6758 7856
rect 7563 7832 7605 7841
rect 7563 7792 7564 7832
rect 7604 7792 7605 7832
rect 7563 7783 7605 7792
rect 8314 7832 8372 7833
rect 8314 7792 8323 7832
rect 8363 7792 8372 7832
rect 8314 7791 8372 7792
rect 8763 7832 8805 7841
rect 8763 7792 8764 7832
rect 8804 7792 8805 7832
rect 8763 7783 8805 7792
rect 9757 7832 9799 7841
rect 9757 7792 9758 7832
rect 9798 7792 9799 7832
rect 9757 7783 9799 7792
rect 10827 7832 10869 7841
rect 10827 7792 10828 7832
rect 10868 7792 10869 7832
rect 10827 7783 10869 7792
rect 14619 7832 14661 7841
rect 14619 7792 14620 7832
rect 14660 7792 14661 7832
rect 14619 7783 14661 7792
rect 19323 7832 19365 7841
rect 19323 7792 19324 7832
rect 19364 7792 19365 7832
rect 19323 7783 19365 7792
rect 25611 7832 25653 7841
rect 25611 7792 25612 7832
rect 25652 7792 25653 7832
rect 25611 7783 25653 7792
rect 32475 7832 32517 7841
rect 32475 7792 32476 7832
rect 32516 7792 32517 7832
rect 32475 7783 32517 7792
rect 44763 7832 44805 7841
rect 44763 7792 44764 7832
rect 44804 7792 44805 7832
rect 44763 7783 44805 7792
rect 1467 7748 1509 7757
rect 1467 7708 1468 7748
rect 1508 7708 1509 7748
rect 1467 7699 1509 7708
rect 1851 7748 1893 7757
rect 1851 7708 1852 7748
rect 1892 7708 1893 7748
rect 1851 7699 1893 7708
rect 4971 7748 5013 7757
rect 4971 7708 4972 7748
rect 5012 7708 5013 7748
rect 4971 7699 5013 7708
rect 7371 7748 7413 7757
rect 7371 7708 7372 7748
rect 7412 7708 7413 7748
rect 7371 7699 7413 7708
rect 8859 7748 8901 7757
rect 8859 7708 8860 7748
rect 8900 7708 8901 7748
rect 8859 7699 8901 7708
rect 9370 7748 9428 7749
rect 9370 7708 9379 7748
rect 9419 7708 9428 7748
rect 9370 7707 9428 7708
rect 9850 7748 9908 7749
rect 9850 7708 9859 7748
rect 9899 7708 9908 7748
rect 9850 7707 9908 7708
rect 9963 7748 10005 7757
rect 9963 7708 9964 7748
rect 10004 7708 10005 7748
rect 9963 7699 10005 7708
rect 10522 7748 10580 7749
rect 10522 7708 10531 7748
rect 10571 7708 10580 7748
rect 10522 7707 10580 7708
rect 11259 7748 11301 7757
rect 11259 7708 11260 7748
rect 11300 7708 11301 7748
rect 11259 7699 11301 7708
rect 12699 7748 12741 7757
rect 12699 7708 12700 7748
rect 12740 7708 12741 7748
rect 12699 7699 12741 7708
rect 13275 7748 13317 7757
rect 13275 7708 13276 7748
rect 13316 7708 13317 7748
rect 13275 7699 13317 7708
rect 15483 7748 15525 7757
rect 15483 7708 15484 7748
rect 15524 7708 15525 7748
rect 15483 7699 15525 7708
rect 16155 7748 16197 7757
rect 16155 7708 16156 7748
rect 16196 7708 16197 7748
rect 16155 7699 16197 7708
rect 16539 7748 16581 7757
rect 16539 7708 16540 7748
rect 16580 7708 16581 7748
rect 16539 7699 16581 7708
rect 18123 7748 18165 7757
rect 18123 7708 18124 7748
rect 18164 7708 18165 7748
rect 18123 7699 18165 7708
rect 18555 7748 18597 7757
rect 18555 7708 18556 7748
rect 18596 7708 18597 7748
rect 18555 7699 18597 7708
rect 18939 7748 18981 7757
rect 18939 7708 18940 7748
rect 18980 7708 18981 7748
rect 18939 7699 18981 7708
rect 19995 7748 20037 7757
rect 19995 7708 19996 7748
rect 20036 7708 20037 7748
rect 19995 7699 20037 7708
rect 20571 7748 20613 7757
rect 20571 7708 20572 7748
rect 20612 7708 20613 7748
rect 20571 7699 20613 7708
rect 22155 7748 22197 7757
rect 22155 7708 22156 7748
rect 22196 7708 22197 7748
rect 22155 7699 22197 7708
rect 24027 7748 24069 7757
rect 24027 7708 24028 7748
rect 24068 7708 24069 7748
rect 24027 7699 24069 7708
rect 28827 7748 28869 7757
rect 28827 7708 28828 7748
rect 28868 7708 28869 7748
rect 28827 7699 28869 7708
rect 29211 7748 29253 7757
rect 29211 7708 29212 7748
rect 29252 7708 29253 7748
rect 29211 7699 29253 7708
rect 29595 7748 29637 7757
rect 29595 7708 29596 7748
rect 29636 7708 29637 7748
rect 29595 7699 29637 7708
rect 32571 7748 32613 7757
rect 32571 7708 32572 7748
rect 32612 7708 32613 7748
rect 32571 7699 32613 7708
rect 36411 7748 36453 7757
rect 36411 7708 36412 7748
rect 36452 7708 36453 7748
rect 36411 7699 36453 7708
rect 39723 7748 39765 7757
rect 39723 7708 39724 7748
rect 39764 7708 39765 7748
rect 39723 7699 39765 7708
rect 41547 7748 41589 7757
rect 41547 7708 41548 7748
rect 41588 7708 41589 7748
rect 41547 7699 41589 7708
rect 43419 7748 43461 7757
rect 43419 7708 43420 7748
rect 43460 7708 43461 7748
rect 43419 7699 43461 7708
rect 45147 7748 45189 7757
rect 45147 7708 45148 7748
rect 45188 7708 45189 7748
rect 45147 7699 45189 7708
rect 1152 7580 45216 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 45216 7580
rect 1152 7516 45216 7540
rect 5979 7412 6021 7421
rect 5979 7372 5980 7412
rect 6020 7372 6021 7412
rect 5979 7363 6021 7372
rect 6298 7412 6356 7413
rect 6298 7372 6307 7412
rect 6347 7372 6356 7412
rect 6298 7371 6356 7372
rect 6795 7412 6837 7421
rect 6795 7372 6796 7412
rect 6836 7372 6837 7412
rect 6795 7363 6837 7372
rect 8506 7412 8564 7413
rect 8506 7372 8515 7412
rect 8555 7372 8564 7412
rect 8506 7371 8564 7372
rect 10810 7412 10868 7413
rect 10810 7372 10819 7412
rect 10859 7372 10868 7412
rect 10810 7371 10868 7372
rect 19275 7412 19317 7421
rect 19275 7372 19276 7412
rect 19316 7372 19317 7412
rect 19275 7363 19317 7372
rect 23691 7412 23733 7421
rect 23691 7372 23692 7412
rect 23732 7372 23733 7412
rect 23691 7363 23733 7372
rect 30219 7412 30261 7421
rect 30219 7372 30220 7412
rect 30260 7372 30261 7412
rect 30219 7363 30261 7372
rect 31947 7412 31989 7421
rect 31947 7372 31948 7412
rect 31988 7372 31989 7412
rect 31947 7363 31989 7372
rect 33147 7412 33189 7421
rect 33147 7372 33148 7412
rect 33188 7372 33189 7412
rect 33147 7363 33189 7372
rect 37083 7412 37125 7421
rect 37083 7372 37084 7412
rect 37124 7372 37125 7412
rect 37083 7363 37125 7372
rect 43995 7412 44037 7421
rect 43995 7372 43996 7412
rect 44036 7372 44037 7412
rect 43995 7363 44037 7372
rect 7083 7328 7125 7337
rect 7083 7288 7084 7328
rect 7124 7288 7125 7328
rect 7083 7279 7125 7288
rect 8619 7328 8661 7337
rect 8619 7288 8620 7328
rect 8660 7288 8661 7328
rect 8619 7279 8661 7288
rect 9867 7328 9909 7337
rect 27147 7328 27189 7337
rect 9867 7288 9868 7328
rect 9908 7288 9909 7328
rect 9867 7279 9909 7288
rect 10626 7319 10672 7328
rect 10626 7279 10627 7319
rect 10667 7279 10672 7319
rect 27147 7288 27148 7328
rect 27188 7288 27189 7328
rect 10626 7270 10672 7279
rect 21946 7277 22004 7282
rect 27147 7279 27189 7288
rect 2187 7244 2229 7253
rect 3819 7244 3861 7253
rect 6123 7244 6165 7253
rect 2187 7204 2188 7244
rect 2228 7204 2229 7244
rect 2187 7195 2229 7204
rect 3435 7235 3477 7244
rect 3435 7195 3436 7235
rect 3476 7195 3477 7235
rect 3819 7204 3820 7244
rect 3860 7204 3861 7244
rect 3819 7195 3861 7204
rect 5067 7235 5109 7244
rect 5067 7195 5068 7235
rect 5108 7195 5109 7235
rect 6123 7204 6124 7244
rect 6164 7204 6165 7244
rect 6123 7195 6165 7204
rect 6315 7244 6357 7253
rect 6315 7204 6316 7244
rect 6356 7204 6357 7244
rect 6315 7195 6357 7204
rect 6507 7244 6549 7253
rect 6507 7204 6508 7244
rect 6548 7204 6549 7244
rect 6507 7195 6549 7204
rect 6641 7244 6699 7245
rect 6641 7204 6650 7244
rect 6690 7204 6699 7244
rect 6641 7203 6699 7204
rect 7179 7244 7221 7253
rect 7179 7204 7180 7244
rect 7220 7204 7221 7244
rect 7179 7195 7221 7204
rect 7408 7244 7466 7245
rect 7408 7204 7417 7244
rect 7457 7204 7466 7244
rect 7408 7203 7466 7204
rect 7642 7244 7700 7245
rect 7642 7204 7651 7244
rect 7691 7204 7700 7244
rect 7642 7203 7700 7204
rect 8410 7244 8468 7245
rect 8410 7204 8419 7244
rect 8459 7204 8468 7244
rect 8410 7203 8468 7204
rect 8729 7244 8771 7253
rect 8729 7204 8730 7244
rect 8770 7204 8771 7244
rect 8729 7195 8771 7204
rect 9003 7244 9045 7253
rect 9232 7244 9290 7245
rect 9003 7204 9004 7244
rect 9044 7204 9045 7244
rect 9003 7195 9045 7204
rect 9138 7235 9184 7244
rect 9138 7195 9139 7235
rect 9179 7195 9184 7235
rect 9232 7204 9241 7244
rect 9281 7204 9290 7244
rect 9232 7203 9290 7204
rect 9483 7244 9525 7253
rect 9483 7204 9484 7244
rect 9524 7204 9525 7244
rect 9483 7195 9525 7204
rect 9754 7244 9812 7245
rect 9754 7204 9763 7244
rect 9803 7204 9812 7244
rect 9754 7203 9812 7204
rect 10330 7244 10388 7245
rect 10722 7244 10780 7245
rect 10330 7204 10339 7244
rect 10379 7204 10388 7244
rect 10330 7203 10388 7204
rect 10443 7235 10485 7244
rect 10443 7195 10444 7235
rect 10484 7195 10485 7235
rect 10722 7204 10731 7244
rect 10771 7204 10780 7244
rect 11062 7244 11104 7253
rect 10722 7203 10780 7204
rect 10848 7233 10890 7242
rect 3435 7186 3477 7195
rect 5067 7186 5109 7195
rect 9138 7186 9184 7195
rect 10443 7186 10485 7195
rect 10848 7193 10849 7233
rect 10889 7193 10890 7233
rect 11062 7204 11063 7244
rect 11103 7204 11104 7244
rect 11062 7195 11104 7204
rect 11307 7244 11349 7253
rect 11307 7204 11308 7244
rect 11348 7204 11349 7244
rect 11307 7195 11349 7204
rect 11595 7244 11637 7253
rect 13707 7244 13749 7253
rect 15531 7244 15573 7253
rect 17530 7244 17588 7245
rect 11595 7204 11596 7244
rect 11636 7204 11637 7244
rect 11595 7195 11637 7204
rect 12843 7235 12885 7244
rect 12843 7195 12844 7235
rect 12884 7195 12885 7235
rect 13707 7204 13708 7244
rect 13748 7204 13749 7244
rect 13707 7195 13749 7204
rect 14955 7235 14997 7244
rect 14955 7195 14956 7235
rect 14996 7195 14997 7235
rect 15531 7204 15532 7244
rect 15572 7204 15573 7244
rect 15531 7195 15573 7204
rect 16779 7235 16821 7244
rect 16779 7195 16780 7235
rect 16820 7195 16821 7235
rect 17530 7204 17539 7244
rect 17579 7204 17588 7244
rect 17530 7203 17588 7204
rect 17643 7244 17685 7253
rect 17643 7204 17644 7244
rect 17684 7204 17685 7244
rect 17643 7195 17685 7204
rect 18027 7244 18069 7253
rect 19546 7244 19604 7245
rect 18027 7204 18028 7244
rect 18068 7204 18069 7244
rect 18027 7195 18069 7204
rect 18603 7235 18645 7244
rect 18603 7195 18604 7235
rect 18644 7195 18645 7235
rect 10848 7184 10890 7193
rect 12843 7186 12885 7195
rect 14955 7186 14997 7195
rect 16779 7186 16821 7195
rect 18603 7186 18645 7195
rect 19083 7235 19125 7244
rect 19083 7195 19084 7235
rect 19124 7195 19125 7235
rect 19546 7204 19555 7244
rect 19595 7204 19604 7244
rect 19546 7203 19604 7204
rect 19659 7244 19701 7253
rect 19659 7204 19660 7244
rect 19700 7204 19701 7244
rect 19659 7195 19701 7204
rect 20043 7244 20085 7253
rect 20043 7204 20044 7244
rect 20084 7204 20085 7244
rect 20043 7195 20085 7204
rect 20619 7235 20661 7244
rect 20619 7195 20620 7235
rect 20660 7195 20661 7235
rect 19083 7186 19125 7195
rect 20619 7186 20661 7195
rect 21099 7235 21141 7244
rect 21946 7237 21955 7277
rect 21995 7237 22004 7277
rect 21946 7236 22004 7237
rect 22059 7244 22101 7253
rect 21099 7195 21100 7235
rect 21140 7195 21141 7235
rect 22059 7204 22060 7244
rect 22100 7204 22101 7244
rect 22059 7195 22101 7204
rect 22443 7244 22485 7253
rect 25515 7244 25557 7253
rect 28587 7244 28629 7253
rect 22443 7204 22444 7244
rect 22484 7204 22485 7244
rect 22443 7195 22485 7204
rect 23019 7235 23061 7244
rect 23019 7195 23020 7235
rect 23060 7195 23061 7235
rect 21099 7186 21141 7195
rect 23019 7186 23061 7195
rect 23499 7235 23541 7244
rect 23499 7195 23500 7235
rect 23540 7195 23541 7235
rect 23499 7186 23541 7195
rect 24267 7235 24309 7244
rect 24267 7195 24268 7235
rect 24308 7195 24309 7235
rect 25515 7204 25516 7244
rect 25556 7204 25557 7244
rect 25515 7195 25557 7204
rect 27339 7235 27381 7244
rect 27339 7195 27340 7235
rect 27380 7195 27381 7235
rect 28587 7204 28588 7244
rect 28628 7204 28629 7244
rect 28587 7195 28629 7204
rect 28779 7244 28821 7253
rect 30507 7244 30549 7253
rect 34731 7244 34773 7253
rect 39531 7244 39573 7253
rect 28779 7204 28780 7244
rect 28820 7204 28821 7244
rect 28779 7195 28821 7204
rect 30027 7235 30069 7244
rect 30027 7195 30028 7235
rect 30068 7195 30069 7235
rect 30507 7204 30508 7244
rect 30548 7204 30549 7244
rect 30507 7195 30549 7204
rect 31755 7235 31797 7244
rect 31755 7195 31756 7235
rect 31796 7195 31797 7235
rect 24267 7186 24309 7195
rect 27339 7186 27381 7195
rect 30027 7186 30069 7195
rect 31755 7186 31797 7195
rect 33483 7235 33525 7244
rect 33483 7195 33484 7235
rect 33524 7195 33525 7235
rect 34731 7204 34732 7244
rect 34772 7204 34773 7244
rect 34731 7195 34773 7204
rect 38283 7235 38325 7244
rect 38283 7195 38284 7235
rect 38324 7195 38325 7235
rect 39531 7204 39532 7244
rect 39572 7204 39573 7244
rect 39531 7195 39573 7204
rect 40282 7244 40340 7245
rect 40282 7204 40291 7244
rect 40331 7204 40340 7244
rect 40282 7203 40340 7204
rect 40395 7244 40437 7253
rect 40395 7204 40396 7244
rect 40436 7204 40437 7244
rect 40395 7195 40437 7204
rect 40779 7244 40821 7253
rect 40779 7204 40780 7244
rect 40820 7204 40821 7244
rect 40779 7195 40821 7204
rect 41355 7235 41397 7244
rect 41355 7195 41356 7235
rect 41396 7195 41397 7235
rect 33483 7186 33525 7195
rect 38283 7186 38325 7195
rect 41355 7186 41397 7195
rect 41835 7235 41877 7244
rect 41835 7195 41836 7235
rect 41876 7195 41877 7235
rect 41835 7186 41877 7195
rect 1227 7160 1269 7169
rect 1227 7120 1228 7160
rect 1268 7120 1269 7160
rect 1227 7111 1269 7120
rect 1611 7160 1653 7169
rect 1611 7120 1612 7160
rect 1652 7120 1653 7160
rect 1611 7111 1653 7120
rect 5739 7160 5781 7169
rect 5739 7120 5740 7160
rect 5780 7120 5781 7160
rect 5739 7111 5781 7120
rect 7298 7160 7340 7169
rect 7298 7120 7299 7160
rect 7339 7120 7340 7160
rect 7298 7111 7340 7120
rect 8043 7160 8085 7169
rect 8043 7120 8044 7160
rect 8084 7120 8085 7160
rect 8043 7111 8085 7120
rect 8283 7160 8325 7169
rect 8283 7120 8284 7160
rect 8324 7120 8325 7160
rect 8283 7111 8325 7120
rect 8907 7160 8949 7169
rect 8907 7120 8908 7160
rect 8948 7120 8949 7160
rect 8907 7111 8949 7120
rect 11194 7160 11252 7161
rect 11194 7120 11203 7160
rect 11243 7120 11252 7160
rect 11194 7119 11252 7120
rect 11403 7160 11445 7169
rect 11403 7120 11404 7160
rect 11444 7120 11445 7160
rect 11403 7111 11445 7120
rect 13323 7160 13365 7169
rect 13323 7120 13324 7160
rect 13364 7120 13365 7160
rect 13323 7111 13365 7120
rect 18123 7160 18165 7169
rect 18123 7120 18124 7160
rect 18164 7120 18165 7160
rect 18123 7111 18165 7120
rect 20139 7160 20181 7169
rect 20139 7120 20140 7160
rect 20180 7120 20181 7160
rect 20139 7111 20181 7120
rect 21322 7160 21380 7161
rect 21322 7120 21331 7160
rect 21371 7120 21380 7160
rect 21322 7119 21380 7120
rect 21483 7160 21525 7169
rect 21483 7120 21484 7160
rect 21524 7120 21525 7160
rect 21483 7111 21525 7120
rect 22539 7160 22581 7169
rect 22539 7120 22540 7160
rect 22580 7120 22581 7160
rect 22539 7111 22581 7120
rect 26187 7160 26229 7169
rect 26187 7120 26188 7160
rect 26228 7120 26229 7160
rect 26187 7111 26229 7120
rect 32331 7160 32373 7169
rect 32331 7120 32332 7160
rect 32372 7120 32373 7160
rect 32331 7111 32373 7120
rect 32715 7160 32757 7169
rect 32715 7120 32716 7160
rect 32756 7120 32757 7160
rect 32715 7111 32757 7120
rect 32907 7160 32949 7169
rect 32907 7120 32908 7160
rect 32948 7120 32949 7160
rect 32907 7111 32949 7120
rect 34923 7160 34965 7169
rect 34923 7120 34924 7160
rect 34964 7120 34965 7160
rect 34923 7111 34965 7120
rect 36459 7160 36501 7169
rect 36459 7120 36460 7160
rect 36500 7120 36501 7160
rect 36459 7111 36501 7120
rect 36843 7160 36885 7169
rect 36843 7120 36844 7160
rect 36884 7120 36885 7160
rect 36843 7111 36885 7120
rect 37419 7160 37461 7169
rect 37419 7120 37420 7160
rect 37460 7120 37461 7160
rect 37419 7111 37461 7120
rect 40011 7160 40053 7169
rect 40011 7120 40012 7160
rect 40052 7120 40053 7160
rect 40011 7111 40053 7120
rect 40875 7160 40917 7169
rect 40875 7120 40876 7160
rect 40916 7120 40917 7160
rect 40875 7111 40917 7120
rect 42058 7160 42116 7161
rect 42058 7120 42067 7160
rect 42107 7120 42116 7160
rect 42058 7119 42116 7120
rect 42411 7160 42453 7169
rect 42411 7120 42412 7160
rect 42452 7120 42453 7160
rect 42411 7111 42453 7120
rect 43371 7160 43413 7169
rect 43371 7120 43372 7160
rect 43412 7120 43413 7160
rect 43371 7111 43413 7120
rect 43755 7160 43797 7169
rect 43755 7120 43756 7160
rect 43796 7120 43797 7160
rect 43755 7111 43797 7120
rect 44139 7160 44181 7169
rect 44139 7120 44140 7160
rect 44180 7120 44181 7160
rect 44139 7111 44181 7120
rect 44523 7160 44565 7169
rect 44523 7120 44524 7160
rect 44564 7120 44565 7160
rect 44523 7111 44565 7120
rect 44907 7160 44949 7169
rect 44907 7120 44908 7160
rect 44948 7120 44949 7160
rect 44907 7111 44949 7120
rect 45147 7160 45189 7169
rect 45147 7120 45148 7160
rect 45188 7120 45189 7160
rect 45147 7111 45189 7120
rect 3627 7076 3669 7085
rect 3627 7036 3628 7076
rect 3668 7036 3669 7076
rect 3627 7027 3669 7036
rect 7622 7076 7664 7085
rect 7622 7036 7623 7076
rect 7663 7036 7664 7076
rect 7622 7027 7664 7036
rect 10155 7076 10197 7085
rect 10155 7036 10156 7076
rect 10196 7036 10197 7076
rect 10155 7027 10197 7036
rect 15147 7076 15189 7085
rect 15147 7036 15148 7076
rect 15188 7036 15189 7076
rect 15147 7027 15189 7036
rect 16971 7076 17013 7085
rect 16971 7036 16972 7076
rect 17012 7036 17013 7076
rect 16971 7027 17013 7036
rect 21723 7076 21765 7085
rect 21723 7036 21724 7076
rect 21764 7036 21765 7076
rect 21723 7027 21765 7036
rect 33291 7076 33333 7085
rect 33291 7036 33292 7076
rect 33332 7036 33333 7076
rect 33291 7027 33333 7036
rect 42171 7076 42213 7085
rect 42171 7036 42172 7076
rect 42212 7036 42213 7076
rect 42171 7027 42213 7036
rect 43611 7076 43653 7085
rect 43611 7036 43612 7076
rect 43652 7036 43653 7076
rect 43611 7027 43653 7036
rect 44379 7076 44421 7085
rect 44379 7036 44380 7076
rect 44420 7036 44421 7076
rect 44379 7027 44421 7036
rect 1467 6992 1509 7001
rect 1467 6952 1468 6992
rect 1508 6952 1509 6992
rect 1467 6943 1509 6952
rect 1851 6992 1893 7001
rect 1851 6952 1852 6992
rect 1892 6952 1893 6992
rect 1851 6943 1893 6952
rect 5259 6992 5301 7001
rect 5259 6952 5260 6992
rect 5300 6952 5301 6992
rect 5259 6943 5301 6952
rect 7834 6992 7892 6993
rect 7834 6952 7843 6992
rect 7883 6952 7892 6992
rect 7834 6951 7892 6952
rect 13035 6992 13077 7001
rect 13035 6952 13036 6992
rect 13076 6952 13077 6992
rect 13035 6943 13077 6952
rect 13563 6992 13605 7001
rect 13563 6952 13564 6992
rect 13604 6952 13605 6992
rect 13563 6943 13605 6952
rect 24075 6992 24117 7001
rect 24075 6952 24076 6992
rect 24116 6952 24117 6992
rect 24075 6943 24117 6952
rect 25947 6992 25989 7001
rect 25947 6952 25948 6992
rect 25988 6952 25989 6992
rect 25947 6943 25989 6952
rect 32091 6992 32133 7001
rect 32091 6952 32092 6992
rect 32132 6952 32133 6992
rect 32091 6943 32133 6952
rect 32475 6992 32517 7001
rect 32475 6952 32476 6992
rect 32516 6952 32517 6992
rect 32475 6943 32517 6952
rect 35163 6992 35205 7001
rect 35163 6952 35164 6992
rect 35204 6952 35205 6992
rect 35163 6943 35205 6952
rect 36699 6992 36741 7001
rect 36699 6952 36700 6992
rect 36740 6952 36741 6992
rect 36699 6943 36741 6952
rect 37179 6992 37221 7001
rect 37179 6952 37180 6992
rect 37220 6952 37221 6992
rect 37179 6943 37221 6952
rect 38091 6992 38133 7001
rect 38091 6952 38092 6992
rect 38132 6952 38133 6992
rect 38091 6943 38133 6952
rect 39771 6992 39813 7001
rect 39771 6952 39772 6992
rect 39812 6952 39813 6992
rect 39771 6943 39813 6952
rect 44763 6992 44805 7001
rect 44763 6952 44764 6992
rect 44804 6952 44805 6992
rect 44763 6943 44805 6952
rect 1152 6824 45216 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 45216 6824
rect 1152 6760 45216 6784
rect 6538 6656 6596 6657
rect 6538 6616 6547 6656
rect 6587 6616 6596 6656
rect 6538 6615 6596 6616
rect 8410 6656 8468 6657
rect 8410 6616 8419 6656
rect 8459 6616 8468 6656
rect 8410 6615 8468 6616
rect 16491 6656 16533 6665
rect 16491 6616 16492 6656
rect 16532 6616 16533 6656
rect 16491 6607 16533 6616
rect 23691 6656 23733 6665
rect 23691 6616 23692 6656
rect 23732 6616 23733 6656
rect 23691 6607 23733 6616
rect 26763 6656 26805 6665
rect 26763 6616 26764 6656
rect 26804 6616 26805 6656
rect 26763 6607 26805 6616
rect 28347 6656 28389 6665
rect 28347 6616 28348 6656
rect 28388 6616 28389 6656
rect 28347 6607 28389 6616
rect 29019 6656 29061 6665
rect 29019 6616 29020 6656
rect 29060 6616 29061 6656
rect 29019 6607 29061 6616
rect 30363 6656 30405 6665
rect 30363 6616 30364 6656
rect 30404 6616 30405 6656
rect 30363 6607 30405 6616
rect 40395 6656 40437 6665
rect 40395 6616 40396 6656
rect 40436 6616 40437 6656
rect 40395 6607 40437 6616
rect 44379 6656 44421 6665
rect 44379 6616 44380 6656
rect 44420 6616 44421 6656
rect 44379 6607 44421 6616
rect 1467 6572 1509 6581
rect 1467 6532 1468 6572
rect 1508 6532 1509 6572
rect 1467 6523 1509 6532
rect 7467 6572 7509 6581
rect 7467 6532 7468 6572
rect 7508 6532 7509 6572
rect 7467 6523 7509 6532
rect 17307 6572 17349 6581
rect 17307 6532 17308 6572
rect 17348 6532 17349 6572
rect 17307 6523 17349 6532
rect 20955 6572 20997 6581
rect 20955 6532 20956 6572
rect 20996 6532 20997 6572
rect 20955 6523 20997 6532
rect 40683 6572 40725 6581
rect 40683 6532 40684 6572
rect 40724 6532 40725 6572
rect 40683 6523 40725 6532
rect 1227 6488 1269 6497
rect 1227 6448 1228 6488
rect 1268 6448 1269 6488
rect 1227 6439 1269 6448
rect 1611 6488 1653 6497
rect 1611 6448 1612 6488
rect 1652 6448 1653 6488
rect 1611 6439 1653 6448
rect 1995 6488 2037 6497
rect 1995 6448 1996 6488
rect 2036 6448 2037 6488
rect 1995 6439 2037 6448
rect 4491 6488 4533 6497
rect 4491 6448 4492 6488
rect 4532 6448 4533 6488
rect 4491 6439 4533 6448
rect 5259 6488 5301 6497
rect 5259 6448 5260 6488
rect 5300 6448 5301 6488
rect 5259 6439 5301 6448
rect 9291 6488 9333 6497
rect 9291 6448 9292 6488
rect 9332 6448 9333 6488
rect 9291 6439 9333 6448
rect 9483 6488 9525 6497
rect 9483 6448 9484 6488
rect 9524 6448 9525 6488
rect 9483 6439 9525 6448
rect 10522 6488 10580 6489
rect 10522 6448 10531 6488
rect 10571 6448 10580 6488
rect 10522 6447 10580 6448
rect 10731 6488 10773 6497
rect 10731 6448 10732 6488
rect 10772 6448 10773 6488
rect 10731 6439 10773 6448
rect 16683 6488 16725 6497
rect 16683 6448 16684 6488
rect 16724 6448 16725 6488
rect 16683 6439 16725 6448
rect 17067 6488 17109 6497
rect 17067 6448 17068 6488
rect 17108 6448 17109 6488
rect 17067 6439 17109 6448
rect 17547 6488 17589 6497
rect 17547 6448 17548 6488
rect 17588 6448 17589 6488
rect 17547 6439 17589 6448
rect 17787 6488 17829 6497
rect 17787 6448 17788 6488
rect 17828 6448 17829 6488
rect 17787 6439 17829 6448
rect 18507 6488 18549 6497
rect 18507 6448 18508 6488
rect 18548 6448 18549 6488
rect 18507 6439 18549 6448
rect 19786 6488 19844 6489
rect 19786 6448 19795 6488
rect 19835 6448 19844 6488
rect 19786 6447 19844 6448
rect 19947 6488 19989 6497
rect 19947 6448 19948 6488
rect 19988 6448 19989 6488
rect 19947 6439 19989 6448
rect 20523 6488 20565 6497
rect 20523 6448 20524 6488
rect 20564 6448 20565 6488
rect 20523 6439 20565 6448
rect 20715 6488 20757 6497
rect 20715 6448 20716 6488
rect 20756 6448 20757 6488
rect 20715 6439 20757 6448
rect 21435 6488 21477 6497
rect 21435 6448 21436 6488
rect 21476 6448 21477 6488
rect 21435 6439 21477 6448
rect 21675 6488 21717 6497
rect 21675 6448 21676 6488
rect 21716 6448 21717 6488
rect 21675 6439 21717 6448
rect 21867 6488 21909 6497
rect 21867 6448 21868 6488
rect 21908 6448 21909 6488
rect 21867 6439 21909 6448
rect 25707 6488 25749 6497
rect 25707 6448 25708 6488
rect 25748 6448 25749 6488
rect 25707 6439 25749 6448
rect 28587 6488 28629 6497
rect 28587 6448 28588 6488
rect 28628 6448 28629 6488
rect 28587 6439 28629 6448
rect 28779 6488 28821 6497
rect 28779 6448 28780 6488
rect 28820 6448 28821 6488
rect 28779 6439 28821 6448
rect 29355 6488 29397 6497
rect 29355 6448 29356 6488
rect 29396 6448 29397 6488
rect 29355 6439 29397 6448
rect 29739 6488 29781 6497
rect 29739 6448 29740 6488
rect 29780 6448 29781 6488
rect 29739 6439 29781 6448
rect 30123 6488 30165 6497
rect 30123 6448 30124 6488
rect 30164 6448 30165 6488
rect 30123 6439 30165 6448
rect 38379 6488 38421 6497
rect 38379 6448 38380 6488
rect 38420 6448 38421 6488
rect 38379 6439 38421 6448
rect 44139 6488 44181 6497
rect 44139 6448 44140 6488
rect 44180 6448 44181 6488
rect 44139 6439 44181 6448
rect 44523 6488 44565 6497
rect 44523 6448 44524 6488
rect 44564 6448 44565 6488
rect 44523 6439 44565 6448
rect 44907 6488 44949 6497
rect 44907 6448 44908 6488
rect 44948 6448 44949 6488
rect 44907 6439 44949 6448
rect 45147 6488 45189 6497
rect 45147 6448 45148 6488
rect 45188 6448 45189 6488
rect 45147 6439 45189 6448
rect 7675 6415 7717 6424
rect 2667 6404 2709 6413
rect 2667 6364 2668 6404
rect 2708 6364 2709 6404
rect 2667 6355 2709 6364
rect 3907 6404 3965 6405
rect 3907 6364 3916 6404
rect 3956 6364 3965 6404
rect 3907 6363 3965 6364
rect 4762 6404 4820 6405
rect 4762 6364 4771 6404
rect 4811 6364 4820 6404
rect 4762 6363 4820 6364
rect 4875 6404 4917 6413
rect 4875 6364 4876 6404
rect 4916 6364 4917 6404
rect 4875 6355 4917 6364
rect 5355 6404 5397 6413
rect 5355 6364 5356 6404
rect 5396 6364 5397 6404
rect 5355 6355 5397 6364
rect 5827 6404 5885 6405
rect 5827 6364 5836 6404
rect 5876 6364 5885 6404
rect 5827 6363 5885 6364
rect 6346 6404 6404 6405
rect 6346 6364 6355 6404
rect 6395 6364 6404 6404
rect 6346 6363 6404 6364
rect 6795 6404 6837 6413
rect 6795 6364 6796 6404
rect 6836 6364 6837 6404
rect 6795 6355 6837 6364
rect 7066 6404 7124 6405
rect 7066 6364 7075 6404
rect 7115 6364 7124 6404
rect 7675 6375 7676 6415
rect 7716 6375 7717 6415
rect 7675 6366 7717 6375
rect 7834 6404 7892 6405
rect 7066 6363 7124 6364
rect 7834 6364 7843 6404
rect 7883 6364 7892 6404
rect 7834 6363 7892 6364
rect 7978 6404 8036 6405
rect 7978 6364 7987 6404
rect 8027 6364 8036 6404
rect 7978 6363 8036 6364
rect 8118 6404 8176 6405
rect 8118 6364 8127 6404
rect 8167 6364 8176 6404
rect 8118 6363 8176 6364
rect 8224 6404 8282 6405
rect 8224 6364 8233 6404
rect 8273 6364 8282 6404
rect 8224 6363 8282 6364
rect 8707 6404 8765 6405
rect 8707 6364 8716 6404
rect 8756 6364 8765 6404
rect 8707 6363 8765 6364
rect 9579 6404 9621 6413
rect 9579 6364 9580 6404
rect 9620 6364 9621 6404
rect 9579 6355 9621 6364
rect 9698 6404 9740 6413
rect 9698 6364 9699 6404
rect 9739 6364 9740 6404
rect 9698 6355 9740 6364
rect 9808 6404 9866 6405
rect 9808 6364 9817 6404
rect 9857 6364 9866 6404
rect 9808 6363 9866 6364
rect 10107 6404 10165 6405
rect 10107 6364 10116 6404
rect 10156 6364 10165 6404
rect 10107 6363 10165 6364
rect 10251 6404 10293 6413
rect 10251 6364 10252 6404
rect 10292 6364 10293 6404
rect 10251 6355 10293 6364
rect 10390 6404 10432 6413
rect 10390 6364 10391 6404
rect 10431 6364 10432 6404
rect 10390 6355 10432 6364
rect 10635 6404 10677 6413
rect 10635 6364 10636 6404
rect 10676 6364 10677 6404
rect 10635 6355 10677 6364
rect 10923 6404 10965 6413
rect 10923 6364 10924 6404
rect 10964 6364 10965 6404
rect 10923 6355 10965 6364
rect 11057 6404 11115 6405
rect 11057 6364 11066 6404
rect 11106 6364 11115 6404
rect 11057 6363 11115 6364
rect 11779 6404 11837 6405
rect 11779 6364 11788 6404
rect 11828 6364 11837 6404
rect 11779 6363 11837 6364
rect 13035 6404 13077 6413
rect 13035 6364 13036 6404
rect 13076 6364 13077 6404
rect 13035 6355 13077 6364
rect 13419 6404 13461 6413
rect 13419 6364 13420 6404
rect 13460 6364 13461 6404
rect 13419 6355 13461 6364
rect 14659 6404 14717 6405
rect 14659 6364 14668 6404
rect 14708 6364 14717 6404
rect 14659 6363 14717 6364
rect 15051 6404 15093 6413
rect 15051 6364 15052 6404
rect 15092 6364 15093 6404
rect 15051 6355 15093 6364
rect 16291 6404 16349 6405
rect 16291 6364 16300 6404
rect 16340 6364 16349 6404
rect 16291 6363 16349 6364
rect 18010 6404 18068 6405
rect 18010 6364 18019 6404
rect 18059 6364 18068 6404
rect 18010 6363 18068 6364
rect 18123 6404 18165 6413
rect 18123 6364 18124 6404
rect 18164 6364 18165 6404
rect 18123 6355 18165 6364
rect 18603 6404 18645 6413
rect 18603 6364 18604 6404
rect 18644 6364 18645 6404
rect 18603 6355 18645 6364
rect 19075 6404 19133 6405
rect 19075 6364 19084 6404
rect 19124 6364 19133 6404
rect 19075 6363 19133 6364
rect 19594 6404 19652 6405
rect 19594 6364 19603 6404
rect 19643 6364 19652 6404
rect 19594 6363 19652 6364
rect 22251 6404 22293 6413
rect 22251 6364 22252 6404
rect 22292 6364 22293 6404
rect 22251 6355 22293 6364
rect 23491 6404 23549 6405
rect 23491 6364 23500 6404
rect 23540 6364 23549 6404
rect 23491 6363 23549 6364
rect 26943 6404 27001 6405
rect 26943 6364 26952 6404
rect 26992 6364 27001 6404
rect 26943 6363 27001 6364
rect 28203 6404 28245 6413
rect 28203 6364 28204 6404
rect 28244 6364 28245 6404
rect 28203 6355 28245 6364
rect 30883 6404 30941 6405
rect 30883 6364 30892 6404
rect 30932 6364 30941 6404
rect 30883 6363 30941 6364
rect 32139 6404 32181 6413
rect 32139 6364 32140 6404
rect 32180 6364 32181 6404
rect 32139 6355 32181 6364
rect 32515 6404 32573 6405
rect 32515 6364 32524 6404
rect 32564 6364 32573 6404
rect 32515 6363 32573 6364
rect 33771 6404 33813 6413
rect 33771 6364 33772 6404
rect 33812 6364 33813 6404
rect 33771 6355 33813 6364
rect 33963 6404 34005 6413
rect 33963 6364 33964 6404
rect 34004 6364 34005 6404
rect 33963 6355 34005 6364
rect 35203 6404 35261 6405
rect 35203 6364 35212 6404
rect 35252 6364 35261 6404
rect 35203 6363 35261 6364
rect 35595 6404 35637 6413
rect 35595 6364 35596 6404
rect 35636 6364 35637 6404
rect 35595 6355 35637 6364
rect 36835 6404 36893 6405
rect 36835 6364 36844 6404
rect 36884 6364 36893 6404
rect 36835 6363 36893 6364
rect 38955 6404 38997 6413
rect 38955 6364 38956 6404
rect 38996 6364 38997 6404
rect 38955 6355 38997 6364
rect 40195 6404 40253 6405
rect 40195 6364 40204 6404
rect 40244 6364 40253 6404
rect 40195 6363 40253 6364
rect 4107 6320 4149 6329
rect 4107 6280 4108 6320
rect 4148 6280 4149 6320
rect 4107 6271 4149 6280
rect 7179 6320 7221 6329
rect 7179 6280 7180 6320
rect 7220 6280 7221 6320
rect 7179 6271 7221 6280
rect 8413 6320 8455 6329
rect 8413 6280 8414 6320
rect 8454 6280 8455 6320
rect 8413 6271 8455 6280
rect 9051 6320 9093 6329
rect 9051 6280 9052 6320
rect 9092 6280 9093 6320
rect 9051 6271 9093 6280
rect 16923 6320 16965 6329
rect 16923 6280 16924 6320
rect 16964 6280 16965 6320
rect 16923 6271 16965 6280
rect 20187 6320 20229 6329
rect 20187 6280 20188 6320
rect 20228 6280 20229 6320
rect 20187 6271 20229 6280
rect 22107 6320 22149 6329
rect 22107 6280 22108 6320
rect 22148 6280 22149 6320
rect 22107 6271 22149 6280
rect 29115 6320 29157 6329
rect 29115 6280 29116 6320
rect 29156 6280 29157 6320
rect 29115 6271 29157 6280
rect 1851 6236 1893 6245
rect 1851 6196 1852 6236
rect 1892 6196 1893 6236
rect 1851 6187 1893 6196
rect 2235 6236 2277 6245
rect 2235 6196 2236 6236
rect 2276 6196 2277 6236
rect 2235 6187 2277 6196
rect 4251 6236 4293 6245
rect 4251 6196 4252 6236
rect 4292 6196 4293 6236
rect 4251 6187 4293 6196
rect 7738 6236 7796 6237
rect 7738 6196 7747 6236
rect 7787 6196 7796 6236
rect 7738 6195 7796 6196
rect 8619 6236 8661 6245
rect 8619 6196 8620 6236
rect 8660 6196 8661 6236
rect 8619 6187 8661 6196
rect 9946 6236 10004 6237
rect 9946 6196 9955 6236
rect 9995 6196 10004 6236
rect 9946 6195 10004 6196
rect 11211 6236 11253 6245
rect 11211 6196 11212 6236
rect 11252 6196 11253 6236
rect 11211 6187 11253 6196
rect 11595 6236 11637 6245
rect 11595 6196 11596 6236
rect 11636 6196 11637 6236
rect 11595 6187 11637 6196
rect 14859 6236 14901 6245
rect 14859 6196 14860 6236
rect 14900 6196 14901 6236
rect 14859 6187 14901 6196
rect 20283 6236 20325 6245
rect 20283 6196 20284 6236
rect 20324 6196 20325 6236
rect 20283 6187 20325 6196
rect 25947 6236 25989 6245
rect 25947 6196 25948 6236
rect 25988 6196 25989 6236
rect 25947 6187 25989 6196
rect 29499 6236 29541 6245
rect 29499 6196 29500 6236
rect 29540 6196 29541 6236
rect 29499 6187 29541 6196
rect 30699 6236 30741 6245
rect 30699 6196 30700 6236
rect 30740 6196 30741 6236
rect 30699 6187 30741 6196
rect 32331 6236 32373 6245
rect 32331 6196 32332 6236
rect 32372 6196 32373 6236
rect 32331 6187 32373 6196
rect 35403 6236 35445 6245
rect 35403 6196 35404 6236
rect 35444 6196 35445 6236
rect 35403 6187 35445 6196
rect 37035 6236 37077 6245
rect 37035 6196 37036 6236
rect 37076 6196 37077 6236
rect 37035 6187 37077 6196
rect 38619 6236 38661 6245
rect 38619 6196 38620 6236
rect 38660 6196 38661 6236
rect 38619 6187 38661 6196
rect 44763 6236 44805 6245
rect 44763 6196 44764 6236
rect 44804 6196 44805 6236
rect 44763 6187 44805 6196
rect 1152 6068 45216 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 45216 6068
rect 1152 6004 45216 6028
rect 5355 5900 5397 5909
rect 5355 5860 5356 5900
rect 5396 5860 5397 5900
rect 5355 5851 5397 5860
rect 11691 5900 11733 5909
rect 11691 5860 11692 5900
rect 11732 5860 11733 5900
rect 11691 5851 11733 5860
rect 16971 5900 17013 5909
rect 16971 5860 16972 5900
rect 17012 5860 17013 5900
rect 16971 5851 17013 5860
rect 35595 5900 35637 5909
rect 35595 5860 35596 5900
rect 35636 5860 35637 5900
rect 35595 5851 35637 5860
rect 1467 5816 1509 5825
rect 1467 5776 1468 5816
rect 1508 5776 1509 5816
rect 1467 5767 1509 5776
rect 6843 5816 6885 5825
rect 6843 5776 6844 5816
rect 6884 5776 6885 5816
rect 6843 5767 6885 5776
rect 11115 5816 11157 5825
rect 11115 5776 11116 5816
rect 11156 5776 11157 5816
rect 11115 5767 11157 5776
rect 36459 5816 36501 5825
rect 36459 5776 36460 5816
rect 36500 5776 36501 5816
rect 36459 5767 36501 5776
rect 39706 5816 39764 5817
rect 39706 5776 39715 5816
rect 39755 5776 39764 5816
rect 39706 5775 39764 5776
rect 45147 5816 45189 5825
rect 45147 5776 45148 5816
rect 45188 5776 45189 5816
rect 45147 5767 45189 5776
rect 2283 5732 2325 5741
rect 3915 5732 3957 5741
rect 5643 5732 5685 5741
rect 2283 5692 2284 5732
rect 2324 5692 2325 5732
rect 2283 5683 2325 5692
rect 3531 5723 3573 5732
rect 3531 5683 3532 5723
rect 3572 5683 3573 5723
rect 3915 5692 3916 5732
rect 3956 5692 3957 5732
rect 3915 5683 3957 5692
rect 5163 5723 5205 5732
rect 5163 5683 5164 5723
rect 5204 5683 5205 5723
rect 5643 5692 5644 5732
rect 5684 5692 5685 5732
rect 5643 5683 5685 5692
rect 5874 5732 5916 5741
rect 5874 5692 5875 5732
rect 5915 5692 5916 5732
rect 5874 5683 5916 5692
rect 5986 5732 6044 5733
rect 5986 5692 5995 5732
rect 6035 5692 6044 5732
rect 5986 5691 6044 5692
rect 6219 5732 6261 5741
rect 6219 5692 6220 5732
rect 6260 5692 6261 5732
rect 6219 5683 6261 5692
rect 6507 5732 6549 5741
rect 6507 5692 6508 5732
rect 6548 5692 6549 5732
rect 6507 5683 6549 5692
rect 6646 5732 6688 5741
rect 6646 5692 6647 5732
rect 6687 5692 6688 5732
rect 6646 5683 6688 5692
rect 7162 5732 7220 5733
rect 8139 5732 8181 5741
rect 7162 5692 7171 5732
rect 7211 5692 7220 5732
rect 7162 5691 7220 5692
rect 7659 5723 7701 5732
rect 7659 5683 7660 5723
rect 7700 5683 7701 5723
rect 8139 5692 8140 5732
rect 8180 5692 8181 5732
rect 8139 5683 8181 5692
rect 8619 5732 8661 5741
rect 8619 5692 8620 5732
rect 8660 5692 8661 5732
rect 8619 5683 8661 5692
rect 8720 5732 8762 5741
rect 8720 5692 8721 5732
rect 8761 5692 8762 5732
rect 8720 5683 8762 5692
rect 10731 5732 10773 5741
rect 10731 5692 10732 5732
rect 10772 5692 10773 5732
rect 10731 5683 10773 5692
rect 10998 5732 11056 5733
rect 13131 5732 13173 5741
rect 10998 5692 11007 5732
rect 11047 5692 11056 5732
rect 10998 5691 11056 5692
rect 11883 5723 11925 5732
rect 11883 5683 11884 5723
rect 11924 5683 11925 5723
rect 13131 5692 13132 5732
rect 13172 5692 13173 5732
rect 13131 5683 13173 5692
rect 13323 5732 13365 5741
rect 15226 5732 15284 5733
rect 13323 5692 13324 5732
rect 13364 5692 13365 5732
rect 13323 5683 13365 5692
rect 14571 5723 14613 5732
rect 14571 5683 14572 5723
rect 14612 5683 14613 5723
rect 15226 5692 15235 5732
rect 15275 5692 15284 5732
rect 15226 5691 15284 5692
rect 15339 5732 15381 5741
rect 15339 5692 15340 5732
rect 15380 5692 15381 5732
rect 15339 5683 15381 5692
rect 15723 5732 15765 5741
rect 17163 5732 17205 5741
rect 18891 5732 18933 5741
rect 23403 5732 23445 5741
rect 15723 5692 15724 5732
rect 15764 5692 15765 5732
rect 15723 5683 15765 5692
rect 16299 5723 16341 5732
rect 16299 5683 16300 5723
rect 16340 5683 16341 5723
rect 3531 5674 3573 5683
rect 5163 5674 5205 5683
rect 7659 5674 7701 5683
rect 11883 5674 11925 5683
rect 14571 5674 14613 5683
rect 16299 5674 16341 5683
rect 16779 5723 16821 5732
rect 16779 5683 16780 5723
rect 16820 5683 16821 5723
rect 17163 5692 17164 5732
rect 17204 5692 17205 5732
rect 17163 5683 17205 5692
rect 18411 5723 18453 5732
rect 18411 5683 18412 5723
rect 18452 5683 18453 5723
rect 18891 5692 18892 5732
rect 18932 5692 18933 5732
rect 18891 5683 18933 5692
rect 22155 5723 22197 5732
rect 20139 5690 20197 5691
rect 16779 5674 16821 5683
rect 18411 5674 18453 5683
rect 1227 5648 1269 5657
rect 1227 5608 1228 5648
rect 1268 5608 1269 5648
rect 1227 5599 1269 5608
rect 1611 5648 1653 5657
rect 1611 5608 1612 5648
rect 1652 5608 1653 5648
rect 1611 5599 1653 5608
rect 5547 5648 5589 5657
rect 6106 5648 6164 5649
rect 5547 5608 5548 5648
rect 5588 5608 5589 5648
rect 5547 5599 5589 5608
rect 5778 5639 5824 5648
rect 5778 5599 5779 5639
rect 5819 5599 5824 5639
rect 6106 5608 6115 5648
rect 6155 5608 6164 5648
rect 6106 5607 6164 5608
rect 6315 5648 6357 5657
rect 6315 5608 6316 5648
rect 6356 5608 6357 5648
rect 6315 5599 6357 5608
rect 8235 5648 8277 5657
rect 8235 5608 8236 5648
rect 8276 5608 8277 5648
rect 8235 5599 8277 5608
rect 9291 5648 9333 5657
rect 9291 5608 9292 5648
rect 9332 5608 9333 5648
rect 9291 5599 9333 5608
rect 9483 5648 9525 5657
rect 9483 5608 9484 5648
rect 9524 5608 9525 5648
rect 9483 5599 9525 5608
rect 10059 5648 10101 5657
rect 10059 5608 10060 5648
rect 10100 5608 10101 5648
rect 10059 5599 10101 5608
rect 10491 5648 10533 5657
rect 10491 5608 10492 5648
rect 10532 5608 10533 5648
rect 10491 5599 10533 5608
rect 15819 5648 15861 5657
rect 20139 5650 20148 5690
rect 20188 5650 20197 5690
rect 22155 5683 22156 5723
rect 22196 5683 22197 5723
rect 23403 5692 23404 5732
rect 23444 5692 23445 5732
rect 23403 5683 23445 5692
rect 23595 5732 23637 5741
rect 25402 5732 25460 5733
rect 23595 5692 23596 5732
rect 23636 5692 23637 5732
rect 23595 5683 23637 5692
rect 24843 5723 24885 5732
rect 24843 5683 24844 5723
rect 24884 5683 24885 5723
rect 25402 5692 25411 5732
rect 25451 5692 25460 5732
rect 25402 5691 25460 5692
rect 25515 5732 25557 5741
rect 25515 5692 25516 5732
rect 25556 5692 25557 5732
rect 25515 5683 25557 5692
rect 25899 5732 25941 5741
rect 30586 5732 30644 5733
rect 25899 5692 25900 5732
rect 25940 5692 25941 5732
rect 25899 5683 25941 5692
rect 26475 5723 26517 5732
rect 26475 5683 26476 5723
rect 26516 5683 26517 5723
rect 22155 5674 22197 5683
rect 24843 5674 24885 5683
rect 26475 5674 26517 5683
rect 26955 5723 26997 5732
rect 26955 5683 26956 5723
rect 26996 5683 26997 5723
rect 30586 5692 30595 5732
rect 30635 5692 30644 5732
rect 30586 5691 30644 5692
rect 30699 5732 30741 5741
rect 30699 5692 30700 5732
rect 30740 5692 30741 5732
rect 30699 5683 30741 5692
rect 31083 5732 31125 5741
rect 33850 5732 33908 5733
rect 31083 5692 31084 5732
rect 31124 5692 31125 5732
rect 31083 5683 31125 5692
rect 31659 5723 31701 5732
rect 31659 5683 31660 5723
rect 31700 5683 31701 5723
rect 26955 5674 26997 5683
rect 31659 5674 31701 5683
rect 32139 5723 32181 5732
rect 32139 5683 32140 5723
rect 32180 5683 32181 5723
rect 33850 5692 33859 5732
rect 33899 5692 33908 5732
rect 33850 5691 33908 5692
rect 33963 5732 34005 5741
rect 33963 5692 33964 5732
rect 34004 5692 34005 5732
rect 33963 5683 34005 5692
rect 34347 5732 34389 5741
rect 36075 5732 36117 5741
rect 34347 5692 34348 5732
rect 34388 5692 34389 5732
rect 34347 5683 34389 5692
rect 34923 5723 34965 5732
rect 34923 5683 34924 5723
rect 34964 5683 34965 5723
rect 32139 5674 32181 5683
rect 34923 5674 34965 5683
rect 35403 5723 35445 5732
rect 35403 5683 35404 5723
rect 35444 5683 35445 5723
rect 36075 5692 36076 5732
rect 36116 5692 36117 5732
rect 36075 5683 36117 5692
rect 36346 5732 36404 5733
rect 36346 5692 36355 5732
rect 36395 5692 36404 5732
rect 36346 5691 36404 5692
rect 36939 5732 36981 5741
rect 40090 5732 40148 5733
rect 36939 5692 36940 5732
rect 36980 5692 36981 5732
rect 36939 5683 36981 5692
rect 38187 5723 38229 5732
rect 38187 5683 38188 5723
rect 38228 5683 38229 5723
rect 40090 5692 40099 5732
rect 40139 5692 40148 5732
rect 40090 5691 40148 5692
rect 35403 5674 35445 5683
rect 38187 5674 38229 5683
rect 20139 5649 20197 5650
rect 15819 5608 15820 5648
rect 15860 5608 15861 5648
rect 15819 5599 15861 5608
rect 20523 5648 20565 5657
rect 20523 5608 20524 5648
rect 20564 5608 20565 5648
rect 20523 5599 20565 5608
rect 21195 5648 21237 5657
rect 21195 5608 21196 5648
rect 21236 5608 21237 5648
rect 21195 5599 21237 5608
rect 21579 5648 21621 5657
rect 21579 5608 21580 5648
rect 21620 5608 21621 5648
rect 21579 5599 21621 5608
rect 21946 5648 22004 5649
rect 21946 5608 21955 5648
rect 21995 5608 22004 5648
rect 21946 5607 22004 5608
rect 25995 5648 26037 5657
rect 25995 5608 25996 5648
rect 26036 5608 26037 5648
rect 25995 5599 26037 5608
rect 27723 5648 27765 5657
rect 27723 5608 27724 5648
rect 27764 5608 27765 5648
rect 27723 5599 27765 5608
rect 27915 5648 27957 5657
rect 27915 5608 27916 5648
rect 27956 5608 27957 5648
rect 27915 5599 27957 5608
rect 28491 5648 28533 5657
rect 28491 5608 28492 5648
rect 28532 5608 28533 5648
rect 28491 5599 28533 5608
rect 28875 5648 28917 5657
rect 28875 5608 28876 5648
rect 28916 5608 28917 5648
rect 28875 5599 28917 5608
rect 29259 5648 29301 5657
rect 29259 5608 29260 5648
rect 29300 5608 29301 5648
rect 29259 5599 29301 5608
rect 29643 5648 29685 5657
rect 29643 5608 29644 5648
rect 29684 5608 29685 5648
rect 29643 5599 29685 5608
rect 30219 5648 30261 5657
rect 30219 5608 30220 5648
rect 30260 5608 30261 5648
rect 30219 5599 30261 5608
rect 31179 5648 31221 5657
rect 31179 5608 31180 5648
rect 31220 5608 31221 5648
rect 31179 5599 31221 5608
rect 32523 5648 32565 5657
rect 32523 5608 32524 5648
rect 32564 5608 32565 5648
rect 32523 5599 32565 5608
rect 33099 5648 33141 5657
rect 33099 5608 33100 5648
rect 33140 5608 33141 5648
rect 33099 5599 33141 5608
rect 33483 5648 33525 5657
rect 33483 5608 33484 5648
rect 33524 5608 33525 5648
rect 33483 5599 33525 5608
rect 34443 5648 34485 5657
rect 34443 5608 34444 5648
rect 34484 5608 34485 5648
rect 34443 5599 34485 5608
rect 38763 5648 38805 5657
rect 38763 5608 38764 5648
rect 38804 5608 38805 5648
rect 38763 5599 38805 5608
rect 38955 5648 38997 5657
rect 38955 5608 38956 5648
rect 38996 5608 38997 5648
rect 38955 5599 38997 5608
rect 44523 5648 44565 5657
rect 44523 5608 44524 5648
rect 44564 5608 44565 5648
rect 44523 5599 44565 5608
rect 44907 5648 44949 5657
rect 44907 5608 44908 5648
rect 44948 5608 44949 5648
rect 44907 5599 44949 5608
rect 5778 5590 5824 5599
rect 3723 5564 3765 5573
rect 3723 5524 3724 5564
rect 3764 5524 3765 5564
rect 3723 5515 3765 5524
rect 9723 5564 9765 5573
rect 9723 5524 9724 5564
rect 9764 5524 9765 5564
rect 9723 5515 9765 5524
rect 25035 5564 25077 5573
rect 25035 5524 25036 5564
rect 25076 5524 25077 5564
rect 25035 5515 25077 5524
rect 27195 5564 27237 5573
rect 27195 5524 27196 5564
rect 27236 5524 27237 5564
rect 27195 5515 27237 5524
rect 28155 5564 28197 5573
rect 28155 5524 28156 5564
rect 28196 5524 28197 5564
rect 28155 5515 28197 5524
rect 32379 5564 32421 5573
rect 32379 5524 32380 5564
rect 32420 5524 32421 5564
rect 32379 5515 32421 5524
rect 32859 5564 32901 5573
rect 32859 5524 32860 5564
rect 32900 5524 32901 5564
rect 32859 5515 32901 5524
rect 36747 5564 36789 5573
rect 36747 5524 36748 5564
rect 36788 5524 36789 5564
rect 36747 5515 36789 5524
rect 42027 5564 42069 5573
rect 42027 5524 42028 5564
rect 42068 5524 42069 5564
rect 42027 5515 42069 5524
rect 44763 5564 44805 5573
rect 44763 5524 44764 5564
rect 44804 5524 44805 5564
rect 44763 5515 44805 5524
rect 1851 5480 1893 5489
rect 1851 5440 1852 5480
rect 1892 5440 1893 5480
rect 1851 5431 1893 5440
rect 6939 5480 6981 5489
rect 6939 5440 6940 5480
rect 6980 5440 6981 5480
rect 6939 5431 6981 5440
rect 9051 5480 9093 5489
rect 9051 5440 9052 5480
rect 9092 5440 9093 5480
rect 9051 5431 9093 5440
rect 9819 5480 9861 5489
rect 9819 5440 9820 5480
rect 9860 5440 9861 5480
rect 9819 5431 9861 5440
rect 10203 5480 10245 5489
rect 10203 5440 10204 5480
rect 10244 5440 10245 5480
rect 10203 5431 10245 5440
rect 11403 5480 11445 5489
rect 11403 5440 11404 5480
rect 11444 5440 11445 5480
rect 11403 5431 11445 5440
rect 14763 5480 14805 5489
rect 14763 5440 14764 5480
rect 14804 5440 14805 5480
rect 14763 5431 14805 5440
rect 18603 5480 18645 5489
rect 18603 5440 18604 5480
rect 18644 5440 18645 5480
rect 18603 5431 18645 5440
rect 20331 5480 20373 5489
rect 20331 5440 20332 5480
rect 20372 5440 20373 5480
rect 20331 5431 20373 5440
rect 20763 5480 20805 5489
rect 20763 5440 20764 5480
rect 20804 5440 20805 5480
rect 20763 5431 20805 5440
rect 21435 5480 21477 5489
rect 21435 5440 21436 5480
rect 21476 5440 21477 5480
rect 21435 5431 21477 5440
rect 21819 5480 21861 5489
rect 21819 5440 21820 5480
rect 21860 5440 21861 5480
rect 21819 5431 21861 5440
rect 27483 5480 27525 5489
rect 27483 5440 27484 5480
rect 27524 5440 27525 5480
rect 27483 5431 27525 5440
rect 28251 5480 28293 5489
rect 28251 5440 28252 5480
rect 28292 5440 28293 5480
rect 28251 5431 28293 5440
rect 28635 5480 28677 5489
rect 28635 5440 28636 5480
rect 28676 5440 28677 5480
rect 28635 5431 28677 5440
rect 29019 5480 29061 5489
rect 29019 5440 29020 5480
rect 29060 5440 29061 5480
rect 29019 5431 29061 5440
rect 29403 5480 29445 5489
rect 29403 5440 29404 5480
rect 29444 5440 29445 5480
rect 29403 5431 29445 5440
rect 29979 5480 30021 5489
rect 29979 5440 29980 5480
rect 30020 5440 30021 5480
rect 29979 5431 30021 5440
rect 32763 5480 32805 5489
rect 32763 5440 32764 5480
rect 32804 5440 32805 5480
rect 32763 5431 32805 5440
rect 33243 5480 33285 5489
rect 33243 5440 33244 5480
rect 33284 5440 33285 5480
rect 33243 5431 33285 5440
rect 38379 5480 38421 5489
rect 38379 5440 38380 5480
rect 38420 5440 38421 5480
rect 38379 5431 38421 5440
rect 38523 5480 38565 5489
rect 38523 5440 38524 5480
rect 38564 5440 38565 5480
rect 38523 5431 38565 5440
rect 39195 5480 39237 5489
rect 39195 5440 39196 5480
rect 39236 5440 39237 5480
rect 39195 5431 39237 5440
rect 1152 5312 45216 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 45216 5312
rect 1152 5248 45216 5272
rect 1851 5144 1893 5153
rect 1851 5104 1852 5144
rect 1892 5104 1893 5144
rect 1851 5095 1893 5104
rect 3195 5144 3237 5153
rect 3195 5104 3196 5144
rect 3236 5104 3237 5144
rect 3195 5095 3237 5104
rect 5547 5144 5589 5153
rect 5547 5104 5548 5144
rect 5588 5104 5589 5144
rect 5547 5095 5589 5104
rect 6603 5144 6645 5153
rect 6603 5104 6604 5144
rect 6644 5104 6645 5144
rect 6603 5095 6645 5104
rect 11434 5144 11492 5145
rect 11434 5104 11443 5144
rect 11483 5104 11492 5144
rect 11434 5103 11492 5104
rect 12411 5144 12453 5153
rect 12411 5104 12412 5144
rect 12452 5104 12453 5144
rect 12411 5095 12453 5104
rect 26955 5144 26997 5153
rect 26955 5104 26956 5144
rect 26996 5104 26997 5144
rect 26955 5095 26997 5104
rect 30058 5144 30116 5145
rect 30058 5104 30067 5144
rect 30107 5104 30116 5144
rect 30058 5103 30116 5104
rect 31659 5144 31701 5153
rect 31659 5104 31660 5144
rect 31700 5104 31701 5144
rect 31659 5095 31701 5104
rect 34059 5144 34101 5153
rect 34059 5104 34060 5144
rect 34100 5104 34101 5144
rect 34059 5095 34101 5104
rect 39291 5144 39333 5153
rect 39291 5104 39292 5144
rect 39332 5104 39333 5144
rect 39291 5095 39333 5104
rect 45147 5144 45189 5153
rect 45147 5104 45148 5144
rect 45188 5104 45189 5144
rect 45147 5095 45189 5104
rect 18411 5060 18453 5069
rect 18411 5020 18412 5060
rect 18452 5020 18453 5060
rect 18411 5011 18453 5020
rect 23115 5060 23157 5069
rect 23115 5020 23116 5060
rect 23156 5020 23157 5060
rect 23115 5011 23157 5020
rect 1227 4976 1269 4985
rect 1227 4936 1228 4976
rect 1268 4936 1269 4976
rect 1227 4927 1269 4936
rect 1611 4976 1653 4985
rect 1611 4936 1612 4976
rect 1652 4936 1653 4976
rect 1611 4927 1653 4936
rect 2571 4976 2613 4985
rect 2571 4936 2572 4976
rect 2612 4936 2613 4976
rect 2571 4927 2613 4936
rect 2955 4976 2997 4985
rect 2955 4936 2956 4976
rect 2996 4936 2997 4976
rect 2955 4927 2997 4936
rect 6219 4976 6261 4985
rect 6219 4936 6220 4976
rect 6260 4936 6261 4976
rect 6219 4927 6261 4936
rect 8715 4976 8757 4985
rect 8715 4936 8716 4976
rect 8756 4936 8757 4976
rect 8715 4927 8757 4936
rect 10155 4976 10197 4985
rect 10155 4936 10156 4976
rect 10196 4936 10197 4976
rect 10155 4927 10197 4936
rect 11787 4976 11829 4985
rect 11787 4936 11788 4976
rect 11828 4936 11829 4976
rect 11787 4927 11829 4936
rect 12171 4976 12213 4985
rect 12171 4936 12172 4976
rect 12212 4936 12213 4976
rect 12171 4927 12213 4936
rect 13131 4976 13173 4985
rect 13131 4936 13132 4976
rect 13172 4936 13173 4976
rect 13131 4927 13173 4936
rect 15339 4976 15381 4985
rect 15339 4936 15340 4976
rect 15380 4936 15381 4976
rect 15339 4927 15381 4936
rect 19179 4976 19221 4985
rect 19179 4936 19180 4976
rect 19220 4936 19221 4976
rect 19179 4927 19221 4936
rect 23499 4976 23541 4985
rect 23499 4936 23500 4976
rect 23540 4936 23541 4976
rect 23499 4927 23541 4936
rect 27339 4976 27381 4985
rect 27339 4936 27340 4976
rect 27380 4936 27381 4976
rect 27339 4927 27381 4936
rect 27723 4976 27765 4985
rect 27723 4936 27724 4976
rect 27764 4936 27765 4976
rect 27723 4927 27765 4936
rect 28779 4976 28821 4985
rect 28779 4936 28780 4976
rect 28820 4936 28821 4976
rect 28779 4927 28821 4936
rect 32043 4976 32085 4985
rect 32043 4936 32044 4976
rect 32084 4936 32085 4976
rect 32043 4927 32085 4936
rect 32427 4976 32469 4985
rect 32427 4936 32428 4976
rect 32468 4936 32469 4976
rect 32427 4927 32469 4936
rect 36171 4976 36213 4985
rect 36171 4936 36172 4976
rect 36212 4936 36213 4976
rect 36171 4927 36213 4936
rect 36363 4976 36405 4985
rect 36363 4936 36364 4976
rect 36404 4936 36405 4976
rect 36363 4927 36405 4936
rect 36939 4976 36981 4985
rect 36939 4936 36940 4976
rect 36980 4936 36981 4976
rect 36939 4927 36981 4936
rect 37899 4976 37941 4985
rect 37899 4936 37900 4976
rect 37940 4936 37941 4976
rect 37899 4927 37941 4936
rect 39178 4976 39236 4977
rect 39178 4936 39187 4976
rect 39227 4936 39236 4976
rect 39178 4935 39236 4936
rect 39531 4976 39573 4985
rect 39531 4936 39532 4976
rect 39572 4936 39573 4976
rect 39531 4927 39573 4936
rect 44523 4976 44565 4985
rect 44523 4936 44524 4976
rect 44564 4936 44565 4976
rect 44523 4927 44565 4936
rect 44907 4976 44949 4985
rect 44907 4936 44908 4976
rect 44948 4936 44949 4976
rect 44907 4927 44949 4936
rect 3723 4892 3765 4901
rect 3723 4852 3724 4892
rect 3764 4852 3765 4892
rect 3723 4843 3765 4852
rect 3915 4892 3957 4901
rect 3915 4852 3916 4892
rect 3956 4852 3957 4892
rect 3915 4843 3957 4852
rect 4107 4892 4149 4901
rect 4107 4852 4108 4892
rect 4148 4852 4149 4892
rect 4107 4843 4149 4852
rect 5347 4892 5405 4893
rect 5347 4852 5356 4892
rect 5396 4852 5405 4892
rect 5347 4851 5405 4852
rect 5835 4892 5877 4901
rect 5835 4852 5836 4892
rect 5876 4852 5877 4892
rect 5835 4843 5877 4852
rect 5954 4892 5996 4901
rect 5954 4852 5955 4892
rect 5995 4852 5996 4892
rect 5954 4843 5996 4852
rect 6064 4892 6122 4893
rect 6064 4852 6073 4892
rect 6113 4852 6122 4892
rect 6064 4851 6122 4852
rect 6891 4892 6933 4901
rect 7275 4892 7317 4901
rect 6891 4852 6892 4892
rect 6932 4852 6933 4892
rect 6891 4843 6933 4852
rect 7026 4883 7072 4892
rect 7026 4843 7027 4883
rect 7067 4843 7072 4883
rect 7275 4852 7276 4892
rect 7316 4852 7317 4892
rect 7275 4843 7317 4852
rect 7738 4892 7796 4893
rect 7738 4852 7747 4892
rect 7787 4852 7796 4892
rect 7738 4851 7796 4852
rect 8227 4892 8285 4893
rect 8227 4852 8236 4892
rect 8276 4852 8285 4892
rect 8227 4851 8285 4852
rect 8811 4892 8853 4901
rect 8811 4852 8812 4892
rect 8852 4852 8853 4892
rect 8811 4843 8853 4852
rect 9195 4892 9237 4901
rect 9195 4852 9196 4892
rect 9236 4852 9237 4892
rect 9195 4843 9237 4852
rect 9296 4891 9338 4900
rect 9296 4851 9297 4891
rect 9337 4851 9338 4891
rect 9658 4892 9716 4893
rect 9658 4852 9667 4892
rect 9707 4852 9716 4892
rect 9658 4851 9716 4852
rect 9771 4892 9813 4901
rect 9771 4852 9772 4892
rect 9812 4852 9813 4892
rect 7026 4834 7072 4843
rect 9296 4842 9338 4851
rect 9771 4843 9813 4852
rect 10251 4892 10293 4901
rect 10251 4852 10252 4892
rect 10292 4852 10293 4892
rect 10251 4843 10293 4852
rect 10723 4892 10781 4893
rect 10723 4852 10732 4892
rect 10772 4852 10781 4892
rect 10723 4851 10781 4852
rect 11211 4892 11269 4893
rect 11211 4852 11220 4892
rect 11260 4852 11269 4892
rect 11211 4851 11269 4852
rect 12634 4892 12692 4893
rect 12634 4852 12643 4892
rect 12683 4852 12692 4892
rect 12634 4851 12692 4852
rect 12747 4892 12789 4901
rect 12747 4852 12748 4892
rect 12788 4852 12789 4892
rect 12747 4843 12789 4852
rect 13227 4892 13269 4901
rect 13227 4852 13228 4892
rect 13268 4852 13269 4892
rect 13227 4843 13269 4852
rect 13699 4892 13757 4893
rect 13699 4852 13708 4892
rect 13748 4852 13757 4892
rect 13699 4851 13757 4852
rect 14218 4892 14276 4893
rect 14218 4852 14227 4892
rect 14267 4852 14276 4892
rect 14218 4851 14276 4852
rect 14842 4892 14900 4893
rect 14842 4852 14851 4892
rect 14891 4852 14900 4892
rect 14842 4851 14900 4852
rect 14955 4892 14997 4901
rect 14955 4852 14956 4892
rect 14996 4852 14997 4892
rect 14955 4843 14997 4852
rect 15435 4892 15477 4901
rect 15435 4852 15436 4892
rect 15476 4852 15477 4892
rect 15435 4843 15477 4852
rect 15907 4892 15965 4893
rect 15907 4852 15916 4892
rect 15956 4852 15965 4892
rect 15907 4851 15965 4852
rect 16395 4892 16453 4893
rect 16395 4852 16404 4892
rect 16444 4852 16453 4892
rect 16395 4851 16453 4852
rect 16971 4892 17013 4901
rect 16971 4852 16972 4892
rect 17012 4852 17013 4892
rect 16971 4843 17013 4852
rect 18211 4892 18269 4893
rect 18211 4852 18220 4892
rect 18260 4852 18269 4892
rect 18211 4851 18269 4852
rect 18682 4892 18740 4893
rect 18682 4852 18691 4892
rect 18731 4852 18740 4892
rect 18682 4851 18740 4852
rect 18795 4892 18837 4901
rect 18795 4852 18796 4892
rect 18836 4852 18837 4892
rect 18795 4843 18837 4852
rect 19275 4892 19317 4901
rect 19275 4852 19276 4892
rect 19316 4852 19317 4892
rect 19275 4843 19317 4852
rect 19747 4892 19805 4893
rect 19747 4852 19756 4892
rect 19796 4852 19805 4892
rect 19747 4851 19805 4852
rect 20266 4892 20324 4893
rect 20266 4852 20275 4892
rect 20315 4852 20324 4892
rect 20266 4851 20324 4852
rect 20458 4892 20516 4893
rect 20458 4852 20467 4892
rect 20507 4852 20516 4892
rect 20458 4851 20516 4852
rect 20715 4892 20757 4901
rect 20715 4852 20716 4892
rect 20756 4852 20757 4892
rect 20715 4843 20757 4852
rect 21955 4892 22013 4893
rect 21955 4852 21964 4892
rect 22004 4852 22013 4892
rect 21955 4851 22013 4852
rect 22443 4892 22485 4901
rect 22443 4852 22444 4892
rect 22484 4852 22485 4892
rect 22443 4843 22485 4852
rect 22714 4892 22772 4893
rect 22714 4852 22723 4892
rect 22763 4852 22772 4892
rect 22714 4851 22772 4852
rect 23971 4892 24029 4893
rect 23971 4852 23980 4892
rect 24020 4852 24029 4892
rect 23971 4851 24029 4852
rect 25227 4892 25269 4901
rect 25227 4852 25228 4892
rect 25268 4852 25269 4892
rect 25227 4843 25269 4852
rect 25515 4892 25557 4901
rect 25515 4852 25516 4892
rect 25556 4852 25557 4892
rect 25515 4843 25557 4852
rect 26755 4892 26813 4893
rect 26755 4852 26764 4892
rect 26804 4852 26813 4892
rect 26755 4851 26813 4852
rect 28282 4892 28340 4893
rect 28282 4852 28291 4892
rect 28331 4852 28340 4892
rect 28282 4851 28340 4852
rect 28395 4892 28437 4901
rect 28395 4852 28396 4892
rect 28436 4852 28437 4892
rect 28395 4843 28437 4852
rect 28875 4892 28917 4901
rect 28875 4852 28876 4892
rect 28916 4852 28917 4892
rect 28875 4843 28917 4852
rect 29347 4892 29405 4893
rect 29347 4852 29356 4892
rect 29396 4852 29405 4892
rect 29347 4851 29405 4852
rect 29866 4892 29924 4893
rect 29866 4852 29875 4892
rect 29915 4852 29924 4892
rect 29866 4851 29924 4852
rect 30219 4892 30261 4901
rect 30219 4852 30220 4892
rect 30260 4852 30261 4892
rect 30219 4843 30261 4852
rect 31467 4892 31525 4893
rect 31467 4852 31476 4892
rect 31516 4852 31525 4892
rect 31467 4851 31525 4852
rect 32619 4892 32661 4901
rect 32619 4852 32620 4892
rect 32660 4852 32661 4892
rect 32619 4843 32661 4852
rect 33859 4892 33917 4893
rect 33859 4852 33868 4892
rect 33908 4852 33917 4892
rect 33859 4851 33917 4852
rect 34347 4892 34389 4901
rect 34347 4852 34348 4892
rect 34388 4852 34389 4892
rect 34347 4843 34389 4852
rect 35595 4892 35653 4893
rect 35595 4852 35604 4892
rect 35644 4852 35653 4892
rect 35595 4851 35653 4852
rect 37402 4892 37460 4893
rect 37402 4852 37411 4892
rect 37451 4852 37460 4892
rect 37402 4851 37460 4852
rect 37515 4892 37557 4901
rect 37515 4852 37516 4892
rect 37556 4852 37557 4892
rect 37515 4843 37557 4852
rect 37995 4892 38037 4901
rect 37995 4852 37996 4892
rect 38036 4852 38037 4892
rect 37995 4843 38037 4852
rect 38467 4892 38525 4893
rect 38467 4852 38476 4892
rect 38516 4852 38525 4892
rect 38467 4851 38525 4852
rect 38955 4892 39013 4893
rect 38955 4852 38964 4892
rect 39004 4852 39013 4892
rect 38955 4851 39013 4852
rect 40282 4892 40340 4893
rect 40282 4852 40291 4892
rect 40331 4852 40340 4892
rect 40282 4851 40340 4852
rect 7546 4808 7604 4809
rect 7546 4768 7555 4808
rect 7595 4768 7604 4808
rect 7546 4767 7604 4768
rect 22155 4808 22197 4817
rect 22155 4768 22156 4808
rect 22196 4768 22197 4808
rect 22155 4759 22197 4768
rect 22827 4808 22869 4817
rect 22827 4768 22828 4808
rect 22868 4768 22869 4808
rect 22827 4759 22869 4768
rect 23787 4808 23829 4817
rect 23787 4768 23788 4808
rect 23828 4768 23829 4808
rect 23787 4759 23829 4768
rect 32187 4808 32229 4817
rect 32187 4768 32188 4808
rect 32228 4768 32229 4808
rect 32187 4759 32229 4768
rect 35787 4808 35829 4817
rect 35787 4768 35788 4808
rect 35828 4768 35829 4808
rect 35787 4759 35829 4768
rect 36603 4808 36645 4817
rect 36603 4768 36604 4808
rect 36644 4768 36645 4808
rect 36603 4759 36645 4768
rect 39898 4808 39956 4809
rect 39898 4768 39907 4808
rect 39947 4768 39956 4808
rect 39898 4767 39956 4768
rect 44763 4808 44805 4817
rect 44763 4768 44764 4808
rect 44804 4768 44805 4808
rect 44763 4759 44805 4768
rect 1467 4724 1509 4733
rect 1467 4684 1468 4724
rect 1508 4684 1509 4724
rect 1467 4675 1509 4684
rect 2811 4724 2853 4733
rect 2811 4684 2812 4724
rect 2852 4684 2853 4724
rect 2811 4675 2853 4684
rect 3898 4724 3956 4725
rect 3898 4684 3907 4724
rect 3947 4684 3956 4724
rect 3898 4683 3956 4684
rect 5739 4724 5781 4733
rect 5739 4684 5740 4724
rect 5780 4684 5781 4724
rect 5739 4675 5781 4684
rect 6459 4724 6501 4733
rect 6459 4684 6460 4724
rect 6500 4684 6501 4724
rect 6459 4675 6501 4684
rect 12027 4724 12069 4733
rect 12027 4684 12028 4724
rect 12068 4684 12069 4724
rect 12027 4675 12069 4684
rect 14379 4724 14421 4733
rect 14379 4684 14380 4724
rect 14420 4684 14421 4724
rect 14379 4675 14421 4684
rect 16587 4724 16629 4733
rect 16587 4684 16588 4724
rect 16628 4684 16629 4724
rect 16587 4675 16629 4684
rect 23259 4724 23301 4733
rect 23259 4684 23260 4724
rect 23300 4684 23301 4724
rect 23259 4675 23301 4684
rect 27099 4724 27141 4733
rect 27099 4684 27100 4724
rect 27140 4684 27141 4724
rect 27099 4675 27141 4684
rect 27483 4724 27525 4733
rect 27483 4684 27484 4724
rect 27524 4684 27525 4724
rect 27483 4675 27525 4684
rect 31803 4724 31845 4733
rect 31803 4684 31804 4724
rect 31844 4684 31845 4724
rect 31803 4675 31845 4684
rect 35931 4724 35973 4733
rect 35931 4684 35932 4724
rect 35972 4684 35973 4724
rect 35931 4675 35973 4684
rect 36699 4724 36741 4733
rect 36699 4684 36700 4724
rect 36740 4684 36741 4724
rect 36699 4675 36741 4684
rect 42219 4724 42261 4733
rect 42219 4684 42220 4724
rect 42260 4684 42261 4724
rect 42219 4675 42261 4684
rect 1152 4556 45216 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 45216 4556
rect 1152 4492 45216 4516
rect 5818 4388 5876 4389
rect 5818 4348 5827 4388
rect 5867 4348 5876 4388
rect 5818 4347 5876 4348
rect 6490 4388 6548 4389
rect 6490 4348 6499 4388
rect 6539 4348 6548 4388
rect 6490 4347 6548 4348
rect 7275 4388 7317 4397
rect 7275 4348 7276 4388
rect 7316 4348 7317 4388
rect 7275 4339 7317 4348
rect 11307 4388 11349 4397
rect 11307 4348 11308 4388
rect 11348 4348 11349 4388
rect 11307 4339 11349 4348
rect 14667 4388 14709 4397
rect 14667 4348 14668 4388
rect 14708 4348 14709 4388
rect 14667 4339 14709 4348
rect 16299 4388 16341 4397
rect 16299 4348 16300 4388
rect 16340 4348 16341 4388
rect 16299 4339 16341 4348
rect 22971 4388 23013 4397
rect 22971 4348 22972 4388
rect 23012 4348 23013 4388
rect 22971 4339 23013 4348
rect 25659 4388 25701 4397
rect 25659 4348 25660 4388
rect 25700 4348 25701 4388
rect 25659 4339 25701 4348
rect 28107 4388 28149 4397
rect 28107 4348 28108 4388
rect 28148 4348 28149 4388
rect 28107 4339 28149 4348
rect 30027 4388 30069 4397
rect 30027 4348 30028 4388
rect 30068 4348 30069 4388
rect 30027 4339 30069 4348
rect 33003 4388 33045 4397
rect 33003 4348 33004 4388
rect 33044 4348 33045 4388
rect 33003 4339 33045 4348
rect 37899 4388 37941 4397
rect 37899 4348 37900 4388
rect 37940 4348 37941 4388
rect 37899 4339 37941 4348
rect 38043 4388 38085 4397
rect 38043 4348 38044 4388
rect 38084 4348 38085 4388
rect 38043 4339 38085 4348
rect 2523 4304 2565 4313
rect 2523 4264 2524 4304
rect 2564 4264 2565 4304
rect 2523 4255 2565 4264
rect 5259 4304 5301 4313
rect 5259 4264 5260 4304
rect 5300 4264 5301 4304
rect 5259 4255 5301 4264
rect 6106 4304 6164 4305
rect 6106 4264 6115 4304
rect 6155 4264 6164 4304
rect 6106 4263 6164 4264
rect 6219 4304 6261 4313
rect 6219 4264 6220 4304
rect 6260 4264 6261 4304
rect 6219 4255 6261 4264
rect 9322 4304 9380 4305
rect 9322 4264 9331 4304
rect 9371 4264 9380 4304
rect 9322 4263 9380 4264
rect 11931 4304 11973 4313
rect 11931 4264 11932 4304
rect 11972 4264 11973 4304
rect 11931 4255 11973 4264
rect 18027 4304 18069 4313
rect 18027 4264 18028 4304
rect 18068 4264 18069 4304
rect 18027 4255 18069 4264
rect 38427 4304 38469 4313
rect 38427 4264 38428 4304
rect 38468 4264 38469 4304
rect 38427 4255 38469 4264
rect 40155 4304 40197 4313
rect 40155 4264 40156 4304
rect 40196 4264 40197 4304
rect 40155 4255 40197 4264
rect 45147 4304 45189 4313
rect 45147 4264 45148 4304
rect 45188 4264 45189 4304
rect 45147 4255 45189 4264
rect 3051 4220 3093 4229
rect 5050 4220 5108 4221
rect 3051 4180 3052 4220
rect 3092 4180 3093 4220
rect 3051 4171 3093 4180
rect 4299 4211 4341 4220
rect 4299 4171 4300 4211
rect 4340 4171 4341 4211
rect 5050 4180 5059 4220
rect 5099 4180 5108 4220
rect 5050 4179 5108 4180
rect 5355 4220 5397 4229
rect 5355 4180 5356 4220
rect 5396 4180 5397 4220
rect 5355 4171 5397 4180
rect 5494 4220 5536 4229
rect 5494 4180 5495 4220
rect 5535 4180 5536 4220
rect 5494 4171 5536 4180
rect 5626 4220 5684 4221
rect 5626 4180 5635 4220
rect 5675 4180 5684 4220
rect 5626 4179 5684 4180
rect 5739 4220 5781 4229
rect 5739 4180 5740 4220
rect 5780 4180 5781 4220
rect 5739 4171 5781 4180
rect 6016 4220 6058 4229
rect 6651 4220 6709 4221
rect 6016 4180 6017 4220
rect 6057 4180 6058 4220
rect 6016 4171 6058 4180
rect 6315 4211 6357 4220
rect 6315 4171 6316 4211
rect 6356 4171 6357 4211
rect 6651 4180 6660 4220
rect 6700 4180 6709 4220
rect 6651 4179 6709 4180
rect 6795 4220 6837 4229
rect 6795 4180 6796 4220
rect 6836 4180 6837 4220
rect 6795 4171 6837 4180
rect 7018 4220 7076 4221
rect 7018 4180 7027 4220
rect 7067 4180 7076 4220
rect 7018 4179 7076 4180
rect 7121 4220 7179 4221
rect 7121 4180 7130 4220
rect 7170 4180 7179 4220
rect 7121 4179 7179 4180
rect 7546 4220 7604 4221
rect 7546 4180 7555 4220
rect 7595 4180 7604 4220
rect 7546 4179 7604 4180
rect 7659 4220 7701 4229
rect 7659 4180 7660 4220
rect 7700 4180 7701 4220
rect 7659 4171 7701 4180
rect 8043 4220 8085 4229
rect 9562 4220 9620 4221
rect 8043 4180 8044 4220
rect 8084 4180 8085 4220
rect 8043 4171 8085 4180
rect 8619 4211 8661 4220
rect 8619 4171 8620 4211
rect 8660 4171 8661 4211
rect 4299 4162 4341 4171
rect 6315 4162 6357 4171
rect 8619 4162 8661 4171
rect 9099 4211 9141 4220
rect 9099 4171 9100 4211
rect 9140 4171 9141 4211
rect 9562 4180 9571 4220
rect 9611 4180 9620 4220
rect 9562 4179 9620 4180
rect 9680 4220 9722 4229
rect 9680 4180 9681 4220
rect 9721 4180 9722 4220
rect 9680 4171 9722 4180
rect 10059 4220 10101 4229
rect 13227 4220 13269 4229
rect 14859 4220 14901 4229
rect 10059 4180 10060 4220
rect 10100 4180 10101 4220
rect 10059 4171 10101 4180
rect 10635 4211 10677 4220
rect 10635 4171 10636 4211
rect 10676 4171 10677 4211
rect 9099 4162 9141 4171
rect 10635 4162 10677 4171
rect 11115 4211 11157 4220
rect 11115 4171 11116 4211
rect 11156 4171 11157 4211
rect 13227 4180 13228 4220
rect 13268 4180 13269 4220
rect 13227 4171 13269 4180
rect 14475 4211 14517 4220
rect 14475 4171 14476 4211
rect 14516 4171 14517 4211
rect 14859 4180 14860 4220
rect 14900 4180 14901 4220
rect 16587 4220 16629 4229
rect 18586 4220 18644 4221
rect 14859 4171 14901 4180
rect 16107 4199 16149 4208
rect 11115 4162 11157 4171
rect 14475 4162 14517 4171
rect 16107 4159 16108 4199
rect 16148 4159 16149 4199
rect 16587 4180 16588 4220
rect 16628 4180 16629 4220
rect 16587 4171 16629 4180
rect 17835 4211 17877 4220
rect 17835 4171 17836 4211
rect 17876 4171 17877 4211
rect 18586 4180 18595 4220
rect 18635 4180 18644 4220
rect 18586 4179 18644 4180
rect 18699 4220 18741 4229
rect 18699 4180 18700 4220
rect 18740 4180 18741 4220
rect 18699 4171 18741 4180
rect 19083 4220 19125 4229
rect 20794 4220 20852 4221
rect 19083 4180 19084 4220
rect 19124 4180 19125 4220
rect 19083 4171 19125 4180
rect 19659 4211 19701 4220
rect 19659 4171 19660 4211
rect 19700 4171 19701 4211
rect 17835 4162 17877 4171
rect 19659 4162 19701 4171
rect 20139 4211 20181 4220
rect 20139 4171 20140 4211
rect 20180 4171 20181 4211
rect 20794 4180 20803 4220
rect 20843 4180 20852 4220
rect 20794 4179 20852 4180
rect 20907 4220 20949 4229
rect 20907 4180 20908 4220
rect 20948 4180 20949 4220
rect 20907 4171 20949 4180
rect 21291 4220 21333 4229
rect 22378 4220 22436 4221
rect 21291 4180 21292 4220
rect 21332 4180 21333 4220
rect 21291 4171 21333 4180
rect 21867 4211 21909 4220
rect 21867 4171 21868 4211
rect 21908 4171 21909 4211
rect 22378 4180 22387 4220
rect 22427 4180 22436 4220
rect 22378 4179 22436 4180
rect 22570 4220 22628 4221
rect 22570 4180 22579 4220
rect 22619 4180 22628 4220
rect 22570 4179 22628 4180
rect 26667 4220 26709 4229
rect 28587 4220 28629 4229
rect 31258 4220 31316 4221
rect 26667 4180 26668 4220
rect 26708 4180 26709 4220
rect 26667 4171 26709 4180
rect 27915 4211 27957 4220
rect 27915 4171 27916 4211
rect 27956 4171 27957 4211
rect 28587 4180 28588 4220
rect 28628 4180 28629 4220
rect 28587 4171 28629 4180
rect 29835 4211 29877 4220
rect 29835 4171 29836 4211
rect 29876 4171 29877 4211
rect 31258 4180 31267 4220
rect 31307 4180 31316 4220
rect 31258 4179 31316 4180
rect 31371 4220 31413 4229
rect 31371 4180 31372 4220
rect 31412 4180 31413 4220
rect 31371 4171 31413 4180
rect 31755 4220 31797 4229
rect 33750 4220 33808 4221
rect 31755 4180 31756 4220
rect 31796 4180 31797 4220
rect 31755 4171 31797 4180
rect 32331 4211 32373 4220
rect 32331 4171 32332 4211
rect 32372 4171 32373 4211
rect 20139 4162 20181 4171
rect 21867 4162 21909 4171
rect 27915 4162 27957 4171
rect 29835 4162 29877 4171
rect 32331 4162 32373 4171
rect 32811 4211 32853 4220
rect 32811 4171 32812 4211
rect 32852 4171 32853 4211
rect 33750 4180 33759 4220
rect 33799 4180 33808 4220
rect 33750 4179 33808 4180
rect 33867 4220 33909 4229
rect 33867 4180 33868 4220
rect 33908 4180 33909 4220
rect 33867 4171 33909 4180
rect 34251 4220 34293 4229
rect 36459 4220 36501 4229
rect 34251 4180 34252 4220
rect 34292 4180 34293 4220
rect 34251 4171 34293 4180
rect 34827 4211 34869 4220
rect 34827 4171 34828 4211
rect 34868 4171 34869 4211
rect 32811 4162 32853 4171
rect 34827 4162 34869 4171
rect 35307 4211 35349 4220
rect 35307 4171 35308 4211
rect 35348 4171 35349 4211
rect 36459 4180 36460 4220
rect 36500 4180 36501 4220
rect 36459 4171 36501 4180
rect 37707 4211 37749 4220
rect 37707 4171 37708 4211
rect 37748 4171 37749 4211
rect 35307 4162 35349 4171
rect 37707 4162 37749 4171
rect 16107 4150 16149 4159
rect 1227 4136 1269 4145
rect 1227 4096 1228 4136
rect 1268 4096 1269 4136
rect 1227 4087 1269 4096
rect 1611 4136 1653 4145
rect 1611 4096 1612 4136
rect 1652 4096 1653 4136
rect 1611 4087 1653 4096
rect 2283 4136 2325 4145
rect 2283 4096 2284 4136
rect 2324 4096 2325 4136
rect 2283 4087 2325 4096
rect 2667 4136 2709 4145
rect 2667 4096 2668 4136
rect 2708 4096 2709 4136
rect 2667 4087 2709 4096
rect 4683 4136 4725 4145
rect 4683 4096 4684 4136
rect 4724 4096 4725 4136
rect 4683 4087 4725 4096
rect 8139 4136 8181 4145
rect 8139 4096 8140 4136
rect 8180 4096 8181 4136
rect 8139 4087 8181 4096
rect 10155 4136 10197 4145
rect 10155 4096 10156 4136
rect 10196 4096 10197 4136
rect 10155 4087 10197 4096
rect 11691 4136 11733 4145
rect 11691 4096 11692 4136
rect 11732 4096 11733 4136
rect 11691 4087 11733 4096
rect 12075 4136 12117 4145
rect 12075 4096 12076 4136
rect 12116 4096 12117 4136
rect 12075 4087 12117 4096
rect 12459 4136 12501 4145
rect 12459 4096 12460 4136
rect 12500 4096 12501 4136
rect 12459 4087 12501 4096
rect 12874 4136 12932 4137
rect 12874 4096 12883 4136
rect 12923 4096 12932 4136
rect 12874 4095 12932 4096
rect 19179 4136 19221 4145
rect 19179 4096 19180 4136
rect 19220 4096 19221 4136
rect 19179 4087 19221 4096
rect 21387 4136 21429 4145
rect 21387 4096 21388 4136
rect 21428 4096 21429 4136
rect 21387 4087 21429 4096
rect 22731 4136 22773 4145
rect 22731 4096 22732 4136
rect 22772 4096 22773 4136
rect 22731 4087 22773 4096
rect 23307 4136 23349 4145
rect 23307 4096 23308 4136
rect 23348 4096 23349 4136
rect 23307 4087 23349 4096
rect 23787 4136 23829 4145
rect 23787 4096 23788 4136
rect 23828 4096 23829 4136
rect 23787 4087 23829 4096
rect 24171 4136 24213 4145
rect 24171 4096 24172 4136
rect 24212 4096 24213 4136
rect 24171 4087 24213 4096
rect 24843 4136 24885 4145
rect 24843 4096 24844 4136
rect 24884 4096 24885 4136
rect 24843 4087 24885 4096
rect 25035 4136 25077 4145
rect 25035 4096 25036 4136
rect 25076 4096 25077 4136
rect 25035 4087 25077 4096
rect 25419 4136 25461 4145
rect 25419 4096 25420 4136
rect 25460 4096 25461 4136
rect 25419 4087 25461 4096
rect 25995 4136 26037 4145
rect 25995 4096 25996 4136
rect 26036 4096 26037 4136
rect 25995 4087 26037 4096
rect 26379 4136 26421 4145
rect 26379 4096 26380 4136
rect 26420 4096 26421 4136
rect 26379 4087 26421 4096
rect 30411 4136 30453 4145
rect 30411 4096 30412 4136
rect 30452 4096 30453 4136
rect 30411 4087 30453 4096
rect 30795 4136 30837 4145
rect 30795 4096 30796 4136
rect 30836 4096 30837 4136
rect 30795 4087 30837 4096
rect 31851 4136 31893 4145
rect 31851 4096 31852 4136
rect 31892 4096 31893 4136
rect 31851 4087 31893 4096
rect 33387 4136 33429 4145
rect 33387 4096 33388 4136
rect 33428 4096 33429 4136
rect 33387 4087 33429 4096
rect 34347 4136 34389 4145
rect 34347 4096 34348 4136
rect 34388 4096 34389 4136
rect 34347 4087 34389 4096
rect 35883 4136 35925 4145
rect 35883 4096 35884 4136
rect 35924 4096 35925 4136
rect 35883 4087 35925 4096
rect 36267 4136 36309 4145
rect 36267 4096 36268 4136
rect 36308 4096 36309 4136
rect 36267 4087 36309 4096
rect 38283 4136 38325 4145
rect 38283 4096 38284 4136
rect 38324 4096 38325 4136
rect 38283 4087 38325 4096
rect 38667 4136 38709 4145
rect 38667 4096 38668 4136
rect 38708 4096 38709 4136
rect 38667 4087 38709 4096
rect 38859 4136 38901 4145
rect 38859 4096 38860 4136
rect 38900 4096 38901 4136
rect 38859 4087 38901 4096
rect 39723 4136 39765 4145
rect 39723 4096 39724 4136
rect 39764 4096 39765 4136
rect 39723 4087 39765 4096
rect 40395 4136 40437 4145
rect 40395 4096 40396 4136
rect 40436 4096 40437 4136
rect 40395 4087 40437 4096
rect 44139 4136 44181 4145
rect 44139 4096 44140 4136
rect 44180 4096 44181 4136
rect 44139 4087 44181 4096
rect 44523 4136 44565 4145
rect 44523 4096 44524 4136
rect 44564 4096 44565 4136
rect 44523 4087 44565 4096
rect 44907 4136 44949 4145
rect 44907 4096 44908 4136
rect 44948 4096 44949 4136
rect 44907 4087 44949 4096
rect 4491 4052 4533 4061
rect 4491 4012 4492 4052
rect 4532 4012 4533 4052
rect 4491 4003 4533 4012
rect 12315 4052 12357 4061
rect 12315 4012 12316 4052
rect 12356 4012 12357 4052
rect 12315 4003 12357 4012
rect 13083 4052 13125 4061
rect 13083 4012 13084 4052
rect 13124 4012 13125 4052
rect 13083 4003 13125 4012
rect 25275 4052 25317 4061
rect 25275 4012 25276 4052
rect 25316 4012 25317 4052
rect 25275 4003 25317 4012
rect 33147 4052 33189 4061
rect 33147 4012 33148 4052
rect 33188 4012 33189 4052
rect 33147 4003 33189 4012
rect 35547 4052 35589 4061
rect 35547 4012 35548 4052
rect 35588 4012 35589 4052
rect 35547 4003 35589 4012
rect 39099 4052 39141 4061
rect 39099 4012 39100 4052
rect 39140 4012 39141 4052
rect 39099 4003 39141 4012
rect 40971 4052 41013 4061
rect 40971 4012 40972 4052
rect 41012 4012 41013 4052
rect 40971 4003 41013 4012
rect 44763 4052 44805 4061
rect 44763 4012 44764 4052
rect 44804 4012 44805 4052
rect 44763 4003 44805 4012
rect 1467 3968 1509 3977
rect 1467 3928 1468 3968
rect 1508 3928 1509 3968
rect 1467 3919 1509 3928
rect 1851 3968 1893 3977
rect 1851 3928 1852 3968
rect 1892 3928 1893 3968
rect 1851 3919 1893 3928
rect 2907 3968 2949 3977
rect 2907 3928 2908 3968
rect 2948 3928 2949 3968
rect 2907 3919 2949 3928
rect 4923 3968 4965 3977
rect 4923 3928 4924 3968
rect 4964 3928 4965 3968
rect 4923 3919 4965 3928
rect 12699 3968 12741 3977
rect 12699 3928 12700 3968
rect 12740 3928 12741 3968
rect 12699 3919 12741 3928
rect 20362 3968 20420 3969
rect 20362 3928 20371 3968
rect 20411 3928 20420 3968
rect 20362 3927 20420 3928
rect 23067 3968 23109 3977
rect 23067 3928 23068 3968
rect 23108 3928 23109 3968
rect 23067 3919 23109 3928
rect 23547 3968 23589 3977
rect 23547 3928 23548 3968
rect 23588 3928 23589 3968
rect 23547 3919 23589 3928
rect 23931 3968 23973 3977
rect 23931 3928 23932 3968
rect 23972 3928 23973 3968
rect 23931 3919 23973 3928
rect 24603 3968 24645 3977
rect 24603 3928 24604 3968
rect 24644 3928 24645 3968
rect 24603 3919 24645 3928
rect 25755 3968 25797 3977
rect 25755 3928 25756 3968
rect 25796 3928 25797 3968
rect 25755 3919 25797 3928
rect 26139 3968 26181 3977
rect 26139 3928 26140 3968
rect 26180 3928 26181 3968
rect 26139 3919 26181 3928
rect 30171 3968 30213 3977
rect 30171 3928 30172 3968
rect 30212 3928 30213 3968
rect 30171 3919 30213 3928
rect 30555 3968 30597 3977
rect 30555 3928 30556 3968
rect 30596 3928 30597 3968
rect 30555 3919 30597 3928
rect 35643 3968 35685 3977
rect 35643 3928 35644 3968
rect 35684 3928 35685 3968
rect 35643 3919 35685 3928
rect 36027 3968 36069 3977
rect 36027 3928 36028 3968
rect 36068 3928 36069 3968
rect 36027 3919 36069 3928
rect 39963 3968 40005 3977
rect 39963 3928 39964 3968
rect 40004 3928 40005 3968
rect 39963 3919 40005 3928
rect 44379 3968 44421 3977
rect 44379 3928 44380 3968
rect 44420 3928 44421 3968
rect 44379 3919 44421 3928
rect 1152 3800 45216 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 45216 3800
rect 1152 3736 45216 3760
rect 3099 3632 3141 3641
rect 3099 3592 3100 3632
rect 3140 3592 3141 3632
rect 3099 3583 3141 3592
rect 8475 3632 8517 3641
rect 8475 3592 8476 3632
rect 8516 3592 8517 3632
rect 8475 3583 8517 3592
rect 9147 3632 9189 3641
rect 9147 3592 9148 3632
rect 9188 3592 9189 3632
rect 9147 3583 9189 3592
rect 9531 3632 9573 3641
rect 9531 3592 9532 3632
rect 9572 3592 9573 3632
rect 9531 3583 9573 3592
rect 19899 3632 19941 3641
rect 19899 3592 19900 3632
rect 19940 3592 19941 3632
rect 19899 3583 19941 3592
rect 23931 3632 23973 3641
rect 23931 3592 23932 3632
rect 23972 3592 23973 3632
rect 23931 3583 23973 3592
rect 32139 3632 32181 3641
rect 32139 3592 32140 3632
rect 32180 3592 32181 3632
rect 32139 3583 32181 3592
rect 33771 3632 33813 3641
rect 33771 3592 33772 3632
rect 33812 3592 33813 3632
rect 33771 3583 33813 3592
rect 35835 3632 35877 3641
rect 35835 3592 35836 3632
rect 35876 3592 35877 3632
rect 35835 3583 35877 3592
rect 36603 3632 36645 3641
rect 36603 3592 36604 3632
rect 36644 3592 36645 3632
rect 36603 3583 36645 3592
rect 39051 3632 39093 3641
rect 39051 3592 39052 3632
rect 39092 3592 39093 3632
rect 39051 3583 39093 3592
rect 45147 3632 45189 3641
rect 45147 3592 45148 3632
rect 45188 3592 45189 3632
rect 45147 3583 45189 3592
rect 15291 3548 15333 3557
rect 15291 3508 15292 3548
rect 15332 3508 15333 3548
rect 15291 3499 15333 3508
rect 18363 3548 18405 3557
rect 18363 3508 18364 3548
rect 18404 3508 18405 3548
rect 18363 3499 18405 3508
rect 26955 3548 26997 3557
rect 26955 3508 26956 3548
rect 26996 3508 26997 3548
rect 26955 3499 26997 3508
rect 37131 3548 37173 3557
rect 37131 3508 37132 3548
rect 37172 3508 37173 3548
rect 37131 3499 37173 3508
rect 41451 3548 41493 3557
rect 41451 3508 41452 3548
rect 41492 3508 41493 3548
rect 41451 3499 41493 3508
rect 1227 3464 1269 3473
rect 1227 3424 1228 3464
rect 1268 3424 1269 3464
rect 1227 3415 1269 3424
rect 1467 3464 1509 3473
rect 1467 3424 1468 3464
rect 1508 3424 1509 3464
rect 1467 3415 1509 3424
rect 1642 3464 1700 3465
rect 1642 3424 1651 3464
rect 1691 3424 1700 3464
rect 1642 3423 1700 3424
rect 1995 3464 2037 3473
rect 1995 3424 1996 3464
rect 2036 3424 2037 3464
rect 1995 3415 2037 3424
rect 2379 3464 2421 3473
rect 2379 3424 2380 3464
rect 2420 3424 2421 3464
rect 2379 3415 2421 3424
rect 2859 3464 2901 3473
rect 7083 3464 7125 3473
rect 2859 3424 2860 3464
rect 2900 3424 2901 3464
rect 2859 3415 2901 3424
rect 5202 3455 5248 3464
rect 5202 3415 5203 3455
rect 5243 3415 5248 3455
rect 5202 3406 5248 3415
rect 5682 3455 5728 3464
rect 5682 3415 5683 3455
rect 5723 3415 5728 3455
rect 7083 3424 7084 3464
rect 7124 3424 7125 3464
rect 7083 3415 7125 3424
rect 8139 3464 8181 3473
rect 8139 3424 8140 3464
rect 8180 3424 8181 3464
rect 8139 3415 8181 3424
rect 8715 3464 8757 3473
rect 8715 3424 8716 3464
rect 8756 3424 8757 3464
rect 8715 3415 8757 3424
rect 8907 3464 8949 3473
rect 8907 3424 8908 3464
rect 8948 3424 8949 3464
rect 8907 3415 8949 3424
rect 9291 3464 9333 3473
rect 9291 3424 9292 3464
rect 9332 3424 9333 3464
rect 9291 3415 9333 3424
rect 10827 3464 10869 3473
rect 10827 3424 10828 3464
rect 10868 3424 10869 3464
rect 10827 3415 10869 3424
rect 12267 3464 12309 3473
rect 12267 3424 12268 3464
rect 12308 3424 12309 3464
rect 12267 3415 12309 3424
rect 13899 3464 13941 3473
rect 13899 3424 13900 3464
rect 13940 3424 13941 3464
rect 13899 3415 13941 3424
rect 14283 3464 14325 3473
rect 14283 3424 14284 3464
rect 14324 3424 14325 3464
rect 14283 3415 14325 3424
rect 14667 3464 14709 3473
rect 14667 3424 14668 3464
rect 14708 3424 14709 3464
rect 14667 3415 14709 3424
rect 15051 3464 15093 3473
rect 15051 3424 15052 3464
rect 15092 3424 15093 3464
rect 15051 3415 15093 3424
rect 17355 3464 17397 3473
rect 17355 3424 17356 3464
rect 17396 3424 17397 3464
rect 17355 3415 17397 3424
rect 17931 3464 17973 3473
rect 17931 3424 17932 3464
rect 17972 3424 17973 3464
rect 17931 3415 17973 3424
rect 18123 3464 18165 3473
rect 18123 3424 18124 3464
rect 18164 3424 18165 3464
rect 18123 3415 18165 3424
rect 18507 3464 18549 3473
rect 18507 3424 18508 3464
rect 18548 3424 18549 3464
rect 18507 3415 18549 3424
rect 18891 3464 18933 3473
rect 18891 3424 18892 3464
rect 18932 3424 18933 3464
rect 18891 3415 18933 3424
rect 19306 3464 19364 3465
rect 19306 3424 19315 3464
rect 19355 3424 19364 3464
rect 19306 3423 19364 3424
rect 19659 3464 19701 3473
rect 19659 3424 19660 3464
rect 19700 3424 19701 3464
rect 19659 3415 19701 3424
rect 20043 3464 20085 3473
rect 20043 3424 20044 3464
rect 20084 3424 20085 3464
rect 20043 3415 20085 3424
rect 23691 3464 23733 3473
rect 23691 3424 23692 3464
rect 23732 3424 23733 3464
rect 23691 3415 23733 3424
rect 24555 3464 24597 3473
rect 24555 3424 24556 3464
rect 24596 3424 24597 3464
rect 24555 3415 24597 3424
rect 26667 3464 26709 3473
rect 26667 3424 26668 3464
rect 26708 3424 26709 3464
rect 26667 3415 26709 3424
rect 28779 3464 28821 3473
rect 28779 3424 28780 3464
rect 28820 3424 28821 3464
rect 28779 3415 28821 3424
rect 36075 3464 36117 3473
rect 36075 3424 36076 3464
rect 36116 3424 36117 3464
rect 36075 3415 36117 3424
rect 36459 3464 36501 3473
rect 36459 3424 36460 3464
rect 36500 3424 36501 3464
rect 36459 3415 36501 3424
rect 36843 3464 36885 3473
rect 36843 3424 36844 3464
rect 36884 3424 36885 3464
rect 36843 3415 36885 3424
rect 41595 3464 41637 3473
rect 41595 3424 41596 3464
rect 41636 3424 41637 3464
rect 41595 3415 41637 3424
rect 41835 3464 41877 3473
rect 41835 3424 41836 3464
rect 41876 3424 41877 3464
rect 41835 3415 41877 3424
rect 44523 3464 44565 3473
rect 44523 3424 44524 3464
rect 44564 3424 44565 3464
rect 44523 3415 44565 3424
rect 44907 3464 44949 3473
rect 44907 3424 44908 3464
rect 44948 3424 44949 3464
rect 44907 3415 44949 3424
rect 5682 3406 5728 3415
rect 3243 3380 3285 3389
rect 3243 3340 3244 3380
rect 3284 3340 3285 3380
rect 3243 3331 3285 3340
rect 4483 3380 4541 3381
rect 4483 3340 4492 3380
rect 4532 3340 4541 3380
rect 4483 3339 4541 3340
rect 5067 3380 5109 3389
rect 5067 3340 5068 3380
rect 5108 3340 5109 3380
rect 5067 3331 5109 3340
rect 5296 3380 5354 3381
rect 5296 3340 5305 3380
rect 5345 3340 5354 3380
rect 5296 3339 5354 3340
rect 5547 3380 5589 3389
rect 5547 3340 5548 3380
rect 5588 3340 5589 3380
rect 5547 3331 5589 3340
rect 5776 3380 5834 3381
rect 5776 3340 5785 3380
rect 5825 3340 5834 3380
rect 5776 3339 5834 3340
rect 6106 3380 6164 3381
rect 6106 3340 6115 3380
rect 6155 3340 6164 3380
rect 6106 3339 6164 3340
rect 6595 3380 6653 3381
rect 6595 3340 6604 3380
rect 6644 3340 6653 3380
rect 6595 3339 6653 3340
rect 7179 3380 7221 3389
rect 7179 3340 7180 3380
rect 7220 3340 7221 3380
rect 7179 3331 7221 3340
rect 7563 3380 7605 3389
rect 7563 3340 7564 3380
rect 7604 3340 7605 3380
rect 7563 3331 7605 3340
rect 7673 3380 7731 3381
rect 7673 3340 7682 3380
rect 7722 3340 7731 3380
rect 7673 3339 7731 3340
rect 9850 3380 9908 3381
rect 9850 3340 9859 3380
rect 9899 3340 9908 3380
rect 9850 3339 9908 3340
rect 10339 3380 10397 3381
rect 10339 3340 10348 3380
rect 10388 3340 10397 3380
rect 10339 3339 10397 3340
rect 10923 3380 10965 3389
rect 10923 3340 10924 3380
rect 10964 3340 10965 3380
rect 10923 3331 10965 3340
rect 11307 3380 11349 3389
rect 11307 3340 11308 3380
rect 11348 3340 11349 3380
rect 11307 3331 11349 3340
rect 11417 3380 11475 3381
rect 11417 3340 11426 3380
rect 11466 3340 11475 3380
rect 11417 3339 11475 3340
rect 11770 3380 11828 3381
rect 11770 3340 11779 3380
rect 11819 3340 11828 3380
rect 11770 3339 11828 3340
rect 11883 3380 11925 3389
rect 11883 3340 11884 3380
rect 11924 3340 11925 3380
rect 11883 3331 11925 3340
rect 12363 3380 12405 3389
rect 12363 3340 12364 3380
rect 12404 3340 12405 3380
rect 12363 3331 12405 3340
rect 12835 3380 12893 3381
rect 12835 3340 12844 3380
rect 12884 3340 12893 3380
rect 12835 3339 12893 3340
rect 13354 3380 13412 3381
rect 13354 3340 13363 3380
rect 13403 3340 13412 3380
rect 13354 3339 13412 3340
rect 15435 3380 15477 3389
rect 15435 3340 15436 3380
rect 15476 3340 15477 3380
rect 15435 3331 15477 3340
rect 16675 3380 16733 3381
rect 16675 3340 16684 3380
rect 16724 3340 16733 3380
rect 16675 3339 16733 3340
rect 20427 3380 20469 3389
rect 20427 3340 20428 3380
rect 20468 3340 20469 3380
rect 20427 3331 20469 3340
rect 21667 3380 21725 3381
rect 21667 3340 21676 3380
rect 21716 3340 21725 3380
rect 21667 3339 21725 3340
rect 22059 3380 22101 3389
rect 22059 3340 22060 3380
rect 22100 3340 22101 3380
rect 22059 3331 22101 3340
rect 23299 3380 23357 3381
rect 23299 3340 23308 3380
rect 23348 3340 23357 3380
rect 23299 3339 23357 3340
rect 24843 3380 24885 3389
rect 24843 3340 24844 3380
rect 24884 3340 24885 3380
rect 24843 3331 24885 3340
rect 26083 3380 26141 3381
rect 26083 3340 26092 3380
rect 26132 3340 26141 3380
rect 26083 3339 26141 3340
rect 27139 3380 27197 3381
rect 27139 3340 27148 3380
rect 27188 3340 27197 3380
rect 27139 3339 27197 3340
rect 28395 3380 28437 3389
rect 28395 3340 28396 3380
rect 28436 3340 28437 3380
rect 28395 3331 28437 3340
rect 29067 3380 29109 3389
rect 29067 3340 29068 3380
rect 29108 3340 29109 3380
rect 29067 3331 29109 3340
rect 30307 3380 30365 3381
rect 30307 3340 30316 3380
rect 30356 3340 30365 3380
rect 30307 3339 30365 3340
rect 30699 3380 30741 3389
rect 30699 3340 30700 3380
rect 30740 3340 30741 3380
rect 30699 3331 30741 3340
rect 31939 3380 31997 3381
rect 31939 3340 31948 3380
rect 31988 3340 31997 3380
rect 31939 3339 31997 3340
rect 32331 3380 32373 3389
rect 32331 3340 32332 3380
rect 32372 3340 32373 3380
rect 32331 3331 32373 3340
rect 33571 3380 33629 3381
rect 33571 3340 33580 3380
rect 33620 3340 33629 3380
rect 33571 3339 33629 3340
rect 34275 3380 34333 3381
rect 34275 3340 34284 3380
rect 34324 3340 34333 3380
rect 34275 3339 34333 3340
rect 35491 3380 35549 3381
rect 35491 3340 35500 3380
rect 35540 3340 35549 3380
rect 35491 3339 35549 3340
rect 37315 3380 37373 3381
rect 37315 3340 37324 3380
rect 37364 3340 37373 3380
rect 37315 3339 37373 3340
rect 38571 3380 38613 3389
rect 38571 3340 38572 3380
rect 38612 3340 38613 3380
rect 38571 3331 38613 3340
rect 39235 3380 39293 3381
rect 39235 3340 39244 3380
rect 39284 3340 39293 3380
rect 39235 3339 39293 3340
rect 40491 3380 40533 3389
rect 40491 3340 40492 3380
rect 40532 3340 40533 3380
rect 40491 3331 40533 3340
rect 40779 3380 40821 3389
rect 40779 3340 40780 3380
rect 40820 3340 40821 3380
rect 40779 3331 40821 3340
rect 41050 3380 41108 3381
rect 41050 3340 41059 3380
rect 41099 3340 41108 3380
rect 41050 3339 41108 3340
rect 1851 3296 1893 3305
rect 1851 3256 1852 3296
rect 1892 3256 1893 3296
rect 1851 3247 1893 3256
rect 2619 3296 2661 3305
rect 2619 3256 2620 3296
rect 2660 3256 2661 3296
rect 2619 3247 2661 3256
rect 4683 3296 4725 3305
rect 4683 3256 4684 3296
rect 4724 3256 4725 3296
rect 4683 3247 4725 3256
rect 5451 3296 5493 3305
rect 5451 3256 5452 3296
rect 5492 3256 5493 3296
rect 5451 3247 5493 3256
rect 8379 3296 8421 3305
rect 8379 3256 8380 3296
rect 8420 3256 8421 3296
rect 8379 3247 8421 3256
rect 9658 3296 9716 3297
rect 9658 3256 9667 3296
rect 9707 3256 9716 3296
rect 9658 3255 9716 3256
rect 17595 3296 17637 3305
rect 17595 3256 17596 3296
rect 17636 3256 17637 3296
rect 17595 3247 17637 3256
rect 23499 3296 23541 3305
rect 23499 3256 23500 3296
rect 23540 3256 23541 3296
rect 23499 3247 23541 3256
rect 41163 3296 41205 3305
rect 41163 3256 41164 3296
rect 41204 3256 41205 3296
rect 41163 3247 41205 3256
rect 2235 3212 2277 3221
rect 2235 3172 2236 3212
rect 2276 3172 2277 3212
rect 2235 3163 2277 3172
rect 4971 3212 5013 3221
rect 4971 3172 4972 3212
rect 5012 3172 5013 3212
rect 4971 3163 5013 3172
rect 5931 3212 5973 3221
rect 5931 3172 5932 3212
rect 5972 3172 5973 3212
rect 5931 3163 5973 3172
rect 13515 3212 13557 3221
rect 13515 3172 13516 3212
rect 13556 3172 13557 3212
rect 13515 3163 13557 3172
rect 14139 3212 14181 3221
rect 14139 3172 14140 3212
rect 14180 3172 14181 3212
rect 14139 3163 14181 3172
rect 14523 3212 14565 3221
rect 14523 3172 14524 3212
rect 14564 3172 14565 3212
rect 14523 3163 14565 3172
rect 14907 3212 14949 3221
rect 14907 3172 14908 3212
rect 14948 3172 14949 3212
rect 14907 3163 14949 3172
rect 16875 3212 16917 3221
rect 16875 3172 16876 3212
rect 16916 3172 16917 3212
rect 16875 3163 16917 3172
rect 17691 3212 17733 3221
rect 17691 3172 17692 3212
rect 17732 3172 17733 3212
rect 17691 3163 17733 3172
rect 18747 3212 18789 3221
rect 18747 3172 18748 3212
rect 18788 3172 18789 3212
rect 18747 3163 18789 3172
rect 19131 3212 19173 3221
rect 19131 3172 19132 3212
rect 19172 3172 19173 3212
rect 19131 3163 19173 3172
rect 19515 3212 19557 3221
rect 19515 3172 19516 3212
rect 19556 3172 19557 3212
rect 19515 3163 19557 3172
rect 20283 3212 20325 3221
rect 20283 3172 20284 3212
rect 20324 3172 20325 3212
rect 20283 3163 20325 3172
rect 21867 3212 21909 3221
rect 21867 3172 21868 3212
rect 21908 3172 21909 3212
rect 21867 3163 21909 3172
rect 24315 3212 24357 3221
rect 24315 3172 24316 3212
rect 24356 3172 24357 3212
rect 24315 3163 24357 3172
rect 26283 3212 26325 3221
rect 26283 3172 26284 3212
rect 26324 3172 26325 3212
rect 26283 3163 26325 3172
rect 26427 3212 26469 3221
rect 26427 3172 26428 3212
rect 26468 3172 26469 3212
rect 26427 3163 26469 3172
rect 28539 3212 28581 3221
rect 28539 3172 28540 3212
rect 28580 3172 28581 3212
rect 28539 3163 28581 3172
rect 30507 3212 30549 3221
rect 30507 3172 30508 3212
rect 30548 3172 30549 3212
rect 30507 3163 30549 3172
rect 35691 3212 35733 3221
rect 35691 3172 35692 3212
rect 35732 3172 35733 3212
rect 35691 3163 35733 3172
rect 36219 3212 36261 3221
rect 36219 3172 36220 3212
rect 36260 3172 36261 3212
rect 36219 3163 36261 3172
rect 44763 3212 44805 3221
rect 44763 3172 44764 3212
rect 44804 3172 44805 3212
rect 44763 3163 44805 3172
rect 1152 3044 45216 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 45216 3044
rect 1152 2980 45216 3004
rect 2331 2876 2373 2885
rect 2331 2836 2332 2876
rect 2372 2836 2373 2876
rect 2331 2827 2373 2836
rect 2715 2876 2757 2885
rect 2715 2836 2716 2876
rect 2756 2836 2757 2876
rect 2715 2827 2757 2836
rect 3483 2876 3525 2885
rect 3483 2836 3484 2876
rect 3524 2836 3525 2876
rect 3483 2827 3525 2836
rect 6682 2876 6740 2877
rect 6682 2836 6691 2876
rect 6731 2836 6740 2876
rect 6682 2835 6740 2836
rect 7179 2876 7221 2885
rect 7179 2836 7180 2876
rect 7220 2836 7221 2876
rect 7179 2827 7221 2836
rect 10635 2876 10677 2885
rect 10635 2836 10636 2876
rect 10676 2836 10677 2876
rect 10635 2827 10677 2836
rect 13707 2876 13749 2885
rect 13707 2836 13708 2876
rect 13748 2836 13749 2876
rect 13707 2827 13749 2836
rect 17355 2876 17397 2885
rect 17355 2836 17356 2876
rect 17396 2836 17397 2876
rect 17355 2827 17397 2836
rect 20139 2876 20181 2885
rect 20139 2836 20140 2876
rect 20180 2836 20181 2876
rect 20139 2827 20181 2836
rect 23211 2876 23253 2885
rect 23211 2836 23212 2876
rect 23252 2836 23253 2876
rect 23211 2827 23253 2836
rect 25803 2876 25845 2885
rect 25803 2836 25804 2876
rect 25844 2836 25845 2876
rect 25803 2827 25845 2836
rect 29835 2876 29877 2885
rect 29835 2836 29836 2876
rect 29876 2836 29877 2876
rect 29835 2827 29877 2836
rect 31947 2876 31989 2885
rect 31947 2836 31948 2876
rect 31988 2836 31989 2876
rect 31947 2827 31989 2836
rect 35787 2876 35829 2885
rect 35787 2836 35788 2876
rect 35828 2836 35829 2876
rect 35787 2827 35829 2836
rect 38043 2876 38085 2885
rect 38043 2836 38044 2876
rect 38084 2836 38085 2876
rect 38043 2827 38085 2836
rect 40251 2876 40293 2885
rect 40251 2836 40252 2876
rect 40292 2836 40293 2876
rect 40251 2827 40293 2836
rect 40923 2876 40965 2885
rect 40923 2836 40924 2876
rect 40964 2836 40965 2876
rect 40923 2827 40965 2836
rect 8811 2792 8853 2801
rect 8811 2752 8812 2792
rect 8852 2752 8853 2792
rect 8811 2743 8853 2752
rect 10443 2792 10485 2801
rect 10443 2752 10444 2792
rect 10484 2752 10485 2792
rect 10443 2743 10485 2752
rect 15339 2792 15381 2801
rect 15339 2752 15340 2792
rect 15380 2752 15381 2792
rect 15339 2743 15381 2752
rect 17787 2792 17829 2801
rect 17787 2752 17788 2792
rect 17828 2752 17829 2792
rect 17787 2743 17829 2752
rect 27819 2792 27861 2801
rect 27819 2752 27820 2792
rect 27860 2752 27861 2792
rect 27819 2743 27861 2752
rect 36459 2792 36501 2801
rect 36459 2752 36460 2792
rect 36500 2752 36501 2792
rect 36459 2743 36501 2752
rect 40107 2792 40149 2801
rect 40107 2752 40108 2792
rect 40148 2752 40149 2792
rect 40107 2743 40149 2752
rect 45147 2792 45189 2801
rect 45147 2752 45148 2792
rect 45188 2752 45189 2792
rect 45147 2743 45189 2752
rect 4779 2708 4821 2717
rect 6358 2708 6400 2717
rect 4779 2668 4780 2708
rect 4820 2668 4821 2708
rect 4779 2659 4821 2668
rect 6027 2699 6069 2708
rect 6027 2659 6028 2699
rect 6068 2659 6069 2699
rect 6358 2668 6359 2708
rect 6399 2668 6400 2708
rect 6358 2659 6400 2668
rect 6603 2708 6645 2717
rect 6603 2668 6604 2708
rect 6644 2668 6645 2708
rect 6603 2659 6645 2668
rect 6891 2708 6933 2717
rect 6891 2668 6892 2708
rect 6932 2668 6933 2708
rect 6891 2659 6933 2668
rect 7025 2708 7083 2709
rect 7025 2668 7034 2708
rect 7074 2668 7083 2708
rect 7025 2667 7083 2668
rect 7371 2708 7413 2717
rect 9003 2708 9045 2717
rect 12035 2708 12077 2717
rect 7371 2668 7372 2708
rect 7412 2668 7413 2708
rect 7371 2659 7413 2668
rect 8619 2699 8661 2708
rect 8619 2659 8620 2699
rect 8660 2659 8661 2699
rect 9003 2668 9004 2708
rect 9044 2668 9045 2708
rect 9003 2659 9045 2668
rect 10251 2699 10293 2708
rect 10251 2659 10252 2699
rect 10292 2659 10293 2699
rect 6027 2650 6069 2659
rect 8619 2650 8661 2659
rect 10251 2650 10293 2659
rect 10827 2699 10869 2708
rect 10827 2659 10828 2699
rect 10868 2659 10869 2699
rect 12035 2668 12036 2708
rect 12076 2668 12077 2708
rect 12035 2659 12077 2668
rect 12255 2708 12297 2717
rect 13899 2708 13941 2717
rect 15610 2708 15668 2709
rect 12255 2668 12256 2708
rect 12296 2668 12297 2708
rect 12255 2659 12297 2668
rect 13515 2699 13557 2708
rect 13515 2659 13516 2699
rect 13556 2659 13557 2699
rect 13899 2668 13900 2708
rect 13940 2668 13941 2708
rect 13899 2659 13941 2668
rect 15147 2699 15189 2708
rect 15147 2659 15148 2699
rect 15188 2659 15189 2699
rect 15610 2668 15619 2708
rect 15659 2668 15668 2708
rect 15610 2667 15668 2668
rect 15723 2708 15765 2717
rect 15723 2668 15724 2708
rect 15764 2668 15765 2708
rect 15723 2659 15765 2668
rect 16107 2708 16149 2717
rect 18394 2708 18452 2709
rect 16107 2668 16108 2708
rect 16148 2668 16149 2708
rect 16107 2659 16149 2668
rect 16683 2699 16725 2708
rect 16683 2659 16684 2699
rect 16724 2659 16725 2699
rect 10827 2650 10869 2659
rect 13515 2650 13557 2659
rect 15147 2650 15189 2659
rect 16683 2650 16725 2659
rect 17163 2699 17205 2708
rect 17163 2659 17164 2699
rect 17204 2659 17205 2699
rect 18394 2668 18403 2708
rect 18443 2668 18452 2708
rect 18394 2667 18452 2668
rect 18507 2708 18549 2717
rect 18507 2668 18508 2708
rect 18548 2668 18549 2708
rect 18507 2659 18549 2668
rect 18891 2708 18933 2717
rect 21466 2708 21524 2709
rect 18891 2668 18892 2708
rect 18932 2668 18933 2708
rect 18891 2659 18933 2668
rect 19467 2699 19509 2708
rect 19467 2659 19468 2699
rect 19508 2659 19509 2699
rect 17163 2650 17205 2659
rect 19467 2650 19509 2659
rect 19947 2699 19989 2708
rect 19947 2659 19948 2699
rect 19988 2659 19989 2699
rect 21466 2668 21475 2708
rect 21515 2668 21524 2708
rect 21466 2667 21524 2668
rect 21579 2708 21621 2717
rect 21579 2668 21580 2708
rect 21620 2668 21621 2708
rect 21579 2659 21621 2668
rect 21963 2708 22005 2717
rect 24058 2708 24116 2709
rect 21963 2668 21964 2708
rect 22004 2668 22005 2708
rect 21963 2659 22005 2668
rect 22539 2699 22581 2708
rect 22539 2659 22540 2699
rect 22580 2659 22581 2699
rect 19947 2650 19989 2659
rect 22539 2650 22581 2659
rect 23019 2699 23061 2708
rect 23019 2659 23020 2699
rect 23060 2659 23061 2699
rect 24058 2668 24067 2708
rect 24107 2668 24116 2708
rect 24058 2667 24116 2668
rect 24171 2708 24213 2717
rect 24171 2668 24172 2708
rect 24212 2668 24213 2708
rect 24171 2659 24213 2668
rect 24555 2708 24597 2717
rect 26379 2708 26421 2717
rect 28090 2708 28148 2709
rect 24555 2668 24556 2708
rect 24596 2668 24597 2708
rect 24555 2659 24597 2668
rect 25131 2699 25173 2708
rect 25131 2659 25132 2699
rect 25172 2659 25173 2699
rect 23019 2650 23061 2659
rect 25131 2650 25173 2659
rect 25611 2699 25653 2708
rect 25611 2659 25612 2699
rect 25652 2659 25653 2699
rect 26379 2668 26380 2708
rect 26420 2668 26421 2708
rect 26379 2659 26421 2668
rect 27627 2699 27669 2708
rect 27627 2659 27628 2699
rect 27668 2659 27669 2699
rect 28090 2668 28099 2708
rect 28139 2668 28148 2708
rect 28090 2667 28148 2668
rect 28203 2708 28245 2717
rect 28203 2668 28204 2708
rect 28244 2668 28245 2708
rect 28203 2659 28245 2668
rect 28587 2708 28629 2717
rect 30202 2708 30260 2709
rect 28587 2668 28588 2708
rect 28628 2668 28629 2708
rect 28587 2659 28629 2668
rect 29163 2699 29205 2708
rect 29163 2659 29164 2699
rect 29204 2659 29205 2699
rect 25611 2650 25653 2659
rect 27627 2650 27669 2659
rect 29163 2650 29205 2659
rect 29643 2699 29685 2708
rect 29643 2659 29644 2699
rect 29684 2659 29685 2699
rect 30202 2668 30211 2708
rect 30251 2668 30260 2708
rect 30202 2667 30260 2668
rect 30315 2708 30357 2717
rect 30315 2668 30316 2708
rect 30356 2668 30357 2708
rect 30315 2659 30357 2668
rect 30699 2708 30741 2717
rect 32331 2708 32373 2717
rect 30699 2668 30700 2708
rect 30740 2668 30741 2708
rect 31755 2699 31797 2708
rect 30699 2659 30741 2668
rect 31275 2666 31317 2675
rect 29643 2650 29685 2659
rect 1227 2624 1269 2633
rect 1227 2584 1228 2624
rect 1268 2584 1269 2624
rect 1227 2575 1269 2584
rect 1611 2624 1653 2633
rect 1611 2584 1612 2624
rect 1652 2584 1653 2624
rect 1611 2575 1653 2584
rect 1851 2624 1893 2633
rect 1851 2584 1852 2624
rect 1892 2584 1893 2624
rect 1851 2575 1893 2584
rect 2091 2624 2133 2633
rect 2091 2584 2092 2624
rect 2132 2584 2133 2624
rect 2091 2575 2133 2584
rect 2475 2624 2517 2633
rect 2475 2584 2476 2624
rect 2516 2584 2517 2624
rect 2475 2575 2517 2584
rect 2859 2624 2901 2633
rect 2859 2584 2860 2624
rect 2900 2584 2901 2624
rect 2859 2575 2901 2584
rect 3243 2624 3285 2633
rect 3243 2584 3244 2624
rect 3284 2584 3285 2624
rect 3243 2575 3285 2584
rect 3627 2624 3669 2633
rect 3627 2584 3628 2624
rect 3668 2584 3669 2624
rect 3627 2575 3669 2584
rect 4011 2624 4053 2633
rect 4011 2584 4012 2624
rect 4052 2584 4053 2624
rect 4011 2575 4053 2584
rect 4395 2624 4437 2633
rect 4395 2584 4396 2624
rect 4436 2584 4437 2624
rect 4395 2575 4437 2584
rect 6490 2624 6548 2625
rect 6490 2584 6499 2624
rect 6539 2584 6548 2624
rect 6490 2583 6548 2584
rect 16203 2624 16245 2633
rect 16203 2584 16204 2624
rect 16244 2584 16245 2624
rect 16203 2575 16245 2584
rect 17547 2624 17589 2633
rect 17547 2584 17548 2624
rect 17588 2584 17589 2624
rect 17547 2575 17589 2584
rect 17931 2624 17973 2633
rect 17931 2584 17932 2624
rect 17972 2584 17973 2624
rect 17931 2575 17973 2584
rect 18987 2624 19029 2633
rect 18987 2584 18988 2624
rect 19028 2584 19029 2624
rect 18987 2575 19029 2584
rect 20619 2624 20661 2633
rect 20619 2584 20620 2624
rect 20660 2584 20661 2624
rect 20619 2575 20661 2584
rect 21003 2624 21045 2633
rect 21003 2584 21004 2624
rect 21044 2584 21045 2624
rect 21003 2575 21045 2584
rect 22059 2624 22101 2633
rect 22059 2584 22060 2624
rect 22100 2584 22101 2624
rect 22059 2575 22101 2584
rect 23595 2624 23637 2633
rect 23595 2584 23596 2624
rect 23636 2584 23637 2624
rect 23595 2575 23637 2584
rect 24651 2624 24693 2633
rect 24651 2584 24652 2624
rect 24692 2584 24693 2624
rect 24651 2575 24693 2584
rect 26187 2624 26229 2633
rect 26187 2584 26188 2624
rect 26228 2584 26229 2624
rect 26187 2575 26229 2584
rect 28683 2624 28725 2633
rect 28683 2584 28684 2624
rect 28724 2584 28725 2624
rect 28683 2575 28725 2584
rect 30795 2624 30837 2633
rect 30795 2584 30796 2624
rect 30836 2584 30837 2624
rect 31275 2626 31276 2666
rect 31316 2626 31317 2666
rect 31755 2659 31756 2699
rect 31796 2659 31797 2699
rect 32331 2668 32332 2708
rect 32372 2668 32373 2708
rect 32331 2659 32373 2668
rect 33579 2708 33637 2709
rect 33579 2668 33588 2708
rect 33628 2668 33637 2708
rect 33579 2667 33637 2668
rect 34042 2708 34100 2709
rect 34042 2668 34051 2708
rect 34091 2668 34100 2708
rect 34042 2667 34100 2668
rect 34155 2708 34197 2717
rect 34155 2668 34156 2708
rect 34196 2668 34197 2708
rect 34155 2659 34197 2668
rect 34539 2708 34581 2717
rect 37899 2708 37941 2717
rect 34539 2668 34540 2708
rect 34580 2668 34581 2708
rect 34539 2659 34581 2668
rect 35115 2699 35157 2708
rect 35115 2659 35116 2699
rect 35156 2659 35157 2699
rect 31755 2650 31797 2659
rect 35115 2650 35157 2659
rect 35595 2699 35637 2708
rect 35595 2659 35596 2699
rect 35636 2659 35637 2699
rect 35595 2650 35637 2659
rect 36651 2699 36693 2708
rect 36651 2659 36652 2699
rect 36692 2659 36693 2699
rect 37899 2668 37900 2708
rect 37940 2668 37941 2708
rect 37899 2659 37941 2668
rect 38667 2708 38709 2717
rect 38667 2668 38668 2708
rect 38708 2668 38709 2708
rect 38667 2659 38709 2668
rect 39915 2699 39957 2708
rect 39915 2659 39916 2699
rect 39956 2659 39957 2699
rect 36651 2650 36693 2659
rect 39915 2650 39957 2659
rect 31275 2617 31317 2626
rect 34635 2624 34677 2633
rect 30795 2575 30837 2584
rect 34635 2584 34636 2624
rect 34676 2584 34677 2624
rect 34635 2575 34677 2584
rect 36171 2624 36213 2633
rect 36171 2584 36172 2624
rect 36212 2584 36213 2624
rect 36171 2575 36213 2584
rect 38283 2624 38325 2633
rect 38283 2584 38284 2624
rect 38324 2584 38325 2624
rect 38283 2575 38325 2584
rect 40491 2624 40533 2633
rect 40491 2584 40492 2624
rect 40532 2584 40533 2624
rect 40491 2575 40533 2584
rect 40683 2624 40725 2633
rect 40683 2584 40684 2624
rect 40724 2584 40725 2624
rect 40683 2575 40725 2584
rect 44139 2624 44181 2633
rect 44139 2584 44140 2624
rect 44180 2584 44181 2624
rect 44139 2575 44181 2584
rect 44523 2624 44565 2633
rect 44523 2584 44524 2624
rect 44564 2584 44565 2624
rect 44523 2575 44565 2584
rect 44907 2624 44949 2633
rect 44907 2584 44908 2624
rect 44948 2584 44949 2624
rect 44907 2575 44949 2584
rect 1467 2540 1509 2549
rect 1467 2500 1468 2540
rect 1508 2500 1509 2540
rect 1467 2491 1509 2500
rect 3867 2540 3909 2549
rect 3867 2500 3868 2540
rect 3908 2500 3909 2540
rect 3867 2491 3909 2500
rect 6219 2540 6261 2549
rect 6219 2500 6220 2540
rect 6260 2500 6261 2540
rect 6219 2491 6261 2500
rect 20859 2540 20901 2549
rect 20859 2500 20860 2540
rect 20900 2500 20901 2540
rect 20859 2491 20901 2500
rect 44763 2540 44805 2549
rect 44763 2500 44764 2540
rect 44804 2500 44805 2540
rect 44763 2491 44805 2500
rect 3099 2456 3141 2465
rect 3099 2416 3100 2456
rect 3140 2416 3141 2456
rect 3099 2407 3141 2416
rect 4251 2456 4293 2465
rect 4251 2416 4252 2456
rect 4292 2416 4293 2456
rect 4251 2407 4293 2416
rect 4635 2456 4677 2465
rect 4635 2416 4636 2456
rect 4676 2416 4677 2456
rect 4635 2407 4677 2416
rect 18171 2456 18213 2465
rect 18171 2416 18172 2456
rect 18212 2416 18213 2456
rect 18171 2407 18213 2416
rect 21243 2456 21285 2465
rect 21243 2416 21244 2456
rect 21284 2416 21285 2456
rect 21243 2407 21285 2416
rect 23835 2456 23877 2465
rect 23835 2416 23836 2456
rect 23876 2416 23877 2456
rect 23835 2407 23877 2416
rect 25947 2456 25989 2465
rect 25947 2416 25948 2456
rect 25988 2416 25989 2456
rect 25947 2407 25989 2416
rect 33771 2456 33813 2465
rect 33771 2416 33772 2456
rect 33812 2416 33813 2456
rect 33771 2407 33813 2416
rect 35931 2456 35973 2465
rect 35931 2416 35932 2456
rect 35972 2416 35973 2456
rect 35931 2407 35973 2416
rect 44379 2456 44421 2465
rect 44379 2416 44380 2456
rect 44420 2416 44421 2456
rect 44379 2407 44421 2416
rect 1152 2288 45216 2312
rect 1152 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 45216 2288
rect 1152 2224 45216 2248
rect 1467 2120 1509 2129
rect 1467 2080 1468 2120
rect 1508 2080 1509 2120
rect 1467 2071 1509 2080
rect 2235 2120 2277 2129
rect 2235 2080 2236 2120
rect 2276 2080 2277 2120
rect 2235 2071 2277 2080
rect 3291 2120 3333 2129
rect 3291 2080 3292 2120
rect 3332 2080 3333 2120
rect 3291 2071 3333 2080
rect 4443 2120 4485 2129
rect 4443 2080 4444 2120
rect 4484 2080 4485 2120
rect 4443 2071 4485 2080
rect 4827 2120 4869 2129
rect 4827 2080 4828 2120
rect 4868 2080 4869 2120
rect 4827 2071 4869 2080
rect 6411 2120 6453 2129
rect 6411 2080 6412 2120
rect 6452 2080 6453 2120
rect 6411 2071 6453 2080
rect 6939 2120 6981 2129
rect 6939 2080 6940 2120
rect 6980 2080 6981 2120
rect 6939 2071 6981 2080
rect 7611 2120 7653 2129
rect 7611 2080 7612 2120
rect 7652 2080 7653 2120
rect 7611 2071 7653 2080
rect 12075 2120 12117 2129
rect 12075 2080 12076 2120
rect 12116 2080 12117 2120
rect 12075 2071 12117 2080
rect 12891 2120 12933 2129
rect 12891 2080 12892 2120
rect 12932 2080 12933 2120
rect 12891 2071 12933 2080
rect 13275 2120 13317 2129
rect 13275 2080 13276 2120
rect 13316 2080 13317 2120
rect 13275 2071 13317 2080
rect 13659 2120 13701 2129
rect 13659 2080 13660 2120
rect 13700 2080 13701 2120
rect 13659 2071 13701 2080
rect 15243 2120 15285 2129
rect 15243 2080 15244 2120
rect 15284 2080 15285 2120
rect 15243 2071 15285 2080
rect 15675 2120 15717 2129
rect 15675 2080 15676 2120
rect 15716 2080 15717 2120
rect 15675 2071 15717 2080
rect 16059 2120 16101 2129
rect 16059 2080 16060 2120
rect 16100 2080 16101 2120
rect 16059 2071 16101 2080
rect 16443 2120 16485 2129
rect 16443 2080 16444 2120
rect 16484 2080 16485 2120
rect 16443 2071 16485 2080
rect 18411 2120 18453 2129
rect 18411 2080 18412 2120
rect 18452 2080 18453 2120
rect 18411 2071 18453 2080
rect 20043 2120 20085 2129
rect 20043 2080 20044 2120
rect 20084 2080 20085 2120
rect 20043 2071 20085 2080
rect 20667 2120 20709 2129
rect 20667 2080 20668 2120
rect 20708 2080 20709 2120
rect 20667 2071 20709 2080
rect 23019 2120 23061 2129
rect 23019 2080 23020 2120
rect 23060 2080 23061 2120
rect 23019 2071 23061 2080
rect 26698 2120 26756 2121
rect 26698 2080 26707 2120
rect 26747 2080 26756 2120
rect 26698 2079 26756 2080
rect 29163 2120 29205 2129
rect 29163 2080 29164 2120
rect 29204 2080 29205 2120
rect 29163 2071 29205 2080
rect 32043 2120 32085 2129
rect 32043 2080 32044 2120
rect 32084 2080 32085 2120
rect 32043 2071 32085 2080
rect 36010 2120 36068 2121
rect 36010 2080 36019 2120
rect 36059 2080 36068 2120
rect 36010 2079 36068 2080
rect 38763 2120 38805 2129
rect 38763 2080 38764 2120
rect 38804 2080 38805 2120
rect 38763 2071 38805 2080
rect 45147 2120 45189 2129
rect 45147 2080 45148 2120
rect 45188 2080 45189 2120
rect 45147 2071 45189 2080
rect 1851 2036 1893 2045
rect 1851 1996 1852 2036
rect 1892 1996 1893 2036
rect 1851 1987 1893 1996
rect 6555 2036 6597 2045
rect 6555 1996 6556 2036
rect 6596 1996 6597 2036
rect 6555 1987 6597 1996
rect 7995 2036 8037 2045
rect 7995 1996 7996 2036
rect 8036 1996 8037 2036
rect 7995 1987 8037 1996
rect 10491 2036 10533 2045
rect 10491 1996 10492 2036
rect 10532 1996 10533 2036
rect 10491 1987 10533 1996
rect 1227 1952 1269 1961
rect 1227 1912 1228 1952
rect 1268 1912 1269 1952
rect 1227 1903 1269 1912
rect 1611 1952 1653 1961
rect 1611 1912 1612 1952
rect 1652 1912 1653 1952
rect 1611 1903 1653 1912
rect 1995 1952 2037 1961
rect 1995 1912 1996 1952
rect 2036 1912 2037 1952
rect 1995 1903 2037 1912
rect 2667 1952 2709 1961
rect 2667 1912 2668 1952
rect 2708 1912 2709 1952
rect 2667 1903 2709 1912
rect 3051 1952 3093 1961
rect 3051 1912 3052 1952
rect 3092 1912 3093 1952
rect 3051 1903 3093 1912
rect 3435 1952 3477 1961
rect 3435 1912 3436 1952
rect 3476 1912 3477 1952
rect 3435 1903 3477 1912
rect 3819 1952 3861 1961
rect 3819 1912 3820 1952
rect 3860 1912 3861 1952
rect 3819 1903 3861 1912
rect 4203 1952 4245 1961
rect 4203 1912 4204 1952
rect 4244 1912 4245 1952
rect 4203 1903 4245 1912
rect 4618 1952 4676 1953
rect 4618 1912 4627 1952
rect 4667 1912 4676 1952
rect 4618 1911 4676 1912
rect 6795 1952 6837 1961
rect 6795 1912 6796 1952
rect 6836 1912 6837 1952
rect 6795 1903 6837 1912
rect 7179 1952 7221 1961
rect 7179 1912 7180 1952
rect 7220 1912 7221 1952
rect 7179 1903 7221 1912
rect 7371 1952 7413 1961
rect 7371 1912 7372 1952
rect 7412 1912 7413 1952
rect 7371 1903 7413 1912
rect 7755 1952 7797 1961
rect 7755 1912 7756 1952
rect 7796 1912 7797 1952
rect 7755 1903 7797 1912
rect 8139 1952 8181 1961
rect 8139 1912 8140 1952
rect 8180 1912 8181 1952
rect 8139 1903 8181 1912
rect 10251 1952 10293 1961
rect 10251 1912 10252 1952
rect 10292 1912 10293 1952
rect 10251 1903 10293 1912
rect 12267 1952 12309 1961
rect 12267 1912 12268 1952
rect 12308 1912 12309 1952
rect 12267 1903 12309 1912
rect 12507 1952 12549 1961
rect 12507 1912 12508 1952
rect 12548 1912 12549 1952
rect 12507 1903 12549 1912
rect 12651 1952 12693 1961
rect 12651 1912 12652 1952
rect 12692 1912 12693 1952
rect 12651 1903 12693 1912
rect 13035 1952 13077 1961
rect 13035 1912 13036 1952
rect 13076 1912 13077 1952
rect 13035 1903 13077 1912
rect 13419 1952 13461 1961
rect 13419 1912 13420 1952
rect 13460 1912 13461 1952
rect 13419 1903 13461 1912
rect 15435 1952 15477 1961
rect 15435 1912 15436 1952
rect 15476 1912 15477 1952
rect 15435 1903 15477 1912
rect 15819 1952 15861 1961
rect 15819 1912 15820 1952
rect 15860 1912 15861 1952
rect 15819 1903 15861 1912
rect 16203 1952 16245 1961
rect 16203 1912 16204 1952
rect 16244 1912 16245 1952
rect 16203 1903 16245 1912
rect 16587 1952 16629 1961
rect 16587 1912 16588 1952
rect 16628 1912 16629 1952
rect 16587 1903 16629 1912
rect 20427 1952 20469 1961
rect 20427 1912 20428 1952
rect 20468 1912 20469 1952
rect 20427 1903 20469 1912
rect 20811 1952 20853 1961
rect 20811 1912 20812 1952
rect 20852 1912 20853 1952
rect 20811 1903 20853 1912
rect 21195 1952 21237 1961
rect 21195 1912 21196 1952
rect 21236 1912 21237 1952
rect 21195 1903 21237 1912
rect 25419 1952 25461 1961
rect 25419 1912 25420 1952
rect 25460 1912 25461 1952
rect 25419 1903 25461 1912
rect 27051 1952 27093 1961
rect 27051 1912 27052 1952
rect 27092 1912 27093 1952
rect 27051 1903 27093 1912
rect 27435 1952 27477 1961
rect 27435 1912 27436 1952
rect 27476 1912 27477 1952
rect 27435 1903 27477 1912
rect 29307 1952 29349 1961
rect 29307 1912 29308 1952
rect 29348 1912 29349 1952
rect 29307 1903 29349 1912
rect 29547 1952 29589 1961
rect 29547 1912 29548 1952
rect 29588 1912 29589 1952
rect 29547 1903 29589 1912
rect 29931 1952 29973 1961
rect 29931 1912 29932 1952
rect 29972 1912 29973 1952
rect 29931 1903 29973 1912
rect 30315 1952 30357 1961
rect 30315 1912 30316 1952
rect 30356 1912 30357 1952
rect 30315 1903 30357 1912
rect 32427 1952 32469 1961
rect 32427 1912 32428 1952
rect 32468 1912 32469 1952
rect 32427 1903 32469 1912
rect 32811 1952 32853 1961
rect 32811 1912 32812 1952
rect 32852 1912 32853 1952
rect 32811 1903 32853 1912
rect 33195 1952 33237 1961
rect 33195 1912 33196 1952
rect 33236 1912 33237 1952
rect 33195 1903 33237 1912
rect 33579 1952 33621 1961
rect 33579 1912 33580 1952
rect 33620 1912 33621 1952
rect 33579 1903 33621 1912
rect 33963 1952 34005 1961
rect 33963 1912 33964 1952
rect 34004 1912 34005 1952
rect 33963 1903 34005 1912
rect 34827 1952 34869 1961
rect 34827 1912 34828 1952
rect 34868 1912 34869 1952
rect 34827 1903 34869 1912
rect 38283 1952 38325 1961
rect 38283 1912 38284 1952
rect 38324 1912 38325 1952
rect 38283 1903 38325 1912
rect 43755 1952 43797 1961
rect 43755 1912 43756 1952
rect 43796 1912 43797 1952
rect 43755 1903 43797 1912
rect 44139 1952 44181 1961
rect 44139 1912 44140 1952
rect 44180 1912 44181 1952
rect 44139 1903 44181 1912
rect 44523 1952 44565 1961
rect 44523 1912 44524 1952
rect 44564 1912 44565 1952
rect 44523 1903 44565 1912
rect 44907 1952 44949 1961
rect 44907 1912 44908 1952
rect 44948 1912 44949 1952
rect 44907 1903 44949 1912
rect 4971 1868 5013 1877
rect 4971 1828 4972 1868
rect 5012 1828 5013 1868
rect 4971 1819 5013 1828
rect 6211 1868 6269 1869
rect 6211 1828 6220 1868
rect 6260 1828 6269 1868
rect 6211 1827 6269 1828
rect 8523 1868 8565 1877
rect 8523 1828 8524 1868
rect 8564 1828 8565 1868
rect 8523 1819 8565 1828
rect 9763 1868 9821 1869
rect 9763 1828 9772 1868
rect 9812 1828 9821 1868
rect 9763 1827 9821 1828
rect 10635 1868 10677 1877
rect 10635 1828 10636 1868
rect 10676 1828 10677 1868
rect 10635 1819 10677 1828
rect 11875 1868 11933 1869
rect 11875 1828 11884 1868
rect 11924 1828 11933 1868
rect 11875 1827 11933 1828
rect 13803 1868 13845 1877
rect 13803 1828 13804 1868
rect 13844 1828 13845 1868
rect 13803 1819 13845 1828
rect 15043 1868 15101 1869
rect 15043 1828 15052 1868
rect 15092 1828 15101 1868
rect 15043 1827 15101 1828
rect 16971 1868 17013 1877
rect 16971 1828 16972 1868
rect 17012 1828 17013 1868
rect 16971 1819 17013 1828
rect 18211 1868 18269 1869
rect 18211 1828 18220 1868
rect 18260 1828 18269 1868
rect 18211 1827 18269 1828
rect 18603 1868 18645 1877
rect 18603 1828 18604 1868
rect 18644 1828 18645 1868
rect 18603 1819 18645 1828
rect 19843 1868 19901 1869
rect 19843 1828 19852 1868
rect 19892 1828 19901 1868
rect 19843 1827 19901 1828
rect 21579 1868 21621 1877
rect 21579 1828 21580 1868
rect 21620 1828 21621 1868
rect 21579 1819 21621 1828
rect 22819 1868 22877 1869
rect 22819 1828 22828 1868
rect 22868 1828 22877 1868
rect 22819 1827 22877 1828
rect 23211 1868 23253 1877
rect 23211 1828 23212 1868
rect 23252 1828 23253 1868
rect 23211 1819 23253 1828
rect 24451 1868 24509 1869
rect 24451 1828 24460 1868
rect 24500 1828 24509 1868
rect 24451 1827 24509 1828
rect 24922 1868 24980 1869
rect 24922 1828 24931 1868
rect 24971 1828 24980 1868
rect 24922 1827 24980 1828
rect 25035 1868 25077 1877
rect 25035 1828 25036 1868
rect 25076 1828 25077 1868
rect 25035 1819 25077 1828
rect 25515 1868 25557 1877
rect 25515 1828 25516 1868
rect 25556 1828 25557 1868
rect 25515 1819 25557 1828
rect 25987 1868 26045 1869
rect 25987 1828 25996 1868
rect 26036 1828 26045 1868
rect 25987 1827 26045 1828
rect 26475 1868 26533 1869
rect 26475 1828 26484 1868
rect 26524 1828 26533 1868
rect 26475 1827 26533 1828
rect 27723 1868 27765 1877
rect 27723 1828 27724 1868
rect 27764 1828 27765 1868
rect 27723 1819 27765 1828
rect 28963 1868 29021 1869
rect 28963 1828 28972 1868
rect 29012 1828 29021 1868
rect 28963 1827 29021 1828
rect 30603 1868 30645 1877
rect 30603 1828 30604 1868
rect 30644 1828 30645 1868
rect 30603 1819 30645 1828
rect 31843 1868 31901 1869
rect 31843 1828 31852 1868
rect 31892 1828 31901 1868
rect 31843 1827 31901 1828
rect 34234 1868 34292 1869
rect 34234 1828 34243 1868
rect 34283 1828 34292 1868
rect 34234 1827 34292 1828
rect 34347 1868 34389 1877
rect 34347 1828 34348 1868
rect 34388 1828 34389 1868
rect 34347 1819 34389 1828
rect 34731 1868 34773 1877
rect 34731 1828 34732 1868
rect 34772 1828 34773 1868
rect 34731 1819 34773 1828
rect 35299 1868 35357 1869
rect 35299 1828 35308 1868
rect 35348 1828 35357 1868
rect 35299 1827 35357 1828
rect 35818 1868 35876 1869
rect 35818 1828 35827 1868
rect 35867 1828 35876 1868
rect 35818 1827 35876 1828
rect 36643 1868 36701 1869
rect 36643 1828 36652 1868
rect 36692 1828 36701 1868
rect 36643 1827 36701 1828
rect 37899 1868 37941 1877
rect 37899 1828 37900 1868
rect 37940 1828 37941 1868
rect 37899 1819 37941 1828
rect 38947 1868 39005 1869
rect 38947 1828 38956 1868
rect 38996 1828 39005 1868
rect 38947 1827 39005 1828
rect 40203 1868 40245 1877
rect 40203 1828 40204 1868
rect 40244 1828 40245 1868
rect 40203 1819 40245 1828
rect 2907 1784 2949 1793
rect 2907 1744 2908 1784
rect 2948 1744 2949 1784
rect 2907 1735 2949 1744
rect 9963 1784 10005 1793
rect 9963 1744 9964 1784
rect 10004 1744 10005 1784
rect 9963 1735 10005 1744
rect 24651 1784 24693 1793
rect 24651 1744 24652 1784
rect 24692 1744 24693 1784
rect 24651 1735 24693 1744
rect 36459 1784 36501 1793
rect 36459 1744 36460 1784
rect 36500 1744 36501 1784
rect 36459 1735 36501 1744
rect 43995 1784 44037 1793
rect 43995 1744 43996 1784
rect 44036 1744 44037 1784
rect 43995 1735 44037 1744
rect 44763 1784 44805 1793
rect 44763 1744 44764 1784
rect 44804 1744 44805 1784
rect 44763 1735 44805 1744
rect 3675 1700 3717 1709
rect 3675 1660 3676 1700
rect 3716 1660 3717 1700
rect 3675 1651 3717 1660
rect 4059 1700 4101 1709
rect 4059 1660 4060 1700
rect 4100 1660 4101 1700
rect 4059 1651 4101 1660
rect 8379 1700 8421 1709
rect 8379 1660 8380 1700
rect 8420 1660 8421 1700
rect 8379 1651 8421 1660
rect 16827 1700 16869 1709
rect 16827 1660 16828 1700
rect 16868 1660 16869 1700
rect 16827 1651 16869 1660
rect 21051 1700 21093 1709
rect 21051 1660 21052 1700
rect 21092 1660 21093 1700
rect 21051 1651 21093 1660
rect 21435 1700 21477 1709
rect 21435 1660 21436 1700
rect 21476 1660 21477 1700
rect 21435 1651 21477 1660
rect 26811 1700 26853 1709
rect 26811 1660 26812 1700
rect 26852 1660 26853 1700
rect 26811 1651 26853 1660
rect 27195 1700 27237 1709
rect 27195 1660 27196 1700
rect 27236 1660 27237 1700
rect 27195 1651 27237 1660
rect 29691 1700 29733 1709
rect 29691 1660 29692 1700
rect 29732 1660 29733 1700
rect 29691 1651 29733 1660
rect 30075 1700 30117 1709
rect 30075 1660 30076 1700
rect 30116 1660 30117 1700
rect 30075 1651 30117 1660
rect 32187 1700 32229 1709
rect 32187 1660 32188 1700
rect 32228 1660 32229 1700
rect 32187 1651 32229 1660
rect 32571 1700 32613 1709
rect 32571 1660 32572 1700
rect 32612 1660 32613 1700
rect 32571 1651 32613 1660
rect 32955 1700 32997 1709
rect 32955 1660 32956 1700
rect 32996 1660 32997 1700
rect 32955 1651 32997 1660
rect 33339 1700 33381 1709
rect 33339 1660 33340 1700
rect 33380 1660 33381 1700
rect 33339 1651 33381 1660
rect 33723 1700 33765 1709
rect 33723 1660 33724 1700
rect 33764 1660 33765 1700
rect 33723 1651 33765 1660
rect 38043 1700 38085 1709
rect 38043 1660 38044 1700
rect 38084 1660 38085 1700
rect 38043 1651 38085 1660
rect 44379 1700 44421 1709
rect 44379 1660 44380 1700
rect 44420 1660 44421 1700
rect 44379 1651 44421 1660
rect 1152 1532 45216 1556
rect 1152 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 45216 1532
rect 1152 1468 45216 1492
<< via1 >>
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 1468 10396 1508 10436
rect 3004 10396 3044 10436
rect 3868 10396 3908 10436
rect 5308 10396 5348 10436
rect 5884 10396 5924 10436
rect 7804 10396 7844 10436
rect 8092 10396 8132 10436
rect 9148 10396 9188 10436
rect 11356 10396 11396 10436
rect 11740 10396 11780 10436
rect 16732 10396 16772 10436
rect 17404 10396 17444 10436
rect 19708 10396 19748 10436
rect 24028 10396 24068 10436
rect 27388 10396 27428 10436
rect 27772 10396 27812 10436
rect 29884 10396 29924 10436
rect 32284 10396 32324 10436
rect 34684 10396 34724 10436
rect 36796 10396 36836 10436
rect 37564 10396 37604 10436
rect 38140 10396 38180 10436
rect 38812 10396 38852 10436
rect 40588 10396 40628 10436
rect 42556 10396 42596 10436
rect 42940 10396 42980 10436
rect 44092 10396 44132 10436
rect 44476 10396 44516 10436
rect 8764 10312 8804 10352
rect 32668 10312 32708 10352
rect 38956 10312 38996 10352
rect 42172 10312 42212 10352
rect 44860 10312 44900 10352
rect 6796 10228 6836 10268
rect 6940 10228 6980 10268
rect 7084 10228 7124 10268
rect 7206 10228 7246 10268
rect 7333 10228 7373 10268
rect 9292 10228 9332 10268
rect 10540 10219 10580 10259
rect 11884 10228 11924 10268
rect 13132 10219 13172 10259
rect 13516 10228 13556 10268
rect 14764 10219 14804 10259
rect 15148 10228 15188 10268
rect 16396 10219 16436 10259
rect 17548 10228 17588 10268
rect 18796 10219 18836 10259
rect 20236 10219 20276 10259
rect 21484 10228 21524 10268
rect 21868 10228 21908 10268
rect 23116 10219 23156 10259
rect 24172 10228 24212 10268
rect 25420 10219 25460 10259
rect 25804 10228 25844 10268
rect 27052 10219 27092 10259
rect 28300 10228 28340 10268
rect 29548 10219 29588 10259
rect 30316 10228 30356 10268
rect 31572 10228 31612 10268
rect 33100 10228 33140 10268
rect 34348 10219 34388 10259
rect 35212 10228 35252 10268
rect 36460 10219 36500 10259
rect 39148 10219 39188 10259
rect 40396 10228 40436 10268
rect 40780 10219 40820 10259
rect 42028 10228 42068 10268
rect 1228 10144 1268 10184
rect 1612 10144 1652 10184
rect 1996 10144 2036 10184
rect 2380 10144 2420 10184
rect 2764 10144 2804 10184
rect 3628 10144 3668 10184
rect 4972 10144 5012 10184
rect 5548 10144 5588 10184
rect 6124 10144 6164 10184
rect 7564 10144 7604 10184
rect 8332 10144 8372 10184
rect 8524 10144 8564 10184
rect 8908 10144 8948 10184
rect 11116 10144 11156 10184
rect 11500 10144 11540 10184
rect 16972 10144 17012 10184
rect 17164 10144 17204 10184
rect 19468 10144 19508 10184
rect 23788 10144 23828 10184
rect 27628 10144 27668 10184
rect 28012 10144 28052 10184
rect 30124 10144 30164 10184
rect 31948 10144 31988 10184
rect 32188 10144 32228 10184
rect 32524 10144 32564 10184
rect 32908 10144 32948 10184
rect 34924 10144 34964 10184
rect 37036 10144 37076 10184
rect 37228 10144 37268 10184
rect 37804 10144 37844 10184
rect 38380 10144 38420 10184
rect 38572 10144 38612 10184
rect 42412 10144 42452 10184
rect 42796 10144 42836 10184
rect 43180 10144 43220 10184
rect 43564 10144 43604 10184
rect 43708 10144 43748 10184
rect 43948 10144 43988 10184
rect 44332 10144 44372 10184
rect 44716 10144 44756 10184
rect 45100 10144 45140 10184
rect 2236 10060 2276 10100
rect 5212 10060 5252 10100
rect 7180 10060 7220 10100
rect 16588 10060 16628 10100
rect 25612 10060 25652 10100
rect 27244 10060 27284 10100
rect 37468 10060 37508 10100
rect 43324 10060 43364 10100
rect 1852 9976 1892 10016
rect 2620 9976 2660 10016
rect 10732 9976 10772 10016
rect 13324 9976 13364 10016
rect 14956 9976 14996 10016
rect 18988 9976 19028 10016
rect 20044 9976 20084 10016
rect 23308 9976 23348 10016
rect 29740 9976 29780 10016
rect 31756 9976 31796 10016
rect 34540 9976 34580 10016
rect 36652 9976 36692 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 5740 9640 5780 9680
rect 7372 9640 7412 9680
rect 13948 9640 13988 9680
rect 14812 9640 14852 9680
rect 18172 9640 18212 9680
rect 20764 9640 20804 9680
rect 26236 9640 26276 9680
rect 33148 9640 33188 9680
rect 33916 9640 33956 9680
rect 44188 9640 44228 9680
rect 44572 9640 44612 9680
rect 21436 9556 21476 9596
rect 43036 9556 43076 9596
rect 1228 9472 1268 9512
rect 1612 9472 1652 9512
rect 1996 9472 2036 9512
rect 2236 9472 2276 9512
rect 8140 9472 8180 9512
rect 8524 9472 8564 9512
rect 9004 9472 9044 9512
rect 11980 9472 12020 9512
rect 13267 9472 13307 9512
rect 13420 9472 13460 9512
rect 14188 9472 14228 9512
rect 14572 9472 14612 9512
rect 15532 9472 15572 9512
rect 16972 9472 17012 9512
rect 17932 9472 17972 9512
rect 18892 9472 18932 9512
rect 20179 9472 20219 9512
rect 20332 9472 20372 9512
rect 21004 9472 21044 9512
rect 21235 9472 21275 9512
rect 22156 9472 22196 9512
rect 23443 9472 23483 9512
rect 23596 9472 23636 9512
rect 24844 9472 24884 9512
rect 26476 9472 26516 9512
rect 26707 9472 26747 9512
rect 26908 9472 26948 9512
rect 27820 9472 27860 9512
rect 29251 9472 29291 9512
rect 31756 9472 31796 9512
rect 33388 9472 33428 9512
rect 33772 9472 33812 9512
rect 34156 9472 34196 9512
rect 35020 9472 35060 9512
rect 36556 9472 36596 9512
rect 42028 9472 42068 9512
rect 42652 9472 42692 9512
rect 42892 9472 42932 9512
rect 43276 9472 43316 9512
rect 43660 9472 43700 9512
rect 44044 9472 44084 9512
rect 44428 9472 44468 9512
rect 44812 9472 44852 9512
rect 4300 9388 4340 9428
rect 5548 9388 5588 9428
rect 5932 9388 5972 9428
rect 7180 9388 7220 9428
rect 7660 9388 7700 9428
rect 7779 9388 7819 9428
rect 7891 9388 7931 9428
rect 9676 9388 9716 9428
rect 10924 9388 10964 9428
rect 11470 9388 11510 9428
rect 11587 9360 11627 9400
rect 12076 9388 12116 9428
rect 12556 9388 12596 9428
rect 13075 9388 13115 9428
rect 15022 9388 15062 9428
rect 15148 9388 15188 9428
rect 15628 9388 15668 9428
rect 16108 9388 16148 9428
rect 16596 9388 16636 9428
rect 18403 9388 18443 9428
rect 18508 9388 18548 9428
rect 18988 9388 19028 9428
rect 19468 9388 19508 9428
rect 19987 9388 20027 9428
rect 21667 9388 21707 9428
rect 21772 9388 21812 9428
rect 22252 9388 22292 9428
rect 22732 9388 22772 9428
rect 23251 9388 23291 9428
rect 24355 9388 24395 9428
rect 24460 9388 24500 9428
rect 24940 9388 24980 9428
rect 25420 9388 25460 9428
rect 25908 9388 25948 9428
rect 27331 9388 27371 9428
rect 27436 9388 27476 9428
rect 27916 9388 27956 9428
rect 28396 9388 28436 9428
rect 28915 9388 28955 9428
rect 29452 9388 29492 9428
rect 30700 9388 30740 9428
rect 31267 9388 31307 9428
rect 31372 9388 31412 9428
rect 31852 9388 31892 9428
rect 32332 9388 32372 9428
rect 32820 9388 32860 9428
rect 34527 9388 34567 9428
rect 34636 9388 34676 9428
rect 35116 9388 35156 9428
rect 35596 9388 35636 9428
rect 36115 9388 36155 9428
rect 37132 9388 37172 9428
rect 38380 9388 38420 9428
rect 38764 9388 38804 9428
rect 40012 9388 40052 9428
rect 40401 9388 40441 9428
rect 41644 9388 41684 9428
rect 7564 9304 7604 9344
rect 20572 9304 20612 9344
rect 36940 9304 36980 9344
rect 43804 9304 43844 9344
rect 1468 9220 1508 9260
rect 1852 9220 1892 9260
rect 7372 9220 7412 9260
rect 8380 9220 8420 9260
rect 8764 9220 8804 9260
rect 9244 9220 9284 9260
rect 11116 9220 11156 9260
rect 13660 9220 13700 9260
rect 16780 9220 16820 9260
rect 17212 9220 17252 9260
rect 23836 9220 23876 9260
rect 26092 9220 26132 9260
rect 29068 9220 29108 9260
rect 33004 9220 33044 9260
rect 33532 9220 33572 9260
rect 36268 9220 36308 9260
rect 36796 9220 36836 9260
rect 40204 9220 40244 9260
rect 41836 9220 41876 9260
rect 42268 9220 42308 9260
rect 43420 9220 43460 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 1852 8884 1892 8924
rect 12460 8884 12500 8924
rect 12652 8884 12692 8924
rect 15724 8884 15764 8924
rect 17356 8884 17396 8924
rect 19372 8884 19412 8924
rect 19708 8884 19748 8924
rect 21676 8884 21716 8924
rect 22108 8884 22148 8924
rect 24268 8884 24308 8924
rect 31756 8884 31796 8924
rect 33388 8884 33428 8924
rect 44476 8884 44516 8924
rect 9676 8800 9716 8840
rect 10492 8800 10532 8840
rect 29404 8800 29444 8840
rect 36220 8800 36260 8840
rect 42172 8800 42212 8840
rect 43036 8800 43076 8840
rect 4300 8716 4340 8756
rect 5548 8707 5588 8747
rect 5932 8716 5972 8756
rect 7180 8707 7220 8747
rect 7719 8716 7759 8756
rect 7837 8696 7877 8736
rect 7939 8716 7979 8756
rect 8236 8716 8276 8756
rect 9484 8707 9524 8747
rect 10723 8716 10763 8756
rect 10828 8716 10868 8756
rect 11212 8716 11252 8756
rect 11788 8707 11828 8747
rect 12268 8707 12308 8747
rect 12836 8716 12876 8756
rect 14092 8716 14132 8756
rect 14284 8716 14324 8756
rect 15532 8707 15572 8747
rect 15916 8716 15956 8756
rect 17164 8707 17204 8747
rect 17635 8716 17675 8756
rect 17740 8716 17780 8756
rect 18124 8716 18164 8756
rect 18700 8707 18740 8747
rect 19180 8707 19220 8747
rect 20236 8716 20276 8756
rect 21484 8707 21524 8747
rect 22828 8716 22868 8756
rect 24076 8707 24116 8747
rect 25228 8716 25268 8756
rect 26476 8707 26516 8747
rect 27052 8716 27092 8756
rect 28300 8707 28340 8747
rect 30019 8716 30059 8756
rect 30124 8716 30164 8756
rect 30508 8716 30548 8756
rect 31084 8707 31124 8747
rect 31564 8707 31604 8747
rect 31948 8716 31988 8756
rect 33196 8707 33236 8747
rect 34339 8716 34379 8756
rect 34444 8716 34484 8756
rect 34828 8716 34868 8756
rect 35404 8707 35444 8747
rect 35884 8707 35924 8747
rect 36748 8716 36788 8756
rect 37996 8707 38036 8747
rect 38380 8716 38420 8756
rect 39628 8707 39668 8747
rect 40291 8716 40331 8756
rect 40393 8716 40433 8756
rect 40780 8716 40820 8756
rect 41356 8707 41396 8747
rect 41836 8707 41876 8747
rect 1228 8632 1268 8672
rect 1612 8632 1652 8672
rect 2572 8632 2612 8672
rect 2812 8632 2852 8672
rect 3916 8632 3956 8672
rect 4156 8632 4196 8672
rect 10252 8632 10292 8672
rect 11308 8632 11348 8672
rect 18220 8632 18260 8672
rect 19948 8632 19988 8672
rect 21868 8632 21908 8672
rect 29116 8632 29156 8672
rect 29548 8632 29588 8672
rect 30604 8632 30644 8672
rect 34924 8632 34964 8672
rect 36115 8632 36155 8672
rect 36460 8632 36500 8672
rect 40876 8632 40916 8672
rect 42067 8632 42107 8672
rect 42412 8632 42452 8672
rect 42796 8632 42836 8672
rect 43372 8632 43412 8672
rect 43756 8632 43796 8672
rect 44092 8632 44132 8672
rect 44332 8632 44372 8672
rect 44716 8632 44756 8672
rect 44908 8632 44948 8672
rect 45148 8632 45188 8672
rect 7372 8548 7412 8588
rect 43996 8548 44036 8588
rect 1468 8464 1508 8504
rect 5740 8464 5780 8504
rect 7564 8464 7604 8504
rect 26668 8464 26708 8504
rect 28492 8464 28532 8504
rect 29788 8464 29828 8504
rect 38188 8464 38228 8504
rect 39820 8464 39860 8504
rect 43132 8464 43172 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 11644 8128 11684 8168
rect 12028 8128 12068 8168
rect 13756 8128 13796 8168
rect 15388 8128 15428 8168
rect 23164 8128 23204 8168
rect 34444 8128 34484 8168
rect 36268 8128 36308 8168
rect 37084 8128 37124 8168
rect 41692 8128 41732 8168
rect 42556 8128 42596 8168
rect 42940 8128 42980 8168
rect 43324 8128 43364 8168
rect 4204 8044 4244 8084
rect 10300 8035 10340 8075
rect 15004 8044 15044 8084
rect 26572 8044 26612 8084
rect 44092 8044 44132 8084
rect 1228 7960 1268 8000
rect 1612 7960 1652 8000
rect 6124 7960 6164 8000
rect 7779 7960 7819 8000
rect 8131 7960 8171 8000
rect 8524 7960 8564 8000
rect 11500 7960 11540 8000
rect 11884 7960 11924 8000
rect 12268 7960 12308 8000
rect 12460 7960 12500 8000
rect 13036 7960 13076 8000
rect 13516 7960 13556 8000
rect 13996 7960 14036 8000
rect 14236 7960 14276 8000
rect 14380 7960 14420 8000
rect 14764 7960 14804 8000
rect 15148 7960 15188 8000
rect 15724 7960 15764 8000
rect 15916 7960 15956 8000
rect 16300 7960 16340 8000
rect 18316 7960 18356 8000
rect 18700 7960 18740 8000
rect 19084 7960 19124 8000
rect 19756 7960 19796 8000
rect 20332 7960 20372 8000
rect 23404 7960 23444 8000
rect 23788 7960 23828 8000
rect 27436 7960 27476 8000
rect 28723 7960 28763 8000
rect 29068 7960 29108 8000
rect 29452 7960 29492 8000
rect 29836 7960 29876 8000
rect 30796 7960 30836 8000
rect 32083 7960 32123 8000
rect 32236 7960 32276 8000
rect 32812 7960 32852 8000
rect 36652 7960 36692 8000
rect 36844 7960 36884 8000
rect 38572 7960 38612 8000
rect 41932 7960 41972 8000
rect 42316 7960 42356 8000
rect 42700 7960 42740 8000
rect 43084 7960 43124 8000
rect 43660 7960 43700 8000
rect 44332 7960 44372 8000
rect 44524 7960 44564 8000
rect 44908 7960 44948 8000
rect 2764 7876 2804 7916
rect 4012 7876 4052 7916
rect 5155 7876 5195 7916
rect 5644 7876 5684 7916
rect 6220 7876 6260 7916
rect 6604 7876 6644 7916
rect 6717 7856 6757 7896
rect 6993 7876 7033 7916
rect 7110 7876 7150 7916
rect 7225 7909 7265 7949
rect 7324 7876 7364 7916
rect 7660 7876 7700 7916
rect 7891 7876 7931 7916
rect 7996 7876 8036 7916
rect 8236 7876 8276 7916
rect 9004 7876 9044 7916
rect 9292 7876 9332 7916
rect 9580 7876 9620 7916
rect 10060 7876 10100 7916
rect 10339 7876 10379 7916
rect 10732 7876 10772 7916
rect 10924 7876 10964 7916
rect 16684 7876 16724 7916
rect 17932 7876 17972 7916
rect 20716 7876 20756 7916
rect 21964 7876 22004 7916
rect 24172 7876 24212 7916
rect 25420 7876 25460 7916
rect 25900 7876 25940 7916
rect 26155 7876 26195 7916
rect 26275 7876 26315 7916
rect 26947 7876 26987 7916
rect 27052 7876 27092 7916
rect 27532 7876 27572 7916
rect 28012 7876 28052 7916
rect 28500 7876 28540 7916
rect 30307 7876 30347 7916
rect 30412 7876 30452 7916
rect 30892 7876 30932 7916
rect 31372 7876 31412 7916
rect 31891 7876 31931 7916
rect 33004 7876 33044 7916
rect 34252 7876 34292 7916
rect 34828 7876 34868 7916
rect 36076 7876 36116 7916
rect 37987 7876 38027 7916
rect 38092 7876 38132 7916
rect 38469 7876 38509 7916
rect 39052 7876 39092 7916
rect 39571 7876 39611 7916
rect 40108 7876 40148 7916
rect 41356 7876 41396 7916
rect 7564 7792 7604 7832
rect 8323 7792 8363 7832
rect 8764 7792 8804 7832
rect 9758 7792 9798 7832
rect 10828 7792 10868 7832
rect 14620 7792 14660 7832
rect 19324 7792 19364 7832
rect 25612 7792 25652 7832
rect 32476 7792 32516 7832
rect 44764 7792 44804 7832
rect 1468 7708 1508 7748
rect 1852 7708 1892 7748
rect 4972 7708 5012 7748
rect 7372 7708 7412 7748
rect 8860 7708 8900 7748
rect 9379 7708 9419 7748
rect 9859 7708 9899 7748
rect 9964 7708 10004 7748
rect 10531 7708 10571 7748
rect 11260 7708 11300 7748
rect 12700 7708 12740 7748
rect 13276 7708 13316 7748
rect 15484 7708 15524 7748
rect 16156 7708 16196 7748
rect 16540 7708 16580 7748
rect 18124 7708 18164 7748
rect 18556 7708 18596 7748
rect 18940 7708 18980 7748
rect 19996 7708 20036 7748
rect 20572 7708 20612 7748
rect 22156 7708 22196 7748
rect 24028 7708 24068 7748
rect 28828 7708 28868 7748
rect 29212 7708 29252 7748
rect 29596 7708 29636 7748
rect 32572 7708 32612 7748
rect 36412 7708 36452 7748
rect 39724 7708 39764 7748
rect 41548 7708 41588 7748
rect 43420 7708 43460 7748
rect 45148 7708 45188 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 5980 7372 6020 7412
rect 6307 7372 6347 7412
rect 6796 7372 6836 7412
rect 8515 7372 8555 7412
rect 10819 7372 10859 7412
rect 19276 7372 19316 7412
rect 23692 7372 23732 7412
rect 30220 7372 30260 7412
rect 31948 7372 31988 7412
rect 33148 7372 33188 7412
rect 37084 7372 37124 7412
rect 43996 7372 44036 7412
rect 7084 7288 7124 7328
rect 8620 7288 8660 7328
rect 9868 7288 9908 7328
rect 10627 7279 10667 7319
rect 27148 7288 27188 7328
rect 2188 7204 2228 7244
rect 3436 7195 3476 7235
rect 3820 7204 3860 7244
rect 5068 7195 5108 7235
rect 6124 7204 6164 7244
rect 6316 7204 6356 7244
rect 6508 7204 6548 7244
rect 6650 7204 6690 7244
rect 7180 7204 7220 7244
rect 7417 7204 7457 7244
rect 7651 7204 7691 7244
rect 8419 7204 8459 7244
rect 8730 7204 8770 7244
rect 9004 7204 9044 7244
rect 9139 7195 9179 7235
rect 9241 7204 9281 7244
rect 9484 7204 9524 7244
rect 9763 7204 9803 7244
rect 10339 7204 10379 7244
rect 10444 7195 10484 7235
rect 10731 7204 10771 7244
rect 10849 7193 10889 7233
rect 11063 7204 11103 7244
rect 11308 7204 11348 7244
rect 11596 7204 11636 7244
rect 12844 7195 12884 7235
rect 13708 7204 13748 7244
rect 14956 7195 14996 7235
rect 15532 7204 15572 7244
rect 16780 7195 16820 7235
rect 17539 7204 17579 7244
rect 17644 7204 17684 7244
rect 18028 7204 18068 7244
rect 18604 7195 18644 7235
rect 19084 7195 19124 7235
rect 19555 7204 19595 7244
rect 19660 7204 19700 7244
rect 20044 7204 20084 7244
rect 20620 7195 20660 7235
rect 21955 7237 21995 7277
rect 21100 7195 21140 7235
rect 22060 7204 22100 7244
rect 22444 7204 22484 7244
rect 23020 7195 23060 7235
rect 23500 7195 23540 7235
rect 24268 7195 24308 7235
rect 25516 7204 25556 7244
rect 27340 7195 27380 7235
rect 28588 7204 28628 7244
rect 28780 7204 28820 7244
rect 30028 7195 30068 7235
rect 30508 7204 30548 7244
rect 31756 7195 31796 7235
rect 33484 7195 33524 7235
rect 34732 7204 34772 7244
rect 38284 7195 38324 7235
rect 39532 7204 39572 7244
rect 40291 7204 40331 7244
rect 40396 7204 40436 7244
rect 40780 7204 40820 7244
rect 41356 7195 41396 7235
rect 41836 7195 41876 7235
rect 1228 7120 1268 7160
rect 1612 7120 1652 7160
rect 5740 7120 5780 7160
rect 7299 7120 7339 7160
rect 8044 7120 8084 7160
rect 8284 7120 8324 7160
rect 8908 7120 8948 7160
rect 11203 7120 11243 7160
rect 11404 7120 11444 7160
rect 13324 7120 13364 7160
rect 18124 7120 18164 7160
rect 20140 7120 20180 7160
rect 21331 7120 21371 7160
rect 21484 7120 21524 7160
rect 22540 7120 22580 7160
rect 26188 7120 26228 7160
rect 32332 7120 32372 7160
rect 32716 7120 32756 7160
rect 32908 7120 32948 7160
rect 34924 7120 34964 7160
rect 36460 7120 36500 7160
rect 36844 7120 36884 7160
rect 37420 7120 37460 7160
rect 40012 7120 40052 7160
rect 40876 7120 40916 7160
rect 42067 7120 42107 7160
rect 42412 7120 42452 7160
rect 43372 7120 43412 7160
rect 43756 7120 43796 7160
rect 44140 7120 44180 7160
rect 44524 7120 44564 7160
rect 44908 7120 44948 7160
rect 45148 7120 45188 7160
rect 3628 7036 3668 7076
rect 7623 7036 7663 7076
rect 10156 7036 10196 7076
rect 15148 7036 15188 7076
rect 16972 7036 17012 7076
rect 21724 7036 21764 7076
rect 33292 7036 33332 7076
rect 42172 7036 42212 7076
rect 43612 7036 43652 7076
rect 44380 7036 44420 7076
rect 1468 6952 1508 6992
rect 1852 6952 1892 6992
rect 5260 6952 5300 6992
rect 7843 6952 7883 6992
rect 13036 6952 13076 6992
rect 13564 6952 13604 6992
rect 24076 6952 24116 6992
rect 25948 6952 25988 6992
rect 32092 6952 32132 6992
rect 32476 6952 32516 6992
rect 35164 6952 35204 6992
rect 36700 6952 36740 6992
rect 37180 6952 37220 6992
rect 38092 6952 38132 6992
rect 39772 6952 39812 6992
rect 44764 6952 44804 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 6547 6616 6587 6656
rect 8419 6616 8459 6656
rect 16492 6616 16532 6656
rect 23692 6616 23732 6656
rect 26764 6616 26804 6656
rect 28348 6616 28388 6656
rect 29020 6616 29060 6656
rect 30364 6616 30404 6656
rect 40396 6616 40436 6656
rect 44380 6616 44420 6656
rect 1468 6532 1508 6572
rect 7468 6532 7508 6572
rect 17308 6532 17348 6572
rect 20956 6532 20996 6572
rect 40684 6532 40724 6572
rect 1228 6448 1268 6488
rect 1612 6448 1652 6488
rect 1996 6448 2036 6488
rect 4492 6448 4532 6488
rect 5260 6448 5300 6488
rect 9292 6448 9332 6488
rect 9484 6448 9524 6488
rect 10531 6448 10571 6488
rect 10732 6448 10772 6488
rect 16684 6448 16724 6488
rect 17068 6448 17108 6488
rect 17548 6448 17588 6488
rect 17788 6448 17828 6488
rect 18508 6448 18548 6488
rect 19795 6448 19835 6488
rect 19948 6448 19988 6488
rect 20524 6448 20564 6488
rect 20716 6448 20756 6488
rect 21436 6448 21476 6488
rect 21676 6448 21716 6488
rect 21868 6448 21908 6488
rect 25708 6448 25748 6488
rect 28588 6448 28628 6488
rect 28780 6448 28820 6488
rect 29356 6448 29396 6488
rect 29740 6448 29780 6488
rect 30124 6448 30164 6488
rect 38380 6448 38420 6488
rect 44140 6448 44180 6488
rect 44524 6448 44564 6488
rect 44908 6448 44948 6488
rect 45148 6448 45188 6488
rect 2668 6364 2708 6404
rect 3916 6364 3956 6404
rect 4771 6364 4811 6404
rect 4876 6364 4916 6404
rect 5356 6364 5396 6404
rect 5836 6364 5876 6404
rect 6355 6364 6395 6404
rect 6796 6364 6836 6404
rect 7075 6364 7115 6404
rect 7676 6375 7716 6415
rect 7843 6364 7883 6404
rect 7987 6364 8027 6404
rect 8127 6364 8167 6404
rect 8233 6364 8273 6404
rect 8716 6364 8756 6404
rect 9580 6364 9620 6404
rect 9699 6364 9739 6404
rect 9817 6364 9857 6404
rect 10116 6364 10156 6404
rect 10252 6364 10292 6404
rect 10391 6364 10431 6404
rect 10636 6364 10676 6404
rect 10924 6364 10964 6404
rect 11066 6364 11106 6404
rect 11788 6364 11828 6404
rect 13036 6364 13076 6404
rect 13420 6364 13460 6404
rect 14668 6364 14708 6404
rect 15052 6364 15092 6404
rect 16300 6364 16340 6404
rect 18019 6364 18059 6404
rect 18124 6364 18164 6404
rect 18604 6364 18644 6404
rect 19084 6364 19124 6404
rect 19603 6364 19643 6404
rect 22252 6364 22292 6404
rect 23500 6364 23540 6404
rect 26952 6364 26992 6404
rect 28204 6364 28244 6404
rect 30892 6364 30932 6404
rect 32140 6364 32180 6404
rect 32524 6364 32564 6404
rect 33772 6364 33812 6404
rect 33964 6364 34004 6404
rect 35212 6364 35252 6404
rect 35596 6364 35636 6404
rect 36844 6364 36884 6404
rect 38956 6364 38996 6404
rect 40204 6364 40244 6404
rect 4108 6280 4148 6320
rect 7180 6280 7220 6320
rect 8414 6280 8454 6320
rect 9052 6280 9092 6320
rect 16924 6280 16964 6320
rect 20188 6280 20228 6320
rect 22108 6280 22148 6320
rect 29116 6280 29156 6320
rect 1852 6196 1892 6236
rect 2236 6196 2276 6236
rect 4252 6196 4292 6236
rect 7747 6196 7787 6236
rect 8620 6196 8660 6236
rect 9955 6196 9995 6236
rect 11212 6196 11252 6236
rect 11596 6196 11636 6236
rect 14860 6196 14900 6236
rect 20284 6196 20324 6236
rect 25948 6196 25988 6236
rect 29500 6196 29540 6236
rect 30700 6196 30740 6236
rect 32332 6196 32372 6236
rect 35404 6196 35444 6236
rect 37036 6196 37076 6236
rect 38620 6196 38660 6236
rect 44764 6196 44804 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 5356 5860 5396 5900
rect 11692 5860 11732 5900
rect 16972 5860 17012 5900
rect 35596 5860 35636 5900
rect 1468 5776 1508 5816
rect 6844 5776 6884 5816
rect 11116 5776 11156 5816
rect 36460 5776 36500 5816
rect 39715 5776 39755 5816
rect 45148 5776 45188 5816
rect 2284 5692 2324 5732
rect 3532 5683 3572 5723
rect 3916 5692 3956 5732
rect 5164 5683 5204 5723
rect 5644 5692 5684 5732
rect 5875 5692 5915 5732
rect 5995 5692 6035 5732
rect 6220 5692 6260 5732
rect 6508 5692 6548 5732
rect 6647 5692 6687 5732
rect 7171 5692 7211 5732
rect 7660 5683 7700 5723
rect 8140 5692 8180 5732
rect 8620 5692 8660 5732
rect 8721 5692 8761 5732
rect 10732 5692 10772 5732
rect 11007 5692 11047 5732
rect 11884 5683 11924 5723
rect 13132 5692 13172 5732
rect 13324 5692 13364 5732
rect 14572 5683 14612 5723
rect 15235 5692 15275 5732
rect 15340 5692 15380 5732
rect 15724 5692 15764 5732
rect 16300 5683 16340 5723
rect 16780 5683 16820 5723
rect 17164 5692 17204 5732
rect 18412 5683 18452 5723
rect 18892 5692 18932 5732
rect 1228 5608 1268 5648
rect 1612 5608 1652 5648
rect 5548 5608 5588 5648
rect 5779 5599 5819 5639
rect 6115 5608 6155 5648
rect 6316 5608 6356 5648
rect 8236 5608 8276 5648
rect 9292 5608 9332 5648
rect 9484 5608 9524 5648
rect 10060 5608 10100 5648
rect 10492 5608 10532 5648
rect 20148 5650 20188 5690
rect 22156 5683 22196 5723
rect 23404 5692 23444 5732
rect 23596 5692 23636 5732
rect 24844 5683 24884 5723
rect 25411 5692 25451 5732
rect 25516 5692 25556 5732
rect 25900 5692 25940 5732
rect 26476 5683 26516 5723
rect 26956 5683 26996 5723
rect 30595 5692 30635 5732
rect 30700 5692 30740 5732
rect 31084 5692 31124 5732
rect 31660 5683 31700 5723
rect 32140 5683 32180 5723
rect 33859 5692 33899 5732
rect 33964 5692 34004 5732
rect 34348 5692 34388 5732
rect 34924 5683 34964 5723
rect 35404 5683 35444 5723
rect 36076 5692 36116 5732
rect 36355 5692 36395 5732
rect 36940 5692 36980 5732
rect 38188 5683 38228 5723
rect 40099 5692 40139 5732
rect 15820 5608 15860 5648
rect 20524 5608 20564 5648
rect 21196 5608 21236 5648
rect 21580 5608 21620 5648
rect 21955 5608 21995 5648
rect 25996 5608 26036 5648
rect 27724 5608 27764 5648
rect 27916 5608 27956 5648
rect 28492 5608 28532 5648
rect 28876 5608 28916 5648
rect 29260 5608 29300 5648
rect 29644 5608 29684 5648
rect 30220 5608 30260 5648
rect 31180 5608 31220 5648
rect 32524 5608 32564 5648
rect 33100 5608 33140 5648
rect 33484 5608 33524 5648
rect 34444 5608 34484 5648
rect 38764 5608 38804 5648
rect 38956 5608 38996 5648
rect 44524 5608 44564 5648
rect 44908 5608 44948 5648
rect 3724 5524 3764 5564
rect 9724 5524 9764 5564
rect 25036 5524 25076 5564
rect 27196 5524 27236 5564
rect 28156 5524 28196 5564
rect 32380 5524 32420 5564
rect 32860 5524 32900 5564
rect 36748 5524 36788 5564
rect 42028 5524 42068 5564
rect 44764 5524 44804 5564
rect 1852 5440 1892 5480
rect 6940 5440 6980 5480
rect 9052 5440 9092 5480
rect 9820 5440 9860 5480
rect 10204 5440 10244 5480
rect 11404 5440 11444 5480
rect 14764 5440 14804 5480
rect 18604 5440 18644 5480
rect 20332 5440 20372 5480
rect 20764 5440 20804 5480
rect 21436 5440 21476 5480
rect 21820 5440 21860 5480
rect 27484 5440 27524 5480
rect 28252 5440 28292 5480
rect 28636 5440 28676 5480
rect 29020 5440 29060 5480
rect 29404 5440 29444 5480
rect 29980 5440 30020 5480
rect 32764 5440 32804 5480
rect 33244 5440 33284 5480
rect 38380 5440 38420 5480
rect 38524 5440 38564 5480
rect 39196 5440 39236 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 1852 5104 1892 5144
rect 3196 5104 3236 5144
rect 5548 5104 5588 5144
rect 6604 5104 6644 5144
rect 11443 5104 11483 5144
rect 12412 5104 12452 5144
rect 26956 5104 26996 5144
rect 30067 5104 30107 5144
rect 31660 5104 31700 5144
rect 34060 5104 34100 5144
rect 39292 5104 39332 5144
rect 45148 5104 45188 5144
rect 18412 5020 18452 5060
rect 23116 5020 23156 5060
rect 1228 4936 1268 4976
rect 1612 4936 1652 4976
rect 2572 4936 2612 4976
rect 2956 4936 2996 4976
rect 6220 4936 6260 4976
rect 8716 4936 8756 4976
rect 10156 4936 10196 4976
rect 11788 4936 11828 4976
rect 12172 4936 12212 4976
rect 13132 4936 13172 4976
rect 15340 4936 15380 4976
rect 19180 4936 19220 4976
rect 23500 4936 23540 4976
rect 27340 4936 27380 4976
rect 27724 4936 27764 4976
rect 28780 4936 28820 4976
rect 32044 4936 32084 4976
rect 32428 4936 32468 4976
rect 36172 4936 36212 4976
rect 36364 4936 36404 4976
rect 36940 4936 36980 4976
rect 37900 4936 37940 4976
rect 39187 4936 39227 4976
rect 39532 4936 39572 4976
rect 44524 4936 44564 4976
rect 44908 4936 44948 4976
rect 3724 4852 3764 4892
rect 3916 4852 3956 4892
rect 4108 4852 4148 4892
rect 5356 4852 5396 4892
rect 5836 4852 5876 4892
rect 5955 4852 5995 4892
rect 6073 4852 6113 4892
rect 6892 4852 6932 4892
rect 7027 4843 7067 4883
rect 7276 4852 7316 4892
rect 7747 4852 7787 4892
rect 8236 4852 8276 4892
rect 8812 4852 8852 4892
rect 9196 4852 9236 4892
rect 9297 4851 9337 4891
rect 9667 4852 9707 4892
rect 9772 4852 9812 4892
rect 10252 4852 10292 4892
rect 10732 4852 10772 4892
rect 11220 4852 11260 4892
rect 12643 4852 12683 4892
rect 12748 4852 12788 4892
rect 13228 4852 13268 4892
rect 13708 4852 13748 4892
rect 14227 4852 14267 4892
rect 14851 4852 14891 4892
rect 14956 4852 14996 4892
rect 15436 4852 15476 4892
rect 15916 4852 15956 4892
rect 16404 4852 16444 4892
rect 16972 4852 17012 4892
rect 18220 4852 18260 4892
rect 18691 4852 18731 4892
rect 18796 4852 18836 4892
rect 19276 4852 19316 4892
rect 19756 4852 19796 4892
rect 20275 4852 20315 4892
rect 20467 4852 20507 4892
rect 20716 4852 20756 4892
rect 21964 4852 22004 4892
rect 22444 4852 22484 4892
rect 22723 4852 22763 4892
rect 23980 4852 24020 4892
rect 25228 4852 25268 4892
rect 25516 4852 25556 4892
rect 26764 4852 26804 4892
rect 28291 4852 28331 4892
rect 28396 4852 28436 4892
rect 28876 4852 28916 4892
rect 29356 4852 29396 4892
rect 29875 4852 29915 4892
rect 30220 4852 30260 4892
rect 31476 4852 31516 4892
rect 32620 4852 32660 4892
rect 33868 4852 33908 4892
rect 34348 4852 34388 4892
rect 35604 4852 35644 4892
rect 37411 4852 37451 4892
rect 37516 4852 37556 4892
rect 37996 4852 38036 4892
rect 38476 4852 38516 4892
rect 38964 4852 39004 4892
rect 40291 4852 40331 4892
rect 7555 4768 7595 4808
rect 22156 4768 22196 4808
rect 22828 4768 22868 4808
rect 23788 4768 23828 4808
rect 32188 4768 32228 4808
rect 35788 4768 35828 4808
rect 36604 4768 36644 4808
rect 39907 4768 39947 4808
rect 44764 4768 44804 4808
rect 1468 4684 1508 4724
rect 2812 4684 2852 4724
rect 3907 4684 3947 4724
rect 5740 4684 5780 4724
rect 6460 4684 6500 4724
rect 12028 4684 12068 4724
rect 14380 4684 14420 4724
rect 16588 4684 16628 4724
rect 23260 4684 23300 4724
rect 27100 4684 27140 4724
rect 27484 4684 27524 4724
rect 31804 4684 31844 4724
rect 35932 4684 35972 4724
rect 36700 4684 36740 4724
rect 42220 4684 42260 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 5827 4348 5867 4388
rect 6499 4348 6539 4388
rect 7276 4348 7316 4388
rect 11308 4348 11348 4388
rect 14668 4348 14708 4388
rect 16300 4348 16340 4388
rect 22972 4348 23012 4388
rect 25660 4348 25700 4388
rect 28108 4348 28148 4388
rect 30028 4348 30068 4388
rect 33004 4348 33044 4388
rect 37900 4348 37940 4388
rect 38044 4348 38084 4388
rect 2524 4264 2564 4304
rect 5260 4264 5300 4304
rect 6115 4264 6155 4304
rect 6220 4264 6260 4304
rect 9331 4264 9371 4304
rect 11932 4264 11972 4304
rect 18028 4264 18068 4304
rect 38428 4264 38468 4304
rect 40156 4264 40196 4304
rect 45148 4264 45188 4304
rect 3052 4180 3092 4220
rect 4300 4171 4340 4211
rect 5059 4180 5099 4220
rect 5356 4180 5396 4220
rect 5495 4180 5535 4220
rect 5635 4180 5675 4220
rect 5740 4180 5780 4220
rect 6017 4180 6057 4220
rect 6316 4171 6356 4211
rect 6660 4180 6700 4220
rect 6796 4180 6836 4220
rect 7027 4180 7067 4220
rect 7130 4180 7170 4220
rect 7555 4180 7595 4220
rect 7660 4180 7700 4220
rect 8044 4180 8084 4220
rect 8620 4171 8660 4211
rect 9100 4171 9140 4211
rect 9571 4180 9611 4220
rect 9681 4180 9721 4220
rect 10060 4180 10100 4220
rect 10636 4171 10676 4211
rect 11116 4171 11156 4211
rect 13228 4180 13268 4220
rect 14476 4171 14516 4211
rect 14860 4180 14900 4220
rect 16108 4159 16148 4199
rect 16588 4180 16628 4220
rect 17836 4171 17876 4211
rect 18595 4180 18635 4220
rect 18700 4180 18740 4220
rect 19084 4180 19124 4220
rect 19660 4171 19700 4211
rect 20140 4171 20180 4211
rect 20803 4180 20843 4220
rect 20908 4180 20948 4220
rect 21292 4180 21332 4220
rect 21868 4171 21908 4211
rect 22387 4180 22427 4220
rect 22579 4180 22619 4220
rect 26668 4180 26708 4220
rect 27916 4171 27956 4211
rect 28588 4180 28628 4220
rect 29836 4171 29876 4211
rect 31267 4180 31307 4220
rect 31372 4180 31412 4220
rect 31756 4180 31796 4220
rect 32332 4171 32372 4211
rect 32812 4171 32852 4211
rect 33759 4180 33799 4220
rect 33868 4180 33908 4220
rect 34252 4180 34292 4220
rect 34828 4171 34868 4211
rect 35308 4171 35348 4211
rect 36460 4180 36500 4220
rect 37708 4171 37748 4211
rect 1228 4096 1268 4136
rect 1612 4096 1652 4136
rect 2284 4096 2324 4136
rect 2668 4096 2708 4136
rect 4684 4096 4724 4136
rect 8140 4096 8180 4136
rect 10156 4096 10196 4136
rect 11692 4096 11732 4136
rect 12076 4096 12116 4136
rect 12460 4096 12500 4136
rect 12883 4096 12923 4136
rect 19180 4096 19220 4136
rect 21388 4096 21428 4136
rect 22732 4096 22772 4136
rect 23308 4096 23348 4136
rect 23788 4096 23828 4136
rect 24172 4096 24212 4136
rect 24844 4096 24884 4136
rect 25036 4096 25076 4136
rect 25420 4096 25460 4136
rect 25996 4096 26036 4136
rect 26380 4096 26420 4136
rect 30412 4096 30452 4136
rect 30796 4096 30836 4136
rect 31852 4096 31892 4136
rect 33388 4096 33428 4136
rect 34348 4096 34388 4136
rect 35884 4096 35924 4136
rect 36268 4096 36308 4136
rect 38284 4096 38324 4136
rect 38668 4096 38708 4136
rect 38860 4096 38900 4136
rect 39724 4096 39764 4136
rect 40396 4096 40436 4136
rect 44140 4096 44180 4136
rect 44524 4096 44564 4136
rect 44908 4096 44948 4136
rect 4492 4012 4532 4052
rect 12316 4012 12356 4052
rect 13084 4012 13124 4052
rect 25276 4012 25316 4052
rect 33148 4012 33188 4052
rect 35548 4012 35588 4052
rect 39100 4012 39140 4052
rect 40972 4012 41012 4052
rect 44764 4012 44804 4052
rect 1468 3928 1508 3968
rect 1852 3928 1892 3968
rect 2908 3928 2948 3968
rect 4924 3928 4964 3968
rect 12700 3928 12740 3968
rect 20371 3928 20411 3968
rect 23068 3928 23108 3968
rect 23548 3928 23588 3968
rect 23932 3928 23972 3968
rect 24604 3928 24644 3968
rect 25756 3928 25796 3968
rect 26140 3928 26180 3968
rect 30172 3928 30212 3968
rect 30556 3928 30596 3968
rect 35644 3928 35684 3968
rect 36028 3928 36068 3968
rect 39964 3928 40004 3968
rect 44380 3928 44420 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 3100 3592 3140 3632
rect 8476 3592 8516 3632
rect 9148 3592 9188 3632
rect 9532 3592 9572 3632
rect 19900 3592 19940 3632
rect 23932 3592 23972 3632
rect 32140 3592 32180 3632
rect 33772 3592 33812 3632
rect 35836 3592 35876 3632
rect 36604 3592 36644 3632
rect 39052 3592 39092 3632
rect 45148 3592 45188 3632
rect 15292 3508 15332 3548
rect 18364 3508 18404 3548
rect 26956 3508 26996 3548
rect 37132 3508 37172 3548
rect 41452 3508 41492 3548
rect 1228 3424 1268 3464
rect 1468 3424 1508 3464
rect 1651 3424 1691 3464
rect 1996 3424 2036 3464
rect 2380 3424 2420 3464
rect 2860 3424 2900 3464
rect 5203 3415 5243 3455
rect 5683 3415 5723 3455
rect 7084 3424 7124 3464
rect 8140 3424 8180 3464
rect 8716 3424 8756 3464
rect 8908 3424 8948 3464
rect 9292 3424 9332 3464
rect 10828 3424 10868 3464
rect 12268 3424 12308 3464
rect 13900 3424 13940 3464
rect 14284 3424 14324 3464
rect 14668 3424 14708 3464
rect 15052 3424 15092 3464
rect 17356 3424 17396 3464
rect 17932 3424 17972 3464
rect 18124 3424 18164 3464
rect 18508 3424 18548 3464
rect 18892 3424 18932 3464
rect 19315 3424 19355 3464
rect 19660 3424 19700 3464
rect 20044 3424 20084 3464
rect 23692 3424 23732 3464
rect 24556 3424 24596 3464
rect 26668 3424 26708 3464
rect 28780 3424 28820 3464
rect 36076 3424 36116 3464
rect 36460 3424 36500 3464
rect 36844 3424 36884 3464
rect 41596 3424 41636 3464
rect 41836 3424 41876 3464
rect 44524 3424 44564 3464
rect 44908 3424 44948 3464
rect 3244 3340 3284 3380
rect 4492 3340 4532 3380
rect 5068 3340 5108 3380
rect 5305 3340 5345 3380
rect 5548 3340 5588 3380
rect 5785 3340 5825 3380
rect 6115 3340 6155 3380
rect 6604 3340 6644 3380
rect 7180 3340 7220 3380
rect 7564 3340 7604 3380
rect 7682 3340 7722 3380
rect 9859 3340 9899 3380
rect 10348 3340 10388 3380
rect 10924 3340 10964 3380
rect 11308 3340 11348 3380
rect 11426 3340 11466 3380
rect 11779 3340 11819 3380
rect 11884 3340 11924 3380
rect 12364 3340 12404 3380
rect 12844 3340 12884 3380
rect 13363 3340 13403 3380
rect 15436 3340 15476 3380
rect 16684 3340 16724 3380
rect 20428 3340 20468 3380
rect 21676 3340 21716 3380
rect 22060 3340 22100 3380
rect 23308 3340 23348 3380
rect 24844 3340 24884 3380
rect 26092 3340 26132 3380
rect 27148 3340 27188 3380
rect 28396 3340 28436 3380
rect 29068 3340 29108 3380
rect 30316 3340 30356 3380
rect 30700 3340 30740 3380
rect 31948 3340 31988 3380
rect 32332 3340 32372 3380
rect 33580 3340 33620 3380
rect 34284 3340 34324 3380
rect 35500 3340 35540 3380
rect 37324 3340 37364 3380
rect 38572 3340 38612 3380
rect 39244 3340 39284 3380
rect 40492 3340 40532 3380
rect 40780 3340 40820 3380
rect 41059 3340 41099 3380
rect 1852 3256 1892 3296
rect 2620 3256 2660 3296
rect 4684 3256 4724 3296
rect 5452 3256 5492 3296
rect 8380 3256 8420 3296
rect 9667 3256 9707 3296
rect 17596 3256 17636 3296
rect 23500 3256 23540 3296
rect 41164 3256 41204 3296
rect 2236 3172 2276 3212
rect 4972 3172 5012 3212
rect 5932 3172 5972 3212
rect 13516 3172 13556 3212
rect 14140 3172 14180 3212
rect 14524 3172 14564 3212
rect 14908 3172 14948 3212
rect 16876 3172 16916 3212
rect 17692 3172 17732 3212
rect 18748 3172 18788 3212
rect 19132 3172 19172 3212
rect 19516 3172 19556 3212
rect 20284 3172 20324 3212
rect 21868 3172 21908 3212
rect 24316 3172 24356 3212
rect 26284 3172 26324 3212
rect 26428 3172 26468 3212
rect 28540 3172 28580 3212
rect 30508 3172 30548 3212
rect 35692 3172 35732 3212
rect 36220 3172 36260 3212
rect 44764 3172 44804 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 2332 2836 2372 2876
rect 2716 2836 2756 2876
rect 3484 2836 3524 2876
rect 6691 2836 6731 2876
rect 7180 2836 7220 2876
rect 10636 2836 10676 2876
rect 13708 2836 13748 2876
rect 17356 2836 17396 2876
rect 20140 2836 20180 2876
rect 23212 2836 23252 2876
rect 25804 2836 25844 2876
rect 29836 2836 29876 2876
rect 31948 2836 31988 2876
rect 35788 2836 35828 2876
rect 38044 2836 38084 2876
rect 40252 2836 40292 2876
rect 40924 2836 40964 2876
rect 8812 2752 8852 2792
rect 10444 2752 10484 2792
rect 15340 2752 15380 2792
rect 17788 2752 17828 2792
rect 27820 2752 27860 2792
rect 36460 2752 36500 2792
rect 40108 2752 40148 2792
rect 45148 2752 45188 2792
rect 4780 2668 4820 2708
rect 6028 2659 6068 2699
rect 6359 2668 6399 2708
rect 6604 2668 6644 2708
rect 6892 2668 6932 2708
rect 7034 2668 7074 2708
rect 7372 2668 7412 2708
rect 8620 2659 8660 2699
rect 9004 2668 9044 2708
rect 10252 2659 10292 2699
rect 10828 2659 10868 2699
rect 12036 2668 12076 2708
rect 12256 2668 12296 2708
rect 13516 2659 13556 2699
rect 13900 2668 13940 2708
rect 15148 2659 15188 2699
rect 15619 2668 15659 2708
rect 15724 2668 15764 2708
rect 16108 2668 16148 2708
rect 16684 2659 16724 2699
rect 17164 2659 17204 2699
rect 18403 2668 18443 2708
rect 18508 2668 18548 2708
rect 18892 2668 18932 2708
rect 19468 2659 19508 2699
rect 19948 2659 19988 2699
rect 21475 2668 21515 2708
rect 21580 2668 21620 2708
rect 21964 2668 22004 2708
rect 22540 2659 22580 2699
rect 23020 2659 23060 2699
rect 24067 2668 24107 2708
rect 24172 2668 24212 2708
rect 24556 2668 24596 2708
rect 25132 2659 25172 2699
rect 25612 2659 25652 2699
rect 26380 2668 26420 2708
rect 27628 2659 27668 2699
rect 28099 2668 28139 2708
rect 28204 2668 28244 2708
rect 28588 2668 28628 2708
rect 29164 2659 29204 2699
rect 29644 2659 29684 2699
rect 30211 2668 30251 2708
rect 30316 2668 30356 2708
rect 30700 2668 30740 2708
rect 1228 2584 1268 2624
rect 1612 2584 1652 2624
rect 1852 2584 1892 2624
rect 2092 2584 2132 2624
rect 2476 2584 2516 2624
rect 2860 2584 2900 2624
rect 3244 2584 3284 2624
rect 3628 2584 3668 2624
rect 4012 2584 4052 2624
rect 4396 2584 4436 2624
rect 6499 2584 6539 2624
rect 16204 2584 16244 2624
rect 17548 2584 17588 2624
rect 17932 2584 17972 2624
rect 18988 2584 19028 2624
rect 20620 2584 20660 2624
rect 21004 2584 21044 2624
rect 22060 2584 22100 2624
rect 23596 2584 23636 2624
rect 24652 2584 24692 2624
rect 26188 2584 26228 2624
rect 28684 2584 28724 2624
rect 30796 2584 30836 2624
rect 31276 2626 31316 2666
rect 31756 2659 31796 2699
rect 32332 2668 32372 2708
rect 33588 2668 33628 2708
rect 34051 2668 34091 2708
rect 34156 2668 34196 2708
rect 34540 2668 34580 2708
rect 35116 2659 35156 2699
rect 35596 2659 35636 2699
rect 36652 2659 36692 2699
rect 37900 2668 37940 2708
rect 38668 2668 38708 2708
rect 39916 2659 39956 2699
rect 34636 2584 34676 2624
rect 36172 2584 36212 2624
rect 38284 2584 38324 2624
rect 40492 2584 40532 2624
rect 40684 2584 40724 2624
rect 44140 2584 44180 2624
rect 44524 2584 44564 2624
rect 44908 2584 44948 2624
rect 1468 2500 1508 2540
rect 3868 2500 3908 2540
rect 6220 2500 6260 2540
rect 20860 2500 20900 2540
rect 44764 2500 44804 2540
rect 3100 2416 3140 2456
rect 4252 2416 4292 2456
rect 4636 2416 4676 2456
rect 18172 2416 18212 2456
rect 21244 2416 21284 2456
rect 23836 2416 23876 2456
rect 25948 2416 25988 2456
rect 33772 2416 33812 2456
rect 35932 2416 35972 2456
rect 44380 2416 44420 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 1468 2080 1508 2120
rect 2236 2080 2276 2120
rect 3292 2080 3332 2120
rect 4444 2080 4484 2120
rect 4828 2080 4868 2120
rect 6412 2080 6452 2120
rect 6940 2080 6980 2120
rect 7612 2080 7652 2120
rect 12076 2080 12116 2120
rect 12892 2080 12932 2120
rect 13276 2080 13316 2120
rect 13660 2080 13700 2120
rect 15244 2080 15284 2120
rect 15676 2080 15716 2120
rect 16060 2080 16100 2120
rect 16444 2080 16484 2120
rect 18412 2080 18452 2120
rect 20044 2080 20084 2120
rect 20668 2080 20708 2120
rect 23020 2080 23060 2120
rect 26707 2080 26747 2120
rect 29164 2080 29204 2120
rect 32044 2080 32084 2120
rect 36019 2080 36059 2120
rect 38764 2080 38804 2120
rect 45148 2080 45188 2120
rect 1852 1996 1892 2036
rect 6556 1996 6596 2036
rect 7996 1996 8036 2036
rect 10492 1996 10532 2036
rect 1228 1912 1268 1952
rect 1612 1912 1652 1952
rect 1996 1912 2036 1952
rect 2668 1912 2708 1952
rect 3052 1912 3092 1952
rect 3436 1912 3476 1952
rect 3820 1912 3860 1952
rect 4204 1912 4244 1952
rect 4627 1912 4667 1952
rect 6796 1912 6836 1952
rect 7180 1912 7220 1952
rect 7372 1912 7412 1952
rect 7756 1912 7796 1952
rect 8140 1912 8180 1952
rect 10252 1912 10292 1952
rect 12268 1912 12308 1952
rect 12508 1912 12548 1952
rect 12652 1912 12692 1952
rect 13036 1912 13076 1952
rect 13420 1912 13460 1952
rect 15436 1912 15476 1952
rect 15820 1912 15860 1952
rect 16204 1912 16244 1952
rect 16588 1912 16628 1952
rect 20428 1912 20468 1952
rect 20812 1912 20852 1952
rect 21196 1912 21236 1952
rect 25420 1912 25460 1952
rect 27052 1912 27092 1952
rect 27436 1912 27476 1952
rect 29308 1912 29348 1952
rect 29548 1912 29588 1952
rect 29932 1912 29972 1952
rect 30316 1912 30356 1952
rect 32428 1912 32468 1952
rect 32812 1912 32852 1952
rect 33196 1912 33236 1952
rect 33580 1912 33620 1952
rect 33964 1912 34004 1952
rect 34828 1912 34868 1952
rect 38284 1912 38324 1952
rect 43756 1912 43796 1952
rect 44140 1912 44180 1952
rect 44524 1912 44564 1952
rect 44908 1912 44948 1952
rect 4972 1828 5012 1868
rect 6220 1828 6260 1868
rect 8524 1828 8564 1868
rect 9772 1828 9812 1868
rect 10636 1828 10676 1868
rect 11884 1828 11924 1868
rect 13804 1828 13844 1868
rect 15052 1828 15092 1868
rect 16972 1828 17012 1868
rect 18220 1828 18260 1868
rect 18604 1828 18644 1868
rect 19852 1828 19892 1868
rect 21580 1828 21620 1868
rect 22828 1828 22868 1868
rect 23212 1828 23252 1868
rect 24460 1828 24500 1868
rect 24931 1828 24971 1868
rect 25036 1828 25076 1868
rect 25516 1828 25556 1868
rect 25996 1828 26036 1868
rect 26484 1828 26524 1868
rect 27724 1828 27764 1868
rect 28972 1828 29012 1868
rect 30604 1828 30644 1868
rect 31852 1828 31892 1868
rect 34243 1828 34283 1868
rect 34348 1828 34388 1868
rect 34732 1828 34772 1868
rect 35308 1828 35348 1868
rect 35827 1828 35867 1868
rect 36652 1828 36692 1868
rect 37900 1828 37940 1868
rect 38956 1828 38996 1868
rect 40204 1828 40244 1868
rect 2908 1744 2948 1784
rect 9964 1744 10004 1784
rect 24652 1744 24692 1784
rect 36460 1744 36500 1784
rect 43996 1744 44036 1784
rect 44764 1744 44804 1784
rect 3676 1660 3716 1700
rect 4060 1660 4100 1700
rect 8380 1660 8420 1700
rect 16828 1660 16868 1700
rect 21052 1660 21092 1700
rect 21436 1660 21476 1700
rect 26812 1660 26852 1700
rect 27196 1660 27236 1700
rect 29692 1660 29732 1700
rect 30076 1660 30116 1700
rect 32188 1660 32228 1700
rect 32572 1660 32612 1700
rect 32956 1660 32996 1700
rect 33340 1660 33380 1700
rect 33724 1660 33764 1700
rect 38044 1660 38084 1700
rect 44380 1660 44420 1700
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
<< metal2 >>
rect 32515 11656 32524 11696
rect 32564 11656 42508 11696
rect 42548 11656 42557 11696
rect 35587 11572 35596 11612
rect 35636 11572 42316 11612
rect 42356 11572 42365 11612
rect 37507 11488 37516 11528
rect 37556 11488 44524 11528
rect 44564 11488 44573 11528
rect 35683 11404 35692 11444
rect 35732 11404 44716 11444
rect 44756 11404 44765 11444
rect 32611 11320 32620 11360
rect 32660 11320 39092 11360
rect 39052 11276 39092 11320
rect 42412 11320 44332 11360
rect 44372 11320 44381 11360
rect 42412 11276 42452 11320
rect 16963 11236 16972 11276
rect 17012 11236 38956 11276
rect 38996 11236 39005 11276
rect 39052 11236 42452 11276
rect 0 11192 90 11212
rect 46278 11192 46368 11212
rect 0 11152 76 11192
rect 116 11152 125 11192
rect 34915 11152 34924 11192
rect 34964 11152 43700 11192
rect 44995 11152 45004 11192
rect 45044 11152 46368 11192
rect 0 11132 90 11152
rect 43660 11108 43700 11152
rect 46278 11132 46368 11152
rect 1987 11068 1996 11108
rect 2036 11068 14476 11108
rect 14516 11068 14525 11108
rect 37795 11068 37804 11108
rect 37844 11068 42124 11108
rect 42164 11068 42173 11108
rect 42307 11068 42316 11108
rect 42356 11068 43564 11108
rect 43604 11068 43613 11108
rect 43660 11068 45100 11108
rect 45140 11068 45149 11108
rect 11491 10984 11500 11024
rect 11540 10984 28012 11024
rect 28052 10984 28061 11024
rect 29251 10984 29260 11024
rect 29300 10984 35020 11024
rect 35060 10984 38764 11024
rect 38804 10984 38813 11024
rect 12940 10900 18412 10940
rect 18452 10900 18461 10940
rect 32899 10900 32908 10940
rect 32948 10900 40300 10940
rect 40340 10900 40349 10940
rect 0 10856 90 10876
rect 0 10816 1324 10856
rect 1364 10816 1373 10856
rect 3043 10816 3052 10856
rect 3092 10816 9676 10856
rect 9716 10816 9725 10856
rect 0 10796 90 10816
rect 12940 10772 12980 10900
rect 46278 10856 46368 10876
rect 14563 10816 14572 10856
rect 14612 10816 40588 10856
rect 40628 10816 40637 10856
rect 43843 10816 43852 10856
rect 43892 10816 46368 10856
rect 46278 10796 46368 10816
rect 4492 10732 12980 10772
rect 14755 10732 14764 10772
rect 14804 10732 21484 10772
rect 21524 10732 28052 10772
rect 28099 10732 28108 10772
rect 28148 10732 37652 10772
rect 38371 10732 38380 10772
rect 38420 10732 42988 10772
rect 43028 10732 43037 10772
rect 67 10648 76 10688
rect 116 10648 2804 10688
rect 0 10520 90 10540
rect 0 10480 2420 10520
rect 0 10460 90 10480
rect 1459 10396 1468 10436
rect 1508 10396 1996 10436
rect 2036 10396 2045 10436
rect 1036 10228 2036 10268
rect 0 10184 90 10204
rect 1036 10184 1076 10228
rect 1996 10184 2036 10228
rect 2380 10184 2420 10480
rect 2764 10184 2804 10648
rect 4492 10436 4532 10732
rect 28012 10688 28052 10732
rect 37612 10688 37652 10732
rect 5548 10648 8236 10688
rect 8276 10648 8285 10688
rect 12940 10648 19564 10688
rect 19604 10648 19613 10688
rect 19948 10648 27532 10688
rect 27572 10648 27581 10688
rect 28012 10648 29260 10688
rect 29300 10648 29309 10688
rect 29443 10648 29452 10688
rect 29492 10648 37516 10688
rect 37556 10648 37565 10688
rect 37612 10648 44428 10688
rect 44468 10648 44477 10688
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 2921 10396 3004 10436
rect 3044 10396 3052 10436
rect 3092 10396 3101 10436
rect 3859 10396 3868 10436
rect 3908 10396 4532 10436
rect 4675 10396 4684 10436
rect 4724 10396 5308 10436
rect 5348 10396 5357 10436
rect 5548 10184 5588 10648
rect 12940 10604 12980 10648
rect 7852 10564 12980 10604
rect 7852 10436 7892 10564
rect 9667 10480 9676 10520
rect 9716 10480 15284 10520
rect 16387 10480 16396 10520
rect 16436 10480 17684 10520
rect 5827 10396 5836 10436
rect 5876 10396 5884 10436
rect 5924 10396 6007 10436
rect 6883 10396 6892 10436
rect 6932 10396 7412 10436
rect 7795 10396 7804 10436
rect 7844 10396 7892 10436
rect 8009 10396 8092 10436
rect 8132 10396 8140 10436
rect 8180 10396 8189 10436
rect 9139 10396 9148 10436
rect 9188 10396 10444 10436
rect 10484 10396 10493 10436
rect 11347 10396 11356 10436
rect 11396 10396 11596 10436
rect 11636 10396 11645 10436
rect 11731 10396 11740 10436
rect 11780 10396 12748 10436
rect 12788 10396 12797 10436
rect 7372 10352 7412 10396
rect 15244 10352 15284 10480
rect 16195 10396 16204 10436
rect 16244 10396 16732 10436
rect 16772 10396 16781 10436
rect 17347 10396 17356 10436
rect 17396 10396 17404 10436
rect 17444 10396 17527 10436
rect 17644 10352 17684 10480
rect 19948 10436 19988 10648
rect 20039 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20425 10604
rect 23692 10564 25612 10604
rect 25652 10564 25661 10604
rect 28003 10564 28012 10604
rect 28052 10564 34732 10604
rect 34772 10564 34781 10604
rect 35159 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 35545 10604
rect 35596 10564 39052 10604
rect 39092 10564 39101 10604
rect 19699 10396 19708 10436
rect 19748 10396 19988 10436
rect 20131 10396 20140 10436
rect 20180 10396 20716 10436
rect 20756 10396 20765 10436
rect 7180 10312 7276 10352
rect 7316 10312 7325 10352
rect 7372 10312 8564 10352
rect 8755 10312 8764 10352
rect 8804 10312 9292 10352
rect 9332 10312 9341 10352
rect 12940 10312 15188 10352
rect 15244 10312 17588 10352
rect 17644 10312 23060 10352
rect 7180 10268 7220 10312
rect 6665 10228 6796 10268
rect 6836 10228 6845 10268
rect 6924 10228 6940 10268
rect 6980 10228 7084 10268
rect 7124 10228 7133 10268
rect 7180 10228 7206 10268
rect 7246 10228 7255 10268
rect 7324 10228 7333 10268
rect 7373 10228 7660 10268
rect 7700 10228 7709 10268
rect 8524 10184 8564 10312
rect 12940 10268 12980 10312
rect 15148 10268 15188 10312
rect 17548 10268 17588 10312
rect 23020 10268 23060 10312
rect 23692 10268 23732 10564
rect 35596 10520 35636 10564
rect 46278 10520 46368 10540
rect 9283 10228 9292 10268
rect 9332 10228 9341 10268
rect 10540 10259 10924 10268
rect 0 10144 1076 10184
rect 1123 10144 1132 10184
rect 1172 10144 1228 10184
rect 1268 10144 1303 10184
rect 1603 10144 1612 10184
rect 1652 10144 1661 10184
rect 1987 10144 1996 10184
rect 2036 10144 2045 10184
rect 2371 10144 2380 10184
rect 2420 10144 2429 10184
rect 2755 10144 2764 10184
rect 2804 10144 2813 10184
rect 3497 10144 3532 10184
rect 3572 10144 3628 10184
rect 3668 10144 3677 10184
rect 4963 10144 4972 10184
rect 5012 10144 5492 10184
rect 5539 10144 5548 10184
rect 5588 10144 5597 10184
rect 6115 10144 6124 10184
rect 6164 10144 6700 10184
rect 6740 10144 6749 10184
rect 6979 10144 6988 10184
rect 7028 10144 7564 10184
rect 7604 10144 7613 10184
rect 8323 10144 8332 10184
rect 8372 10144 8381 10184
rect 8515 10144 8524 10184
rect 8564 10144 8573 10184
rect 8777 10144 8908 10184
rect 8948 10144 8957 10184
rect 0 10124 90 10144
rect 0 9848 90 9868
rect 1612 9848 1652 10144
rect 5452 10100 5492 10144
rect 8332 10100 8372 10144
rect 9292 10100 9332 10228
rect 10580 10228 10924 10259
rect 10964 10228 10973 10268
rect 11683 10228 11692 10268
rect 11732 10228 11884 10268
rect 11924 10228 11933 10268
rect 11980 10228 12980 10268
rect 13132 10259 13172 10268
rect 10540 10210 10580 10219
rect 10985 10144 11116 10184
rect 11156 10144 11165 10184
rect 11491 10144 11500 10184
rect 11540 10144 11671 10184
rect 11980 10100 12020 10228
rect 13507 10228 13516 10268
rect 13556 10228 14476 10268
rect 14516 10228 14525 10268
rect 14729 10259 14860 10268
rect 14729 10228 14764 10259
rect 13132 10184 13172 10219
rect 14804 10228 14860 10259
rect 14900 10228 14909 10268
rect 15139 10228 15148 10268
rect 15188 10228 15197 10268
rect 16265 10228 16396 10268
rect 16436 10228 16445 10268
rect 16492 10228 17204 10268
rect 17539 10228 17548 10268
rect 17588 10228 17597 10268
rect 18796 10259 20140 10268
rect 14764 10184 14804 10219
rect 16396 10210 16436 10219
rect 12844 10144 14380 10184
rect 14420 10144 14429 10184
rect 14572 10144 14804 10184
rect 12844 10100 12884 10144
rect 2227 10060 2236 10100
rect 2276 10060 2284 10100
rect 2324 10060 2407 10100
rect 5203 10060 5212 10100
rect 5252 10060 5356 10100
rect 5396 10060 5405 10100
rect 5452 10060 5740 10100
rect 5780 10060 5789 10100
rect 6211 10060 6220 10100
rect 6260 10060 6932 10100
rect 7049 10060 7180 10100
rect 7220 10060 7229 10100
rect 7276 10060 8372 10100
rect 8419 10060 8428 10100
rect 8468 10060 12020 10100
rect 12835 10060 12844 10100
rect 12884 10060 12893 10100
rect 6892 10016 6932 10060
rect 7276 10016 7316 10060
rect 14572 10016 14612 10144
rect 16492 10100 16532 10228
rect 17164 10184 17204 10228
rect 18836 10228 20140 10259
rect 20180 10228 20189 10268
rect 20236 10259 21292 10268
rect 18796 10210 18836 10219
rect 20276 10228 21292 10259
rect 21332 10228 21341 10268
rect 21475 10228 21484 10268
rect 21524 10228 21655 10268
rect 21859 10228 21868 10268
rect 21908 10228 22039 10268
rect 23020 10259 23732 10268
rect 23020 10228 23116 10259
rect 20236 10210 20276 10219
rect 23156 10228 23732 10259
rect 23788 10480 34348 10520
rect 34388 10480 34397 10520
rect 34924 10480 35636 10520
rect 35692 10480 43220 10520
rect 43267 10480 43276 10520
rect 43316 10480 44276 10520
rect 23116 10210 23156 10219
rect 23788 10184 23828 10480
rect 24019 10396 24028 10436
rect 24068 10396 24268 10436
rect 24308 10396 24317 10436
rect 26563 10396 26572 10436
rect 26612 10396 27388 10436
rect 27428 10396 27437 10436
rect 27715 10396 27724 10436
rect 27764 10396 27772 10436
rect 27812 10396 27895 10436
rect 28867 10396 28876 10436
rect 28916 10396 29884 10436
rect 29924 10396 29933 10436
rect 30019 10396 30028 10436
rect 30068 10396 32284 10436
rect 32324 10396 32333 10436
rect 34627 10396 34636 10436
rect 34676 10396 34684 10436
rect 34724 10396 34807 10436
rect 26851 10312 26860 10352
rect 26900 10312 28340 10352
rect 31171 10312 31180 10352
rect 31220 10312 32668 10352
rect 32708 10312 32717 10352
rect 32908 10312 33580 10352
rect 33620 10312 34252 10352
rect 34292 10312 34301 10352
rect 28300 10268 28340 10312
rect 32908 10268 32948 10312
rect 24041 10228 24172 10268
rect 24212 10228 24221 10268
rect 25027 10228 25036 10268
rect 25076 10259 25460 10268
rect 25076 10228 25420 10259
rect 25673 10228 25804 10268
rect 25844 10228 25853 10268
rect 27052 10259 27572 10268
rect 25420 10210 25460 10219
rect 27092 10228 27572 10259
rect 27052 10210 27092 10219
rect 16841 10144 16972 10184
rect 17012 10144 17021 10184
rect 17155 10144 17164 10184
rect 17204 10144 17213 10184
rect 19337 10144 19468 10184
rect 19508 10144 19517 10184
rect 23779 10144 23788 10184
rect 23828 10144 23837 10184
rect 27532 10100 27572 10228
rect 27628 10228 28108 10268
rect 28148 10228 28157 10268
rect 28291 10228 28300 10268
rect 28340 10228 28349 10268
rect 29513 10259 29644 10268
rect 29513 10228 29548 10259
rect 27628 10184 27668 10228
rect 29588 10228 29644 10259
rect 29684 10228 30260 10268
rect 30307 10228 30316 10268
rect 30356 10228 30700 10268
rect 30740 10228 30749 10268
rect 31563 10228 31572 10268
rect 31612 10228 32948 10268
rect 33036 10228 33100 10268
rect 33140 10228 33196 10268
rect 33236 10228 33271 10268
rect 34348 10259 34828 10268
rect 29548 10210 29588 10219
rect 30220 10184 30260 10228
rect 32188 10184 32228 10228
rect 34388 10228 34828 10259
rect 34868 10228 34877 10268
rect 34348 10210 34388 10219
rect 34924 10184 34964 10480
rect 35011 10228 35020 10268
rect 35060 10228 35212 10268
rect 35252 10228 35261 10268
rect 27619 10144 27628 10184
rect 27668 10144 27677 10184
rect 28003 10144 28012 10184
rect 28052 10144 29452 10184
rect 29492 10144 29501 10184
rect 30115 10144 30124 10184
rect 30164 10144 30173 10184
rect 30220 10144 31468 10184
rect 31508 10144 31517 10184
rect 31651 10144 31660 10184
rect 31700 10144 31948 10184
rect 31988 10144 31997 10184
rect 32179 10144 32188 10184
rect 32228 10144 32237 10184
rect 32515 10144 32524 10184
rect 32564 10144 32695 10184
rect 32777 10144 32908 10184
rect 32948 10144 32957 10184
rect 34915 10144 34924 10184
rect 34964 10144 34973 10184
rect 30124 10100 30164 10144
rect 35692 10100 35732 10480
rect 43180 10436 43220 10480
rect 44236 10436 44276 10480
rect 45388 10480 46368 10520
rect 35779 10396 35788 10436
rect 35828 10396 36796 10436
rect 36836 10396 36845 10436
rect 36931 10396 36940 10436
rect 36980 10396 37564 10436
rect 37604 10396 37613 10436
rect 38083 10396 38092 10436
rect 38132 10396 38140 10436
rect 38180 10396 38263 10436
rect 38803 10396 38812 10436
rect 38852 10396 39244 10436
rect 39284 10396 39293 10436
rect 40457 10396 40588 10436
rect 40628 10396 40637 10436
rect 41539 10396 41548 10436
rect 41588 10396 42556 10436
rect 42596 10396 42605 10436
rect 42691 10396 42700 10436
rect 42740 10396 42940 10436
rect 42980 10396 42989 10436
rect 43180 10396 44092 10436
rect 44132 10396 44141 10436
rect 44236 10396 44476 10436
rect 44516 10396 44525 10436
rect 38825 10312 38956 10352
rect 38996 10312 39005 10352
rect 40387 10312 40396 10352
rect 40436 10312 42172 10352
rect 42212 10312 42221 10352
rect 42796 10312 43180 10352
rect 43220 10312 43229 10352
rect 43363 10312 43372 10352
rect 43412 10312 44860 10352
rect 44900 10312 44909 10352
rect 35779 10228 35788 10268
rect 35828 10259 36500 10268
rect 35828 10228 36460 10259
rect 36460 10210 36500 10219
rect 37036 10228 39092 10268
rect 37036 10184 37076 10228
rect 37027 10144 37036 10184
rect 37076 10144 37085 10184
rect 37219 10144 37228 10184
rect 37268 10144 37277 10184
rect 37673 10144 37804 10184
rect 37844 10144 37853 10184
rect 38249 10144 38380 10184
rect 38420 10144 38429 10184
rect 38563 10144 38572 10184
rect 38612 10144 38621 10184
rect 37228 10100 37268 10144
rect 38572 10100 38612 10144
rect 39052 10100 39092 10228
rect 39148 10259 39188 10268
rect 39235 10228 39244 10268
rect 39284 10228 40396 10268
rect 40436 10228 40445 10268
rect 40780 10259 40820 10268
rect 39148 10184 39188 10219
rect 41897 10228 42028 10268
rect 42068 10228 42077 10268
rect 40780 10184 40820 10219
rect 42796 10184 42836 10312
rect 42883 10228 42892 10268
rect 42932 10228 43988 10268
rect 43948 10184 43988 10228
rect 39139 10144 39148 10184
rect 39188 10144 40820 10184
rect 42403 10144 42412 10184
rect 42452 10144 42461 10184
rect 42787 10144 42796 10184
rect 42836 10144 42845 10184
rect 43171 10144 43180 10184
rect 43220 10144 43276 10184
rect 43316 10144 43351 10184
rect 43433 10144 43564 10184
rect 43604 10144 43613 10184
rect 43699 10144 43708 10184
rect 43748 10144 43756 10184
rect 43796 10144 43879 10184
rect 43939 10144 43948 10184
rect 43988 10144 43997 10184
rect 44201 10144 44332 10184
rect 44372 10144 44381 10184
rect 44585 10144 44716 10184
rect 44756 10144 44765 10184
rect 44969 10144 45100 10184
rect 45140 10144 45149 10184
rect 42412 10100 42452 10144
rect 45388 10100 45428 10480
rect 46278 10460 46368 10480
rect 46278 10184 46368 10204
rect 45475 10144 45484 10184
rect 45524 10144 46368 10184
rect 46278 10124 46368 10144
rect 14659 10060 14668 10100
rect 14708 10060 15092 10100
rect 15139 10060 15148 10100
rect 15188 10060 16532 10100
rect 16579 10060 16588 10100
rect 16628 10060 17452 10100
rect 17492 10060 17501 10100
rect 17740 10060 19948 10100
rect 19988 10060 25556 10100
rect 25603 10060 25612 10100
rect 25652 10060 25900 10100
rect 25940 10060 25949 10100
rect 27235 10060 27244 10100
rect 27284 10060 27340 10100
rect 27380 10060 27415 10100
rect 27532 10060 27628 10100
rect 27668 10060 27677 10100
rect 30124 10060 35732 10100
rect 36259 10060 36268 10100
rect 36308 10060 37268 10100
rect 37459 10060 37468 10100
rect 37508 10060 38284 10100
rect 38324 10060 38333 10100
rect 38572 10060 38996 10100
rect 39052 10060 41740 10100
rect 41780 10060 41789 10100
rect 42412 10060 43324 10100
rect 43364 10060 43373 10100
rect 44227 10060 44236 10100
rect 44276 10060 45428 10100
rect 15052 10016 15092 10060
rect 1843 9976 1852 10016
rect 1892 9976 1901 10016
rect 2611 9976 2620 10016
rect 2660 9976 2956 10016
rect 2996 9976 3005 10016
rect 6892 9976 7316 10016
rect 10601 9976 10732 10016
rect 10772 9976 10781 10016
rect 13193 9976 13324 10016
rect 13364 9976 13373 10016
rect 13507 9976 13516 10016
rect 13556 9976 14612 10016
rect 14825 9976 14956 10016
rect 14996 9976 15005 10016
rect 15052 9976 17644 10016
rect 17684 9976 17693 10016
rect 0 9808 1652 9848
rect 0 9788 90 9808
rect 1852 9764 1892 9976
rect 17740 9932 17780 10060
rect 25516 10016 25556 10060
rect 38956 10016 38996 10060
rect 17827 9976 17836 10016
rect 17876 9976 18700 10016
rect 18740 9976 18749 10016
rect 18979 9976 18988 10016
rect 19028 9976 19276 10016
rect 19316 9976 19325 10016
rect 19913 9976 20044 10016
rect 20084 9976 20093 10016
rect 23177 9976 23308 10016
rect 23348 9976 23357 10016
rect 25516 9976 27052 10016
rect 27092 9976 29452 10016
rect 29492 9976 29501 10016
rect 29609 9976 29740 10016
rect 29780 9976 29789 10016
rect 31625 9976 31756 10016
rect 31796 9976 31805 10016
rect 34409 9976 34540 10016
rect 34580 9976 34589 10016
rect 36521 9976 36652 10016
rect 36692 9976 36701 10016
rect 38956 9976 41836 10016
rect 41876 9976 41885 10016
rect 2083 9892 2092 9932
rect 2132 9892 7892 9932
rect 8515 9892 8524 9932
rect 8564 9892 17780 9932
rect 17932 9892 25132 9932
rect 25172 9892 25181 9932
rect 26947 9892 26956 9932
rect 26996 9892 33100 9932
rect 33140 9892 33149 9932
rect 34819 9892 34828 9932
rect 34868 9892 40396 9932
rect 40436 9892 42028 9932
rect 42068 9892 42077 9932
rect 42211 9892 42220 9932
rect 42260 9892 43276 9932
rect 43316 9892 43325 9932
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 7852 9764 7892 9892
rect 17932 9848 17972 9892
rect 46278 9848 46368 9868
rect 10531 9808 10540 9848
rect 10580 9808 17972 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 20428 9808 21868 9848
rect 21908 9808 21917 9848
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 34627 9808 34636 9848
rect 34676 9808 41932 9848
rect 41972 9808 41981 9848
rect 44803 9808 44812 9848
rect 44852 9808 46368 9848
rect 1852 9724 2668 9764
rect 2708 9724 2900 9764
rect 5731 9724 5740 9764
rect 5780 9724 7508 9764
rect 7852 9724 20140 9764
rect 20180 9724 20189 9764
rect 2860 9596 2900 9724
rect 7468 9680 7508 9724
rect 20428 9680 20468 9808
rect 46278 9788 46368 9808
rect 5731 9640 5740 9680
rect 5780 9640 6316 9680
rect 6356 9640 6365 9680
rect 7241 9640 7276 9680
rect 7316 9640 7372 9680
rect 7412 9640 7421 9680
rect 7468 9640 8428 9680
rect 8468 9640 8477 9680
rect 9004 9640 12460 9680
rect 12500 9640 12509 9680
rect 13891 9640 13900 9680
rect 13940 9640 13948 9680
rect 13988 9640 14071 9680
rect 14803 9640 14812 9680
rect 14852 9640 15052 9680
rect 15092 9640 15101 9680
rect 18163 9640 18172 9680
rect 18212 9640 18508 9680
rect 18548 9640 18557 9680
rect 18691 9640 18700 9680
rect 18740 9640 20468 9680
rect 20524 9724 25076 9764
rect 652 9556 1132 9596
rect 1172 9556 1181 9596
rect 1315 9556 1324 9596
rect 1364 9556 2036 9596
rect 2860 9556 8660 9596
rect 0 9512 90 9532
rect 652 9512 692 9556
rect 1996 9512 2036 9556
rect 8140 9512 8180 9556
rect 0 9472 692 9512
rect 1097 9472 1228 9512
rect 1268 9472 1277 9512
rect 1603 9472 1612 9512
rect 1652 9472 1661 9512
rect 1987 9472 1996 9512
rect 2036 9472 2045 9512
rect 2227 9472 2236 9512
rect 2276 9472 2900 9512
rect 0 9452 90 9472
rect 1612 9344 1652 9472
rect 2860 9428 2900 9472
rect 5548 9472 7220 9512
rect 5548 9428 5588 9472
rect 7180 9428 7220 9472
rect 7660 9472 7948 9512
rect 7988 9472 7997 9512
rect 8131 9472 8140 9512
rect 8180 9472 8189 9512
rect 8393 9472 8524 9512
rect 8564 9472 8573 9512
rect 7660 9428 7700 9472
rect 2860 9388 4300 9428
rect 4340 9388 5492 9428
rect 5539 9388 5548 9428
rect 5588 9388 5719 9428
rect 5923 9388 5932 9428
rect 5972 9388 6356 9428
rect 7020 9388 7084 9428
rect 7124 9388 7180 9428
rect 7651 9388 7660 9428
rect 7700 9388 7709 9428
rect 7756 9388 7779 9428
rect 7819 9388 7828 9428
rect 7882 9388 7891 9428
rect 7931 9388 7940 9428
rect 172 9304 1652 9344
rect 0 9176 90 9196
rect 172 9176 212 9304
rect 5452 9260 5492 9388
rect 5548 9379 5588 9388
rect 1459 9220 1468 9260
rect 1508 9220 1517 9260
rect 1843 9220 1852 9260
rect 1892 9220 2188 9260
rect 2228 9220 2237 9260
rect 5452 9220 5740 9260
rect 5780 9220 5789 9260
rect 0 9136 212 9176
rect 0 9116 90 9136
rect 0 8840 90 8860
rect 1468 8840 1508 9220
rect 6316 9092 6356 9388
rect 7180 9379 7220 9388
rect 7267 9304 7276 9344
rect 7316 9304 7564 9344
rect 7604 9304 7613 9344
rect 7660 9260 7700 9388
rect 7363 9220 7372 9260
rect 7412 9220 7700 9260
rect 7756 9176 7796 9388
rect 7891 9344 7931 9388
rect 8524 9344 8564 9472
rect 8620 9428 8660 9556
rect 9004 9512 9044 9640
rect 20524 9596 20564 9724
rect 20681 9640 20764 9680
rect 20804 9640 20812 9680
rect 20852 9640 20861 9680
rect 25036 9596 25076 9724
rect 27436 9724 34444 9764
rect 34484 9724 34493 9764
rect 39043 9724 39052 9764
rect 39092 9724 42796 9764
rect 42836 9724 42845 9764
rect 27436 9680 27476 9724
rect 25411 9640 25420 9680
rect 25460 9640 26236 9680
rect 26276 9640 26285 9680
rect 26380 9640 27476 9680
rect 26380 9596 26420 9640
rect 9388 9556 11788 9596
rect 11828 9556 11837 9596
rect 11980 9556 20564 9596
rect 20620 9556 21380 9596
rect 21427 9556 21436 9596
rect 21476 9556 21964 9596
rect 22004 9556 22013 9596
rect 22147 9556 22156 9596
rect 22196 9556 24940 9596
rect 24980 9556 24989 9596
rect 25036 9556 26420 9596
rect 8873 9472 9004 9512
rect 9044 9472 9053 9512
rect 9388 9428 9428 9556
rect 11980 9512 12020 9556
rect 11299 9472 11308 9512
rect 11348 9472 11980 9512
rect 12020 9472 12029 9512
rect 13258 9472 13267 9512
rect 13307 9472 13420 9512
rect 13460 9472 13469 9512
rect 14057 9472 14092 9512
rect 14132 9472 14188 9512
rect 14228 9472 14237 9512
rect 14441 9472 14572 9512
rect 14612 9472 14621 9512
rect 15401 9472 15532 9512
rect 15572 9472 15581 9512
rect 16963 9472 16972 9512
rect 17012 9472 17143 9512
rect 17801 9472 17836 9512
rect 17876 9472 17932 9512
rect 17972 9472 17981 9512
rect 18028 9472 18892 9512
rect 18932 9472 18941 9512
rect 20170 9472 20179 9512
rect 20219 9472 20332 9512
rect 20372 9472 20381 9512
rect 10924 9428 10964 9437
rect 12556 9428 12596 9437
rect 16108 9428 16148 9437
rect 18028 9428 18068 9472
rect 19468 9428 19508 9437
rect 20620 9428 20660 9556
rect 21340 9512 21380 9556
rect 20995 9472 21004 9512
rect 21044 9472 21175 9512
rect 21226 9472 21235 9512
rect 21275 9472 21284 9512
rect 21340 9472 22004 9512
rect 22147 9472 22156 9512
rect 22196 9472 22252 9512
rect 22292 9472 22327 9512
rect 23434 9472 23443 9512
rect 23483 9472 23596 9512
rect 23636 9472 23645 9512
rect 23692 9472 24844 9512
rect 24884 9472 24893 9512
rect 21244 9428 21284 9472
rect 21964 9428 22004 9472
rect 22732 9428 22772 9437
rect 8620 9388 9428 9428
rect 9545 9388 9676 9428
rect 9716 9388 9725 9428
rect 10793 9388 10924 9428
rect 10964 9388 10973 9428
rect 11452 9388 11470 9428
rect 11510 9388 11519 9428
rect 10924 9379 10964 9388
rect 7843 9304 7852 9344
rect 7892 9304 7931 9344
rect 8140 9304 8564 9344
rect 6787 9136 6796 9176
rect 6836 9136 7756 9176
rect 7796 9136 7805 9176
rect 8140 9092 8180 9304
rect 8371 9220 8380 9260
rect 8420 9220 8620 9260
rect 8660 9220 8669 9260
rect 8755 9220 8764 9260
rect 8804 9220 9100 9260
rect 9140 9220 9149 9260
rect 9235 9220 9244 9260
rect 9284 9220 10060 9260
rect 10100 9220 10109 9260
rect 11107 9220 11116 9260
rect 11156 9220 11212 9260
rect 11252 9220 11287 9260
rect 11452 9092 11492 9388
rect 11578 9360 11587 9400
rect 11636 9360 11767 9400
rect 11945 9388 12076 9428
rect 12116 9388 12125 9428
rect 12596 9388 12748 9428
rect 12788 9388 12797 9428
rect 13066 9388 13075 9428
rect 13115 9388 13324 9428
rect 13364 9388 13373 9428
rect 14891 9388 14956 9428
rect 14996 9388 15022 9428
rect 15062 9388 15071 9428
rect 15139 9388 15148 9428
rect 15188 9388 15197 9428
rect 15427 9388 15436 9428
rect 15476 9388 15628 9428
rect 15668 9388 15677 9428
rect 15811 9388 15820 9428
rect 15860 9388 16108 9428
rect 16579 9388 16588 9428
rect 16636 9388 16759 9428
rect 17731 9388 17740 9428
rect 17780 9388 18068 9428
rect 18115 9388 18124 9428
rect 18164 9388 18403 9428
rect 18443 9388 18452 9428
rect 18499 9388 18508 9428
rect 18548 9388 18679 9428
rect 18857 9388 18988 9428
rect 19028 9388 19037 9428
rect 19913 9388 19987 9428
rect 20027 9388 20044 9428
rect 20084 9388 20093 9428
rect 20140 9388 20660 9428
rect 20899 9388 20908 9428
rect 20948 9388 21284 9428
rect 21475 9388 21484 9428
rect 21524 9388 21667 9428
rect 21707 9388 21716 9428
rect 21763 9388 21772 9428
rect 21812 9388 21859 9428
rect 21964 9388 22252 9428
rect 22292 9388 22301 9428
rect 23177 9388 23251 9428
rect 23291 9388 23308 9428
rect 23348 9388 23357 9428
rect 12556 9344 12596 9388
rect 15148 9344 15188 9388
rect 11875 9304 11884 9344
rect 11924 9304 12596 9344
rect 12643 9304 12652 9344
rect 12692 9304 14668 9344
rect 14708 9304 14717 9344
rect 15043 9304 15052 9344
rect 15092 9304 15188 9344
rect 16108 9344 16148 9388
rect 19468 9344 19508 9388
rect 20140 9344 20180 9388
rect 21772 9344 21812 9388
rect 22732 9344 22772 9388
rect 16108 9304 20180 9344
rect 20563 9304 20572 9344
rect 20612 9304 21580 9344
rect 21620 9304 21629 9344
rect 21763 9304 21772 9344
rect 21812 9304 21821 9344
rect 22051 9304 22060 9344
rect 22100 9304 22732 9344
rect 22772 9304 22781 9344
rect 23692 9260 23732 9472
rect 24317 9388 24355 9428
rect 24395 9388 24404 9428
rect 24451 9388 24460 9428
rect 24500 9388 24509 9428
rect 24643 9388 24652 9428
rect 24692 9388 24940 9428
rect 24980 9388 24989 9428
rect 24364 9344 24404 9388
rect 24460 9344 24500 9388
rect 25036 9344 25076 9556
rect 26467 9472 26476 9512
rect 26516 9472 26647 9512
rect 26698 9472 26707 9512
rect 26747 9472 26756 9512
rect 26825 9472 26908 9512
rect 26948 9472 26956 9512
rect 26996 9472 27005 9512
rect 27293 9472 27340 9512
rect 27380 9472 27389 9512
rect 25420 9428 25460 9437
rect 25289 9388 25420 9428
rect 25460 9388 25469 9428
rect 25891 9388 25900 9428
rect 25948 9388 26071 9428
rect 25420 9379 25460 9388
rect 26716 9344 26756 9472
rect 27340 9428 27380 9472
rect 27436 9428 27476 9640
rect 28492 9640 32276 9680
rect 32323 9640 32332 9680
rect 32372 9640 33148 9680
rect 33188 9640 33197 9680
rect 33475 9640 33484 9680
rect 33524 9640 33916 9680
rect 33956 9640 33965 9680
rect 40291 9640 40300 9680
rect 40340 9640 44188 9680
rect 44228 9640 44237 9680
rect 44419 9640 44428 9680
rect 44468 9640 44572 9680
rect 44612 9640 44621 9680
rect 27689 9472 27820 9512
rect 27860 9472 27869 9512
rect 28396 9428 28436 9437
rect 28492 9428 28532 9640
rect 32236 9596 32276 9640
rect 32236 9556 32372 9596
rect 29242 9472 29251 9512
rect 29291 9472 29300 9512
rect 29539 9472 29548 9512
rect 29588 9472 30740 9512
rect 31625 9472 31660 9512
rect 31700 9472 31756 9512
rect 31796 9472 31805 9512
rect 29260 9428 29300 9472
rect 27322 9388 27331 9428
rect 27371 9388 27380 9428
rect 27427 9388 27436 9428
rect 27476 9388 27485 9428
rect 27907 9388 27916 9428
rect 27956 9388 27965 9428
rect 28387 9388 28396 9428
rect 28436 9388 28567 9428
rect 28906 9388 28915 9428
rect 28955 9388 29300 9428
rect 29452 9428 29492 9437
rect 30700 9428 30740 9472
rect 32332 9428 32372 9556
rect 33388 9556 38956 9596
rect 38996 9556 39005 9596
rect 39235 9556 39244 9596
rect 39284 9556 41548 9596
rect 41588 9556 41597 9596
rect 41731 9556 41740 9596
rect 41780 9556 43036 9596
rect 43076 9556 43085 9596
rect 43180 9556 44468 9596
rect 33388 9512 33428 9556
rect 43180 9512 43220 9556
rect 44428 9512 44468 9556
rect 46278 9512 46368 9532
rect 33379 9472 33388 9512
rect 33428 9472 33437 9512
rect 33763 9472 33772 9512
rect 33812 9472 33821 9512
rect 34025 9472 34156 9512
rect 34196 9472 34205 9512
rect 34531 9472 34540 9512
rect 34580 9472 34589 9512
rect 34819 9472 34828 9512
rect 34868 9472 35020 9512
rect 35060 9472 35069 9512
rect 36547 9472 36556 9512
rect 36596 9472 36748 9512
rect 36788 9472 36797 9512
rect 37132 9472 39148 9512
rect 39188 9472 39197 9512
rect 39331 9472 39340 9512
rect 39380 9472 41684 9512
rect 41897 9472 42028 9512
rect 42068 9472 42077 9512
rect 42499 9472 42508 9512
rect 42548 9472 42652 9512
rect 42692 9472 42701 9512
rect 42761 9472 42892 9512
rect 42932 9472 42941 9512
rect 43075 9472 43084 9512
rect 43124 9472 43220 9512
rect 43267 9472 43276 9512
rect 43316 9472 43447 9512
rect 43529 9472 43660 9512
rect 43700 9472 43709 9512
rect 43913 9472 44044 9512
rect 44084 9472 44093 9512
rect 44419 9472 44428 9512
rect 44468 9472 44477 9512
rect 44803 9472 44812 9512
rect 44852 9472 44861 9512
rect 44908 9472 46368 9512
rect 30691 9388 30700 9428
rect 30740 9388 30749 9428
rect 31258 9388 31267 9428
rect 31307 9388 31316 9428
rect 31363 9388 31372 9428
rect 31412 9388 31468 9428
rect 31508 9388 31543 9428
rect 31843 9388 31852 9428
rect 31892 9388 31901 9428
rect 32201 9388 32332 9428
rect 32372 9388 32381 9428
rect 32811 9388 32820 9428
rect 32860 9388 32869 9428
rect 27916 9344 27956 9388
rect 28396 9387 28532 9388
rect 28396 9379 28436 9387
rect 29452 9344 29492 9388
rect 31276 9344 31316 9388
rect 24355 9304 24364 9344
rect 24404 9304 24413 9344
rect 24460 9304 25076 9344
rect 26092 9304 26756 9344
rect 27427 9304 27436 9344
rect 27476 9304 27916 9344
rect 27956 9304 27965 9344
rect 28492 9304 29204 9344
rect 29452 9304 29548 9344
rect 29588 9304 29597 9344
rect 31276 9304 31756 9344
rect 31796 9304 31805 9344
rect 26092 9260 26132 9304
rect 11779 9220 11788 9260
rect 11828 9220 12980 9260
rect 13651 9220 13660 9260
rect 13700 9220 14380 9260
rect 14420 9220 14429 9260
rect 16771 9220 16780 9260
rect 16820 9220 16972 9260
rect 17012 9220 17021 9260
rect 17203 9220 17212 9260
rect 17252 9220 18508 9260
rect 18548 9220 18557 9260
rect 19363 9220 19372 9260
rect 19412 9220 23732 9260
rect 23827 9220 23836 9260
rect 23876 9220 25900 9260
rect 25940 9220 25949 9260
rect 26083 9220 26092 9260
rect 26132 9220 26141 9260
rect 12940 9176 12980 9220
rect 28492 9176 28532 9304
rect 29164 9260 29204 9304
rect 31852 9260 31892 9388
rect 32332 9379 32372 9388
rect 28937 9220 29068 9260
rect 29108 9220 29117 9260
rect 29164 9220 31892 9260
rect 12940 9136 14284 9176
rect 14324 9136 14333 9176
rect 18691 9136 18700 9176
rect 18740 9136 21100 9176
rect 21140 9136 21149 9176
rect 21196 9136 28532 9176
rect 21196 9092 21236 9136
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 6316 9052 8180 9092
rect 8323 9052 8332 9092
rect 8372 9052 11308 9092
rect 11348 9052 11357 9092
rect 11452 9052 12692 9092
rect 15907 9052 15916 9092
rect 15956 9052 18644 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 20611 9052 20620 9092
rect 20660 9052 20908 9092
rect 20948 9052 21236 9092
rect 21763 9052 21772 9092
rect 21812 9052 24748 9092
rect 24788 9052 24797 9092
rect 25123 9052 25132 9092
rect 25172 9052 32716 9092
rect 32756 9052 32765 9092
rect 6316 9008 6356 9052
rect 2860 8968 6356 9008
rect 9955 8968 9964 9008
rect 10004 8968 12364 9008
rect 12404 8968 12413 9008
rect 2860 8924 2900 8968
rect 12652 8924 12692 9052
rect 18604 9008 18644 9052
rect 32812 9008 32852 9388
rect 33772 9344 33812 9472
rect 34540 9428 34580 9472
rect 35596 9428 35636 9437
rect 37132 9428 37172 9472
rect 40012 9428 40052 9472
rect 41644 9428 41684 9472
rect 44812 9428 44852 9472
rect 34493 9388 34527 9428
rect 34567 9388 34580 9428
rect 34627 9388 34636 9428
rect 34676 9388 34724 9428
rect 34915 9388 34924 9428
rect 34964 9388 35116 9428
rect 35156 9388 35165 9428
rect 35636 9388 35884 9428
rect 35924 9388 35933 9428
rect 36106 9388 36115 9428
rect 36155 9388 36652 9428
rect 36692 9388 36701 9428
rect 37123 9388 37132 9428
rect 37172 9388 37303 9428
rect 38249 9388 38380 9428
rect 38420 9388 38429 9428
rect 38633 9388 38764 9428
rect 38804 9388 38813 9428
rect 40052 9388 40128 9428
rect 40270 9388 40396 9428
rect 40441 9388 40450 9428
rect 41731 9388 41740 9428
rect 41780 9388 44852 9428
rect 34684 9344 34724 9388
rect 35596 9379 35636 9388
rect 37132 9379 37172 9388
rect 40012 9379 40052 9388
rect 41644 9379 41684 9388
rect 44908 9344 44948 9472
rect 46278 9452 46368 9472
rect 33100 9304 33812 9344
rect 34435 9304 34444 9344
rect 34484 9304 34724 9344
rect 36809 9304 36940 9344
rect 36980 9304 36989 9344
rect 40195 9304 40204 9344
rect 40244 9304 41356 9344
rect 41396 9304 41405 9344
rect 43276 9304 43804 9344
rect 43844 9304 43853 9344
rect 43939 9304 43948 9344
rect 43988 9304 44948 9344
rect 33100 9260 33140 9304
rect 43276 9260 43316 9304
rect 32995 9220 33004 9260
rect 33044 9220 33140 9260
rect 33379 9220 33388 9260
rect 33428 9220 33532 9260
rect 33572 9220 33581 9260
rect 36137 9220 36268 9260
rect 36308 9220 36317 9260
rect 36787 9220 36796 9260
rect 36836 9220 36844 9260
rect 36884 9220 36967 9260
rect 40195 9220 40204 9260
rect 40244 9220 40396 9260
rect 40436 9220 40445 9260
rect 41827 9220 41836 9260
rect 41876 9220 42028 9260
rect 42068 9220 42077 9260
rect 42259 9220 42268 9260
rect 42308 9220 42548 9260
rect 42787 9220 42796 9260
rect 42836 9220 43316 9260
rect 43363 9220 43372 9260
rect 43412 9220 43420 9260
rect 43460 9220 43543 9260
rect 42508 9176 42548 9220
rect 46278 9176 46368 9196
rect 37411 9136 37420 9176
rect 37460 9136 41452 9176
rect 41492 9136 41501 9176
rect 42508 9136 43276 9176
rect 43316 9136 43325 9176
rect 44611 9136 44620 9176
rect 44660 9136 46368 9176
rect 46278 9116 46368 9136
rect 33283 9052 33292 9092
rect 33332 9052 34964 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 37315 9052 37324 9092
rect 37364 9052 43084 9092
rect 43124 9052 43133 9092
rect 34924 9008 34964 9052
rect 15724 8968 16588 9008
rect 16628 8968 16637 9008
rect 18604 8968 21196 9008
rect 21236 8968 21245 9008
rect 21475 8968 21484 9008
rect 21524 8968 21716 9008
rect 15724 8924 15764 8968
rect 21676 8924 21716 8968
rect 21772 8968 27860 9008
rect 27907 8968 27916 9008
rect 27956 8968 32524 9008
rect 32564 8968 32573 9008
rect 32812 8968 33140 9008
rect 33187 8968 33196 9008
rect 33236 8968 34828 9008
rect 34868 8968 34877 9008
rect 34924 8968 41740 9008
rect 41780 8968 41789 9008
rect 41923 8968 41932 9008
rect 41972 8968 43372 9008
rect 43412 8968 43421 9008
rect 1843 8884 1852 8924
rect 1892 8884 2900 8924
rect 5452 8884 11020 8924
rect 11060 8884 11069 8924
rect 12329 8884 12460 8924
rect 12500 8884 12509 8924
rect 12643 8884 12652 8924
rect 12692 8884 12701 8924
rect 15715 8884 15724 8924
rect 15764 8884 15773 8924
rect 17347 8884 17356 8924
rect 17396 8884 18124 8924
rect 18164 8884 18173 8924
rect 19363 8884 19372 8924
rect 19412 8884 19468 8924
rect 19508 8884 19543 8924
rect 19651 8884 19660 8924
rect 19700 8884 19708 8924
rect 19748 8884 19831 8924
rect 21667 8884 21676 8924
rect 21716 8884 21725 8924
rect 0 8800 1228 8840
rect 1268 8800 1277 8840
rect 1468 8800 3956 8840
rect 0 8780 90 8800
rect 3916 8756 3956 8800
rect 5452 8756 5492 8884
rect 21772 8840 21812 8968
rect 27820 8924 27860 8968
rect 33100 8924 33140 8968
rect 21948 8884 21964 8924
rect 22004 8884 22108 8924
rect 22148 8884 23980 8924
rect 24020 8884 24029 8924
rect 24233 8884 24268 8924
rect 24308 8884 24364 8924
rect 24404 8884 24413 8924
rect 24931 8884 24940 8924
rect 24980 8884 27764 8924
rect 27811 8884 27820 8924
rect 27860 8884 29780 8924
rect 31747 8884 31756 8924
rect 31796 8884 32812 8924
rect 32852 8884 32861 8924
rect 33100 8884 33388 8924
rect 33428 8884 33437 8924
rect 34915 8884 34924 8924
rect 34964 8884 38476 8924
rect 38516 8884 38525 8924
rect 39715 8884 39724 8924
rect 39764 8884 40340 8924
rect 42019 8884 42028 8924
rect 42068 8884 44044 8924
rect 44084 8884 44093 8924
rect 44393 8884 44476 8924
rect 44516 8884 44524 8924
rect 44564 8884 44573 8924
rect 27724 8840 27764 8884
rect 29740 8840 29780 8884
rect 40300 8840 40340 8884
rect 46278 8840 46368 8860
rect 6979 8800 6988 8840
rect 7028 8800 7765 8840
rect 9091 8800 9100 8840
rect 9140 8800 9676 8840
rect 9716 8800 9725 8840
rect 10409 8800 10492 8840
rect 10532 8800 10540 8840
rect 10580 8800 10589 8840
rect 10685 8800 10732 8840
rect 10772 8800 10781 8840
rect 11203 8800 11212 8840
rect 11252 8800 12308 8840
rect 7725 8756 7765 8800
rect 10732 8756 10772 8800
rect 3916 8716 4300 8756
rect 4340 8716 5492 8756
rect 5539 8716 5548 8756
rect 5588 8716 5719 8756
rect 5801 8716 5932 8756
rect 5972 8716 5981 8756
rect 7075 8716 7084 8756
rect 7124 8747 7255 8756
rect 7124 8716 7180 8747
rect 3916 8672 3956 8716
rect 5548 8698 5588 8707
rect 5932 8672 5972 8716
rect 7220 8716 7255 8747
rect 7710 8716 7719 8756
rect 7759 8716 7768 8756
rect 7180 8698 7220 8707
rect 7825 8696 7837 8736
rect 7877 8696 7886 8736
rect 7930 8716 7939 8756
rect 7988 8716 8119 8756
rect 8227 8716 8236 8756
rect 8276 8716 8428 8756
rect 8468 8716 8477 8756
rect 8803 8716 8812 8756
rect 8852 8747 10060 8756
rect 8852 8716 9484 8747
rect 9524 8716 10060 8747
rect 10100 8716 10109 8756
rect 10714 8716 10723 8756
rect 10763 8716 10772 8756
rect 10819 8716 10828 8756
rect 10868 8716 10999 8756
rect 11177 8716 11212 8756
rect 11252 8716 11308 8756
rect 11348 8716 11357 8756
rect 11753 8747 11884 8756
rect 11753 8716 11788 8747
rect 9484 8698 9524 8707
rect 11828 8716 11884 8747
rect 11924 8716 11933 8756
rect 12268 8747 12308 8800
rect 17740 8800 21812 8840
rect 21859 8800 21868 8840
rect 21908 8800 25804 8840
rect 25844 8800 25853 8840
rect 25987 8800 25996 8840
rect 26036 8800 27668 8840
rect 27724 8800 29012 8840
rect 29395 8800 29404 8840
rect 29444 8800 29644 8840
rect 29684 8800 29693 8840
rect 29740 8800 33196 8840
rect 33236 8800 33245 8840
rect 34156 8800 35444 8840
rect 35971 8800 35980 8840
rect 36020 8800 36220 8840
rect 36260 8800 36269 8840
rect 40300 8800 42172 8840
rect 42212 8800 42221 8840
rect 43027 8800 43036 8840
rect 43076 8800 46368 8840
rect 17740 8756 17780 8800
rect 25228 8756 25268 8800
rect 27628 8756 27668 8800
rect 28972 8756 29012 8800
rect 11788 8698 11828 8707
rect 12714 8716 12836 8756
rect 12884 8716 12894 8756
rect 14083 8716 14092 8756
rect 14132 8716 14228 8756
rect 14275 8716 14284 8756
rect 14324 8716 14455 8756
rect 14851 8716 14860 8756
rect 14900 8747 15572 8756
rect 14900 8716 15532 8747
rect 12268 8698 12308 8707
rect 7825 8672 7865 8696
rect 14188 8672 14228 8716
rect 15785 8716 15916 8756
rect 15956 8716 15965 8756
rect 17164 8747 17204 8756
rect 15532 8698 15572 8707
rect 17443 8716 17452 8756
rect 17492 8716 17635 8756
rect 17675 8716 17684 8756
rect 17731 8716 17740 8756
rect 17780 8716 17911 8756
rect 18115 8716 18124 8756
rect 18164 8716 18295 8756
rect 18499 8716 18508 8756
rect 18548 8747 18740 8756
rect 18548 8716 18700 8747
rect 17164 8672 17204 8707
rect 19145 8747 19276 8756
rect 19145 8716 19180 8747
rect 18700 8698 18740 8707
rect 19220 8716 19276 8747
rect 19316 8716 19325 8756
rect 19939 8716 19948 8756
rect 19988 8716 20236 8756
rect 20276 8716 20285 8756
rect 20803 8716 20812 8756
rect 20852 8747 21524 8756
rect 20852 8716 21484 8747
rect 19180 8698 19220 8707
rect 21667 8716 21676 8756
rect 21716 8716 22828 8756
rect 22868 8716 22877 8756
rect 23945 8716 24076 8756
rect 24116 8716 24125 8756
rect 24643 8716 24652 8756
rect 24692 8716 24940 8756
rect 24980 8716 24989 8756
rect 25219 8716 25228 8756
rect 25268 8716 25277 8756
rect 25699 8716 25708 8756
rect 25748 8747 26516 8756
rect 25748 8716 26476 8747
rect 21484 8698 21524 8707
rect 24076 8698 24116 8707
rect 26921 8716 27052 8756
rect 27092 8716 27101 8756
rect 27628 8716 28012 8756
rect 28052 8716 28061 8756
rect 28169 8716 28300 8756
rect 28340 8716 28349 8756
rect 28972 8716 29684 8756
rect 29731 8716 29740 8756
rect 29780 8716 30019 8756
rect 30059 8716 30068 8756
rect 30115 8716 30124 8756
rect 30164 8716 30220 8756
rect 30260 8716 30295 8756
rect 30377 8716 30508 8756
rect 30548 8716 30557 8756
rect 30953 8716 31084 8756
rect 31124 8716 31133 8756
rect 31433 8716 31564 8756
rect 31604 8716 31613 8756
rect 31817 8716 31852 8756
rect 31892 8716 31948 8756
rect 31988 8716 31997 8756
rect 32044 8716 33140 8756
rect 26476 8698 26516 8707
rect 28300 8698 28340 8707
rect 29644 8672 29684 8716
rect 31084 8698 31124 8707
rect 31564 8698 31604 8707
rect 32044 8672 32084 8716
rect 1097 8632 1228 8672
rect 1268 8632 1277 8672
rect 1603 8632 1612 8672
rect 1652 8632 1661 8672
rect 1987 8632 1996 8672
rect 2036 8632 2572 8672
rect 2612 8632 2621 8672
rect 2681 8632 2764 8672
rect 2804 8632 2812 8672
rect 2852 8632 2861 8672
rect 3907 8632 3916 8672
rect 3956 8632 3965 8672
rect 4147 8632 4156 8672
rect 4196 8632 4300 8672
rect 4340 8632 4349 8672
rect 5644 8632 5972 8672
rect 7276 8632 7865 8672
rect 10243 8632 10252 8672
rect 10292 8632 10636 8672
rect 10676 8632 10685 8672
rect 11273 8632 11308 8672
rect 11348 8632 11404 8672
rect 11444 8632 11453 8672
rect 13027 8632 13036 8672
rect 13076 8632 13996 8672
rect 14036 8632 14045 8672
rect 14179 8632 14188 8672
rect 14228 8632 14237 8672
rect 17164 8632 17548 8672
rect 17588 8632 17597 8672
rect 18211 8632 18220 8672
rect 18260 8632 18604 8672
rect 18644 8632 18653 8672
rect 19939 8632 19948 8672
rect 19988 8632 21388 8672
rect 21428 8632 21437 8672
rect 21859 8632 21868 8672
rect 21908 8632 22060 8672
rect 22100 8632 22109 8672
rect 29059 8632 29068 8672
rect 29108 8632 29116 8672
rect 29156 8632 29239 8672
rect 29539 8632 29548 8672
rect 29588 8632 29597 8672
rect 29644 8632 30604 8672
rect 30644 8632 30892 8672
rect 30932 8632 30941 8672
rect 31660 8632 32084 8672
rect 32131 8632 32140 8672
rect 32180 8632 33004 8672
rect 33044 8632 33053 8672
rect 1612 8588 1652 8632
rect 844 8548 1652 8588
rect 0 8504 90 8524
rect 844 8504 884 8548
rect 5644 8504 5684 8632
rect 7276 8588 7316 8632
rect 6595 8548 6604 8588
rect 6644 8548 7316 8588
rect 7363 8548 7372 8588
rect 7412 8548 7543 8588
rect 8092 8548 11884 8588
rect 11924 8548 11933 8588
rect 15811 8548 15820 8588
rect 15860 8548 29452 8588
rect 29492 8548 29501 8588
rect 0 8464 884 8504
rect 1459 8464 1468 8504
rect 1508 8464 5684 8504
rect 5731 8464 5740 8504
rect 5780 8464 6796 8504
rect 6836 8464 6845 8504
rect 7433 8464 7468 8504
rect 7508 8464 7564 8504
rect 7604 8464 7613 8504
rect 0 8444 90 8464
rect 8092 8420 8132 8548
rect 29548 8504 29588 8632
rect 31660 8588 31700 8632
rect 30403 8548 30412 8588
rect 30452 8548 31700 8588
rect 33100 8588 33140 8716
rect 33196 8747 33283 8756
rect 33236 8716 33283 8747
rect 33196 8672 33236 8707
rect 34156 8672 34196 8800
rect 34330 8716 34339 8756
rect 34379 8716 34388 8756
rect 34435 8716 34444 8756
rect 34484 8716 34540 8756
rect 34580 8716 34615 8756
rect 34697 8716 34828 8756
rect 34868 8716 34877 8756
rect 35404 8747 35444 8800
rect 46278 8780 46368 8800
rect 33187 8632 33196 8672
rect 33236 8632 33245 8672
rect 33292 8632 34196 8672
rect 34348 8672 34388 8716
rect 35404 8698 35444 8707
rect 35884 8747 36268 8756
rect 35924 8716 36268 8747
rect 36308 8716 36317 8756
rect 36617 8716 36748 8756
rect 36788 8716 36797 8756
rect 37027 8716 37036 8756
rect 37076 8747 38036 8756
rect 37076 8716 37996 8747
rect 35884 8698 35924 8707
rect 38249 8716 38380 8756
rect 38420 8716 38429 8756
rect 38476 8747 39668 8756
rect 38476 8716 39628 8747
rect 37996 8672 38036 8707
rect 38476 8672 38516 8716
rect 40282 8716 40291 8756
rect 40331 8716 40340 8756
rect 40384 8716 40393 8756
rect 40433 8716 40492 8756
rect 40532 8716 40573 8756
rect 40649 8716 40780 8756
rect 40820 8716 40829 8756
rect 41225 8716 41356 8756
rect 41396 8716 41405 8756
rect 41635 8716 41644 8756
rect 41684 8747 41876 8756
rect 41684 8716 41836 8747
rect 39628 8698 39668 8707
rect 40300 8672 40340 8716
rect 41356 8698 41396 8707
rect 41836 8698 41876 8707
rect 41932 8716 44372 8756
rect 34348 8632 34444 8672
rect 34484 8632 34493 8672
rect 34793 8632 34924 8672
rect 34964 8632 34973 8672
rect 36106 8632 36115 8672
rect 36155 8632 36460 8672
rect 36500 8632 36509 8672
rect 37996 8632 38516 8672
rect 38563 8632 38572 8672
rect 38612 8632 39572 8672
rect 40300 8632 40396 8672
rect 40436 8632 40445 8672
rect 40588 8632 40876 8672
rect 40916 8632 40925 8672
rect 33292 8588 33332 8632
rect 39532 8588 39572 8632
rect 40588 8588 40628 8632
rect 41932 8588 41972 8716
rect 44332 8672 44372 8716
rect 42058 8632 42067 8672
rect 42107 8632 42412 8672
rect 42452 8632 42461 8672
rect 42665 8632 42796 8672
rect 42836 8632 42845 8672
rect 42979 8632 42988 8672
rect 43028 8632 43316 8672
rect 43363 8632 43372 8672
rect 43412 8632 43543 8672
rect 43625 8632 43756 8672
rect 43796 8632 43805 8672
rect 43852 8632 44092 8672
rect 44132 8632 44141 8672
rect 44323 8632 44332 8672
rect 44372 8632 44381 8672
rect 44585 8632 44716 8672
rect 44756 8632 44765 8672
rect 44899 8632 44908 8672
rect 44948 8632 45079 8672
rect 45139 8632 45148 8672
rect 45188 8632 46252 8672
rect 46292 8632 46301 8672
rect 33100 8548 33332 8588
rect 34531 8548 34540 8588
rect 34580 8548 38324 8588
rect 39532 8548 40628 8588
rect 41443 8548 41452 8588
rect 41492 8548 41972 8588
rect 43276 8588 43316 8632
rect 43852 8588 43892 8632
rect 43276 8548 43892 8588
rect 43987 8548 43996 8588
rect 44036 8548 45332 8588
rect 9283 8464 9292 8504
rect 9332 8464 13420 8504
rect 13460 8464 13469 8504
rect 13795 8464 13804 8504
rect 13844 8464 24364 8504
rect 24404 8464 24413 8504
rect 26537 8464 26668 8504
rect 26708 8464 26717 8504
rect 28361 8464 28492 8504
rect 28532 8464 28541 8504
rect 29251 8464 29260 8504
rect 29300 8464 29588 8504
rect 29779 8464 29788 8504
rect 29828 8464 29836 8504
rect 29876 8464 29959 8504
rect 30019 8464 30028 8504
rect 30068 8464 37940 8504
rect 38057 8464 38188 8504
rect 38228 8464 38237 8504
rect 5443 8380 5452 8420
rect 5492 8380 8132 8420
rect 9667 8380 9676 8420
rect 9716 8380 11308 8420
rect 11348 8380 11357 8420
rect 14179 8380 14188 8420
rect 14228 8380 22540 8420
rect 22580 8380 22589 8420
rect 23395 8380 23404 8420
rect 23444 8380 35884 8420
rect 35924 8380 35933 8420
rect 37900 8336 37940 8464
rect 38284 8420 38324 8548
rect 45292 8504 45332 8548
rect 46278 8504 46368 8524
rect 39689 8464 39820 8504
rect 39860 8464 39869 8504
rect 41539 8464 41548 8504
rect 41588 8464 43132 8504
rect 43172 8464 43181 8504
rect 45292 8464 46368 8504
rect 46278 8444 46368 8464
rect 38284 8380 41644 8420
rect 41684 8380 41693 8420
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 7651 8296 7660 8336
rect 7700 8296 8524 8336
rect 8564 8296 11500 8336
rect 11540 8296 11549 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 19276 8296 25172 8336
rect 25411 8296 25420 8336
rect 25460 8296 28300 8336
rect 28340 8296 28349 8336
rect 28579 8296 28588 8336
rect 28628 8296 31660 8336
rect 31700 8296 31709 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 37900 8296 38420 8336
rect 19276 8252 19316 8296
rect 9859 8212 9868 8252
rect 9908 8212 11828 8252
rect 11875 8212 11884 8252
rect 11924 8212 14036 8252
rect 0 8168 90 8188
rect 11788 8168 11828 8212
rect 0 8128 1228 8168
rect 1268 8128 1277 8168
rect 4012 8128 6988 8168
rect 7028 8128 7037 8168
rect 7363 8128 7372 8168
rect 7412 8128 7988 8168
rect 10243 8128 10252 8168
rect 10292 8128 11020 8168
rect 11060 8128 11069 8168
rect 11491 8128 11500 8168
rect 11540 8128 11644 8168
rect 11684 8128 11693 8168
rect 11788 8128 12028 8168
rect 12068 8128 13612 8168
rect 13652 8128 13661 8168
rect 13747 8128 13756 8168
rect 13796 8128 13804 8168
rect 13844 8128 13927 8168
rect 0 8108 90 8128
rect 1097 7960 1228 8000
rect 1268 7960 1277 8000
rect 1603 7960 1612 8000
rect 1652 7960 1661 8000
rect 0 7832 90 7852
rect 1612 7832 1652 7960
rect 4012 7916 4052 8128
rect 4195 8044 4204 8084
rect 4244 8044 6836 8084
rect 6115 7960 6124 8000
rect 6164 7960 6508 8000
rect 6548 7960 6557 8000
rect 5644 7916 5684 7925
rect 2563 7876 2572 7916
rect 2612 7876 2764 7916
rect 2804 7876 2813 7916
rect 3427 7876 3436 7916
rect 3476 7876 4012 7916
rect 4291 7876 4300 7916
rect 4340 7876 5155 7916
rect 5195 7876 5204 7916
rect 5684 7876 5932 7916
rect 5972 7876 5981 7916
rect 6211 7876 6220 7916
rect 6260 7876 6269 7916
rect 6473 7876 6604 7916
rect 6644 7876 6653 7916
rect 6796 7896 6836 8044
rect 7228 8044 7468 8084
rect 7508 8044 7517 8084
rect 7651 8044 7660 8084
rect 7700 8044 7709 8084
rect 7228 7958 7268 8044
rect 7660 8000 7700 8044
rect 7948 8000 7988 8128
rect 13996 8084 14036 8212
rect 14380 8212 19316 8252
rect 25132 8252 25172 8296
rect 25132 8212 38092 8252
rect 38132 8212 38141 8252
rect 14380 8168 14420 8212
rect 38380 8168 38420 8296
rect 42604 8296 45004 8336
rect 45044 8296 45053 8336
rect 42604 8168 42644 8296
rect 43180 8212 45484 8252
rect 45524 8212 45533 8252
rect 43180 8168 43220 8212
rect 46278 8168 46368 8188
rect 14284 8128 14420 8168
rect 14668 8128 15244 8168
rect 15284 8128 15293 8168
rect 15379 8128 15388 8168
rect 15428 8128 17740 8168
rect 17780 8128 17789 8168
rect 17923 8128 17932 8168
rect 17972 8128 23060 8168
rect 23107 8128 23116 8168
rect 23156 8128 23164 8168
rect 23204 8128 23287 8168
rect 23404 8128 29876 8168
rect 14284 8084 14324 8128
rect 8035 8044 8044 8084
rect 8084 8044 8468 8084
rect 7660 7960 7779 8000
rect 7819 7960 7828 8000
rect 7948 7960 8036 8000
rect 8122 7960 8131 8000
rect 8180 7960 8311 8000
rect 7225 7949 7268 7958
rect 4012 7867 4052 7876
rect 5644 7867 5684 7876
rect 0 7792 1652 7832
rect 0 7772 90 7792
rect 6220 7748 6260 7876
rect 6708 7856 6717 7896
rect 6757 7856 6836 7896
rect 6984 7876 6993 7916
rect 7033 7876 7042 7916
rect 7101 7876 7110 7916
rect 7150 7915 7159 7916
rect 7150 7876 7172 7915
rect 7265 7918 7268 7949
rect 7996 7916 8036 7960
rect 7225 7900 7265 7909
rect 7315 7876 7324 7916
rect 7364 7876 7372 7916
rect 7412 7876 7495 7916
rect 7651 7876 7660 7916
rect 7700 7876 7831 7916
rect 7882 7876 7891 7916
rect 7931 7876 7940 7916
rect 7987 7876 7996 7916
rect 8036 7876 8045 7916
rect 8092 7876 8236 7916
rect 8276 7876 8285 7916
rect 6988 7832 7028 7876
rect 7119 7875 7172 7876
rect 7132 7832 7172 7875
rect 7891 7832 7931 7876
rect 6955 7792 6988 7832
rect 7028 7792 7037 7832
rect 7132 7792 7276 7832
rect 7316 7792 7325 7832
rect 7468 7792 7564 7832
rect 7604 7792 7613 7832
rect 7852 7792 7931 7832
rect 1459 7708 1468 7748
rect 1508 7708 1708 7748
rect 1748 7708 1757 7748
rect 1843 7708 1852 7748
rect 1892 7708 1901 7748
rect 4963 7708 4972 7748
rect 5012 7708 5143 7748
rect 6220 7708 7084 7748
rect 7124 7708 7133 7748
rect 7180 7708 7372 7748
rect 7412 7708 7421 7748
rect 1852 7664 1892 7708
rect 1852 7624 7124 7664
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 0 7496 90 7516
rect 7084 7496 7124 7624
rect 7180 7580 7220 7708
rect 7468 7664 7508 7792
rect 7852 7664 7892 7792
rect 7267 7624 7276 7664
rect 7316 7624 7508 7664
rect 7843 7624 7852 7664
rect 7892 7624 7901 7664
rect 8092 7580 8132 7876
rect 8428 7832 8468 8044
rect 9580 8075 10772 8084
rect 9580 8044 10300 8075
rect 8515 7960 8524 8000
rect 8564 7960 8716 8000
rect 8756 7960 8765 8000
rect 9580 7916 9620 8044
rect 10340 8044 10772 8075
rect 10300 8026 10340 8035
rect 10060 7916 10100 7925
rect 10732 7916 10772 8044
rect 11500 8044 13708 8084
rect 13748 8044 13757 8084
rect 13996 8044 14324 8084
rect 11500 8000 11540 8044
rect 14668 8000 14708 8128
rect 23020 8084 23060 8128
rect 23404 8084 23444 8128
rect 14995 8044 15004 8084
rect 15044 8044 22924 8084
rect 22964 8044 22973 8084
rect 23020 8044 23444 8084
rect 23491 8044 23500 8084
rect 23540 8044 26132 8084
rect 26179 8044 26188 8084
rect 26228 8044 26572 8084
rect 26612 8044 26621 8084
rect 27340 8044 29780 8084
rect 26092 8000 26132 8044
rect 27340 8000 27380 8044
rect 11491 7960 11500 8000
rect 11540 7960 11549 8000
rect 11875 7960 11884 8000
rect 11924 7960 11933 8000
rect 12259 7960 12268 8000
rect 12308 7960 12317 8000
rect 12451 7960 12460 8000
rect 12500 7960 12631 8000
rect 13001 7960 13036 8000
rect 13076 7960 13132 8000
rect 13172 7960 13181 8000
rect 13385 7960 13516 8000
rect 13556 7960 13565 8000
rect 13987 7960 13996 8000
rect 14036 7960 14045 8000
rect 14105 7960 14188 8000
rect 14228 7960 14236 8000
rect 14276 7960 14285 8000
rect 14371 7960 14380 8000
rect 14420 7960 14708 8000
rect 14755 7960 14764 8000
rect 14804 7960 15092 8000
rect 15139 7960 15148 8000
rect 15188 7960 15197 8000
rect 15619 7960 15628 8000
rect 15668 7960 15724 8000
rect 15764 7960 15799 8000
rect 15907 7960 15916 8000
rect 15956 7960 15965 8000
rect 16291 7960 16300 8000
rect 16340 7960 17260 8000
rect 17300 7960 17309 8000
rect 18185 7960 18316 8000
rect 18356 7960 18365 8000
rect 18691 7960 18700 8000
rect 18740 7960 18749 8000
rect 18953 7960 19084 8000
rect 19124 7960 19133 8000
rect 19625 7960 19756 8000
rect 19796 7960 19805 8000
rect 20323 7960 20332 8000
rect 20372 7960 21772 8000
rect 21812 7960 21821 8000
rect 23273 7960 23404 8000
rect 23444 7960 23453 8000
rect 23657 7960 23788 8000
rect 23828 7960 23837 8000
rect 26092 7960 27380 8000
rect 27427 7960 27436 8000
rect 27476 7960 27607 8000
rect 28012 7960 28588 8000
rect 28628 7960 28637 8000
rect 28714 7960 28723 8000
rect 28763 7960 29068 8000
rect 29108 7960 29117 8000
rect 29321 7960 29452 8000
rect 29492 7960 29501 8000
rect 8515 7876 8524 7916
rect 8564 7876 9004 7916
rect 9044 7876 9053 7916
rect 9161 7876 9292 7916
rect 9332 7876 9341 7916
rect 9475 7876 9484 7916
rect 9524 7876 9580 7916
rect 9620 7876 9655 7916
rect 9929 7876 10060 7916
rect 10100 7876 10109 7916
rect 10217 7876 10339 7916
rect 10388 7876 10397 7916
rect 10723 7876 10732 7916
rect 10772 7876 10781 7916
rect 10915 7876 10924 7916
rect 10964 7876 11788 7916
rect 11828 7876 11837 7916
rect 10060 7867 10100 7876
rect 11884 7832 11924 7960
rect 12268 7916 12308 7960
rect 13996 7916 14036 7960
rect 12268 7876 13900 7916
rect 13940 7876 13949 7916
rect 13996 7876 14764 7916
rect 14804 7876 14813 7916
rect 15052 7832 15092 7960
rect 15148 7916 15188 7960
rect 15148 7876 15860 7916
rect 8314 7792 8323 7832
rect 8363 7792 8468 7832
rect 8755 7792 8764 7832
rect 8804 7792 8908 7832
rect 8948 7792 8957 7832
rect 9676 7792 9758 7832
rect 9798 7792 9807 7832
rect 10348 7792 10828 7832
rect 10868 7792 10877 7832
rect 11884 7792 13804 7832
rect 13844 7792 13853 7832
rect 14611 7792 14620 7832
rect 14660 7792 14956 7832
rect 14996 7792 15005 7832
rect 15052 7792 15628 7832
rect 15668 7792 15677 7832
rect 8851 7708 8860 7748
rect 8900 7708 8909 7748
rect 9370 7708 9379 7748
rect 9419 7708 9580 7748
rect 9620 7708 9629 7748
rect 8860 7580 8900 7708
rect 7180 7540 8132 7580
rect 8716 7540 8900 7580
rect 9676 7580 9716 7792
rect 10348 7748 10388 7792
rect 15820 7748 15860 7876
rect 15916 7832 15956 7960
rect 17932 7916 17972 7925
rect 18700 7916 18740 7960
rect 20332 7916 20372 7960
rect 21964 7916 22004 7925
rect 25420 7916 25460 7925
rect 27340 7916 27380 7960
rect 28012 7916 28052 7960
rect 29740 7916 29780 8044
rect 29836 8000 29876 8128
rect 29932 8128 31604 8168
rect 31651 8128 31660 8168
rect 31700 8128 34156 8168
rect 34196 8128 34205 8168
rect 34313 8128 34444 8168
rect 34484 8128 34493 8168
rect 36137 8128 36268 8168
rect 36308 8128 36317 8168
rect 36643 8128 36652 8168
rect 36692 8128 37084 8168
rect 37124 8128 37132 8168
rect 37172 8128 37181 8168
rect 38380 8128 41692 8168
rect 41732 8128 41741 8168
rect 42547 8128 42556 8168
rect 42596 8128 42644 8168
rect 42931 8128 42940 8168
rect 42980 8128 43220 8168
rect 43315 8128 43324 8168
rect 43364 8128 43948 8168
rect 43988 8128 43997 8168
rect 46243 8128 46252 8168
rect 46292 8128 46368 8168
rect 29827 7960 29836 8000
rect 29876 7960 29885 8000
rect 29932 7916 29972 8128
rect 31564 8084 31604 8128
rect 46278 8108 46368 8128
rect 30499 8044 30508 8084
rect 30548 8044 31468 8084
rect 31508 8044 31517 8084
rect 31564 8044 40780 8084
rect 40820 8044 40829 8084
rect 41827 8044 41836 8084
rect 41876 8044 44092 8084
rect 44132 8044 44141 8084
rect 30796 8000 30836 8044
rect 38572 8000 38612 8044
rect 30787 7960 30796 8000
rect 30836 7960 30845 8000
rect 32074 7960 32083 8000
rect 32123 7960 32236 8000
rect 32276 7960 32285 8000
rect 32681 7960 32812 8000
rect 32852 7960 32861 8000
rect 34252 7960 35828 8000
rect 36521 7960 36652 8000
rect 36692 7960 36701 8000
rect 36835 7960 36844 8000
rect 36884 7960 37015 8000
rect 37996 7960 38188 8000
rect 38228 7960 38237 8000
rect 38563 7960 38572 8000
rect 38612 7960 38621 8000
rect 41452 7960 41932 8000
rect 41972 7960 41981 8000
rect 42185 7960 42316 8000
rect 42356 7960 42365 8000
rect 42569 7960 42700 8000
rect 42740 7960 42749 8000
rect 42953 7960 43084 8000
rect 43124 7960 43133 8000
rect 43363 7960 43372 8000
rect 43412 7960 43660 8000
rect 43700 7960 43709 8000
rect 44323 7960 44332 8000
rect 44372 7960 44381 8000
rect 44515 7960 44524 8000
rect 44564 7960 44695 8000
rect 44899 7960 44908 8000
rect 44948 7960 45079 8000
rect 31372 7916 31412 7925
rect 34252 7916 34292 7960
rect 35788 7916 35828 7960
rect 36076 7916 36116 7925
rect 37996 7916 38036 7960
rect 39052 7916 39092 7925
rect 41356 7916 41396 7925
rect 16553 7876 16684 7916
rect 16724 7876 16733 7916
rect 17972 7876 18220 7916
rect 18260 7876 18269 7916
rect 18403 7876 18412 7916
rect 18452 7876 18740 7916
rect 19651 7876 19660 7916
rect 19700 7876 20372 7916
rect 20707 7876 20716 7916
rect 20756 7876 21004 7916
rect 21044 7876 21053 7916
rect 21833 7876 21964 7916
rect 22004 7876 22013 7916
rect 23107 7876 23116 7916
rect 23156 7876 24172 7916
rect 24212 7876 24221 7916
rect 25289 7876 25420 7916
rect 25460 7876 25469 7916
rect 25612 7876 25900 7916
rect 25940 7876 25949 7916
rect 26033 7876 26092 7916
rect 26132 7876 26155 7916
rect 26195 7876 26213 7916
rect 26266 7876 26275 7916
rect 26324 7876 26455 7916
rect 26659 7876 26668 7916
rect 26708 7876 26947 7916
rect 26987 7876 26996 7916
rect 27043 7876 27052 7916
rect 27092 7876 27101 7916
rect 27340 7876 27532 7916
rect 27572 7876 27581 7916
rect 28483 7876 28492 7916
rect 28540 7876 28663 7916
rect 29740 7876 29972 7916
rect 30298 7876 30307 7916
rect 30347 7876 30356 7916
rect 30403 7876 30412 7916
rect 30452 7876 30583 7916
rect 30761 7876 30892 7916
rect 30932 7876 30941 7916
rect 31075 7876 31084 7916
rect 31124 7876 31372 7916
rect 31412 7876 31660 7916
rect 31700 7876 31709 7916
rect 31882 7876 31891 7916
rect 31931 7876 31948 7916
rect 31988 7876 32071 7916
rect 32140 7876 33004 7916
rect 33044 7876 33053 7916
rect 34121 7876 34252 7916
rect 34292 7876 34301 7916
rect 34793 7876 34828 7916
rect 34868 7876 34924 7916
rect 34964 7876 34973 7916
rect 35779 7876 35788 7916
rect 35828 7876 36076 7916
rect 37978 7876 37987 7916
rect 38027 7876 38036 7916
rect 38083 7876 38092 7916
rect 38132 7876 38263 7916
rect 38345 7876 38469 7916
rect 38516 7876 38525 7916
rect 39562 7876 39571 7916
rect 39611 7876 39820 7916
rect 39860 7876 39869 7916
rect 40099 7876 40108 7916
rect 40148 7876 40157 7916
rect 17932 7867 17972 7876
rect 21964 7867 22004 7876
rect 25420 7867 25460 7876
rect 25612 7832 25652 7876
rect 27052 7832 27092 7876
rect 28012 7832 28052 7876
rect 30316 7832 30356 7876
rect 31372 7867 31412 7876
rect 32140 7832 32180 7876
rect 34252 7867 34292 7876
rect 36076 7867 36116 7876
rect 15916 7792 16780 7832
rect 16820 7792 16829 7832
rect 19315 7792 19324 7832
rect 19364 7792 21908 7832
rect 21868 7748 21908 7792
rect 22060 7792 24652 7832
rect 24692 7792 24701 7832
rect 25603 7792 25612 7832
rect 25652 7792 25661 7832
rect 26467 7792 26476 7832
rect 26516 7792 27092 7832
rect 27139 7792 27148 7832
rect 27188 7792 28052 7832
rect 28108 7792 30028 7832
rect 30068 7792 30077 7832
rect 30307 7792 30316 7832
rect 30356 7792 30403 7832
rect 31747 7792 31756 7832
rect 31796 7792 32180 7832
rect 32345 7792 32428 7832
rect 32468 7792 32476 7832
rect 32516 7792 32525 7832
rect 22060 7748 22100 7792
rect 28108 7748 28148 7792
rect 9850 7708 9859 7748
rect 9899 7708 9908 7748
rect 9955 7708 9964 7748
rect 10004 7708 10388 7748
rect 10522 7708 10531 7748
rect 10571 7708 10580 7748
rect 10819 7708 10828 7748
rect 10868 7708 11260 7748
rect 11300 7708 11309 7748
rect 12691 7708 12700 7748
rect 12740 7708 13132 7748
rect 13172 7708 13181 7748
rect 13267 7708 13276 7748
rect 13316 7708 14188 7748
rect 14228 7708 14237 7748
rect 14764 7708 15340 7748
rect 15380 7708 15484 7748
rect 15524 7708 15533 7748
rect 15820 7708 16012 7748
rect 16052 7708 16061 7748
rect 16147 7708 16156 7748
rect 16196 7708 16300 7748
rect 16340 7708 16349 7748
rect 16531 7708 16540 7748
rect 16580 7708 16972 7748
rect 17012 7708 17021 7748
rect 18115 7708 18124 7748
rect 18164 7708 18173 7748
rect 18547 7708 18556 7748
rect 18596 7708 18605 7748
rect 18931 7708 18940 7748
rect 18980 7708 19372 7748
rect 19412 7708 19421 7748
rect 19865 7708 19948 7748
rect 19988 7708 19996 7748
rect 20036 7708 20045 7748
rect 20563 7708 20572 7748
rect 20612 7708 21580 7748
rect 21620 7708 21629 7748
rect 21868 7708 22100 7748
rect 22147 7708 22156 7748
rect 22196 7708 22327 7748
rect 24019 7708 24028 7748
rect 24068 7708 25900 7748
rect 25940 7708 25949 7748
rect 26275 7708 26284 7748
rect 26324 7708 28148 7748
rect 28195 7708 28204 7748
rect 28244 7708 28828 7748
rect 28868 7708 28877 7748
rect 29059 7708 29068 7748
rect 29108 7708 29212 7748
rect 29252 7708 29261 7748
rect 29443 7708 29452 7748
rect 29492 7708 29596 7748
rect 29636 7708 29645 7748
rect 32035 7708 32044 7748
rect 32084 7708 32572 7748
rect 32612 7708 32621 7748
rect 33763 7708 33772 7748
rect 33812 7708 36412 7748
rect 36452 7708 36461 7748
rect 9868 7664 9908 7708
rect 9868 7624 10348 7664
rect 10388 7624 10397 7664
rect 10540 7580 10580 7708
rect 14764 7664 14804 7708
rect 11011 7624 11020 7664
rect 11060 7624 14804 7664
rect 18124 7580 18164 7708
rect 18556 7664 18596 7708
rect 39052 7664 39092 7876
rect 40108 7832 40148 7876
rect 41356 7832 41396 7876
rect 39619 7792 39628 7832
rect 39668 7792 40148 7832
rect 40195 7792 40204 7832
rect 40244 7792 41396 7832
rect 41452 7748 41492 7960
rect 44332 7916 44372 7960
rect 41635 7876 41644 7916
rect 41684 7876 44372 7916
rect 46278 7832 46368 7852
rect 42115 7792 42124 7832
rect 42164 7792 43220 7832
rect 44755 7792 44764 7832
rect 44804 7792 46368 7832
rect 43180 7748 43220 7792
rect 46278 7772 46368 7792
rect 39715 7708 39724 7748
rect 39764 7708 41492 7748
rect 41539 7708 41548 7748
rect 41588 7708 41836 7748
rect 41876 7708 41885 7748
rect 43180 7708 43420 7748
rect 43460 7708 43469 7748
rect 45139 7708 45148 7748
rect 45188 7708 45197 7748
rect 45148 7664 45188 7708
rect 18556 7624 18988 7664
rect 19028 7624 19037 7664
rect 19084 7624 20716 7664
rect 20756 7624 20765 7664
rect 28291 7624 28300 7664
rect 28340 7624 33964 7664
rect 34004 7624 34013 7664
rect 34147 7624 34156 7664
rect 34196 7624 39052 7664
rect 39092 7624 39101 7664
rect 45148 7624 46252 7664
rect 46292 7624 46301 7664
rect 9676 7540 10252 7580
rect 10292 7540 10301 7580
rect 10540 7540 10676 7580
rect 18115 7540 18124 7580
rect 18164 7540 18173 7580
rect 0 7456 1228 7496
rect 1268 7456 1277 7496
rect 6316 7456 6988 7496
rect 7028 7456 7037 7496
rect 7084 7456 8044 7496
rect 8084 7456 8093 7496
rect 0 7436 90 7456
rect 6316 7412 6356 7456
rect 8716 7412 8756 7540
rect 8908 7456 9428 7496
rect 9763 7456 9772 7496
rect 9812 7456 10540 7496
rect 10580 7456 10589 7496
rect 5897 7372 5980 7412
rect 6020 7372 6028 7412
rect 6068 7372 6077 7412
rect 6298 7372 6307 7412
rect 6347 7372 6356 7412
rect 6787 7372 6796 7412
rect 6836 7372 7660 7412
rect 7700 7372 7709 7412
rect 8506 7372 8515 7412
rect 8555 7372 8716 7412
rect 8756 7372 8765 7412
rect 8908 7328 8948 7456
rect 9388 7412 9428 7456
rect 2188 7288 2668 7328
rect 2708 7288 3860 7328
rect 2188 7244 2228 7288
rect 3820 7244 3860 7288
rect 6124 7288 6699 7328
rect 7075 7288 7084 7328
rect 7124 7288 8140 7328
rect 8180 7288 8189 7328
rect 8611 7288 8620 7328
rect 8660 7288 8948 7328
rect 9004 7372 9196 7412
rect 9236 7372 9245 7412
rect 9388 7372 10388 7412
rect 6124 7244 6164 7288
rect 6659 7244 6699 7288
rect 9004 7244 9044 7372
rect 10348 7328 10388 7372
rect 10636 7328 10676 7540
rect 19084 7412 19124 7624
rect 19171 7540 19180 7580
rect 19220 7540 19508 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 21763 7540 21772 7580
rect 21812 7540 21821 7580
rect 29923 7540 29932 7580
rect 29972 7540 30220 7580
rect 30260 7540 30269 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 19468 7496 19508 7540
rect 21772 7496 21812 7540
rect 46278 7496 46368 7516
rect 19468 7456 21196 7496
rect 21236 7456 21245 7496
rect 21772 7456 22004 7496
rect 10810 7372 10819 7412
rect 10859 7372 10868 7412
rect 13411 7372 13420 7412
rect 13460 7372 15668 7412
rect 17635 7372 17644 7412
rect 17684 7372 19124 7412
rect 19267 7372 19276 7412
rect 19316 7372 19756 7412
rect 19796 7372 19805 7412
rect 20227 7372 20236 7412
rect 20276 7372 21772 7412
rect 21812 7372 21821 7412
rect 9250 7288 9580 7328
rect 9620 7288 9629 7328
rect 9859 7288 9868 7328
rect 9908 7288 9964 7328
rect 10004 7288 10039 7328
rect 10348 7288 10484 7328
rect 9250 7244 9290 7288
rect 2179 7204 2188 7244
rect 2228 7204 2237 7244
rect 3305 7204 3436 7244
rect 3476 7204 3485 7244
rect 3811 7204 3820 7244
rect 3860 7204 3869 7244
rect 4387 7204 4396 7244
rect 4436 7235 5548 7244
rect 4436 7204 5068 7235
rect 3436 7186 3476 7195
rect 5108 7204 5548 7235
rect 5588 7204 5597 7244
rect 6115 7204 6124 7244
rect 6164 7204 6173 7244
rect 6307 7204 6316 7244
rect 6356 7204 6452 7244
rect 6499 7204 6508 7244
rect 6548 7204 6557 7244
rect 6641 7204 6650 7244
rect 6690 7204 6796 7244
rect 6836 7204 6845 7244
rect 7049 7204 7180 7244
rect 7220 7204 7229 7244
rect 7337 7204 7417 7244
rect 7457 7204 7468 7244
rect 7508 7204 7517 7244
rect 7642 7204 7651 7244
rect 7700 7204 7831 7244
rect 8410 7204 8419 7244
rect 8459 7204 8564 7244
rect 8721 7204 8730 7244
rect 8770 7204 8812 7244
rect 8852 7204 8901 7244
rect 8995 7204 9004 7244
rect 9044 7204 9053 7244
rect 9130 7235 9188 7244
rect 5068 7186 5108 7195
rect 0 7160 90 7180
rect 6412 7160 6452 7204
rect 6508 7160 6548 7204
rect 0 7120 1228 7160
rect 1268 7120 1277 7160
rect 1603 7120 1612 7160
rect 1652 7120 1661 7160
rect 5731 7120 5740 7160
rect 5780 7120 5789 7160
rect 6403 7120 6412 7160
rect 6452 7120 6461 7160
rect 6508 7120 7220 7160
rect 7267 7120 7276 7160
rect 7339 7120 7447 7160
rect 7913 7120 8044 7160
rect 8084 7120 8093 7160
rect 8275 7120 8284 7160
rect 8324 7120 8428 7160
rect 8468 7120 8477 7160
rect 0 7100 90 7120
rect 1612 7076 1652 7120
rect 172 7036 1652 7076
rect 3619 7036 3628 7076
rect 3668 7036 4300 7076
rect 4340 7036 4349 7076
rect 0 6824 90 6844
rect 172 6824 212 7036
rect 5740 6992 5780 7120
rect 6508 7076 6548 7120
rect 7180 7076 7220 7120
rect 5827 7036 5836 7076
rect 5876 7036 6548 7076
rect 7171 7036 7180 7076
rect 7220 7036 7229 7076
rect 7614 7036 7623 7076
rect 7663 7036 7756 7076
rect 7796 7036 7805 7076
rect 1459 6952 1468 6992
rect 1508 6952 1612 6992
rect 1652 6952 1661 6992
rect 1843 6952 1852 6992
rect 1892 6952 4780 6992
rect 4820 6952 4829 6992
rect 5251 6952 5260 6992
rect 5300 6952 5309 6992
rect 5740 6952 6124 6992
rect 6164 6952 6173 6992
rect 7834 6952 7843 6992
rect 7883 6952 7948 6992
rect 7988 6952 8023 6992
rect 5260 6908 5300 6952
rect 8524 6908 8564 7204
rect 9130 7195 9139 7235
rect 9179 7195 9188 7235
rect 9232 7204 9241 7244
rect 9281 7204 9290 7244
rect 9475 7204 9484 7244
rect 9524 7204 9572 7244
rect 9737 7204 9763 7244
rect 9803 7204 9868 7244
rect 9908 7204 9917 7244
rect 10156 7204 10339 7244
rect 10379 7204 10388 7244
rect 10444 7235 10484 7288
rect 10618 7319 10676 7328
rect 10618 7279 10627 7319
rect 10667 7279 10676 7319
rect 10828 7328 10868 7372
rect 15628 7328 15668 7372
rect 10828 7288 11060 7328
rect 14275 7288 14284 7328
rect 14324 7288 15572 7328
rect 15628 7288 19220 7328
rect 10618 7278 10676 7279
rect 11020 7244 11060 7288
rect 15532 7244 15572 7288
rect 9130 7194 9188 7195
rect 9148 7160 9188 7194
rect 9532 7160 9572 7204
rect 10156 7160 10196 7204
rect 10722 7204 10731 7244
rect 10771 7204 10780 7244
rect 10444 7186 10484 7195
rect 10732 7160 10772 7204
rect 10828 7193 10849 7233
rect 10889 7193 10898 7233
rect 11020 7204 11063 7244
rect 11103 7204 11112 7244
rect 11203 7204 11212 7244
rect 11252 7204 11308 7244
rect 11348 7204 11383 7244
rect 11561 7204 11596 7244
rect 11636 7204 11692 7244
rect 11732 7204 11741 7244
rect 11875 7204 11884 7244
rect 11924 7235 12884 7244
rect 11924 7204 12844 7235
rect 13411 7204 13420 7244
rect 13460 7204 13708 7244
rect 13748 7204 14572 7244
rect 14612 7204 14621 7244
rect 14825 7204 14956 7244
rect 14996 7204 15005 7244
rect 15523 7204 15532 7244
rect 15572 7204 15581 7244
rect 16387 7204 16396 7244
rect 16436 7235 16820 7244
rect 16436 7204 16780 7235
rect 8899 7120 8908 7160
rect 8948 7120 8957 7160
rect 9148 7120 9196 7160
rect 9236 7120 9245 7160
rect 9475 7120 9484 7160
rect 9524 7120 9572 7160
rect 9667 7120 9676 7160
rect 9716 7120 10156 7160
rect 10196 7120 10205 7160
rect 10693 7120 10732 7160
rect 10772 7120 10781 7160
rect 8908 6992 8948 7120
rect 10828 7076 10868 7193
rect 12844 7186 12884 7195
rect 14956 7186 14996 7195
rect 17530 7204 17539 7244
rect 17579 7204 17588 7244
rect 17635 7204 17644 7244
rect 17684 7204 17815 7244
rect 18019 7204 18028 7244
rect 18068 7204 18260 7244
rect 18473 7204 18508 7244
rect 18548 7235 18644 7244
rect 18548 7204 18604 7235
rect 16780 7186 16820 7195
rect 17548 7160 17588 7204
rect 18220 7160 18260 7204
rect 18691 7204 18700 7244
rect 18740 7235 19124 7244
rect 18740 7204 19084 7235
rect 18604 7186 18644 7195
rect 19084 7186 19124 7195
rect 19180 7160 19220 7288
rect 19564 7288 21292 7328
rect 21332 7288 21341 7328
rect 19564 7244 19604 7288
rect 21964 7286 22004 7456
rect 23596 7456 25804 7496
rect 25844 7456 25853 7496
rect 33148 7456 34252 7496
rect 34292 7456 34301 7496
rect 36940 7456 43372 7496
rect 43412 7456 43421 7496
rect 46243 7456 46252 7496
rect 46292 7456 46368 7496
rect 23596 7412 23636 7456
rect 33148 7412 33188 7456
rect 22339 7372 22348 7412
rect 22388 7372 23636 7412
rect 23683 7372 23692 7412
rect 23732 7372 23788 7412
rect 23828 7372 23863 7412
rect 24451 7372 24460 7412
rect 24500 7372 28204 7412
rect 28244 7372 28253 7412
rect 30185 7372 30220 7412
rect 30260 7372 30316 7412
rect 30356 7372 30365 7412
rect 31817 7372 31948 7412
rect 31988 7372 31997 7412
rect 33139 7372 33148 7412
rect 33188 7372 33197 7412
rect 33484 7372 33772 7412
rect 33812 7372 33821 7412
rect 22627 7288 22636 7328
rect 22676 7288 27148 7328
rect 27188 7288 27197 7328
rect 28780 7288 32908 7328
rect 32948 7288 32957 7328
rect 21954 7277 22004 7286
rect 19546 7204 19555 7244
rect 19595 7204 19604 7244
rect 19651 7204 19660 7244
rect 19700 7204 19709 7244
rect 19900 7204 20044 7244
rect 20084 7204 20093 7244
rect 20227 7204 20236 7244
rect 20276 7235 20660 7244
rect 20276 7204 20620 7235
rect 19660 7160 19700 7204
rect 11011 7120 11020 7160
rect 11060 7120 11203 7160
rect 11243 7120 11252 7160
rect 11299 7120 11308 7160
rect 11348 7120 11404 7160
rect 11444 7120 11479 7160
rect 12940 7120 13324 7160
rect 13364 7120 14860 7160
rect 14900 7120 14909 7160
rect 16972 7120 17588 7160
rect 17644 7120 18124 7160
rect 18164 7120 18173 7160
rect 18220 7120 18412 7160
rect 18452 7120 18461 7160
rect 19180 7120 19700 7160
rect 12940 7076 12980 7120
rect 16972 7076 17012 7120
rect 10147 7036 10156 7076
rect 10196 7036 10868 7076
rect 12835 7036 12844 7076
rect 12884 7036 12980 7076
rect 15017 7036 15148 7076
rect 15188 7036 15197 7076
rect 16963 7036 16972 7076
rect 17012 7036 17021 7076
rect 8908 6952 9676 6992
rect 9716 6952 9725 6992
rect 9772 6952 11692 6992
rect 11732 6952 11741 6992
rect 13027 6952 13036 6992
rect 13076 6952 13207 6992
rect 13555 6952 13564 6992
rect 13604 6952 14380 6992
rect 14420 6952 14429 6992
rect 16195 6952 16204 6992
rect 16244 6952 17452 6992
rect 17492 6952 17501 6992
rect 5260 6868 7276 6908
rect 7316 6868 7325 6908
rect 8524 6868 9484 6908
rect 9524 6868 9533 6908
rect 9772 6824 9812 6952
rect 10723 6868 10732 6908
rect 10772 6868 11500 6908
rect 11540 6868 11549 6908
rect 17644 6824 17684 7120
rect 18124 7076 18164 7120
rect 19900 7076 19940 7204
rect 20620 7186 20660 7195
rect 21100 7235 21484 7244
rect 21140 7204 21484 7235
rect 21524 7204 21533 7244
rect 21954 7237 21955 7277
rect 21995 7237 22004 7277
rect 28780 7244 28820 7288
rect 21954 7228 22004 7237
rect 22051 7204 22060 7244
rect 22100 7204 22231 7244
rect 22313 7204 22444 7244
rect 22484 7204 22493 7244
rect 22723 7204 22732 7244
rect 22772 7235 23060 7244
rect 22772 7204 23020 7235
rect 21100 7186 21140 7195
rect 23369 7204 23500 7244
rect 23540 7204 23549 7244
rect 24268 7235 24500 7244
rect 23020 7186 23060 7195
rect 23500 7186 23540 7195
rect 24308 7204 24500 7235
rect 24547 7204 24556 7244
rect 24596 7204 25516 7244
rect 25556 7204 25565 7244
rect 27209 7204 27340 7244
rect 27380 7204 27389 7244
rect 28579 7204 28588 7244
rect 28628 7204 28724 7244
rect 28771 7204 28780 7244
rect 28820 7204 28951 7244
rect 29897 7204 30028 7244
rect 30068 7204 30077 7244
rect 30377 7204 30508 7244
rect 30548 7204 30557 7244
rect 31756 7235 32948 7244
rect 24268 7186 24308 7195
rect 24460 7160 24500 7204
rect 27340 7186 27380 7195
rect 28684 7160 28724 7204
rect 30028 7160 30068 7195
rect 31796 7204 32948 7235
rect 31756 7160 31796 7195
rect 32908 7160 32948 7204
rect 33484 7235 33524 7372
rect 36940 7328 36980 7456
rect 46278 7436 46368 7456
rect 37075 7372 37084 7412
rect 37124 7372 37132 7412
rect 37172 7372 37255 7412
rect 43987 7372 43996 7412
rect 44036 7372 44812 7412
rect 44852 7372 44861 7412
rect 33571 7288 33580 7328
rect 33620 7288 36980 7328
rect 39043 7288 39052 7328
rect 39092 7288 40916 7328
rect 33859 7204 33868 7244
rect 33908 7204 34732 7244
rect 34772 7204 34781 7244
rect 34915 7204 34924 7244
rect 34964 7204 36940 7244
rect 36980 7204 36989 7244
rect 37507 7204 37516 7244
rect 37556 7235 38324 7244
rect 37556 7204 38284 7235
rect 33484 7186 33524 7195
rect 36460 7160 36500 7204
rect 38371 7204 38380 7244
rect 38420 7204 39532 7244
rect 39572 7204 39581 7244
rect 40282 7204 40291 7244
rect 40331 7204 40340 7244
rect 40387 7204 40396 7244
rect 40436 7204 40492 7244
rect 40532 7204 40567 7244
rect 40771 7204 40780 7244
rect 40820 7204 40829 7244
rect 38284 7160 38324 7195
rect 40300 7160 40340 7204
rect 40780 7160 40820 7204
rect 40876 7160 40916 7288
rect 41225 7204 41356 7244
rect 41396 7204 41405 7244
rect 41705 7204 41836 7244
rect 41876 7204 41885 7244
rect 41356 7186 41396 7195
rect 41836 7186 41876 7195
rect 46278 7160 46368 7180
rect 20009 7120 20140 7160
rect 20180 7120 20189 7160
rect 21322 7120 21331 7160
rect 21371 7120 21484 7160
rect 21524 7120 21533 7160
rect 22243 7120 22252 7160
rect 22292 7120 22540 7160
rect 22580 7120 22589 7160
rect 23116 7120 23404 7160
rect 23444 7120 23453 7160
rect 24460 7120 25708 7160
rect 25748 7120 25757 7160
rect 26057 7120 26188 7160
rect 26228 7120 26237 7160
rect 28675 7120 28684 7160
rect 28724 7120 28733 7160
rect 30028 7120 31796 7160
rect 32201 7120 32236 7160
rect 32276 7120 32332 7160
rect 32372 7120 32381 7160
rect 32707 7120 32716 7160
rect 32756 7120 32765 7160
rect 32899 7120 32908 7160
rect 32948 7120 32957 7160
rect 34531 7120 34540 7160
rect 34580 7120 34924 7160
rect 34964 7120 34973 7160
rect 36451 7120 36460 7160
rect 36500 7120 36509 7160
rect 36835 7120 36844 7160
rect 36884 7120 36893 7160
rect 37123 7120 37132 7160
rect 37172 7120 37420 7160
rect 37460 7120 37469 7160
rect 38284 7120 38900 7160
rect 39139 7120 39148 7160
rect 39188 7120 40012 7160
rect 40052 7120 40061 7160
rect 40300 7120 40396 7160
rect 40436 7120 40445 7160
rect 40579 7120 40588 7160
rect 40628 7120 40820 7160
rect 40867 7120 40876 7160
rect 40916 7120 40925 7160
rect 42058 7120 42067 7160
rect 42107 7120 42412 7160
rect 42452 7120 42461 7160
rect 43241 7120 43372 7160
rect 43412 7120 43421 7160
rect 43625 7120 43756 7160
rect 43796 7120 43805 7160
rect 44009 7120 44044 7160
rect 44084 7120 44140 7160
rect 44180 7120 44189 7160
rect 44515 7120 44524 7160
rect 44564 7120 44573 7160
rect 44777 7120 44908 7160
rect 44948 7120 44957 7160
rect 45139 7120 45148 7160
rect 45188 7120 46368 7160
rect 23116 7076 23156 7120
rect 32716 7076 32756 7120
rect 36844 7076 36884 7120
rect 18124 7036 21484 7076
rect 21524 7036 21533 7076
rect 21715 7036 21724 7076
rect 21764 7036 23156 7076
rect 23203 7036 23212 7076
rect 23252 7036 24212 7076
rect 30787 7036 30796 7076
rect 30836 7036 32228 7076
rect 32419 7036 32428 7076
rect 32468 7036 32756 7076
rect 32803 7036 32812 7076
rect 32852 7036 33292 7076
rect 33332 7036 33341 7076
rect 33763 7036 33772 7076
rect 33812 7036 36884 7076
rect 24172 6992 24212 7036
rect 32188 6992 32228 7036
rect 38860 6992 38900 7120
rect 39811 7036 39820 7076
rect 39860 7036 42172 7076
rect 42212 7036 42221 7076
rect 43603 7036 43612 7076
rect 43652 7036 43852 7076
rect 43892 7036 43901 7076
rect 44297 7036 44380 7076
rect 44420 7036 44428 7076
rect 44468 7036 44477 7076
rect 17827 6952 17836 6992
rect 17876 6952 19412 6992
rect 19651 6952 19660 6992
rect 19700 6952 24076 6992
rect 24116 6952 24125 6992
rect 24172 6952 25948 6992
rect 25988 6952 25997 6992
rect 26851 6952 26860 6992
rect 26900 6952 30412 6992
rect 30452 6952 30461 6992
rect 30595 6952 30604 6992
rect 30644 6952 32092 6992
rect 32132 6952 32141 6992
rect 32188 6952 32476 6992
rect 32516 6952 32525 6992
rect 35155 6952 35164 6992
rect 35204 6952 36500 6992
rect 36617 6952 36700 6992
rect 36740 6952 36748 6992
rect 36788 6952 36797 6992
rect 37123 6952 37132 6992
rect 37172 6952 37180 6992
rect 37220 6952 37303 6992
rect 37961 6952 38092 6992
rect 38132 6952 38141 6992
rect 38860 6952 39244 6992
rect 39284 6952 39772 6992
rect 39812 6952 39821 6992
rect 19372 6908 19412 6952
rect 19372 6868 32236 6908
rect 32276 6868 32285 6908
rect 34915 6868 34924 6908
rect 34964 6868 35692 6908
rect 35732 6868 35741 6908
rect 0 6784 212 6824
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 4675 6784 4684 6824
rect 4724 6784 9812 6824
rect 9859 6784 9868 6824
rect 9908 6784 18508 6824
rect 18548 6784 18557 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 19747 6784 19756 6824
rect 19796 6784 32084 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 0 6764 90 6784
rect 3427 6700 3436 6740
rect 3476 6700 7756 6740
rect 7796 6700 7805 6740
rect 11500 6700 12844 6740
rect 12884 6700 13076 6740
rect 14851 6700 14860 6740
rect 14900 6700 22924 6740
rect 22964 6700 22973 6740
rect 27427 6700 27436 6740
rect 27476 6700 31948 6740
rect 31988 6700 31997 6740
rect 6115 6616 6124 6656
rect 6164 6616 6547 6656
rect 6587 6616 6596 6656
rect 8410 6616 8419 6656
rect 8459 6616 8468 6656
rect 8803 6616 8812 6656
rect 8852 6616 10252 6656
rect 10292 6616 10732 6656
rect 10772 6616 10781 6656
rect 1459 6532 1468 6572
rect 1508 6532 3724 6572
rect 3764 6532 3773 6572
rect 3820 6532 4684 6572
rect 4724 6532 4733 6572
rect 7459 6532 7468 6572
rect 7508 6532 7517 6572
rect 0 6488 90 6508
rect 3820 6488 3860 6532
rect 7468 6488 7508 6532
rect 8428 6488 8468 6616
rect 9187 6532 9196 6572
rect 9236 6532 9524 6572
rect 9484 6488 9524 6532
rect 0 6448 1228 6488
rect 1268 6448 1277 6488
rect 1603 6448 1612 6488
rect 1652 6448 1661 6488
rect 1708 6448 1996 6488
rect 2036 6448 2045 6488
rect 2860 6448 3860 6488
rect 4361 6448 4492 6488
rect 4532 6448 4541 6488
rect 5251 6448 5260 6488
rect 5300 6448 5548 6488
rect 5588 6448 5597 6488
rect 6796 6448 6988 6488
rect 7028 6448 7037 6488
rect 7468 6448 7700 6488
rect 7939 6448 7948 6488
rect 7988 6448 8036 6488
rect 0 6428 90 6448
rect 1612 6320 1652 6448
rect 76 6280 1652 6320
rect 76 6172 116 6280
rect 0 6112 116 6172
rect 0 6092 90 6112
rect 1708 5900 1748 6448
rect 2563 6364 2572 6404
rect 2612 6364 2668 6404
rect 2708 6364 2743 6404
rect 2860 6236 2900 6448
rect 1843 6196 1852 6236
rect 1892 6196 1901 6236
rect 2227 6196 2236 6236
rect 2276 6196 2900 6236
rect 3916 6404 3956 6413
rect 5836 6404 5876 6413
rect 6796 6404 6836 6448
rect 7660 6415 7700 6448
rect 4291 6364 4300 6404
rect 4340 6364 4771 6404
rect 4811 6364 4820 6404
rect 4867 6364 4876 6404
rect 4916 6364 5047 6404
rect 5321 6364 5356 6404
rect 5396 6364 5452 6404
rect 5492 6364 5501 6404
rect 5876 6364 6028 6404
rect 6068 6364 6077 6404
rect 6346 6364 6355 6404
rect 6395 6364 6412 6404
rect 6452 6364 6535 6404
rect 6787 6364 6796 6404
rect 6836 6364 6845 6404
rect 6953 6364 7075 6404
rect 7124 6364 7133 6404
rect 7660 6375 7676 6415
rect 7716 6375 7725 6415
rect 7804 6404 7892 6425
rect 7996 6404 8036 6448
rect 8136 6448 8468 6488
rect 9161 6448 9292 6488
rect 9332 6448 9341 6488
rect 9475 6448 9484 6488
rect 9524 6448 9533 6488
rect 8136 6404 8176 6448
rect 8716 6404 8756 6413
rect 9580 6404 9620 6616
rect 9667 6532 9676 6572
rect 9716 6532 10580 6572
rect 10540 6488 10580 6532
rect 9699 6448 10292 6488
rect 10339 6448 10348 6488
rect 10388 6448 10397 6488
rect 10522 6448 10531 6488
rect 10571 6448 10580 6488
rect 10723 6448 10732 6488
rect 10772 6448 11020 6488
rect 11060 6448 11069 6488
rect 9699 6404 9739 6448
rect 10252 6404 10292 6448
rect 10348 6404 10388 6448
rect 7804 6364 7843 6404
rect 7883 6364 7892 6404
rect 7978 6364 7987 6404
rect 8027 6364 8036 6404
rect 8118 6364 8127 6404
rect 8167 6364 8176 6404
rect 8224 6364 8233 6404
rect 8276 6364 8407 6404
rect 8585 6364 8716 6404
rect 8756 6364 8765 6404
rect 9571 6364 9580 6404
rect 9620 6364 9629 6404
rect 9690 6364 9699 6404
rect 9739 6364 9748 6404
rect 9808 6364 9817 6404
rect 9857 6364 9964 6404
rect 10004 6364 10013 6404
rect 10107 6364 10116 6404
rect 172 5860 1748 5900
rect 0 5816 90 5836
rect 172 5816 212 5860
rect 1852 5816 1892 6196
rect 3916 6152 3956 6364
rect 4099 6280 4108 6320
rect 4148 6280 5740 6320
rect 5780 6280 5789 6320
rect 5836 6236 5876 6364
rect 7804 6320 7844 6364
rect 8716 6355 8756 6364
rect 9699 6320 9739 6364
rect 7049 6280 7180 6320
rect 7220 6280 7229 6320
rect 7804 6280 8044 6320
rect 8084 6280 8414 6320
rect 8454 6280 8463 6320
rect 9043 6280 9052 6320
rect 9092 6280 9484 6320
rect 9524 6280 9739 6320
rect 10156 6320 10196 6404
rect 10243 6364 10252 6404
rect 10292 6364 10301 6404
rect 10348 6364 10391 6404
rect 10431 6364 10440 6404
rect 10627 6364 10636 6404
rect 10676 6364 10924 6404
rect 10964 6364 10973 6404
rect 11057 6364 11066 6404
rect 11106 6364 11404 6404
rect 11444 6364 11453 6404
rect 10636 6320 10676 6364
rect 10156 6280 10292 6320
rect 10339 6280 10348 6320
rect 10388 6280 10676 6320
rect 10252 6236 10292 6280
rect 4195 6196 4204 6236
rect 4244 6196 4252 6236
rect 4292 6196 4375 6236
rect 5347 6196 5356 6236
rect 5396 6196 5876 6236
rect 6019 6196 6028 6236
rect 6068 6196 7747 6236
rect 7787 6196 7796 6236
rect 8489 6196 8620 6236
rect 8660 6196 8669 6236
rect 9929 6196 9955 6236
rect 9995 6196 10060 6236
rect 10100 6196 10109 6236
rect 10243 6196 10252 6236
rect 10292 6196 10301 6236
rect 11081 6196 11212 6236
rect 11252 6196 11261 6236
rect 11500 6152 11540 6700
rect 11788 6404 11828 6413
rect 13036 6404 13076 6700
rect 32044 6656 32084 6784
rect 36460 6740 36500 6952
rect 44524 6908 44564 7120
rect 46278 7100 46368 7120
rect 44755 6952 44764 6992
rect 44804 6952 46252 6992
rect 46292 6952 46301 6992
rect 37219 6868 37228 6908
rect 37268 6868 44564 6908
rect 46278 6824 46368 6844
rect 40291 6784 40300 6824
rect 40340 6784 43468 6824
rect 43508 6784 43517 6824
rect 46243 6784 46252 6824
rect 46292 6784 46368 6824
rect 46278 6764 46368 6784
rect 36460 6700 43564 6740
rect 43604 6700 43613 6740
rect 16483 6616 16492 6656
rect 16532 6616 18700 6656
rect 18740 6616 18749 6656
rect 20140 6616 23308 6656
rect 23348 6616 23357 6656
rect 23491 6616 23500 6656
rect 23540 6616 23692 6656
rect 23732 6616 23741 6656
rect 25795 6616 25804 6656
rect 25844 6616 26764 6656
rect 26804 6616 26813 6656
rect 28003 6616 28012 6656
rect 28052 6616 28348 6656
rect 28388 6616 28397 6656
rect 29011 6616 29020 6656
rect 29060 6616 30028 6656
rect 30068 6616 30077 6656
rect 30355 6616 30364 6656
rect 30404 6616 31372 6656
rect 31412 6616 31421 6656
rect 32044 6616 32428 6656
rect 32468 6616 32477 6656
rect 34339 6616 34348 6656
rect 34388 6616 37132 6656
rect 37172 6616 37181 6656
rect 40265 6616 40396 6656
rect 40436 6616 40445 6656
rect 44227 6616 44236 6656
rect 44276 6616 44380 6656
rect 44420 6616 44429 6656
rect 20140 6572 20180 6616
rect 14467 6532 14476 6572
rect 14516 6532 15092 6572
rect 17299 6532 17308 6572
rect 17348 6532 20180 6572
rect 20899 6532 20908 6572
rect 20948 6532 20956 6572
rect 20996 6532 21079 6572
rect 21379 6532 21388 6572
rect 21428 6532 40012 6572
rect 40052 6532 40061 6572
rect 40553 6532 40684 6572
rect 40724 6532 40733 6572
rect 14668 6404 14708 6413
rect 15052 6404 15092 6532
rect 46278 6488 46368 6508
rect 16553 6448 16588 6488
rect 16628 6448 16684 6488
rect 16724 6448 16733 6488
rect 16937 6448 17068 6488
rect 17108 6448 17117 6488
rect 17443 6448 17452 6488
rect 17492 6448 17548 6488
rect 17588 6448 17623 6488
rect 17705 6448 17788 6488
rect 17828 6448 17836 6488
rect 17876 6448 17885 6488
rect 18028 6448 18124 6488
rect 18164 6448 18173 6488
rect 18377 6448 18508 6488
rect 18548 6448 18557 6488
rect 19786 6448 19795 6488
rect 19835 6448 19948 6488
rect 19988 6448 19997 6488
rect 20515 6448 20524 6488
rect 20564 6448 20573 6488
rect 20707 6448 20716 6488
rect 20756 6448 20887 6488
rect 21427 6448 21436 6488
rect 21476 6448 21485 6488
rect 21667 6448 21676 6488
rect 21716 6448 21868 6488
rect 21908 6448 22060 6488
rect 22100 6448 22109 6488
rect 22156 6448 22348 6488
rect 22388 6448 22397 6488
rect 25577 6448 25708 6488
rect 25748 6448 25757 6488
rect 28579 6448 28588 6488
rect 28628 6448 28780 6488
rect 28820 6448 28829 6488
rect 29347 6448 29356 6488
rect 29396 6448 29588 6488
rect 29635 6448 29644 6488
rect 29684 6448 29740 6488
rect 29780 6448 29815 6488
rect 29932 6448 30124 6488
rect 30164 6448 30508 6488
rect 30548 6448 30557 6488
rect 30892 6448 32564 6488
rect 33187 6448 33196 6488
rect 33236 6448 34540 6488
rect 34580 6448 34589 6488
rect 37132 6448 38380 6488
rect 38420 6448 38429 6488
rect 44009 6448 44140 6488
rect 44180 6448 44189 6488
rect 44323 6448 44332 6488
rect 44372 6448 44524 6488
rect 44564 6448 44573 6488
rect 44707 6448 44716 6488
rect 44756 6448 44908 6488
rect 44948 6448 44957 6488
rect 45139 6448 45148 6488
rect 45188 6448 46368 6488
rect 16300 6404 16340 6413
rect 18028 6404 18068 6448
rect 19084 6404 19124 6413
rect 20524 6404 20564 6448
rect 11753 6364 11788 6404
rect 11828 6364 11884 6404
rect 11924 6364 11933 6404
rect 13027 6364 13036 6404
rect 13076 6364 13085 6404
rect 13289 6364 13420 6404
rect 13460 6364 13469 6404
rect 14508 6364 14572 6404
rect 14612 6364 14668 6404
rect 15043 6364 15052 6404
rect 15092 6364 15101 6404
rect 16265 6364 16300 6404
rect 16340 6364 16396 6404
rect 16436 6364 16445 6404
rect 18010 6364 18019 6404
rect 18059 6364 18068 6404
rect 18115 6364 18124 6404
rect 18164 6364 18173 6404
rect 18473 6364 18604 6404
rect 18644 6364 18653 6404
rect 19124 6364 19276 6404
rect 19316 6364 19325 6404
rect 19594 6364 19603 6404
rect 19643 6364 19660 6404
rect 19700 6364 19783 6404
rect 19843 6364 19852 6404
rect 19892 6364 20564 6404
rect 21436 6404 21476 6448
rect 22156 6404 22196 6448
rect 23500 6404 23540 6413
rect 26952 6404 26992 6413
rect 21436 6364 22196 6404
rect 22243 6364 22252 6404
rect 22292 6364 22924 6404
rect 22964 6364 22973 6404
rect 26371 6364 26380 6404
rect 26420 6364 26952 6404
rect 26992 6364 27340 6404
rect 27380 6364 27389 6404
rect 28073 6364 28204 6404
rect 28244 6364 28253 6404
rect 11788 6355 11828 6364
rect 14668 6320 14708 6364
rect 16300 6355 16340 6364
rect 14668 6280 15820 6320
rect 15860 6280 15869 6320
rect 16915 6280 16924 6320
rect 16964 6280 17740 6320
rect 17780 6280 17789 6320
rect 18124 6236 18164 6364
rect 19084 6355 19124 6364
rect 19276 6320 19316 6364
rect 23500 6320 23540 6364
rect 26952 6355 26992 6364
rect 29548 6320 29588 6448
rect 29932 6404 29972 6448
rect 30892 6404 30932 6448
rect 32524 6404 32564 6448
rect 33964 6404 34004 6448
rect 35212 6404 35252 6413
rect 36844 6404 36884 6413
rect 29731 6364 29740 6404
rect 29780 6364 29972 6404
rect 30019 6364 30028 6404
rect 30068 6364 30892 6404
rect 31939 6364 31948 6404
rect 31988 6364 32140 6404
rect 32180 6364 32189 6404
rect 33475 6364 33484 6404
rect 33524 6364 33772 6404
rect 33812 6364 33821 6404
rect 33955 6364 33964 6404
rect 34004 6364 34013 6404
rect 34819 6364 34828 6404
rect 34868 6364 35212 6404
rect 35395 6364 35404 6404
rect 35444 6364 35596 6404
rect 35636 6364 35645 6404
rect 36713 6364 36844 6404
rect 36884 6364 36893 6404
rect 30892 6355 30932 6364
rect 32524 6355 32564 6364
rect 19276 6280 20044 6320
rect 20084 6280 20093 6320
rect 20179 6280 20188 6320
rect 20228 6280 21196 6320
rect 21236 6280 21245 6320
rect 21475 6280 21484 6320
rect 21524 6280 21620 6320
rect 21955 6280 21964 6320
rect 22004 6280 22108 6320
rect 22148 6280 25036 6320
rect 25076 6280 25085 6320
rect 25804 6280 26860 6320
rect 26900 6280 26909 6320
rect 28291 6280 28300 6320
rect 28340 6280 29116 6320
rect 29156 6280 29165 6320
rect 29548 6280 30260 6320
rect 30307 6280 30316 6320
rect 30356 6280 30836 6320
rect 21580 6236 21620 6280
rect 25804 6236 25844 6280
rect 11587 6196 11596 6236
rect 11636 6196 11767 6236
rect 14729 6196 14860 6236
rect 14900 6196 14909 6236
rect 14956 6196 18164 6236
rect 20275 6196 20284 6236
rect 20324 6196 20524 6236
rect 20564 6196 20573 6236
rect 21580 6196 25844 6236
rect 25939 6196 25948 6236
rect 25988 6196 26284 6236
rect 26324 6196 26333 6236
rect 28483 6196 28492 6236
rect 28532 6196 29500 6236
rect 29540 6196 29549 6236
rect 30115 6196 30124 6236
rect 30164 6196 30173 6236
rect 14956 6152 14996 6196
rect 30124 6152 30164 6196
rect 3916 6112 4396 6152
rect 4436 6112 4445 6152
rect 6115 6112 6124 6152
rect 6164 6112 11540 6152
rect 12835 6112 12844 6152
rect 12884 6112 14996 6152
rect 18499 6112 18508 6152
rect 18548 6112 24308 6152
rect 24355 6112 24364 6152
rect 24404 6112 30164 6152
rect 30220 6152 30260 6280
rect 30796 6236 30836 6280
rect 30988 6280 32468 6320
rect 30988 6236 31028 6280
rect 32428 6236 32468 6280
rect 30569 6196 30700 6236
rect 30740 6196 30749 6236
rect 30796 6196 31028 6236
rect 32131 6196 32140 6236
rect 32180 6196 32332 6236
rect 32372 6196 32381 6236
rect 32428 6196 33004 6236
rect 33044 6196 33053 6236
rect 33772 6152 33812 6364
rect 35212 6355 35252 6364
rect 36844 6355 36884 6364
rect 35395 6196 35404 6236
rect 35444 6196 35596 6236
rect 35636 6196 35645 6236
rect 36067 6196 36076 6236
rect 36116 6196 37036 6236
rect 37076 6196 37085 6236
rect 37132 6152 37172 6448
rect 46278 6428 46368 6448
rect 40204 6404 40244 6413
rect 38825 6364 38956 6404
rect 38996 6364 39005 6404
rect 40073 6364 40204 6404
rect 40244 6364 40253 6404
rect 40204 6320 40244 6364
rect 37603 6280 37612 6320
rect 37652 6280 40244 6320
rect 38611 6196 38620 6236
rect 38660 6196 41068 6236
rect 41108 6196 41117 6236
rect 44755 6196 44764 6236
rect 44804 6196 44813 6236
rect 44764 6152 44804 6196
rect 46278 6152 46368 6172
rect 30220 6112 32908 6152
rect 32948 6112 32957 6152
rect 33772 6112 37172 6152
rect 40291 6112 40300 6152
rect 40340 6112 43948 6152
rect 43988 6112 43997 6152
rect 44764 6112 46368 6152
rect 24268 6068 24308 6112
rect 46278 6092 46368 6112
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 7267 6028 7276 6068
rect 7316 6028 8236 6068
rect 8276 6028 8285 6068
rect 8611 6028 8620 6068
rect 8660 6028 14092 6068
rect 14132 6028 14141 6068
rect 18403 6028 18412 6068
rect 18452 6028 19756 6068
rect 19796 6028 19805 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 22051 6028 22060 6068
rect 22100 6028 24172 6068
rect 24212 6028 24221 6068
rect 24268 6028 27436 6068
rect 27476 6028 27485 6068
rect 27715 6028 27724 6068
rect 27764 6028 28780 6068
rect 28820 6028 30124 6068
rect 30164 6028 30173 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 2092 5944 17588 5984
rect 17923 5944 17932 5984
rect 17972 5944 32812 5984
rect 32852 5944 32861 5984
rect 32908 5944 33772 5984
rect 33812 5944 33821 5984
rect 34723 5944 34732 5984
rect 34772 5944 38764 5984
rect 38804 5944 38813 5984
rect 2092 5900 2132 5944
rect 2083 5860 2092 5900
rect 2132 5860 2141 5900
rect 4483 5860 4492 5900
rect 4532 5860 5356 5900
rect 5396 5860 5405 5900
rect 5740 5860 5836 5900
rect 5876 5860 5885 5900
rect 6019 5860 6028 5900
rect 6068 5860 6077 5900
rect 9283 5860 9292 5900
rect 9332 5860 11692 5900
rect 11732 5860 11741 5900
rect 16963 5860 16972 5900
rect 17012 5860 17068 5900
rect 17108 5860 17143 5900
rect 5740 5816 5780 5860
rect 0 5776 212 5816
rect 1459 5776 1468 5816
rect 1508 5776 1612 5816
rect 1652 5776 1661 5816
rect 1852 5776 5780 5816
rect 5836 5776 5932 5816
rect 5972 5776 5981 5816
rect 0 5756 90 5776
rect 5836 5732 5876 5776
rect 6028 5732 6068 5860
rect 17548 5816 17588 5944
rect 32908 5900 32948 5944
rect 17635 5860 17644 5900
rect 17684 5860 23212 5900
rect 23252 5860 28820 5900
rect 31939 5860 31948 5900
rect 31988 5860 32948 5900
rect 32995 5860 33004 5900
rect 33044 5860 34540 5900
rect 34580 5860 34589 5900
rect 35561 5860 35596 5900
rect 35636 5860 35692 5900
rect 35732 5860 35741 5900
rect 28780 5816 28820 5860
rect 46278 5816 46368 5836
rect 6220 5776 6844 5816
rect 6884 5776 6893 5816
rect 7075 5776 7084 5816
rect 7124 5776 10348 5816
rect 10388 5776 10397 5816
rect 11107 5776 11116 5816
rect 11156 5776 11308 5816
rect 11348 5776 11357 5816
rect 13219 5776 13228 5816
rect 13268 5776 13364 5816
rect 17548 5776 20236 5816
rect 20276 5776 20285 5816
rect 20419 5776 20428 5816
rect 20468 5776 23884 5816
rect 23924 5776 23933 5816
rect 24163 5776 24172 5816
rect 24212 5776 25804 5816
rect 25844 5776 25853 5816
rect 28780 5776 29740 5816
rect 29780 5776 29789 5816
rect 30604 5776 30700 5816
rect 30740 5776 30749 5816
rect 32093 5776 32140 5816
rect 32180 5776 32189 5816
rect 35308 5776 36172 5816
rect 36212 5776 36460 5816
rect 36500 5776 36509 5816
rect 36643 5776 36652 5816
rect 36692 5776 39715 5816
rect 39755 5776 39764 5816
rect 45139 5776 45148 5816
rect 45188 5776 46368 5816
rect 6220 5732 6260 5776
rect 13324 5732 13364 5776
rect 30604 5732 30644 5776
rect 2153 5692 2284 5732
rect 2324 5692 2333 5732
rect 3401 5692 3532 5732
rect 3572 5692 3581 5732
rect 3628 5692 3916 5732
rect 3956 5692 4108 5732
rect 4148 5692 4157 5732
rect 4387 5692 4396 5732
rect 4436 5723 5204 5732
rect 4436 5692 5164 5723
rect 3532 5674 3572 5683
rect 67 5608 76 5648
rect 116 5608 1228 5648
rect 1268 5608 1277 5648
rect 1603 5608 1612 5648
rect 1652 5608 1661 5648
rect 1612 5564 1652 5608
rect 3628 5564 3668 5692
rect 5513 5692 5644 5732
rect 5684 5692 5693 5732
rect 5836 5692 5875 5732
rect 5915 5692 5924 5732
rect 5986 5692 5995 5732
rect 6035 5692 6068 5732
rect 6211 5692 6220 5732
rect 6260 5692 6269 5732
rect 6499 5692 6508 5732
rect 6548 5692 6557 5732
rect 6604 5692 6647 5732
rect 6687 5692 6696 5732
rect 7049 5692 7171 5732
rect 7220 5692 7229 5732
rect 7459 5692 7468 5732
rect 7508 5723 7852 5732
rect 7508 5692 7660 5723
rect 5164 5674 5204 5683
rect 5539 5608 5548 5648
rect 5588 5608 5597 5648
rect 5770 5639 5836 5648
rect 844 5524 1652 5564
rect 2179 5524 2188 5564
rect 2228 5524 3668 5564
rect 3715 5524 3724 5564
rect 3764 5524 4300 5564
rect 4340 5524 4349 5564
rect 0 5480 90 5500
rect 0 5440 76 5480
rect 116 5440 125 5480
rect 0 5420 90 5440
rect 0 5144 90 5164
rect 844 5144 884 5524
rect 5548 5480 5588 5608
rect 5770 5599 5779 5639
rect 5819 5608 5836 5639
rect 5876 5608 5959 5648
rect 6106 5608 6115 5648
rect 6155 5608 6164 5648
rect 6211 5608 6220 5648
rect 6260 5608 6316 5648
rect 6356 5608 6391 5648
rect 5819 5599 5828 5608
rect 5770 5598 5828 5599
rect 6124 5480 6164 5608
rect 1843 5440 1852 5480
rect 1892 5440 2380 5480
rect 2420 5440 2429 5480
rect 2563 5440 2572 5480
rect 2612 5440 5452 5480
rect 5492 5440 5501 5480
rect 5548 5440 6164 5480
rect 6508 5396 6548 5692
rect 6604 5648 6644 5692
rect 7700 5692 7852 5723
rect 7892 5692 7901 5732
rect 8131 5692 8140 5732
rect 8180 5692 8428 5732
rect 8468 5692 8477 5732
rect 8611 5692 8620 5732
rect 8660 5692 8669 5732
rect 8712 5692 8721 5732
rect 8761 5692 8892 5732
rect 9187 5692 9196 5732
rect 9236 5692 10444 5732
rect 10484 5692 10493 5732
rect 10723 5692 10732 5732
rect 10772 5692 10781 5732
rect 10998 5692 11007 5732
rect 11047 5692 11596 5732
rect 11636 5692 11645 5732
rect 11753 5692 11884 5732
rect 11924 5692 11933 5732
rect 12931 5692 12940 5732
rect 12980 5692 13132 5732
rect 13172 5692 13181 5732
rect 13315 5692 13324 5732
rect 13364 5692 13373 5732
rect 13603 5692 13612 5732
rect 13652 5692 14228 5732
rect 7660 5674 7700 5683
rect 8620 5648 8660 5692
rect 10732 5672 10780 5692
rect 11884 5674 11924 5683
rect 10740 5648 10780 5672
rect 6595 5608 6604 5648
rect 6644 5608 6653 5648
rect 8227 5608 8236 5648
rect 8276 5608 8285 5648
rect 8620 5608 8812 5648
rect 8852 5608 8861 5648
rect 9283 5608 9292 5648
rect 9332 5608 9341 5648
rect 9475 5608 9484 5648
rect 9524 5608 9676 5648
rect 9716 5608 9725 5648
rect 10051 5608 10060 5648
rect 10100 5608 10348 5648
rect 10388 5608 10397 5648
rect 10483 5608 10492 5648
rect 10532 5608 10580 5648
rect 10740 5608 11020 5648
rect 11060 5608 11069 5648
rect 13420 5608 14092 5648
rect 14132 5608 14141 5648
rect 8236 5564 8276 5608
rect 7651 5524 7660 5564
rect 7700 5524 8276 5564
rect 9292 5564 9332 5608
rect 10540 5564 10580 5608
rect 13420 5564 13460 5608
rect 9292 5524 9580 5564
rect 9620 5524 9629 5564
rect 9715 5524 9724 5564
rect 9764 5524 9772 5564
rect 9812 5524 9895 5564
rect 10540 5524 13460 5564
rect 14188 5564 14228 5692
rect 14572 5723 14612 5732
rect 14851 5692 14860 5732
rect 14900 5692 15235 5732
rect 15275 5692 15284 5732
rect 15331 5692 15340 5732
rect 15380 5692 15389 5732
rect 15689 5692 15724 5732
rect 15764 5692 15820 5732
rect 15860 5692 15869 5732
rect 16300 5723 16492 5732
rect 14572 5648 14612 5683
rect 14572 5608 15148 5648
rect 15188 5608 15197 5648
rect 15340 5564 15380 5692
rect 16340 5692 16492 5723
rect 16532 5692 16541 5732
rect 16780 5723 16820 5732
rect 16300 5674 16340 5683
rect 17033 5692 17164 5732
rect 17204 5692 17213 5732
rect 17539 5692 17548 5732
rect 17588 5723 18508 5732
rect 17588 5692 18412 5723
rect 15427 5608 15436 5648
rect 15476 5608 15820 5648
rect 15860 5608 15869 5648
rect 14188 5524 15380 5564
rect 16780 5564 16820 5683
rect 18452 5692 18508 5723
rect 18548 5692 18612 5732
rect 18761 5692 18892 5732
rect 18932 5692 18941 5732
rect 20380 5692 20812 5732
rect 20852 5692 20861 5732
rect 21340 5692 22004 5732
rect 22147 5692 22156 5732
rect 22196 5692 22327 5732
rect 23203 5692 23212 5732
rect 23252 5692 23404 5732
rect 23444 5692 23453 5732
rect 23587 5692 23596 5732
rect 23636 5692 23645 5732
rect 24067 5692 24076 5732
rect 24116 5692 24364 5732
rect 24404 5723 24884 5732
rect 24404 5692 24844 5723
rect 18412 5674 18452 5683
rect 20139 5650 20148 5690
rect 20188 5650 20276 5690
rect 20236 5648 20276 5650
rect 20380 5648 20420 5692
rect 20236 5608 20420 5648
rect 20515 5608 20524 5648
rect 20564 5608 20908 5648
rect 20948 5608 20957 5648
rect 21065 5608 21196 5648
rect 21236 5608 21245 5648
rect 21340 5564 21380 5692
rect 21964 5648 22004 5692
rect 22156 5674 22196 5683
rect 23596 5648 23636 5692
rect 24844 5674 24884 5683
rect 25036 5692 25411 5732
rect 25451 5692 25460 5732
rect 25507 5692 25516 5732
rect 25556 5692 25687 5732
rect 25865 5692 25900 5732
rect 25940 5692 25996 5732
rect 26036 5692 26045 5732
rect 26476 5723 26764 5732
rect 21571 5608 21580 5648
rect 21620 5608 21629 5648
rect 21946 5608 21955 5648
rect 21995 5608 22004 5648
rect 22243 5608 22252 5648
rect 22292 5608 23636 5648
rect 16780 5524 20140 5564
rect 20180 5524 20189 5564
rect 20323 5524 20332 5564
rect 20372 5524 21380 5564
rect 21580 5564 21620 5608
rect 25036 5564 25076 5692
rect 26516 5692 26764 5723
rect 26804 5692 26813 5732
rect 26956 5723 26996 5732
rect 26476 5648 26516 5683
rect 25123 5608 25132 5648
rect 25172 5608 25708 5648
rect 25748 5608 25996 5648
rect 26036 5608 26045 5648
rect 26380 5608 26516 5648
rect 26956 5648 26996 5683
rect 28876 5692 30316 5732
rect 30356 5692 30365 5732
rect 30586 5692 30595 5732
rect 30635 5692 30644 5732
rect 30691 5692 30700 5732
rect 30740 5692 30836 5732
rect 30883 5692 30892 5732
rect 30932 5692 31084 5732
rect 31124 5692 31133 5732
rect 31625 5723 31756 5732
rect 31625 5692 31660 5723
rect 28876 5648 28916 5692
rect 30796 5648 30836 5692
rect 31700 5692 31756 5723
rect 31796 5692 31805 5732
rect 32140 5723 32180 5776
rect 35308 5732 35348 5776
rect 46278 5756 46368 5776
rect 31660 5674 31700 5683
rect 32140 5674 32180 5683
rect 33768 5692 33859 5732
rect 33899 5692 33908 5732
rect 33955 5692 33964 5732
rect 34004 5692 34060 5732
rect 34100 5692 34135 5732
rect 34217 5692 34348 5732
rect 34388 5692 34397 5732
rect 34627 5692 34636 5732
rect 34676 5723 35348 5732
rect 34676 5692 34924 5723
rect 26956 5608 27148 5648
rect 27188 5608 27197 5648
rect 27593 5608 27724 5648
rect 27764 5608 27773 5648
rect 27907 5608 27916 5648
rect 27956 5608 27965 5648
rect 28099 5608 28108 5648
rect 28148 5608 28492 5648
rect 28532 5608 28541 5648
rect 28867 5608 28876 5648
rect 28916 5608 28925 5648
rect 29129 5608 29260 5648
rect 29300 5608 29309 5648
rect 29635 5608 29644 5648
rect 29684 5608 29693 5648
rect 30211 5608 30220 5648
rect 30260 5608 30269 5648
rect 30499 5608 30508 5648
rect 30548 5608 30836 5648
rect 31145 5608 31180 5648
rect 31220 5608 31276 5648
rect 31316 5608 31325 5648
rect 32515 5608 32524 5648
rect 32564 5608 32573 5648
rect 32620 5608 33044 5648
rect 33091 5608 33100 5648
rect 33140 5608 33271 5648
rect 33475 5608 33484 5648
rect 33524 5608 33533 5648
rect 26380 5564 26420 5608
rect 27916 5564 27956 5608
rect 29644 5564 29684 5608
rect 21580 5524 24460 5564
rect 24500 5524 24509 5564
rect 25027 5524 25036 5564
rect 25076 5524 25085 5564
rect 25411 5524 25420 5564
rect 25460 5524 26420 5564
rect 27187 5524 27196 5564
rect 27236 5524 27956 5564
rect 28147 5524 28156 5564
rect 28196 5524 29548 5564
rect 29588 5524 29597 5564
rect 29644 5524 30164 5564
rect 6931 5440 6940 5480
rect 6980 5440 7028 5480
rect 7171 5440 7180 5480
rect 7220 5440 8620 5480
rect 8660 5440 8669 5480
rect 8995 5440 9004 5480
rect 9044 5440 9052 5480
rect 9092 5440 9175 5480
rect 9379 5440 9388 5480
rect 9428 5440 9820 5480
rect 9860 5440 9869 5480
rect 10121 5440 10204 5480
rect 10244 5440 10252 5480
rect 10292 5440 11116 5480
rect 11156 5440 11165 5480
rect 11273 5440 11404 5480
rect 11444 5440 11453 5480
rect 11500 5440 14572 5480
rect 14612 5440 14621 5480
rect 14755 5440 14764 5480
rect 14804 5440 14813 5480
rect 18473 5440 18604 5480
rect 18644 5440 18653 5480
rect 20323 5440 20332 5480
rect 20372 5440 20428 5480
rect 20468 5440 20503 5480
rect 20755 5440 20764 5480
rect 20804 5440 21236 5480
rect 21427 5440 21436 5480
rect 21476 5440 21716 5480
rect 21811 5440 21820 5480
rect 21860 5440 21908 5480
rect 23779 5440 23788 5480
rect 23828 5440 27484 5480
rect 27524 5440 27533 5480
rect 27628 5440 28252 5480
rect 28292 5440 28301 5480
rect 28387 5440 28396 5480
rect 28436 5440 28636 5480
rect 28676 5440 28685 5480
rect 28780 5440 29020 5480
rect 29060 5440 29069 5480
rect 29164 5440 29404 5480
rect 29444 5440 29453 5480
rect 29731 5440 29740 5480
rect 29780 5440 29980 5480
rect 30020 5440 30029 5480
rect 5635 5356 5644 5396
rect 5684 5356 6548 5396
rect 6988 5312 7028 5440
rect 11500 5396 11540 5440
rect 9004 5356 11540 5396
rect 9004 5312 9044 5356
rect 14764 5312 14804 5440
rect 18499 5356 18508 5396
rect 18548 5356 20140 5396
rect 20180 5356 20189 5396
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 6883 5272 6892 5312
rect 6932 5272 7028 5312
rect 7084 5272 9044 5312
rect 10060 5272 13420 5312
rect 13460 5272 13469 5312
rect 14275 5272 14284 5312
rect 14324 5272 14804 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 19363 5272 19372 5312
rect 19412 5272 21140 5312
rect 1852 5188 6548 5228
rect 1852 5144 1892 5188
rect 0 5104 884 5144
rect 1843 5104 1852 5144
rect 1892 5104 1901 5144
rect 3113 5104 3196 5144
rect 3236 5104 3244 5144
rect 3284 5104 3293 5144
rect 5539 5104 5548 5144
rect 5588 5104 5644 5144
rect 5684 5104 5719 5144
rect 0 5084 90 5104
rect 6508 5060 6548 5188
rect 6595 5104 6604 5144
rect 6644 5104 6775 5144
rect 7084 5060 7124 5272
rect 10060 5228 10100 5272
rect 7363 5188 7372 5228
rect 7412 5188 10100 5228
rect 11788 5188 16396 5228
rect 16436 5188 16445 5228
rect 18508 5188 20812 5228
rect 20852 5188 20861 5228
rect 8515 5104 8524 5144
rect 8564 5104 10004 5144
rect 11434 5104 11443 5144
rect 11483 5104 11596 5144
rect 11636 5104 11645 5144
rect 9964 5060 10004 5104
rect 2371 5020 2380 5060
rect 2420 5020 3916 5060
rect 3956 5020 3965 5060
rect 4099 5020 4108 5060
rect 4148 5020 6452 5060
rect 6508 5020 7124 5060
rect 7171 5020 7180 5060
rect 7220 5020 8044 5060
rect 8084 5020 8180 5060
rect 8227 5020 8236 5060
rect 8276 5020 9908 5060
rect 6412 4976 6452 5020
rect 67 4936 76 4976
rect 116 4936 1228 4976
rect 1268 4936 1277 4976
rect 1603 4936 1612 4976
rect 1652 4936 1661 4976
rect 2179 4936 2188 4976
rect 2228 4936 2572 4976
rect 2612 4936 2621 4976
rect 2860 4936 2956 4976
rect 2996 4936 4148 4976
rect 1612 4892 1652 4936
rect 2860 4892 2900 4936
rect 4108 4892 4148 4936
rect 5836 4936 6028 4976
rect 6068 4936 6077 4976
rect 6211 4936 6220 4976
rect 6260 4936 6356 4976
rect 6412 4936 7892 4976
rect 5356 4892 5396 4901
rect 5836 4892 5876 4936
rect 172 4852 1652 4892
rect 2275 4852 2284 4892
rect 2324 4852 2900 4892
rect 3593 4852 3724 4892
rect 3764 4852 3773 4892
rect 3907 4852 3916 4892
rect 3956 4852 3965 4892
rect 4099 4852 4108 4892
rect 4148 4852 5300 4892
rect 0 4808 90 4828
rect 0 4768 76 4808
rect 116 4768 125 4808
rect 0 4748 90 4768
rect 0 4472 90 4492
rect 172 4472 212 4852
rect 3916 4808 3956 4852
rect 3916 4768 4204 4808
rect 4244 4768 4253 4808
rect 5260 4724 5300 4852
rect 5396 4852 5452 4892
rect 5492 4852 5527 4892
rect 5705 4852 5740 4892
rect 5780 4852 5836 4892
rect 5876 4852 5885 4892
rect 5946 4852 5955 4892
rect 5995 4852 6013 4892
rect 6064 4852 6073 4892
rect 6113 4852 6124 4892
rect 6164 4852 6253 4892
rect 5356 4843 5396 4852
rect 5973 4808 6013 4852
rect 5973 4768 6220 4808
rect 6260 4768 6269 4808
rect 1459 4684 1468 4724
rect 1508 4684 1517 4724
rect 2729 4684 2812 4724
rect 2852 4684 2860 4724
rect 2900 4684 3012 4724
rect 3898 4684 3907 4724
rect 3947 4684 3956 4724
rect 5260 4684 5492 4724
rect 5731 4684 5740 4724
rect 5780 4684 5911 4724
rect 1468 4556 1508 4684
rect 1468 4516 2900 4556
rect 0 4432 212 4472
rect 0 4412 90 4432
rect 2860 4388 2900 4516
rect 3916 4472 3956 4684
rect 5452 4640 5492 4684
rect 6316 4640 6356 4936
rect 6761 4852 6892 4892
rect 6932 4852 6941 4892
rect 7018 4883 7220 4892
rect 7018 4843 7027 4883
rect 7067 4852 7220 4883
rect 7267 4852 7276 4892
rect 7316 4852 7447 4892
rect 7625 4852 7747 4892
rect 7796 4852 7805 4892
rect 7067 4843 7076 4852
rect 7018 4842 7076 4843
rect 7180 4808 7220 4852
rect 7180 4768 7555 4808
rect 7595 4768 7604 4808
rect 7852 4724 7892 4936
rect 8140 4892 8180 5020
rect 8716 4976 8756 5020
rect 8707 4936 8716 4976
rect 8756 4936 8765 4976
rect 9283 4936 9292 4976
rect 9332 4936 9716 4976
rect 8236 4892 8276 4901
rect 9676 4892 9716 4936
rect 9868 4892 9908 5020
rect 9964 5020 10636 5060
rect 10676 5020 11020 5060
rect 11060 5020 11069 5060
rect 9964 4976 10004 5020
rect 11788 4976 11828 5188
rect 12329 5104 12412 5144
rect 12452 5104 12460 5144
rect 12500 5104 12509 5144
rect 12940 5104 17164 5144
rect 17204 5104 17213 5144
rect 12940 5060 12980 5104
rect 11884 5020 12980 5060
rect 13027 5020 13036 5060
rect 13076 5020 13085 5060
rect 13612 5020 13844 5060
rect 18211 5020 18220 5060
rect 18260 5020 18412 5060
rect 18452 5020 18461 5060
rect 9964 4936 10156 4976
rect 10196 4936 10205 4976
rect 11779 4936 11788 4976
rect 11828 4936 11837 4976
rect 10732 4892 10772 4901
rect 8140 4852 8236 4892
rect 8515 4852 8524 4892
rect 8564 4852 8812 4892
rect 8852 4852 8861 4892
rect 9065 4852 9196 4892
rect 9236 4852 9245 4892
rect 8236 4843 8276 4852
rect 9288 4851 9297 4891
rect 9337 4851 9346 4891
rect 9658 4852 9667 4892
rect 9707 4852 9716 4892
rect 9763 4852 9772 4892
rect 9812 4852 9821 4892
rect 9868 4852 10252 4892
rect 10292 4852 10301 4892
rect 10435 4852 10444 4892
rect 10484 4852 10732 4892
rect 11107 4852 11116 4892
rect 11156 4852 11220 4892
rect 11260 4852 11500 4892
rect 11540 4852 11549 4892
rect 9297 4808 9337 4851
rect 9772 4808 9812 4852
rect 10732 4843 10772 4852
rect 8707 4768 8716 4808
rect 8756 4768 9337 4808
rect 9379 4768 9388 4808
rect 9428 4768 10636 4808
rect 10676 4768 10685 4808
rect 11884 4724 11924 5020
rect 13036 4976 13076 5020
rect 13612 4976 13652 5020
rect 12163 4936 12172 4976
rect 12212 4936 12460 4976
rect 12500 4936 12509 4976
rect 12652 4936 13076 4976
rect 13123 4936 13132 4976
rect 13172 4936 13324 4976
rect 13364 4936 13373 4976
rect 13420 4936 13652 4976
rect 12652 4892 12692 4936
rect 13132 4892 13172 4936
rect 13420 4892 13460 4936
rect 13708 4892 13748 4901
rect 12634 4852 12643 4892
rect 12683 4852 12692 4892
rect 12739 4852 12748 4892
rect 12788 4852 12919 4892
rect 13027 4852 13036 4892
rect 13076 4852 13172 4892
rect 13219 4852 13228 4892
rect 13268 4852 13460 4892
rect 13577 4852 13708 4892
rect 13748 4852 13757 4892
rect 13228 4808 13268 4852
rect 13708 4843 13748 4852
rect 12643 4768 12652 4808
rect 12692 4768 13268 4808
rect 13804 4808 13844 5020
rect 15043 4936 15052 4976
rect 15092 4936 15340 4976
rect 15380 4936 15820 4976
rect 15860 4936 15869 4976
rect 15916 4936 16492 4976
rect 16532 4936 17108 4976
rect 15916 4892 15956 4936
rect 14153 4852 14227 4892
rect 14267 4852 14284 4892
rect 14324 4852 14333 4892
rect 14659 4852 14668 4892
rect 14708 4852 14851 4892
rect 14891 4852 14900 4892
rect 14947 4852 14956 4892
rect 14996 4852 15005 4892
rect 15305 4852 15436 4892
rect 15476 4852 15485 4892
rect 16291 4852 16300 4892
rect 16340 4852 16404 4892
rect 16444 4852 16471 4892
rect 16675 4852 16684 4892
rect 16724 4852 16972 4892
rect 17012 4852 17021 4892
rect 14956 4808 14996 4852
rect 15916 4843 15956 4852
rect 13804 4768 14996 4808
rect 17068 4724 17108 4936
rect 18220 4892 18260 4901
rect 18508 4892 18548 5188
rect 18595 5104 18604 5144
rect 18644 5104 18653 5144
rect 18787 5104 18796 5144
rect 18836 5104 21004 5144
rect 21044 5104 21053 5144
rect 18260 4852 18548 4892
rect 18604 4892 18644 5104
rect 21100 5060 21140 5272
rect 21196 5144 21236 5440
rect 21676 5396 21716 5440
rect 21868 5396 21908 5440
rect 27628 5396 27668 5440
rect 28780 5396 28820 5440
rect 21676 5356 21772 5396
rect 21812 5356 21821 5396
rect 21868 5356 22252 5396
rect 22292 5356 22301 5396
rect 27043 5356 27052 5396
rect 27092 5356 27668 5396
rect 27811 5356 27820 5396
rect 27860 5356 28820 5396
rect 29164 5312 29204 5440
rect 27907 5272 27916 5312
rect 27956 5272 29204 5312
rect 30124 5228 30164 5524
rect 21955 5188 21964 5228
rect 22004 5188 28876 5228
rect 28916 5188 28925 5228
rect 29932 5188 30164 5228
rect 21196 5104 26188 5144
rect 26228 5104 26237 5144
rect 26947 5104 26956 5144
rect 26996 5104 27148 5144
rect 27188 5104 27197 5144
rect 29932 5060 29972 5188
rect 30220 5144 30260 5608
rect 30796 5564 30836 5608
rect 32524 5564 32564 5608
rect 30796 5524 30988 5564
rect 31028 5524 31037 5564
rect 32371 5524 32380 5564
rect 32420 5524 32564 5564
rect 32620 5480 32660 5608
rect 33004 5564 33044 5608
rect 33484 5564 33524 5608
rect 32707 5524 32716 5564
rect 32756 5524 32860 5564
rect 32900 5524 32909 5564
rect 33004 5524 33196 5564
rect 33236 5524 33245 5564
rect 33484 5524 33676 5564
rect 33716 5524 33725 5564
rect 30499 5440 30508 5480
rect 30548 5440 32660 5480
rect 32755 5440 32764 5480
rect 32804 5440 32813 5480
rect 32995 5440 33004 5480
rect 33044 5440 33244 5480
rect 33284 5440 33293 5480
rect 32764 5228 32804 5440
rect 32764 5188 33620 5228
rect 33580 5144 33620 5188
rect 33768 5144 33808 5692
rect 34964 5692 35348 5723
rect 35404 5723 35596 5732
rect 34924 5674 34964 5683
rect 35444 5692 35596 5723
rect 35636 5692 35645 5732
rect 35945 5692 36076 5732
rect 36116 5692 36125 5732
rect 36233 5692 36355 5732
rect 36404 5692 36413 5732
rect 36809 5692 36940 5732
rect 36980 5692 36989 5732
rect 38057 5692 38188 5732
rect 38228 5692 38237 5732
rect 40090 5692 40099 5732
rect 40139 5692 40300 5732
rect 40340 5692 40349 5732
rect 41347 5692 41356 5732
rect 41396 5692 42068 5732
rect 35404 5674 35444 5683
rect 38188 5674 38228 5683
rect 33859 5608 33868 5648
rect 33908 5608 34444 5648
rect 34484 5608 34493 5648
rect 38755 5608 38764 5648
rect 38804 5608 38813 5648
rect 38947 5608 38956 5648
rect 38996 5608 39127 5648
rect 40675 5608 40684 5648
rect 40724 5608 40733 5648
rect 38764 5564 38804 5608
rect 42028 5564 42068 5692
rect 44393 5608 44524 5648
rect 44564 5608 44573 5648
rect 44777 5608 44908 5648
rect 44948 5608 44957 5648
rect 35596 5524 36364 5564
rect 36404 5524 36413 5564
rect 36739 5524 36748 5564
rect 36788 5524 38804 5564
rect 42019 5524 42028 5564
rect 42068 5524 42077 5564
rect 44755 5524 44764 5564
rect 44804 5524 45620 5564
rect 35596 5480 35636 5524
rect 34051 5440 34060 5480
rect 34100 5440 35636 5480
rect 36364 5480 36404 5524
rect 45580 5480 45620 5524
rect 46278 5480 46368 5500
rect 36364 5440 37516 5480
rect 37556 5440 37565 5480
rect 38249 5440 38380 5480
rect 38420 5440 38429 5480
rect 38515 5440 38524 5480
rect 38564 5440 38572 5480
rect 38612 5440 38695 5480
rect 39187 5440 39196 5480
rect 39236 5440 41972 5480
rect 45580 5440 46368 5480
rect 41932 5396 41972 5440
rect 46278 5420 46368 5440
rect 41932 5356 43084 5396
rect 43124 5356 43133 5396
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 46278 5144 46368 5164
rect 30058 5104 30067 5144
rect 30107 5104 30260 5144
rect 30307 5104 30316 5144
rect 30356 5104 31372 5144
rect 31412 5104 31421 5144
rect 31529 5104 31564 5144
rect 31604 5104 31660 5144
rect 31700 5104 31709 5144
rect 32227 5104 32236 5144
rect 32276 5104 32716 5144
rect 32756 5104 32765 5144
rect 33571 5104 33580 5144
rect 33620 5104 33629 5144
rect 33768 5104 34060 5144
rect 34100 5104 34109 5144
rect 36451 5104 36460 5144
rect 36500 5104 38132 5144
rect 38371 5104 38380 5144
rect 38420 5104 38900 5144
rect 39139 5104 39148 5144
rect 39188 5104 39292 5144
rect 39332 5104 39341 5144
rect 45139 5104 45148 5144
rect 45188 5104 46368 5144
rect 38092 5060 38132 5104
rect 19276 5020 20524 5060
rect 20564 5020 20573 5060
rect 21100 5020 21964 5060
rect 22004 5020 22013 5060
rect 22435 5020 22444 5060
rect 22484 5020 23060 5060
rect 23107 5020 23116 5060
rect 23156 5020 23165 5060
rect 23971 5020 23980 5060
rect 24020 5020 26380 5060
rect 26420 5020 26429 5060
rect 28579 5020 28588 5060
rect 28628 5020 29732 5060
rect 29932 5020 33388 5060
rect 33428 5020 33437 5060
rect 38092 5020 38516 5060
rect 18691 4936 18700 4976
rect 18740 4936 19180 4976
rect 19220 4936 19229 4976
rect 19276 4892 19316 5020
rect 19756 4892 19796 4901
rect 21964 4892 22004 4901
rect 23020 4892 23060 5020
rect 23116 4976 23156 5020
rect 29692 4976 29732 5020
rect 23116 4936 23500 4976
rect 23540 4936 23549 4976
rect 24547 4936 24556 4976
rect 24596 4936 25556 4976
rect 27209 4936 27340 4976
rect 27380 4936 27389 4976
rect 27523 4936 27532 4976
rect 27572 4936 27724 4976
rect 27764 4936 27773 4976
rect 28771 4936 28780 4976
rect 28820 4936 28876 4976
rect 28916 4936 28951 4976
rect 29692 4936 30260 4976
rect 31913 4936 32044 4976
rect 32084 4936 32093 4976
rect 32297 4936 32428 4976
rect 32468 4936 32477 4976
rect 32524 4936 33004 4976
rect 33044 4936 33053 4976
rect 33868 4936 34828 4976
rect 34868 4936 34877 4976
rect 35683 4936 35692 4976
rect 35732 4936 36172 4976
rect 36212 4936 36221 4976
rect 36355 4936 36364 4976
rect 36404 4936 36413 4976
rect 36809 4936 36940 4976
rect 36980 4936 36989 4976
rect 37769 4936 37900 4976
rect 37940 4936 37949 4976
rect 23980 4892 24020 4901
rect 25516 4892 25556 4936
rect 26764 4892 26804 4901
rect 29356 4892 29396 4901
rect 30220 4892 30260 4936
rect 32524 4892 32564 4936
rect 33868 4892 33908 4936
rect 36364 4892 36404 4936
rect 38476 4892 38516 5020
rect 38860 4976 38900 5104
rect 46278 5084 46368 5104
rect 43939 5020 43948 5060
rect 43988 5020 44948 5060
rect 44908 4976 44948 5020
rect 38860 4936 38996 4976
rect 39178 4936 39187 4976
rect 39227 4936 39532 4976
rect 39572 4936 39581 4976
rect 40963 4936 40972 4976
rect 41012 4936 41021 4976
rect 43555 4936 43564 4976
rect 43604 4936 44524 4976
rect 44564 4936 44573 4976
rect 44899 4936 44908 4976
rect 44948 4936 44957 4976
rect 38956 4892 38996 4936
rect 18604 4852 18691 4892
rect 18731 4852 18740 4892
rect 18787 4852 18796 4892
rect 18836 4852 18967 4892
rect 19267 4852 19276 4892
rect 19316 4852 19325 4892
rect 19555 4852 19564 4892
rect 19604 4852 19756 4892
rect 20201 4852 20275 4892
rect 20315 4852 20332 4892
rect 20372 4852 20381 4892
rect 20458 4852 20467 4892
rect 20507 4852 20564 4892
rect 20707 4852 20716 4892
rect 20756 4852 21676 4892
rect 21716 4852 21725 4892
rect 21833 4852 21964 4892
rect 22004 4852 22013 4892
rect 22156 4852 22444 4892
rect 22484 4852 22493 4892
rect 22627 4852 22636 4892
rect 22676 4852 22723 4892
rect 22763 4852 22807 4892
rect 23020 4852 23828 4892
rect 23971 4852 23980 4892
rect 24020 4852 24151 4892
rect 25123 4852 25132 4892
rect 25172 4852 25228 4892
rect 25268 4852 25303 4892
rect 25507 4852 25516 4892
rect 25556 4852 25565 4892
rect 26804 4852 27628 4892
rect 27668 4852 27677 4892
rect 28099 4852 28108 4892
rect 28148 4852 28291 4892
rect 28331 4852 28340 4892
rect 28387 4852 28396 4892
rect 28436 4852 28445 4892
rect 28675 4852 28684 4892
rect 28724 4852 28876 4892
rect 28916 4852 28925 4892
rect 29225 4852 29356 4892
rect 29396 4852 29405 4892
rect 29866 4852 29875 4892
rect 29915 4852 30028 4892
rect 30068 4852 30077 4892
rect 30211 4852 30220 4892
rect 30260 4852 30269 4892
rect 31433 4852 31476 4892
rect 31516 4852 31564 4892
rect 31604 4852 31613 4892
rect 31747 4852 31756 4892
rect 31796 4852 32564 4892
rect 32611 4852 32620 4892
rect 32660 4852 32669 4892
rect 34243 4852 34252 4892
rect 34292 4852 34348 4892
rect 34388 4852 34423 4892
rect 35453 4852 35596 4892
rect 35644 4852 35788 4892
rect 35828 4852 35837 4892
rect 35971 4852 35980 4892
rect 36020 4852 36460 4892
rect 36500 4852 36564 4892
rect 37402 4852 37411 4892
rect 37451 4852 37460 4892
rect 37507 4852 37516 4892
rect 37556 4852 37687 4892
rect 37865 4852 37996 4892
rect 38036 4852 38045 4892
rect 38955 4852 38964 4892
rect 39004 4852 39013 4892
rect 40282 4852 40291 4892
rect 40340 4852 40471 4892
rect 18220 4843 18260 4852
rect 19276 4808 19316 4852
rect 19756 4843 19796 4852
rect 20524 4808 20564 4852
rect 21964 4843 22004 4852
rect 22156 4808 22196 4852
rect 23788 4808 23828 4852
rect 23980 4843 24020 4852
rect 26764 4843 26804 4852
rect 18316 4768 19316 4808
rect 19939 4768 19948 4808
rect 19988 4768 20428 4808
rect 20468 4768 20477 4808
rect 20524 4768 20908 4808
rect 20948 4768 20957 4808
rect 22147 4768 22156 4808
rect 22196 4768 22205 4808
rect 22723 4768 22732 4808
rect 22772 4768 22828 4808
rect 22868 4768 23732 4808
rect 23779 4768 23788 4808
rect 23828 4768 23837 4808
rect 18316 4724 18356 4768
rect 23692 4724 23732 4768
rect 6451 4684 6460 4724
rect 6500 4684 7180 4724
rect 7220 4684 7229 4724
rect 7852 4684 11924 4724
rect 12019 4684 12028 4724
rect 12068 4684 14180 4724
rect 14249 4684 14284 4724
rect 14324 4684 14380 4724
rect 14420 4684 14429 4724
rect 14476 4684 16108 4724
rect 16148 4684 16157 4724
rect 16457 4684 16588 4724
rect 16628 4684 16637 4724
rect 17068 4684 18356 4724
rect 20035 4684 20044 4724
rect 20084 4684 23260 4724
rect 23300 4684 23309 4724
rect 23692 4684 25420 4724
rect 25460 4684 25469 4724
rect 25987 4684 25996 4724
rect 26036 4684 27100 4724
rect 27140 4684 27149 4724
rect 27244 4684 27484 4724
rect 27524 4684 27533 4724
rect 14140 4640 14180 4684
rect 14476 4640 14516 4684
rect 27244 4640 27284 4684
rect 4003 4600 4012 4640
rect 4052 4600 5396 4640
rect 5452 4600 6260 4640
rect 6316 4600 6988 4640
rect 7028 4600 7037 4640
rect 7084 4600 12212 4640
rect 14140 4600 14516 4640
rect 18595 4600 18604 4640
rect 18644 4600 19892 4640
rect 5356 4556 5396 4600
rect 6220 4556 6260 4600
rect 7084 4556 7124 4600
rect 12172 4556 12212 4600
rect 19852 4556 19892 4600
rect 19948 4600 21292 4640
rect 21332 4600 21868 4640
rect 21908 4600 21917 4640
rect 26179 4600 26188 4640
rect 26228 4600 27284 4640
rect 19948 4556 19988 4600
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 5356 4516 6164 4556
rect 6220 4516 7124 4556
rect 7372 4516 10732 4556
rect 10772 4516 10781 4556
rect 12172 4516 13364 4556
rect 13411 4516 13420 4556
rect 13460 4516 16820 4556
rect 17443 4516 17452 4556
rect 17492 4516 19660 4556
rect 19700 4516 19709 4556
rect 19852 4516 19988 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 20515 4516 20524 4556
rect 20564 4516 25516 4556
rect 25556 4516 25565 4556
rect 26083 4516 26092 4556
rect 26132 4516 27340 4556
rect 27380 4516 27389 4556
rect 6124 4472 6164 4516
rect 7372 4472 7412 4516
rect 13324 4472 13364 4516
rect 16780 4472 16820 4516
rect 28396 4472 28436 4852
rect 29356 4843 29396 4852
rect 32620 4808 32660 4852
rect 33868 4843 33908 4852
rect 37420 4808 37460 4852
rect 38476 4808 38516 4852
rect 46278 4808 46368 4828
rect 29452 4768 32188 4808
rect 32228 4768 32237 4808
rect 32323 4768 32332 4808
rect 32372 4768 32660 4808
rect 35683 4768 35692 4808
rect 35732 4768 35788 4808
rect 35828 4768 35863 4808
rect 36595 4768 36604 4808
rect 36644 4768 37364 4808
rect 37420 4768 37900 4808
rect 37940 4768 37949 4808
rect 38476 4768 39476 4808
rect 39785 4768 39907 4808
rect 39956 4768 39965 4808
rect 44755 4768 44764 4808
rect 44804 4768 46368 4808
rect 29452 4724 29492 4768
rect 28867 4684 28876 4724
rect 28916 4684 29492 4724
rect 30211 4684 30220 4724
rect 30260 4684 31804 4724
rect 31844 4684 31853 4724
rect 32332 4684 34484 4724
rect 32332 4640 32372 4684
rect 34444 4640 34484 4684
rect 35692 4684 35932 4724
rect 35972 4684 35981 4724
rect 36076 4684 36700 4724
rect 36740 4684 36749 4724
rect 35692 4640 35732 4684
rect 36076 4640 36116 4684
rect 29251 4600 29260 4640
rect 29300 4600 32372 4640
rect 32419 4600 32428 4640
rect 32468 4600 34348 4640
rect 34388 4600 34397 4640
rect 34444 4600 35732 4640
rect 35980 4600 36116 4640
rect 35980 4556 36020 4600
rect 29539 4516 29548 4556
rect 29588 4516 33964 4556
rect 34004 4516 34013 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 35875 4516 35884 4556
rect 35924 4516 36020 4556
rect 37324 4556 37364 4768
rect 39436 4724 39476 4768
rect 46278 4748 46368 4768
rect 39436 4684 42220 4724
rect 42260 4684 42269 4724
rect 37324 4516 44620 4556
rect 44660 4516 44669 4556
rect 46278 4472 46368 4492
rect 3916 4432 5972 4472
rect 6124 4432 7412 4472
rect 7747 4432 7756 4472
rect 7796 4432 9196 4472
rect 9236 4432 9245 4472
rect 9571 4432 9580 4472
rect 9620 4432 11444 4472
rect 13315 4432 13324 4472
rect 13364 4432 16684 4472
rect 16724 4432 16733 4472
rect 16780 4432 28436 4472
rect 28675 4432 28684 4472
rect 28724 4432 31124 4472
rect 31171 4432 31180 4472
rect 31220 4432 40300 4472
rect 40340 4432 40436 4472
rect 5932 4388 5972 4432
rect 11404 4388 11444 4432
rect 31084 4388 31124 4432
rect 2860 4348 5548 4388
rect 5588 4348 5597 4388
rect 5705 4348 5827 4388
rect 5876 4348 5885 4388
rect 5932 4348 6260 4388
rect 6490 4348 6499 4388
rect 6539 4348 6548 4388
rect 6979 4348 6988 4388
rect 7028 4348 7220 4388
rect 7267 4348 7276 4388
rect 7316 4348 7447 4388
rect 7651 4348 7660 4388
rect 7700 4348 10732 4388
rect 10772 4348 10781 4388
rect 11177 4348 11308 4388
rect 11348 4348 11357 4388
rect 11404 4348 13228 4388
rect 13268 4348 13277 4388
rect 14537 4348 14668 4388
rect 14708 4348 14717 4388
rect 16169 4348 16300 4388
rect 16340 4348 16349 4388
rect 18211 4348 18220 4388
rect 18260 4348 20276 4388
rect 22147 4348 22156 4388
rect 22196 4348 22972 4388
rect 23012 4348 23212 4388
rect 23252 4348 23261 4388
rect 25577 4348 25660 4388
rect 25700 4348 25708 4388
rect 25748 4348 25757 4388
rect 26371 4348 26380 4388
rect 26420 4348 27052 4388
rect 27092 4348 27101 4388
rect 27977 4348 28108 4388
rect 28148 4348 28157 4388
rect 28771 4348 28780 4388
rect 28820 4348 29740 4388
rect 29780 4348 29789 4388
rect 29897 4348 30028 4388
rect 30068 4348 30077 4388
rect 31084 4348 31852 4388
rect 31892 4348 32428 4388
rect 32468 4348 32477 4388
rect 32995 4348 33004 4388
rect 33044 4348 33053 4388
rect 33571 4348 33580 4388
rect 33620 4348 36076 4388
rect 36116 4348 36125 4388
rect 37769 4348 37900 4388
rect 37940 4348 37949 4388
rect 38035 4348 38044 4388
rect 38084 4348 38092 4388
rect 38132 4348 38215 4388
rect 6220 4304 6260 4348
rect 2467 4264 2476 4304
rect 2516 4264 2524 4304
rect 2564 4264 2647 4304
rect 5251 4264 5260 4304
rect 5300 4264 5492 4304
rect 5452 4220 5492 4264
rect 5644 4264 5740 4304
rect 5780 4264 5789 4304
rect 5923 4264 5932 4304
rect 5972 4264 6115 4304
rect 6155 4264 6164 4304
rect 6211 4264 6220 4304
rect 6260 4264 6269 4304
rect 5644 4220 5684 4264
rect 6508 4220 6548 4348
rect 7180 4304 7220 4348
rect 6595 4264 6604 4304
rect 6644 4264 6836 4304
rect 7180 4264 9331 4304
rect 9371 4264 9380 4304
rect 6796 4220 6836 4264
rect 10060 4220 10100 4348
rect 10636 4264 11269 4304
rect 11923 4264 11932 4304
rect 11972 4264 12940 4304
rect 12980 4264 12989 4304
rect 14275 4264 14284 4304
rect 14324 4264 15148 4304
rect 15188 4264 15197 4304
rect 16060 4264 16588 4304
rect 16628 4264 16637 4304
rect 18019 4264 18028 4304
rect 18068 4264 18644 4304
rect 10636 4220 10676 4264
rect 11229 4220 11269 4264
rect 16060 4220 16100 4264
rect 18604 4220 18644 4264
rect 19276 4264 20084 4304
rect 19276 4220 19316 4264
rect 2284 4180 3052 4220
rect 3092 4180 3101 4220
rect 3523 4180 3532 4220
rect 3572 4180 4108 4220
rect 4148 4211 4340 4220
rect 4148 4180 4300 4211
rect 0 4136 90 4156
rect 2284 4136 2324 4180
rect 4483 4180 4492 4220
rect 4532 4180 5059 4220
rect 5099 4180 5108 4220
rect 5225 4180 5356 4220
rect 5396 4180 5405 4220
rect 5452 4180 5495 4220
rect 5535 4180 5544 4220
rect 5626 4180 5635 4220
rect 5675 4180 5684 4220
rect 5731 4180 5740 4220
rect 5780 4180 5836 4220
rect 5876 4180 5911 4220
rect 6008 4180 6017 4220
rect 6068 4180 6188 4220
rect 6316 4211 6548 4220
rect 4300 4162 4340 4171
rect 6356 4180 6548 4211
rect 6651 4180 6660 4220
rect 6316 4162 6356 4171
rect 6700 4136 6740 4220
rect 6787 4180 6796 4220
rect 6836 4180 6845 4220
rect 7018 4180 7027 4220
rect 7067 4180 7076 4220
rect 7121 4180 7130 4220
rect 7170 4180 7180 4220
rect 7220 4180 7310 4220
rect 7546 4180 7555 4220
rect 7595 4180 7604 4220
rect 7651 4180 7660 4220
rect 7700 4180 7756 4220
rect 7796 4180 7831 4220
rect 7913 4180 8044 4220
rect 8084 4180 8093 4220
rect 8419 4180 8428 4220
rect 8468 4211 8660 4220
rect 8468 4180 8620 4211
rect 7036 4136 7076 4180
rect 0 4096 1228 4136
rect 1268 4096 1277 4136
rect 1603 4096 1612 4136
rect 1652 4096 1661 4136
rect 2275 4096 2284 4136
rect 2324 4096 2333 4136
rect 2537 4096 2668 4136
rect 2708 4096 2717 4136
rect 4396 4096 4684 4136
rect 4724 4096 4733 4136
rect 6700 4096 6796 4136
rect 6836 4096 6845 4136
rect 6979 4096 6988 4136
rect 7028 4096 7076 4136
rect 0 4076 90 4096
rect 1612 4052 1652 4096
rect 172 4012 1652 4052
rect 0 3800 90 3820
rect 172 3800 212 4012
rect 1459 3928 1468 3968
rect 1508 3928 1517 3968
rect 1843 3928 1852 3968
rect 1892 3928 2380 3968
rect 2420 3928 2429 3968
rect 2899 3928 2908 3968
rect 2948 3928 4300 3968
rect 4340 3928 4349 3968
rect 0 3760 212 3800
rect 0 3740 90 3760
rect 1468 3632 1508 3928
rect 4396 3800 4436 4096
rect 7564 4052 7604 4180
rect 8969 4180 9100 4220
rect 9140 4180 9149 4220
rect 9449 4180 9484 4220
rect 9524 4180 9571 4220
rect 9611 4180 9629 4220
rect 9672 4180 9681 4220
rect 9721 4180 9772 4220
rect 9812 4180 9881 4220
rect 10051 4180 10060 4220
rect 10100 4180 10109 4220
rect 10505 4180 10636 4220
rect 10676 4180 10685 4220
rect 10985 4180 11116 4220
rect 11156 4180 11165 4220
rect 11229 4180 12844 4220
rect 12884 4180 12893 4220
rect 13193 4180 13228 4220
rect 13268 4180 13324 4220
rect 13364 4180 13373 4220
rect 14476 4211 14516 4220
rect 8620 4162 8660 4171
rect 9100 4162 9140 4171
rect 7651 4096 7660 4136
rect 7700 4096 8140 4136
rect 8180 4096 8236 4136
rect 8276 4096 8285 4136
rect 9676 4052 9716 4180
rect 10636 4162 10676 4171
rect 11116 4162 11156 4171
rect 14851 4180 14860 4220
rect 14900 4180 15031 4220
rect 15148 4199 16100 4220
rect 15148 4180 16108 4199
rect 14476 4136 14516 4171
rect 15148 4136 15188 4180
rect 16060 4159 16108 4180
rect 16148 4159 16157 4199
rect 16483 4180 16492 4220
rect 16532 4180 16588 4220
rect 16628 4180 16663 4220
rect 17539 4180 17548 4220
rect 17588 4211 17876 4220
rect 17588 4180 17836 4211
rect 18586 4180 18595 4220
rect 18635 4180 18644 4220
rect 18691 4180 18700 4220
rect 18740 4180 18871 4220
rect 19075 4180 19084 4220
rect 19124 4180 19276 4220
rect 19316 4180 19325 4220
rect 19660 4211 19756 4220
rect 17836 4162 17876 4171
rect 19700 4180 19756 4211
rect 19796 4180 19948 4220
rect 19988 4180 19997 4220
rect 19660 4162 19700 4171
rect 4483 4012 4492 4052
rect 4532 4012 7604 4052
rect 8035 4012 8044 4052
rect 8084 4012 8812 4052
rect 8852 4012 9716 4052
rect 9772 4096 10156 4136
rect 10196 4096 10252 4136
rect 10292 4096 10301 4136
rect 11561 4096 11692 4136
rect 11732 4096 11741 4136
rect 11945 4096 11980 4136
rect 12020 4096 12076 4136
rect 12116 4096 12125 4136
rect 12451 4096 12460 4136
rect 12500 4096 12509 4136
rect 12874 4096 12883 4136
rect 12923 4096 12932 4136
rect 14476 4096 14764 4136
rect 14804 4096 15188 4136
rect 19171 4096 19180 4136
rect 19220 4096 19468 4136
rect 19508 4096 19517 4136
rect 9772 3968 9812 4096
rect 12233 4012 12316 4052
rect 12356 4012 12364 4052
rect 12404 4012 12413 4052
rect 4915 3928 4924 3968
rect 4964 3928 5740 3968
rect 5780 3928 5789 3968
rect 7555 3928 7564 3968
rect 7604 3928 8428 3968
rect 8468 3928 9812 3968
rect 10243 3928 10252 3968
rect 10292 3928 12172 3968
rect 12212 3928 12221 3968
rect 12460 3884 12500 4096
rect 12892 4052 12932 4096
rect 20044 4052 20084 4264
rect 20236 4220 20276 4348
rect 33004 4304 33044 4348
rect 20323 4264 20332 4304
rect 20372 4264 20948 4304
rect 20995 4264 21004 4304
rect 21044 4264 27188 4304
rect 27331 4264 27340 4304
rect 27380 4264 29644 4304
rect 29684 4264 30452 4304
rect 31267 4264 31276 4304
rect 31316 4264 31796 4304
rect 33004 4264 36308 4304
rect 37699 4264 37708 4304
rect 37748 4264 38428 4304
rect 38468 4264 38477 4304
rect 40003 4264 40012 4304
rect 40052 4264 40156 4304
rect 40196 4264 40205 4304
rect 20908 4220 20948 4264
rect 20140 4211 20276 4220
rect 20180 4180 20276 4211
rect 20611 4180 20620 4220
rect 20660 4180 20803 4220
rect 20843 4180 20852 4220
rect 20899 4180 20908 4220
rect 20948 4180 20957 4220
rect 21187 4180 21196 4220
rect 21236 4180 21292 4220
rect 21332 4180 21367 4220
rect 21737 4180 21868 4220
rect 21908 4180 21917 4220
rect 22313 4180 22387 4220
rect 22427 4180 22444 4220
rect 22484 4180 22493 4220
rect 22570 4180 22579 4220
rect 22619 4180 23348 4220
rect 23395 4180 23404 4220
rect 23444 4180 23828 4220
rect 23875 4180 23884 4220
rect 23924 4180 26284 4220
rect 26324 4180 26612 4220
rect 26659 4180 26668 4220
rect 26708 4180 26839 4220
rect 20140 4162 20180 4171
rect 21868 4162 21908 4171
rect 23308 4136 23348 4180
rect 23788 4136 23828 4180
rect 26572 4136 26612 4180
rect 20236 4096 21388 4136
rect 21428 4096 21437 4136
rect 22339 4096 22348 4136
rect 22388 4096 22732 4136
rect 22772 4096 22781 4136
rect 23299 4096 23308 4136
rect 23348 4096 23357 4136
rect 23779 4096 23788 4136
rect 23828 4096 23837 4136
rect 24163 4096 24172 4136
rect 24212 4096 24268 4136
rect 24308 4096 24343 4136
rect 24713 4096 24844 4136
rect 24884 4096 24893 4136
rect 25027 4096 25036 4136
rect 25076 4096 25420 4136
rect 25460 4096 25612 4136
rect 25652 4096 25661 4136
rect 25891 4096 25900 4136
rect 25940 4096 25996 4136
rect 26036 4096 26071 4136
rect 26371 4096 26380 4136
rect 26420 4096 26429 4136
rect 26572 4096 27052 4136
rect 27092 4096 27101 4136
rect 20236 4052 20276 4096
rect 12892 4012 12940 4052
rect 12980 4012 12989 4052
rect 13075 4012 13084 4052
rect 13124 4012 19604 4052
rect 20044 4012 20276 4052
rect 20323 4012 20332 4052
rect 20372 4012 21964 4052
rect 22004 4012 22013 4052
rect 12691 3928 12700 3968
rect 12740 3928 13036 3968
rect 13076 3928 13085 3968
rect 15043 3928 15052 3968
rect 15092 3928 19468 3968
rect 19508 3928 19517 3968
rect 19564 3884 19604 4012
rect 20227 3928 20236 3968
rect 20276 3928 20371 3968
rect 20411 3928 20420 3968
rect 21187 3928 21196 3968
rect 21236 3928 22828 3968
rect 22868 3928 22877 3968
rect 23011 3928 23020 3968
rect 23060 3928 23068 3968
rect 23108 3928 23191 3968
rect 23417 3928 23500 3968
rect 23540 3928 23548 3968
rect 23588 3928 23597 3968
rect 23801 3928 23884 3968
rect 23924 3928 23932 3968
rect 23972 3928 23981 3968
rect 24451 3928 24460 3968
rect 24500 3928 24604 3968
rect 24644 3928 24653 3968
rect 24844 3884 24884 4096
rect 26380 4052 26420 4096
rect 27148 4052 27188 4264
rect 30412 4220 30452 4264
rect 31756 4220 31796 4264
rect 27235 4180 27244 4220
rect 27284 4211 27956 4220
rect 27284 4180 27916 4211
rect 28457 4180 28588 4220
rect 28628 4180 28637 4220
rect 29836 4211 29932 4220
rect 27916 4162 27956 4171
rect 29876 4180 29932 4211
rect 29972 4180 30007 4220
rect 30412 4180 30836 4220
rect 31258 4180 31267 4220
rect 31307 4180 31316 4220
rect 31363 4180 31372 4220
rect 31412 4180 31508 4220
rect 31747 4180 31756 4220
rect 31796 4180 32044 4220
rect 32084 4180 32093 4220
rect 32332 4211 32428 4220
rect 29836 4162 29876 4171
rect 30796 4136 30836 4180
rect 31276 4136 31316 4180
rect 30403 4096 30412 4136
rect 30452 4096 30508 4136
rect 30548 4096 30583 4136
rect 30787 4096 30796 4136
rect 30836 4096 30845 4136
rect 31267 4096 31276 4136
rect 31316 4096 31363 4136
rect 31468 4052 31508 4180
rect 32372 4180 32428 4211
rect 32468 4180 32503 4220
rect 32812 4211 32852 4220
rect 32332 4162 32372 4171
rect 33750 4180 33759 4220
rect 33799 4180 33812 4220
rect 33859 4180 33868 4220
rect 33908 4180 34039 4220
rect 34243 4180 34252 4220
rect 34292 4180 34423 4220
rect 34627 4180 34636 4220
rect 34676 4211 34868 4220
rect 34676 4180 34828 4211
rect 31721 4096 31852 4136
rect 31892 4096 31901 4136
rect 25116 4012 25228 4052
rect 25268 4012 25276 4052
rect 25316 4012 26276 4052
rect 26380 4012 26572 4052
rect 26612 4012 26621 4052
rect 27148 4012 31508 4052
rect 25420 3928 25756 3968
rect 25796 3928 25805 3968
rect 25900 3928 26140 3968
rect 26180 3928 26189 3968
rect 25420 3884 25460 3928
rect 4483 3844 4492 3884
rect 4532 3844 5644 3884
rect 5684 3844 5693 3884
rect 5827 3844 5836 3884
rect 5876 3844 7372 3884
rect 7412 3844 7421 3884
rect 9187 3844 9196 3884
rect 9236 3844 12268 3884
rect 12308 3844 12317 3884
rect 12460 3844 13172 3884
rect 13699 3844 13708 3884
rect 13748 3844 15092 3884
rect 15811 3844 15820 3884
rect 15860 3844 19316 3884
rect 19564 3844 24884 3884
rect 25027 3844 25036 3884
rect 25076 3844 25460 3884
rect 13132 3800 13172 3844
rect 15052 3800 15092 3844
rect 19276 3800 19316 3844
rect 25900 3800 25940 3928
rect 26236 3884 26276 4012
rect 27139 3928 27148 3968
rect 27188 3928 30172 3968
rect 30212 3928 30221 3968
rect 30547 3928 30556 3968
rect 30596 3928 31564 3968
rect 31604 3928 31613 3968
rect 26236 3844 32332 3884
rect 32372 3844 32381 3884
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 4396 3760 11212 3800
rect 11252 3760 11261 3800
rect 13132 3760 14956 3800
rect 14996 3760 15005 3800
rect 15052 3760 16876 3800
rect 16916 3760 16925 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 19276 3760 21004 3800
rect 21044 3760 21053 3800
rect 21292 3760 25172 3800
rect 25219 3760 25228 3800
rect 25268 3760 25940 3800
rect 28675 3760 28684 3800
rect 28724 3760 30220 3800
rect 30260 3760 30269 3800
rect 2860 3676 5164 3716
rect 5204 3676 5213 3716
rect 5260 3676 14860 3716
rect 14900 3676 14909 3716
rect 15052 3676 21196 3716
rect 21236 3676 21245 3716
rect 2860 3632 2900 3676
rect 5260 3632 5300 3676
rect 15052 3632 15092 3676
rect 21292 3632 21332 3760
rect 25132 3716 25172 3760
rect 25132 3676 26092 3716
rect 26132 3676 26141 3716
rect 26467 3676 26476 3716
rect 26516 3676 27052 3716
rect 27092 3676 27101 3716
rect 29827 3676 29836 3716
rect 29876 3676 30508 3716
rect 30548 3676 30557 3716
rect 31952 3676 32332 3716
rect 32372 3676 32381 3716
rect 31952 3632 31992 3676
rect 32812 3632 32852 4171
rect 33772 4136 33812 4180
rect 34828 4162 34868 4171
rect 35308 4211 35692 4220
rect 35348 4180 35692 4211
rect 35732 4180 35741 4220
rect 35308 4162 35348 4171
rect 36268 4136 36308 4264
rect 36451 4180 36460 4220
rect 36500 4180 36631 4220
rect 37603 4180 37612 4220
rect 37652 4211 37783 4220
rect 37652 4180 37708 4211
rect 37748 4180 37783 4211
rect 37708 4162 37748 4171
rect 40396 4136 40436 4432
rect 45148 4432 46368 4472
rect 45148 4304 45188 4432
rect 46278 4412 46368 4432
rect 45139 4264 45148 4304
rect 45188 4264 45197 4304
rect 43267 4180 43276 4220
rect 43316 4180 44564 4220
rect 44524 4136 44564 4180
rect 46278 4136 46368 4156
rect 32995 4096 33004 4136
rect 33044 4096 33388 4136
rect 33428 4096 33437 4136
rect 33571 4096 33580 4136
rect 33620 4096 33812 4136
rect 34217 4096 34348 4136
rect 34388 4096 34397 4136
rect 35404 4096 35884 4136
rect 35924 4096 35933 4136
rect 36259 4096 36268 4136
rect 36308 4096 36317 4136
rect 38275 4096 38284 4136
rect 38324 4096 38333 4136
rect 38537 4096 38668 4136
rect 38708 4096 38717 4136
rect 38851 4096 38860 4136
rect 38900 4096 39031 4136
rect 39619 4096 39628 4136
rect 39668 4096 39724 4136
rect 39764 4096 39799 4136
rect 40387 4096 40396 4136
rect 40436 4096 40445 4136
rect 40684 4096 44140 4136
rect 44180 4096 44189 4136
rect 44515 4096 44524 4136
rect 44564 4096 44573 4136
rect 44620 4096 44908 4136
rect 44948 4096 44957 4136
rect 45676 4096 46368 4136
rect 35404 4052 35444 4096
rect 38284 4052 38324 4096
rect 40684 4052 40724 4096
rect 44620 4052 44660 4096
rect 45676 4052 45716 4096
rect 46278 4076 46368 4096
rect 32899 4012 32908 4052
rect 32948 4012 33148 4052
rect 33188 4012 33197 4052
rect 34531 4012 34540 4052
rect 34580 4012 35444 4052
rect 35539 4012 35548 4052
rect 35588 4012 38324 4052
rect 39091 4012 39100 4052
rect 39140 4012 40724 4052
rect 40841 4012 40972 4052
rect 41012 4012 41021 4052
rect 43180 4012 44660 4052
rect 44755 4012 44764 4052
rect 44804 4012 45716 4052
rect 34435 3928 34444 3968
rect 34484 3928 35644 3968
rect 35684 3928 35693 3968
rect 35779 3928 35788 3968
rect 35828 3928 36028 3968
rect 36068 3928 36077 3968
rect 39955 3928 39964 3968
rect 40004 3928 41644 3968
rect 41684 3928 41693 3968
rect 43180 3884 43220 4012
rect 44371 3928 44380 3968
rect 44420 3928 44564 3968
rect 35107 3844 35116 3884
rect 35156 3844 43220 3884
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 32899 3676 32908 3716
rect 32948 3676 34540 3716
rect 34580 3676 40492 3716
rect 40532 3676 40541 3716
rect 1468 3592 2900 3632
rect 3017 3592 3100 3632
rect 3140 3592 3148 3632
rect 3188 3592 3197 3632
rect 4204 3592 5300 3632
rect 5356 3592 7276 3632
rect 7316 3592 7325 3632
rect 8467 3592 8476 3632
rect 8516 3592 8620 3632
rect 8660 3592 8669 3632
rect 9065 3592 9148 3632
rect 9188 3592 9196 3632
rect 9236 3592 9245 3632
rect 9523 3592 9532 3632
rect 9572 3592 15092 3632
rect 16579 3592 16588 3632
rect 16628 3592 18892 3632
rect 18932 3592 18941 3632
rect 19171 3592 19180 3632
rect 19220 3592 19564 3632
rect 19604 3592 19613 3632
rect 19891 3592 19900 3632
rect 19940 3592 21332 3632
rect 23923 3592 23932 3632
rect 23972 3592 26572 3632
rect 26612 3592 26621 3632
rect 26947 3592 26956 3632
rect 26996 3592 28204 3632
rect 28244 3592 31992 3632
rect 32131 3592 32140 3632
rect 32180 3592 32852 3632
rect 33571 3592 33580 3632
rect 33620 3592 33772 3632
rect 33812 3592 33821 3632
rect 33868 3592 35836 3632
rect 35876 3592 35885 3632
rect 36547 3592 36556 3632
rect 36596 3592 36604 3632
rect 36644 3592 36727 3632
rect 37411 3592 37420 3632
rect 37460 3592 39052 3632
rect 39092 3592 39101 3632
rect 41059 3592 41068 3632
rect 41108 3592 43220 3632
rect 1123 3508 1132 3548
rect 1172 3508 2420 3548
rect 0 3464 90 3484
rect 2380 3464 2420 3508
rect 4204 3464 4244 3592
rect 5356 3464 5396 3592
rect 33868 3548 33908 3592
rect 5932 3508 6316 3548
rect 6356 3508 6365 3548
rect 7363 3508 7372 3548
rect 7412 3508 8180 3548
rect 5932 3464 5972 3508
rect 8140 3464 8180 3508
rect 8716 3508 14668 3548
rect 14708 3508 14717 3548
rect 15283 3508 15292 3548
rect 15332 3508 18220 3548
rect 18260 3508 18269 3548
rect 18355 3508 18364 3548
rect 18404 3508 19364 3548
rect 8716 3464 8756 3508
rect 19324 3464 19364 3508
rect 19660 3508 20236 3548
rect 20276 3508 20285 3548
rect 20332 3508 24364 3548
rect 24404 3508 24413 3548
rect 24547 3508 24556 3548
rect 24596 3508 26956 3548
rect 26996 3508 27005 3548
rect 30115 3508 30124 3548
rect 30164 3508 32084 3548
rect 19660 3464 19700 3508
rect 0 3424 1228 3464
rect 1268 3424 1277 3464
rect 1411 3424 1420 3464
rect 1460 3424 1468 3464
rect 1508 3424 1591 3464
rect 1642 3424 1651 3464
rect 1691 3424 1748 3464
rect 1865 3424 1996 3464
rect 2036 3424 2045 3464
rect 2371 3424 2380 3464
rect 2420 3424 2429 3464
rect 2825 3424 2860 3464
rect 2900 3424 2956 3464
rect 2996 3424 4204 3464
rect 4244 3424 4253 3464
rect 5194 3455 5396 3464
rect 0 3404 90 3424
rect 0 3128 90 3148
rect 1708 3128 1748 3424
rect 5194 3415 5203 3455
rect 5243 3424 5396 3455
rect 5674 3455 5972 3464
rect 5243 3415 5252 3424
rect 5194 3414 5252 3415
rect 5674 3415 5683 3455
rect 5723 3424 5972 3455
rect 6017 3424 6220 3464
rect 6260 3424 6269 3464
rect 7075 3424 7084 3464
rect 7124 3424 7133 3464
rect 7180 3424 7468 3464
rect 7508 3424 7517 3464
rect 8131 3424 8140 3464
rect 8180 3424 8189 3464
rect 8707 3424 8716 3464
rect 8756 3424 8765 3464
rect 8899 3424 8908 3464
rect 8948 3424 8957 3464
rect 9283 3424 9292 3464
rect 9332 3424 9341 3464
rect 10723 3424 10732 3464
rect 10772 3424 10828 3464
rect 10868 3424 10903 3464
rect 11011 3424 11020 3464
rect 11060 3424 11348 3464
rect 5723 3415 5732 3424
rect 5674 3414 5732 3415
rect 4492 3380 4532 3389
rect 6017 3380 6057 3424
rect 6604 3380 6644 3389
rect 3043 3340 3052 3380
rect 3092 3340 3244 3380
rect 3284 3340 3293 3380
rect 4291 3340 4300 3380
rect 4340 3340 4492 3380
rect 5059 3340 5068 3380
rect 5108 3340 5117 3380
rect 5296 3340 5305 3380
rect 5345 3340 5548 3380
rect 5588 3340 5597 3380
rect 5776 3340 5785 3380
rect 5825 3340 6057 3380
rect 6106 3340 6115 3380
rect 6155 3340 6316 3380
rect 6356 3340 6365 3380
rect 6644 3340 6796 3380
rect 6836 3340 6845 3380
rect 4492 3331 4532 3340
rect 5068 3296 5108 3340
rect 6604 3331 6644 3340
rect 1843 3256 1852 3296
rect 1892 3256 2092 3296
rect 2132 3256 2141 3296
rect 2611 3256 2620 3296
rect 2660 3256 4396 3296
rect 4436 3256 4445 3296
rect 4675 3256 4684 3296
rect 4724 3256 5108 3296
rect 5443 3256 5452 3296
rect 5492 3256 5740 3296
rect 5780 3256 5789 3296
rect 5836 3256 6124 3296
rect 6164 3256 6173 3296
rect 5068 3212 5108 3256
rect 5836 3212 5876 3256
rect 7084 3212 7124 3424
rect 7180 3380 7220 3424
rect 8140 3380 8180 3424
rect 7171 3340 7180 3380
rect 7220 3340 7351 3380
rect 7433 3340 7564 3380
rect 7604 3340 7613 3380
rect 7673 3340 7682 3380
rect 7722 3340 7852 3380
rect 7892 3340 7901 3380
rect 8140 3340 8812 3380
rect 8852 3340 8861 3380
rect 8371 3256 8380 3296
rect 8420 3256 8620 3296
rect 8660 3256 8669 3296
rect 2227 3172 2236 3212
rect 2276 3172 2572 3212
rect 2612 3172 2621 3212
rect 4963 3172 4972 3212
rect 5012 3172 5021 3212
rect 5068 3172 5876 3212
rect 5923 3172 5932 3212
rect 5972 3172 6508 3212
rect 6548 3172 6557 3212
rect 7084 3172 8812 3212
rect 8852 3172 8861 3212
rect 0 3088 1748 3128
rect 4972 3128 5012 3172
rect 4972 3088 6796 3128
rect 6836 3088 6845 3128
rect 0 3068 90 3088
rect 8908 3044 8948 3424
rect 9292 3128 9332 3424
rect 10348 3380 10388 3389
rect 11308 3380 11348 3424
rect 11788 3424 12020 3464
rect 12067 3424 12076 3464
rect 12116 3424 12268 3464
rect 12308 3424 12317 3464
rect 13769 3424 13900 3464
rect 13940 3424 13949 3464
rect 14275 3424 14284 3464
rect 14324 3424 14476 3464
rect 14516 3424 14525 3464
rect 14659 3424 14668 3464
rect 14708 3424 14764 3464
rect 14804 3424 14839 3464
rect 14921 3424 15052 3464
rect 15092 3424 15101 3464
rect 16099 3424 16108 3464
rect 16148 3424 16724 3464
rect 17225 3424 17356 3464
rect 17396 3424 17405 3464
rect 17801 3424 17932 3464
rect 17972 3424 17981 3464
rect 18115 3424 18124 3464
rect 18164 3424 18173 3464
rect 18377 3424 18508 3464
rect 18548 3424 18557 3464
rect 18761 3424 18892 3464
rect 18932 3424 18941 3464
rect 19306 3424 19315 3464
rect 19355 3424 19364 3464
rect 19651 3424 19660 3464
rect 19700 3424 19709 3464
rect 20035 3424 20044 3464
rect 20084 3424 20140 3464
rect 20180 3424 20244 3464
rect 11788 3380 11828 3424
rect 9850 3340 9859 3380
rect 9899 3340 10252 3380
rect 10292 3340 10301 3380
rect 10388 3340 10636 3380
rect 10676 3340 10685 3380
rect 10793 3340 10828 3380
rect 10868 3340 10924 3380
rect 10964 3340 10973 3380
rect 11299 3340 11308 3380
rect 11348 3340 11357 3380
rect 11417 3340 11426 3380
rect 11466 3340 11500 3380
rect 11540 3340 11606 3380
rect 11770 3340 11779 3380
rect 11819 3340 11828 3380
rect 11875 3340 11884 3380
rect 11924 3340 11933 3380
rect 10348 3296 10388 3340
rect 9545 3256 9667 3296
rect 9716 3256 9725 3296
rect 9772 3256 10388 3296
rect 11308 3296 11348 3340
rect 11308 3256 11684 3296
rect 9772 3212 9812 3256
rect 11644 3212 11684 3256
rect 11884 3212 11924 3340
rect 11980 3296 12020 3424
rect 12844 3380 12884 3389
rect 16684 3380 16724 3424
rect 18124 3380 18164 3424
rect 20332 3380 20372 3508
rect 32044 3464 32084 3508
rect 33196 3508 33908 3548
rect 35107 3508 35116 3548
rect 35156 3508 37132 3548
rect 37172 3508 37181 3548
rect 41443 3508 41452 3548
rect 41492 3508 41876 3548
rect 33196 3464 33236 3508
rect 41836 3464 41876 3508
rect 43180 3464 43220 3592
rect 44524 3548 44564 3928
rect 46278 3800 46368 3820
rect 45148 3760 46368 3800
rect 45148 3632 45188 3760
rect 46278 3740 46368 3760
rect 45139 3592 45148 3632
rect 45188 3592 45197 3632
rect 44524 3508 45428 3548
rect 45388 3464 45428 3508
rect 46278 3464 46368 3484
rect 23561 3424 23692 3464
rect 23732 3424 23741 3464
rect 24547 3424 24556 3464
rect 24596 3424 24748 3464
rect 24788 3424 24797 3464
rect 26537 3424 26668 3464
rect 26708 3424 26717 3464
rect 27235 3424 27244 3464
rect 27284 3424 28780 3464
rect 28820 3424 28829 3464
rect 29155 3424 29164 3464
rect 29204 3424 30316 3464
rect 30356 3424 30487 3464
rect 32044 3424 33236 3464
rect 34293 3424 34540 3464
rect 34580 3424 34589 3464
rect 35587 3424 35596 3464
rect 35636 3424 35645 3464
rect 35945 3424 36076 3464
rect 36116 3424 36125 3464
rect 36259 3424 36268 3464
rect 36308 3424 36460 3464
rect 36500 3424 36509 3464
rect 36835 3424 36844 3464
rect 36884 3424 36893 3464
rect 40291 3424 40300 3464
rect 40340 3424 41596 3464
rect 41636 3424 41645 3464
rect 41827 3424 41836 3464
rect 41876 3424 41885 3464
rect 43180 3424 44524 3464
rect 44564 3424 44573 3464
rect 44899 3424 44908 3464
rect 44948 3424 44957 3464
rect 45388 3424 46368 3464
rect 21676 3380 21716 3389
rect 23308 3380 23348 3389
rect 26092 3380 26132 3389
rect 27148 3380 27188 3389
rect 30316 3380 30356 3424
rect 31948 3380 31988 3389
rect 33580 3380 33620 3389
rect 34293 3380 34333 3424
rect 12355 3340 12364 3380
rect 12404 3340 12556 3380
rect 12596 3340 12605 3380
rect 12713 3340 12844 3380
rect 12884 3340 12893 3380
rect 13354 3340 13363 3380
rect 13403 3340 13708 3380
rect 13748 3340 13757 3380
rect 14188 3340 15436 3380
rect 15476 3340 16588 3380
rect 16628 3340 16637 3380
rect 16724 3340 17836 3380
rect 17876 3340 17885 3380
rect 18124 3340 18988 3380
rect 19028 3340 19037 3380
rect 19708 3340 20372 3380
rect 20419 3340 20428 3380
rect 20468 3340 20524 3380
rect 20564 3340 20599 3380
rect 21929 3340 21964 3380
rect 22004 3340 22060 3380
rect 22100 3340 22109 3380
rect 23177 3340 23212 3380
rect 23252 3340 23308 3380
rect 24835 3340 24844 3380
rect 24884 3340 25015 3380
rect 25603 3340 25612 3380
rect 25652 3340 26092 3380
rect 27043 3340 27052 3380
rect 27092 3340 27148 3380
rect 27188 3340 27223 3380
rect 28195 3340 28204 3380
rect 28244 3340 28396 3380
rect 28436 3340 28780 3380
rect 28820 3340 28829 3380
rect 29059 3340 29068 3380
rect 29108 3340 29260 3380
rect 29300 3340 29309 3380
rect 30569 3340 30700 3380
rect 30740 3340 30749 3380
rect 32201 3340 32332 3380
rect 32372 3340 32381 3380
rect 34275 3340 34284 3380
rect 34324 3340 34333 3380
rect 35500 3380 35540 3389
rect 35596 3380 35636 3424
rect 36844 3380 36884 3424
rect 35540 3340 35636 3380
rect 35683 3340 35692 3380
rect 35732 3340 36884 3380
rect 37324 3380 37364 3389
rect 39244 3380 39284 3389
rect 44908 3380 44948 3424
rect 46278 3404 46368 3424
rect 37891 3340 37900 3380
rect 37940 3340 38572 3380
rect 38612 3340 38621 3380
rect 38947 3340 38956 3380
rect 38996 3340 39244 3380
rect 39284 3340 39293 3380
rect 40361 3340 40492 3380
rect 40532 3340 40541 3380
rect 40649 3340 40780 3380
rect 40820 3340 40829 3380
rect 40963 3340 40972 3380
rect 41012 3340 41059 3380
rect 41099 3340 41143 3380
rect 41731 3340 41740 3380
rect 41780 3340 44948 3380
rect 12844 3331 12884 3340
rect 14188 3296 14228 3340
rect 16684 3331 16724 3340
rect 19708 3296 19748 3340
rect 21676 3296 21716 3340
rect 23212 3296 23252 3340
rect 23308 3331 23348 3340
rect 26092 3331 26132 3340
rect 27148 3331 27188 3340
rect 30316 3331 30356 3340
rect 31948 3296 31988 3340
rect 11980 3256 12076 3296
rect 12116 3256 12125 3296
rect 13276 3256 14228 3296
rect 14467 3256 14476 3296
rect 14516 3256 16645 3296
rect 17587 3256 17596 3296
rect 17636 3256 19748 3296
rect 19939 3256 19948 3296
rect 19988 3256 21484 3296
rect 21524 3256 21533 3296
rect 21676 3256 22828 3296
rect 22868 3256 23252 3296
rect 23491 3256 23500 3296
rect 23540 3256 24460 3296
rect 24500 3256 24509 3296
rect 30892 3256 31988 3296
rect 33580 3296 33620 3340
rect 35500 3296 35540 3340
rect 37324 3296 37364 3340
rect 39244 3331 39284 3340
rect 33580 3256 36268 3296
rect 36308 3256 36317 3296
rect 36451 3256 36460 3296
rect 36500 3256 36940 3296
rect 36980 3256 37364 3296
rect 39907 3256 39916 3296
rect 39956 3256 41164 3296
rect 41204 3256 41213 3296
rect 13276 3212 13316 3256
rect 9379 3172 9388 3212
rect 9428 3172 9812 3212
rect 9955 3172 9964 3212
rect 10004 3172 11540 3212
rect 11644 3172 11924 3212
rect 12845 3172 13316 3212
rect 13385 3172 13516 3212
rect 13556 3172 13565 3212
rect 13891 3172 13900 3212
rect 13940 3172 14140 3212
rect 14180 3172 14189 3212
rect 14441 3172 14524 3212
rect 14564 3172 14572 3212
rect 14612 3172 14621 3212
rect 14899 3172 14908 3212
rect 14948 3172 16532 3212
rect 11500 3128 11540 3172
rect 12845 3128 12885 3172
rect 9292 3088 11308 3128
rect 11348 3088 11357 3128
rect 11500 3088 12885 3128
rect 12940 3088 14860 3128
rect 14900 3088 14909 3128
rect 12940 3044 12980 3088
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 7660 3004 7756 3044
rect 7796 3004 7805 3044
rect 8908 3004 12980 3044
rect 16492 3044 16532 3172
rect 16605 3128 16645 3256
rect 16867 3172 16876 3212
rect 16916 3172 17164 3212
rect 17204 3172 17213 3212
rect 17539 3172 17548 3212
rect 17588 3172 17692 3212
rect 17732 3172 17741 3212
rect 17827 3172 17836 3212
rect 17876 3172 18508 3212
rect 18548 3172 18557 3212
rect 18739 3172 18748 3212
rect 18788 3172 18796 3212
rect 18836 3172 18919 3212
rect 19123 3172 19132 3212
rect 19172 3172 19181 3212
rect 19507 3172 19516 3212
rect 19556 3172 20180 3212
rect 20275 3172 20284 3212
rect 20324 3172 21620 3212
rect 21737 3172 21868 3212
rect 21908 3172 21917 3212
rect 22147 3172 22156 3212
rect 22196 3172 23060 3212
rect 24185 3172 24268 3212
rect 24308 3172 24316 3212
rect 24356 3172 24365 3212
rect 25699 3172 25708 3212
rect 25748 3172 26036 3212
rect 26153 3172 26284 3212
rect 26324 3172 26333 3212
rect 26419 3172 26428 3212
rect 26468 3172 26476 3212
rect 26516 3172 26599 3212
rect 27427 3172 27436 3212
rect 27476 3172 28540 3212
rect 28580 3172 28589 3212
rect 30377 3172 30508 3212
rect 30548 3172 30557 3212
rect 19132 3128 19172 3172
rect 20140 3128 20180 3172
rect 21580 3128 21620 3172
rect 23020 3128 23060 3172
rect 25996 3128 26036 3172
rect 30892 3128 30932 3256
rect 30979 3172 30988 3212
rect 31028 3172 34348 3212
rect 34388 3172 34397 3212
rect 34540 3172 35116 3212
rect 35156 3172 35165 3212
rect 35683 3172 35692 3212
rect 35732 3172 35884 3212
rect 35924 3172 35933 3212
rect 35980 3172 36220 3212
rect 36260 3172 36269 3212
rect 44755 3172 44764 3212
rect 44804 3172 44813 3212
rect 34540 3128 34580 3172
rect 35980 3128 36020 3172
rect 16605 3088 18700 3128
rect 18740 3088 18749 3128
rect 19132 3088 19364 3128
rect 20140 3088 21524 3128
rect 21580 3088 22540 3128
rect 22580 3088 22589 3128
rect 23020 3088 25900 3128
rect 25940 3088 25949 3128
rect 25996 3088 30932 3128
rect 31267 3088 31276 3128
rect 31316 3088 34580 3128
rect 34636 3088 36020 3128
rect 44764 3128 44804 3172
rect 46278 3128 46368 3148
rect 44764 3088 46368 3128
rect 19324 3044 19364 3088
rect 21484 3044 21524 3088
rect 34636 3044 34676 3088
rect 46278 3068 46368 3088
rect 16492 3004 18412 3044
rect 18452 3004 18461 3044
rect 19324 3004 19756 3044
rect 19796 3004 19805 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 21484 3004 22156 3044
rect 22196 3004 22205 3044
rect 24355 3004 24364 3044
rect 24404 3004 29356 3044
rect 29396 3004 30836 3044
rect 30883 3004 30892 3044
rect 30932 3004 34676 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 35587 3004 35596 3044
rect 35636 3004 35884 3044
rect 35924 3004 35933 3044
rect 7660 2960 7700 3004
rect 30796 2960 30836 3004
rect 2659 2920 2668 2960
rect 2708 2920 5452 2960
rect 5492 2920 5501 2960
rect 5923 2920 5932 2960
rect 5972 2920 7700 2960
rect 9964 2920 10772 2960
rect 11683 2920 11692 2960
rect 11732 2920 16492 2960
rect 16532 2920 16541 2960
rect 17260 2920 17548 2960
rect 17588 2920 18604 2960
rect 18644 2920 18836 2960
rect 18883 2920 18892 2960
rect 18932 2920 21964 2960
rect 22004 2920 22013 2960
rect 23020 2920 26476 2960
rect 26516 2920 26525 2960
rect 29251 2920 29260 2960
rect 29300 2920 30028 2960
rect 30068 2920 30077 2960
rect 30796 2920 31660 2960
rect 31700 2920 31709 2960
rect 31852 2920 33004 2960
rect 33044 2920 33053 2960
rect 34915 2920 34924 2960
rect 34964 2920 35692 2960
rect 35732 2920 35741 2960
rect 37420 2920 38668 2960
rect 38708 2920 38717 2960
rect 2249 2836 2332 2876
rect 2372 2836 2380 2876
rect 2420 2836 2429 2876
rect 2707 2836 2716 2876
rect 2756 2836 2900 2876
rect 0 2792 90 2812
rect 2860 2792 2900 2836
rect 0 2752 1996 2792
rect 2036 2752 2045 2792
rect 2851 2752 2860 2792
rect 2900 2752 2909 2792
rect 0 2732 90 2752
rect 1852 2668 2276 2708
rect 1852 2624 1892 2668
rect 1219 2584 1228 2624
rect 1268 2584 1277 2624
rect 1603 2584 1612 2624
rect 1652 2584 1661 2624
rect 1843 2584 1852 2624
rect 1892 2584 1901 2624
rect 2083 2584 2092 2624
rect 2132 2584 2141 2624
rect 0 2456 90 2476
rect 1228 2456 1268 2584
rect 1385 2500 1468 2540
rect 1508 2500 1516 2540
rect 1556 2500 1565 2540
rect 0 2416 1268 2456
rect 0 2396 90 2416
rect 1612 2204 1652 2584
rect 2092 2456 2132 2584
rect 2236 2540 2276 2668
rect 2956 2624 2996 2920
rect 9964 2876 10004 2920
rect 10732 2876 10772 2920
rect 17260 2876 17300 2920
rect 3427 2836 3436 2876
rect 3476 2836 3484 2876
rect 3524 2836 3607 2876
rect 4195 2836 4204 2876
rect 4244 2836 4253 2876
rect 5932 2836 6220 2876
rect 6260 2836 6269 2876
rect 6569 2836 6691 2876
rect 6740 2836 6749 2876
rect 7171 2836 7180 2876
rect 7220 2836 7229 2876
rect 8716 2836 10004 2876
rect 10243 2836 10252 2876
rect 10292 2836 10636 2876
rect 10676 2836 10685 2876
rect 10732 2836 12652 2876
rect 12692 2836 12701 2876
rect 13577 2836 13708 2876
rect 13748 2836 13757 2876
rect 15427 2836 15436 2876
rect 15476 2836 16148 2876
rect 4204 2792 4244 2836
rect 3331 2752 3340 2792
rect 3380 2752 4108 2792
rect 4148 2752 4157 2792
rect 4204 2752 4820 2792
rect 4780 2708 4820 2752
rect 5932 2708 5972 2836
rect 7180 2792 7220 2836
rect 8716 2792 8756 2836
rect 6659 2752 7220 2792
rect 7267 2752 7276 2792
rect 7316 2752 8756 2792
rect 8803 2752 8812 2792
rect 8852 2752 9484 2792
rect 9524 2752 9533 2792
rect 10435 2752 10444 2792
rect 10484 2752 11500 2792
rect 11540 2752 11549 2792
rect 12076 2752 12404 2792
rect 12547 2752 12556 2792
rect 12596 2752 13420 2792
rect 13460 2752 13469 2792
rect 13516 2752 14284 2792
rect 14324 2752 14333 2792
rect 15331 2752 15340 2792
rect 15380 2752 16052 2792
rect 6659 2708 6699 2752
rect 3427 2668 3436 2708
rect 3476 2668 4724 2708
rect 4771 2668 4780 2708
rect 4820 2668 4972 2708
rect 5012 2668 5021 2708
rect 5443 2668 5452 2708
rect 5492 2699 6068 2708
rect 5492 2668 6028 2699
rect 4684 2624 4724 2668
rect 6115 2668 6124 2708
rect 6164 2668 6359 2708
rect 6399 2668 6408 2708
rect 6595 2668 6604 2708
rect 6644 2668 6699 2708
rect 6761 2668 6796 2708
rect 6836 2668 6892 2708
rect 6932 2668 6941 2708
rect 7025 2668 7034 2708
rect 7074 2668 7084 2708
rect 7124 2668 7214 2708
rect 7363 2668 7372 2708
rect 7412 2668 7543 2708
rect 8620 2699 8660 2708
rect 6028 2650 6068 2659
rect 8873 2668 9004 2708
rect 9044 2668 9053 2708
rect 10060 2699 10868 2708
rect 10060 2668 10252 2699
rect 8620 2624 8660 2659
rect 10060 2624 10100 2668
rect 10292 2668 10828 2699
rect 10252 2650 10292 2659
rect 10915 2668 10924 2708
rect 10964 2668 12036 2708
rect 12076 2668 12116 2752
rect 12158 2668 12256 2708
rect 12296 2687 12308 2708
rect 2345 2584 2476 2624
rect 2516 2584 2525 2624
rect 2851 2584 2860 2624
rect 2900 2584 2996 2624
rect 3113 2584 3244 2624
rect 3284 2584 3293 2624
rect 3619 2584 3628 2624
rect 3668 2584 3677 2624
rect 4003 2584 4012 2624
rect 4052 2584 4204 2624
rect 4244 2584 4253 2624
rect 4387 2584 4396 2624
rect 4436 2584 4567 2624
rect 4684 2584 5972 2624
rect 6377 2584 6499 2624
rect 6548 2584 6557 2624
rect 6691 2584 6700 2624
rect 6740 2584 9676 2624
rect 9716 2584 10100 2624
rect 10828 2624 10868 2659
rect 12259 2647 12268 2668
rect 12308 2647 12317 2687
rect 12364 2624 12404 2752
rect 13516 2708 13556 2752
rect 12739 2668 12748 2708
rect 12788 2699 13556 2708
rect 12788 2668 13516 2699
rect 13891 2668 13900 2708
rect 13940 2668 13949 2708
rect 15017 2668 15148 2708
rect 15188 2668 15197 2708
rect 15610 2668 15619 2708
rect 15659 2668 15668 2708
rect 15715 2668 15724 2708
rect 15764 2668 15820 2708
rect 15860 2668 15895 2708
rect 13516 2650 13556 2659
rect 10828 2584 11884 2624
rect 11924 2584 11933 2624
rect 12364 2584 12980 2624
rect 2236 2500 2956 2540
rect 2996 2500 3005 2540
rect 2092 2416 2900 2456
rect 3091 2416 3100 2456
rect 3140 2416 3148 2456
rect 3188 2416 3271 2456
rect 2860 2372 2900 2416
rect 3628 2372 3668 2584
rect 3859 2500 3868 2540
rect 3908 2500 5644 2540
rect 5684 2500 5693 2540
rect 5932 2456 5972 2584
rect 12940 2540 12980 2584
rect 13900 2540 13940 2668
rect 15148 2650 15188 2659
rect 15628 2540 15668 2668
rect 6019 2500 6028 2540
rect 6068 2500 6220 2540
rect 6260 2500 7852 2540
rect 7892 2500 7901 2540
rect 8131 2500 8140 2540
rect 8180 2500 12556 2540
rect 12596 2500 12605 2540
rect 12940 2500 13804 2540
rect 13844 2500 13940 2540
rect 15139 2500 15148 2540
rect 15188 2500 15668 2540
rect 16012 2540 16052 2752
rect 16108 2708 16148 2836
rect 16204 2836 17300 2876
rect 17347 2836 17356 2876
rect 17396 2836 17836 2876
rect 17876 2836 17885 2876
rect 16099 2668 16108 2708
rect 16148 2668 16157 2708
rect 16204 2624 16244 2836
rect 18796 2792 18836 2920
rect 23020 2876 23060 2920
rect 31852 2876 31892 2920
rect 37420 2876 37460 2920
rect 18979 2836 18988 2876
rect 19028 2836 20140 2876
rect 20180 2836 20189 2876
rect 21484 2836 21868 2876
rect 21908 2836 21917 2876
rect 22723 2836 22732 2876
rect 22772 2836 23060 2876
rect 23203 2836 23212 2876
rect 23252 2836 23692 2876
rect 23732 2836 23741 2876
rect 25795 2836 25804 2876
rect 25844 2836 26668 2876
rect 26708 2836 26717 2876
rect 26764 2836 29644 2876
rect 29684 2836 29693 2876
rect 29827 2836 29836 2876
rect 29876 2836 31892 2876
rect 31939 2836 31948 2876
rect 31988 2836 33964 2876
rect 34004 2836 34013 2876
rect 34339 2836 34348 2876
rect 34388 2836 34676 2876
rect 35779 2836 35788 2876
rect 35828 2836 37460 2876
rect 37507 2836 37516 2876
rect 37556 2836 38044 2876
rect 38084 2836 38093 2876
rect 39523 2836 39532 2876
rect 39572 2836 40252 2876
rect 40292 2836 40301 2876
rect 40915 2836 40924 2876
rect 40964 2836 41740 2876
rect 41780 2836 41789 2876
rect 16684 2752 17452 2792
rect 17492 2752 17501 2792
rect 17548 2752 17788 2792
rect 17828 2752 17837 2792
rect 18220 2752 18316 2792
rect 18356 2752 18365 2792
rect 18499 2752 18508 2792
rect 18548 2752 18644 2792
rect 18796 2752 19508 2792
rect 16684 2699 16724 2752
rect 17548 2708 17588 2752
rect 18220 2708 18260 2752
rect 17033 2668 17164 2708
rect 17204 2668 17213 2708
rect 17347 2668 17356 2708
rect 17396 2668 17588 2708
rect 17635 2668 17644 2708
rect 17684 2668 17693 2708
rect 17827 2668 17836 2708
rect 17876 2668 18260 2708
rect 18365 2668 18403 2708
rect 18443 2668 18452 2708
rect 18499 2668 18508 2708
rect 18548 2668 18557 2708
rect 16684 2650 16724 2659
rect 17164 2650 17204 2659
rect 17644 2624 17684 2668
rect 18412 2624 18452 2668
rect 16195 2584 16204 2624
rect 16244 2584 16253 2624
rect 17417 2584 17548 2624
rect 17588 2584 17597 2624
rect 17644 2584 17932 2624
rect 17972 2584 17981 2624
rect 18403 2584 18412 2624
rect 18452 2584 18461 2624
rect 18508 2540 18548 2668
rect 18604 2624 18644 2752
rect 18883 2668 18892 2708
rect 18932 2668 19180 2708
rect 19220 2668 19229 2708
rect 19468 2699 19508 2752
rect 21484 2708 21524 2836
rect 22435 2752 22444 2792
rect 22484 2752 26420 2792
rect 26380 2708 26420 2752
rect 19468 2650 19508 2659
rect 19948 2699 20236 2708
rect 19988 2668 20236 2699
rect 20276 2668 20285 2708
rect 20620 2668 21100 2708
rect 21140 2668 21149 2708
rect 21466 2668 21475 2708
rect 21515 2668 21524 2708
rect 21571 2668 21580 2708
rect 21620 2668 21676 2708
rect 21716 2668 21751 2708
rect 21833 2668 21964 2708
rect 22004 2668 22013 2708
rect 22540 2699 22924 2708
rect 19948 2650 19988 2659
rect 20620 2624 20660 2668
rect 22580 2668 22924 2699
rect 22964 2668 22973 2708
rect 23020 2699 23060 2708
rect 22540 2650 22580 2659
rect 23107 2668 23116 2708
rect 23156 2668 24067 2708
rect 24107 2668 24116 2708
rect 24163 2668 24172 2708
rect 24212 2668 24221 2708
rect 24425 2668 24556 2708
rect 24596 2668 24605 2708
rect 24835 2668 24844 2708
rect 24884 2699 25324 2708
rect 24884 2668 25132 2699
rect 23020 2624 23060 2659
rect 18604 2584 18988 2624
rect 19028 2584 19276 2624
rect 19316 2584 19325 2624
rect 20611 2584 20620 2624
rect 20660 2584 20669 2624
rect 20716 2584 21004 2624
rect 21044 2584 21053 2624
rect 21283 2584 21292 2624
rect 21332 2584 22060 2624
rect 22100 2584 22109 2624
rect 23020 2584 23156 2624
rect 23299 2584 23308 2624
rect 23348 2584 23596 2624
rect 23636 2584 23645 2624
rect 20716 2540 20756 2584
rect 23116 2540 23156 2584
rect 24172 2540 24212 2668
rect 25172 2668 25324 2699
rect 25364 2668 25373 2708
rect 25481 2668 25612 2708
rect 25652 2668 25661 2708
rect 25891 2668 25900 2708
rect 25940 2668 26324 2708
rect 26371 2668 26380 2708
rect 26420 2668 26429 2708
rect 25132 2650 25172 2659
rect 25612 2650 25652 2659
rect 26284 2624 26324 2668
rect 26764 2624 26804 2836
rect 27811 2752 27820 2792
rect 27860 2752 28148 2792
rect 28108 2708 28148 2752
rect 28204 2708 28244 2836
rect 34636 2792 34676 2836
rect 46278 2792 46368 2812
rect 28579 2752 28588 2792
rect 28628 2752 29780 2792
rect 27497 2668 27628 2708
rect 27668 2668 27677 2708
rect 28090 2668 28099 2708
rect 28139 2668 28148 2708
rect 28195 2668 28204 2708
rect 28244 2668 28253 2708
rect 28387 2668 28396 2708
rect 28436 2668 28588 2708
rect 28628 2668 28637 2708
rect 29033 2668 29164 2708
rect 29204 2668 29213 2708
rect 29347 2668 29356 2708
rect 29396 2699 29684 2708
rect 29396 2668 29644 2699
rect 27628 2650 27668 2659
rect 29164 2650 29204 2659
rect 29644 2650 29684 2659
rect 29740 2624 29780 2752
rect 30220 2752 30508 2792
rect 30548 2752 30557 2792
rect 30604 2752 31084 2792
rect 31124 2752 31133 2792
rect 31180 2752 31660 2792
rect 31700 2752 32428 2792
rect 32468 2752 32477 2792
rect 32611 2752 32620 2792
rect 32660 2752 34196 2792
rect 34636 2752 36460 2792
rect 36500 2752 36509 2792
rect 37795 2752 37804 2792
rect 37844 2752 40052 2792
rect 40099 2752 40108 2792
rect 40148 2752 40780 2792
rect 40820 2752 40829 2792
rect 45139 2752 45148 2792
rect 45188 2752 46368 2792
rect 30220 2708 30260 2752
rect 30604 2708 30644 2752
rect 31180 2708 31220 2752
rect 34156 2708 34196 2752
rect 40012 2708 40052 2752
rect 46278 2732 46368 2752
rect 30202 2668 30211 2708
rect 30251 2668 30260 2708
rect 30307 2668 30316 2708
rect 30356 2668 30644 2708
rect 30691 2668 30700 2708
rect 30740 2668 30871 2708
rect 31084 2668 31220 2708
rect 31756 2699 32044 2708
rect 31084 2624 31124 2668
rect 31267 2626 31276 2666
rect 31316 2626 31447 2666
rect 31796 2668 32044 2699
rect 32084 2668 32093 2708
rect 32323 2668 32332 2708
rect 32372 2668 32908 2708
rect 32948 2668 32957 2708
rect 33579 2668 33588 2708
rect 33628 2668 33868 2708
rect 33908 2668 33917 2708
rect 34042 2668 34051 2708
rect 34091 2668 34100 2708
rect 34147 2668 34156 2708
rect 34196 2668 34327 2708
rect 34531 2668 34540 2708
rect 34580 2668 34732 2708
rect 34772 2668 34781 2708
rect 34985 2668 35116 2708
rect 35156 2668 35165 2708
rect 35465 2668 35596 2708
rect 35636 2668 35645 2708
rect 36259 2668 36268 2708
rect 36308 2699 36692 2708
rect 36308 2668 36652 2699
rect 31756 2650 31796 2659
rect 34060 2624 34100 2668
rect 35116 2650 35156 2659
rect 35596 2650 35636 2659
rect 37769 2668 37900 2708
rect 37940 2668 37949 2708
rect 38537 2668 38668 2708
rect 38708 2668 38717 2708
rect 38947 2668 38956 2708
rect 38996 2699 39956 2708
rect 38996 2668 39916 2699
rect 36652 2650 36692 2659
rect 40012 2668 44948 2708
rect 39916 2650 39956 2659
rect 44908 2624 44948 2668
rect 24643 2584 24652 2624
rect 24692 2584 24748 2624
rect 24788 2584 24823 2624
rect 26179 2584 26188 2624
rect 26228 2584 26237 2624
rect 26284 2584 26804 2624
rect 28579 2584 28588 2624
rect 28628 2584 28684 2624
rect 28724 2584 28759 2624
rect 29740 2584 30508 2624
rect 30548 2584 30557 2624
rect 30787 2584 30796 2624
rect 30836 2584 31124 2624
rect 33580 2584 33964 2624
rect 34004 2584 34013 2624
rect 34060 2584 34348 2624
rect 34388 2584 34397 2624
rect 34531 2584 34540 2624
rect 34580 2584 34636 2624
rect 34676 2584 34711 2624
rect 36163 2584 36172 2624
rect 36212 2584 36221 2624
rect 36739 2584 36748 2624
rect 36788 2584 38284 2624
rect 38324 2584 38333 2624
rect 40483 2584 40492 2624
rect 40532 2584 40541 2624
rect 40675 2584 40684 2624
rect 40724 2584 40855 2624
rect 43075 2584 43084 2624
rect 43124 2584 44140 2624
rect 44180 2584 44189 2624
rect 44515 2584 44524 2624
rect 44564 2584 44573 2624
rect 44899 2584 44908 2624
rect 44948 2584 44957 2624
rect 26188 2540 26228 2584
rect 33580 2540 33620 2584
rect 36172 2540 36212 2584
rect 16012 2500 17740 2540
rect 17780 2500 17789 2540
rect 17836 2500 18548 2540
rect 18787 2500 18796 2540
rect 18836 2500 20756 2540
rect 20851 2500 20860 2540
rect 20900 2500 22732 2540
rect 22772 2500 22781 2540
rect 23107 2500 23116 2540
rect 23156 2500 23165 2540
rect 23596 2500 24212 2540
rect 25699 2500 25708 2540
rect 25748 2500 26132 2540
rect 26188 2500 30220 2540
rect 30260 2500 30269 2540
rect 31948 2500 33620 2540
rect 33676 2500 36212 2540
rect 4243 2416 4252 2456
rect 4292 2416 4532 2456
rect 4627 2416 4636 2456
rect 4676 2416 5740 2456
rect 5780 2416 5789 2456
rect 5932 2416 12268 2456
rect 12308 2416 12317 2456
rect 12451 2416 12460 2456
rect 12500 2416 15436 2456
rect 15476 2416 15485 2456
rect 4492 2372 4532 2416
rect 17836 2372 17876 2500
rect 18163 2416 18172 2456
rect 18212 2416 18220 2456
rect 18260 2416 18343 2456
rect 19267 2416 19276 2456
rect 19316 2416 20524 2456
rect 20564 2416 20573 2456
rect 21235 2416 21244 2456
rect 21284 2416 22924 2456
rect 22964 2416 22973 2456
rect 23596 2372 23636 2500
rect 26092 2456 26132 2500
rect 31948 2456 31988 2500
rect 33676 2456 33716 2500
rect 23827 2416 23836 2456
rect 23876 2416 24460 2456
rect 24500 2416 24509 2456
rect 24556 2416 25948 2456
rect 25988 2416 25997 2456
rect 26092 2416 28780 2456
rect 28820 2416 28829 2456
rect 29155 2416 29164 2456
rect 29204 2416 31988 2456
rect 32323 2416 32332 2456
rect 32372 2416 33716 2456
rect 33763 2416 33772 2456
rect 33812 2416 34540 2456
rect 34580 2416 34589 2456
rect 35923 2416 35932 2456
rect 35972 2416 35981 2456
rect 36067 2416 36076 2456
rect 36116 2416 37420 2456
rect 37460 2416 38188 2456
rect 38228 2416 38237 2456
rect 24556 2372 24596 2416
rect 35932 2372 35972 2416
rect 2860 2332 3340 2372
rect 3380 2332 3389 2372
rect 3628 2332 4396 2372
rect 4436 2332 4445 2372
rect 4492 2332 7660 2372
rect 7700 2332 7709 2372
rect 8716 2332 12556 2372
rect 12596 2332 12605 2372
rect 13411 2332 13420 2372
rect 13460 2332 16204 2372
rect 16244 2332 16253 2372
rect 16867 2332 16876 2372
rect 16916 2332 17876 2372
rect 18700 2332 21388 2372
rect 21428 2332 21437 2372
rect 21571 2332 21580 2372
rect 21620 2332 23636 2372
rect 24067 2332 24076 2372
rect 24116 2332 24596 2372
rect 24643 2332 24652 2372
rect 24692 2332 31660 2372
rect 31700 2332 31709 2372
rect 31756 2332 35972 2372
rect 8716 2288 8756 2332
rect 18700 2288 18740 2332
rect 31756 2288 31796 2332
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 4108 2248 8756 2288
rect 8803 2248 8812 2288
rect 8852 2248 12940 2288
rect 12980 2248 12989 2288
rect 13132 2248 14380 2288
rect 14420 2248 14429 2288
rect 17347 2248 17356 2288
rect 17396 2248 18740 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 20899 2248 20908 2288
rect 20948 2248 29684 2288
rect 30019 2248 30028 2288
rect 30068 2248 30220 2288
rect 30260 2248 30269 2288
rect 31267 2248 31276 2288
rect 31316 2248 31796 2288
rect 31948 2248 32908 2288
rect 32948 2248 32957 2288
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 35107 2248 35116 2288
rect 35156 2248 39916 2288
rect 39956 2248 39965 2288
rect 172 2164 1652 2204
rect 1996 2164 3532 2204
rect 3572 2164 3581 2204
rect 0 2120 90 2140
rect 172 2120 212 2164
rect 1996 2120 2036 2164
rect 0 2080 212 2120
rect 1459 2080 1468 2120
rect 1508 2080 2036 2120
rect 2153 2080 2236 2120
rect 2276 2080 2284 2120
rect 2324 2080 2333 2120
rect 3283 2080 3292 2120
rect 3332 2080 4012 2120
rect 4052 2080 4061 2120
rect 0 2060 90 2080
rect 1843 1996 1852 2036
rect 1892 1996 3532 2036
rect 3572 1996 3581 2036
rect 4108 1952 4148 2248
rect 13132 2204 13172 2248
rect 6124 2164 11980 2204
rect 12020 2164 12029 2204
rect 12892 2164 13172 2204
rect 13228 2164 14476 2204
rect 14516 2164 14525 2204
rect 18499 2164 18508 2204
rect 18548 2164 21676 2204
rect 21716 2164 21725 2204
rect 23011 2164 23020 2204
rect 23060 2164 23069 2204
rect 23203 2164 23212 2204
rect 23252 2164 29164 2204
rect 29204 2164 29213 2204
rect 4361 2080 4444 2120
rect 4484 2080 4492 2120
rect 4532 2080 4541 2120
rect 4819 2080 4828 2120
rect 4868 2080 6028 2120
rect 6068 2080 6077 2120
rect 6124 2036 6164 2164
rect 12892 2120 12932 2164
rect 13228 2120 13268 2164
rect 23020 2120 23060 2164
rect 6281 2080 6412 2120
rect 6452 2080 6461 2120
rect 6883 2080 6892 2120
rect 6932 2080 6940 2120
rect 6980 2080 7063 2120
rect 7603 2080 7612 2120
rect 7652 2080 8428 2120
rect 8468 2080 8477 2120
rect 8611 2080 8620 2120
rect 8660 2080 11788 2120
rect 11828 2080 11837 2120
rect 11945 2080 12076 2120
rect 12116 2080 12125 2120
rect 12172 2080 12748 2120
rect 12788 2080 12797 2120
rect 12883 2080 12892 2120
rect 12932 2080 12941 2120
rect 13228 2080 13276 2120
rect 13316 2080 13325 2120
rect 13651 2080 13660 2120
rect 13700 2080 14188 2120
rect 14228 2080 14237 2120
rect 15139 2080 15148 2120
rect 15188 2080 15244 2120
rect 15284 2080 15319 2120
rect 15523 2080 15532 2120
rect 15572 2080 15676 2120
rect 15716 2080 15725 2120
rect 15907 2080 15916 2120
rect 15956 2080 16060 2120
rect 16100 2080 16109 2120
rect 16435 2080 16444 2120
rect 16484 2080 16684 2120
rect 16724 2080 16733 2120
rect 18403 2080 18412 2120
rect 18452 2080 18604 2120
rect 18644 2080 18653 2120
rect 20035 2080 20044 2120
rect 20084 2080 20236 2120
rect 20276 2080 20285 2120
rect 20659 2080 20668 2120
rect 20708 2080 22484 2120
rect 23011 2080 23020 2120
rect 23060 2080 23107 2120
rect 24739 2080 24748 2120
rect 24788 2080 25708 2120
rect 25748 2080 25757 2120
rect 26698 2080 26707 2120
rect 26747 2080 27244 2120
rect 27284 2080 27293 2120
rect 27340 2080 29108 2120
rect 29155 2080 29164 2120
rect 29204 2080 29356 2120
rect 29396 2080 29405 2120
rect 12172 2036 12212 2080
rect 22444 2036 22484 2080
rect 27340 2036 27380 2080
rect 4204 1996 4300 2036
rect 4340 1996 4349 2036
rect 4492 1996 6164 2036
rect 6547 1996 6556 2036
rect 6596 1996 6988 2036
rect 7028 1996 7037 2036
rect 7987 1996 7996 2036
rect 8036 1996 9772 2036
rect 9812 1996 9821 2036
rect 10483 1996 10492 2036
rect 10532 1996 12212 2036
rect 12268 1996 13268 2036
rect 4204 1952 4244 1996
rect 556 1912 1228 1952
rect 1268 1912 1277 1952
rect 1411 1912 1420 1952
rect 1460 1912 1612 1952
rect 1652 1912 1661 1952
rect 1987 1912 1996 1952
rect 2036 1912 2045 1952
rect 2659 1912 2668 1952
rect 2708 1912 2764 1952
rect 2804 1912 2839 1952
rect 3043 1912 3052 1952
rect 3092 1912 3101 1952
rect 3305 1912 3436 1952
rect 3476 1912 3485 1952
rect 3811 1912 3820 1952
rect 3860 1912 4148 1952
rect 4195 1912 4204 1952
rect 4244 1912 4253 1952
rect 0 1784 90 1804
rect 556 1784 596 1912
rect 1996 1868 2036 1912
rect 643 1828 652 1868
rect 692 1828 2036 1868
rect 3052 1868 3092 1912
rect 4492 1868 4532 1996
rect 12268 1952 12308 1996
rect 3052 1828 4532 1868
rect 4588 1912 4627 1952
rect 4667 1912 4676 1952
rect 4771 1912 4780 1952
rect 4820 1912 6260 1952
rect 6787 1912 6796 1952
rect 6836 1912 6932 1952
rect 7049 1912 7180 1952
rect 7220 1912 7229 1952
rect 7363 1912 7372 1952
rect 7412 1912 7543 1952
rect 7747 1912 7756 1952
rect 7796 1912 7805 1952
rect 8009 1912 8140 1952
rect 8180 1912 8189 1952
rect 10243 1912 10252 1952
rect 10292 1912 10301 1952
rect 12259 1912 12268 1952
rect 12308 1912 12317 1952
rect 12377 1912 12460 1952
rect 12500 1912 12508 1952
rect 12548 1912 12557 1952
rect 12643 1912 12652 1952
rect 12692 1912 12844 1952
rect 12884 1912 12893 1952
rect 13027 1912 13036 1952
rect 13076 1912 13085 1952
rect 0 1744 596 1784
rect 2899 1744 2908 1784
rect 2948 1744 4300 1784
rect 4340 1744 4349 1784
rect 0 1724 90 1744
rect 4588 1700 4628 1912
rect 6220 1868 6260 1912
rect 4841 1828 4972 1868
rect 5012 1828 5021 1868
rect 6220 1819 6260 1828
rect 3667 1660 3676 1700
rect 3716 1660 3956 1700
rect 4051 1660 4060 1700
rect 4100 1660 4492 1700
rect 4532 1660 4541 1700
rect 4588 1660 6740 1700
rect 3916 1532 3956 1660
rect 4195 1576 4204 1616
rect 4244 1576 6644 1616
rect 3916 1492 4588 1532
rect 4628 1492 4637 1532
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 0 1448 90 1468
rect 6604 1448 6644 1576
rect 6700 1532 6740 1660
rect 6892 1616 6932 1912
rect 7756 1784 7796 1912
rect 9772 1868 9812 1877
rect 8227 1828 8236 1868
rect 8276 1828 8524 1868
rect 8564 1828 8620 1868
rect 8660 1828 8724 1868
rect 9667 1828 9676 1868
rect 9716 1828 9772 1868
rect 9812 1828 9847 1868
rect 9772 1819 9812 1828
rect 7756 1744 9716 1784
rect 9929 1744 9964 1784
rect 10004 1744 10060 1784
rect 10100 1744 10109 1784
rect 9676 1700 9716 1744
rect 10252 1700 10292 1912
rect 11884 1868 11924 1877
rect 10505 1828 10540 1868
rect 10580 1828 10636 1868
rect 10676 1828 10685 1868
rect 11753 1828 11884 1868
rect 11924 1828 11933 1868
rect 11884 1819 11924 1828
rect 13036 1700 13076 1912
rect 13228 1868 13268 1996
rect 18604 1996 20180 2036
rect 13411 1912 13420 1952
rect 13460 1912 14476 1952
rect 14516 1912 14525 1952
rect 15427 1912 15436 1952
rect 15476 1912 15485 1952
rect 15811 1912 15820 1952
rect 15860 1912 15916 1952
rect 15956 1912 15991 1952
rect 16195 1912 16204 1952
rect 16244 1912 16253 1952
rect 16579 1912 16588 1952
rect 16628 1912 17068 1952
rect 17108 1912 17117 1952
rect 15052 1868 15092 1877
rect 15436 1868 15476 1912
rect 13228 1828 13556 1868
rect 13673 1828 13804 1868
rect 13844 1828 13853 1868
rect 15092 1828 15340 1868
rect 15380 1828 15389 1868
rect 15436 1828 15724 1868
rect 15764 1828 15773 1868
rect 13516 1700 13556 1828
rect 15052 1819 15092 1828
rect 16204 1784 16244 1912
rect 18220 1868 18260 1877
rect 18604 1868 18644 1996
rect 19852 1868 19892 1877
rect 16841 1828 16972 1868
rect 17012 1828 17021 1868
rect 18211 1828 18220 1868
rect 18260 1828 18391 1868
rect 18595 1828 18604 1868
rect 18644 1828 18775 1868
rect 19363 1828 19372 1868
rect 19412 1828 19852 1868
rect 20140 1868 20180 1996
rect 20428 1996 21004 2036
rect 21044 1996 21053 2036
rect 21100 1996 22348 2036
rect 22388 1996 22397 2036
rect 22444 1996 23116 2036
rect 23156 1996 23165 2036
rect 24547 1996 24556 2036
rect 24596 1996 25172 2036
rect 25411 1996 25420 2036
rect 25460 1996 27380 2036
rect 20428 1952 20468 1996
rect 21100 1952 21140 1996
rect 25132 1952 25172 1996
rect 29068 1952 29108 2080
rect 29644 2036 29684 2248
rect 31948 2204 31988 2248
rect 40492 2204 40532 2584
rect 44524 2540 44564 2584
rect 43459 2500 43468 2540
rect 43508 2500 44564 2540
rect 44755 2500 44764 2540
rect 44804 2500 45812 2540
rect 45772 2456 45812 2500
rect 46278 2456 46368 2476
rect 44371 2416 44380 2456
rect 44420 2416 45292 2456
rect 45332 2416 45341 2456
rect 45772 2416 46368 2456
rect 46278 2396 46368 2416
rect 29827 2164 29836 2204
rect 29876 2164 31988 2204
rect 35116 2164 37996 2204
rect 38036 2164 38045 2204
rect 38188 2164 40532 2204
rect 35116 2120 35156 2164
rect 38188 2120 38228 2164
rect 46278 2120 46368 2140
rect 29923 2080 29932 2120
rect 29972 2080 31564 2120
rect 31604 2080 31613 2120
rect 31913 2080 32044 2120
rect 32084 2080 32093 2120
rect 32428 2080 33716 2120
rect 29155 1996 29164 2036
rect 29204 1996 29588 2036
rect 29644 1996 30356 2036
rect 29548 1952 29588 1996
rect 30316 1952 30356 1996
rect 32428 1952 32468 2080
rect 33676 2036 33716 2080
rect 34060 2080 35156 2120
rect 36010 2080 36019 2120
rect 36059 2080 38228 2120
rect 38633 2080 38764 2120
rect 38804 2080 38813 2120
rect 45139 2080 45148 2120
rect 45188 2080 46368 2120
rect 33100 1996 33332 2036
rect 33676 1996 33964 2036
rect 34004 1996 34013 2036
rect 20419 1912 20428 1952
rect 20468 1912 20477 1952
rect 20803 1912 20812 1952
rect 20852 1912 21140 1952
rect 21187 1912 21196 1952
rect 21236 1912 22060 1952
rect 22100 1912 22109 1952
rect 24460 1912 24940 1952
rect 24980 1912 24989 1952
rect 25132 1912 25420 1952
rect 25460 1912 25469 1952
rect 25996 1912 26708 1952
rect 26921 1912 26956 1952
rect 26996 1912 27052 1952
rect 27092 1912 27101 1952
rect 27305 1912 27436 1952
rect 27476 1912 27485 1952
rect 27619 1912 27628 1952
rect 27668 1912 29012 1952
rect 29068 1912 29308 1952
rect 29348 1912 29357 1952
rect 29539 1912 29548 1952
rect 29588 1912 29597 1952
rect 29731 1912 29740 1952
rect 29780 1912 29932 1952
rect 29972 1912 29981 1952
rect 30307 1912 30316 1952
rect 30356 1912 30365 1952
rect 32419 1912 32428 1952
rect 32468 1912 32477 1952
rect 32803 1912 32812 1952
rect 32852 1912 33004 1952
rect 33044 1912 33053 1952
rect 22828 1868 22868 1877
rect 24460 1868 24500 1912
rect 25996 1868 26036 1912
rect 26668 1868 26708 1912
rect 28972 1868 29012 1912
rect 31852 1868 31892 1877
rect 33100 1868 33140 1996
rect 33187 1912 33196 1952
rect 33236 1912 33245 1952
rect 20140 1828 21580 1868
rect 21620 1828 21629 1868
rect 22697 1828 22828 1868
rect 22868 1828 22877 1868
rect 23177 1828 23212 1868
rect 23252 1828 23308 1868
rect 23348 1828 23357 1868
rect 18220 1819 18260 1828
rect 19852 1819 19892 1828
rect 22828 1819 22868 1828
rect 24460 1819 24500 1828
rect 24652 1828 24931 1868
rect 24971 1828 24980 1868
rect 25027 1828 25036 1868
rect 25076 1828 25085 1868
rect 25507 1828 25516 1868
rect 25556 1828 25708 1868
rect 25748 1828 25757 1868
rect 26275 1828 26284 1868
rect 26324 1828 26484 1868
rect 26524 1828 26533 1868
rect 26668 1828 27532 1868
rect 27572 1828 27581 1868
rect 27715 1828 27724 1868
rect 27764 1828 27895 1868
rect 29012 1828 29932 1868
rect 29972 1828 29981 1868
rect 30403 1828 30412 1868
rect 30452 1828 30604 1868
rect 30644 1828 30653 1868
rect 31555 1828 31564 1868
rect 31604 1828 31852 1868
rect 31892 1828 32044 1868
rect 32084 1828 32093 1868
rect 32419 1828 32428 1868
rect 32468 1828 33140 1868
rect 24652 1784 24692 1828
rect 25036 1784 25076 1828
rect 25996 1784 26036 1828
rect 28972 1819 29012 1828
rect 31852 1819 31892 1828
rect 33196 1784 33236 1912
rect 33292 1868 33332 1996
rect 33449 1912 33484 1952
rect 33524 1912 33580 1952
rect 33620 1912 33629 1952
rect 33763 1912 33772 1952
rect 33812 1912 33964 1952
rect 34004 1912 34013 1952
rect 34060 1868 34100 2080
rect 34723 1996 34732 2036
rect 34772 1996 34781 2036
rect 34732 1952 34772 1996
rect 34252 1912 34540 1952
rect 34580 1912 34589 1952
rect 34636 1912 34772 1952
rect 34819 1912 34828 1952
rect 34868 1912 34924 1952
rect 34964 1912 34999 1952
rect 34252 1868 34292 1912
rect 34636 1868 34676 1912
rect 35116 1868 35156 2080
rect 46278 2060 46368 2080
rect 33292 1828 34100 1868
rect 34234 1828 34243 1868
rect 34283 1828 34292 1868
rect 34339 1828 34348 1868
rect 34388 1828 34676 1868
rect 34723 1828 34732 1868
rect 34772 1828 35156 1868
rect 35212 1996 37268 2036
rect 37769 1996 37900 2036
rect 37940 1996 40244 2036
rect 41635 1996 41644 2036
rect 41684 1996 44564 2036
rect 44611 1996 44620 2036
rect 44660 1996 44669 2036
rect 35212 1784 35252 1996
rect 37228 1952 37268 1996
rect 35308 1912 35884 1952
rect 35924 1912 35933 1952
rect 37228 1912 37844 1952
rect 35308 1868 35348 1912
rect 36652 1868 36692 1877
rect 35818 1828 35827 1868
rect 35867 1828 36500 1868
rect 35308 1819 35348 1828
rect 36460 1784 36500 1828
rect 36692 1828 37420 1868
rect 37460 1828 37469 1868
rect 36652 1819 36692 1828
rect 37804 1784 37844 1912
rect 37900 1868 37940 1996
rect 38153 1912 38284 1952
rect 38324 1912 38333 1952
rect 38956 1868 38996 1877
rect 40204 1868 40244 1996
rect 44524 1952 44564 1996
rect 44620 1952 44660 1996
rect 43747 1912 43756 1952
rect 43796 1912 43805 1952
rect 44009 1912 44140 1952
rect 44180 1912 44189 1952
rect 44515 1912 44524 1952
rect 44564 1912 44573 1952
rect 44620 1912 44908 1952
rect 44948 1912 44957 1952
rect 37891 1828 37900 1868
rect 37940 1828 37949 1868
rect 38825 1828 38956 1868
rect 38996 1828 39005 1868
rect 40195 1828 40204 1868
rect 40244 1828 40253 1868
rect 38956 1819 38996 1828
rect 16204 1744 18028 1784
rect 18068 1744 18077 1784
rect 20035 1744 20044 1784
rect 20084 1744 21484 1784
rect 21524 1744 21533 1784
rect 24643 1744 24652 1784
rect 24692 1744 24701 1784
rect 24931 1744 24940 1784
rect 24980 1744 25076 1784
rect 25315 1744 25324 1784
rect 25364 1744 26036 1784
rect 29251 1744 29260 1784
rect 29300 1744 31276 1784
rect 31316 1744 31325 1784
rect 33196 1744 35252 1784
rect 36451 1744 36460 1784
rect 36500 1744 36509 1784
rect 37804 1744 38900 1784
rect 38860 1700 38900 1744
rect 8371 1660 8380 1700
rect 8420 1660 8620 1700
rect 8660 1660 8669 1700
rect 9676 1660 10156 1700
rect 10196 1660 10205 1700
rect 10252 1660 12940 1700
rect 12980 1660 12989 1700
rect 13036 1660 13364 1700
rect 13516 1660 14572 1700
rect 14612 1660 14621 1700
rect 16819 1660 16828 1700
rect 16868 1660 20948 1700
rect 21043 1660 21052 1700
rect 21092 1660 21332 1700
rect 21427 1660 21436 1700
rect 21476 1660 23692 1700
rect 23732 1660 23741 1700
rect 26188 1660 26812 1700
rect 26852 1660 26861 1700
rect 26956 1660 27196 1700
rect 27236 1660 27245 1700
rect 27340 1660 29692 1700
rect 29732 1660 29741 1700
rect 29836 1660 30076 1700
rect 30116 1660 30125 1700
rect 31651 1660 31660 1700
rect 31700 1660 32188 1700
rect 32228 1660 32237 1700
rect 32419 1660 32428 1700
rect 32468 1660 32572 1700
rect 32612 1660 32621 1700
rect 32812 1660 32956 1700
rect 32996 1660 33005 1700
rect 33187 1660 33196 1700
rect 33236 1660 33340 1700
rect 33380 1660 33389 1700
rect 33475 1660 33484 1700
rect 33524 1660 33724 1700
rect 33764 1660 33773 1700
rect 34732 1660 34964 1700
rect 36163 1660 36172 1700
rect 36212 1660 38044 1700
rect 38084 1660 38093 1700
rect 38860 1660 39724 1700
rect 39764 1660 39773 1700
rect 6892 1576 13172 1616
rect 6700 1492 13036 1532
rect 13076 1492 13085 1532
rect 13132 1448 13172 1576
rect 13324 1532 13364 1660
rect 20908 1616 20948 1660
rect 21292 1616 21332 1660
rect 26188 1616 26228 1660
rect 13699 1576 13708 1616
rect 13748 1576 20716 1616
rect 20756 1576 20765 1616
rect 20908 1576 21196 1616
rect 21236 1576 21245 1616
rect 21292 1576 23308 1616
rect 23348 1576 23357 1616
rect 24643 1576 24652 1616
rect 24692 1576 26228 1616
rect 26956 1532 26996 1660
rect 27340 1532 27380 1660
rect 29836 1616 29876 1660
rect 32812 1616 32852 1660
rect 34732 1616 34772 1660
rect 29539 1576 29548 1616
rect 29588 1576 29876 1616
rect 32428 1576 32852 1616
rect 32899 1576 32908 1616
rect 32948 1576 34772 1616
rect 34924 1616 34964 1660
rect 43756 1616 43796 1912
rect 46278 1784 46368 1804
rect 43987 1744 43996 1784
rect 44036 1744 44620 1784
rect 44660 1744 44669 1784
rect 44755 1744 44764 1784
rect 44804 1744 46368 1784
rect 46278 1724 46368 1744
rect 44371 1660 44380 1700
rect 44420 1660 45388 1700
rect 45428 1660 45437 1700
rect 34924 1576 43796 1616
rect 32428 1532 32468 1576
rect 13324 1492 14900 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 22540 1492 24556 1532
rect 24596 1492 24605 1532
rect 24835 1492 24844 1532
rect 24884 1492 26996 1532
rect 27052 1492 27380 1532
rect 30220 1492 32468 1532
rect 32812 1492 34924 1532
rect 34964 1492 34973 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 35596 1492 39820 1532
rect 39860 1492 39869 1532
rect 0 1408 652 1448
rect 692 1408 701 1448
rect 6604 1408 12172 1448
rect 12212 1408 12221 1448
rect 13132 1408 14284 1448
rect 14324 1408 14333 1448
rect 0 1388 90 1408
rect 14860 1280 14900 1492
rect 22540 1448 22580 1492
rect 27052 1448 27092 1492
rect 30220 1448 30260 1492
rect 15907 1408 15916 1448
rect 15956 1408 20180 1448
rect 21475 1408 21484 1448
rect 21524 1408 22580 1448
rect 25603 1408 25612 1448
rect 25652 1408 27092 1448
rect 27331 1408 27340 1448
rect 27380 1408 30260 1448
rect 20140 1364 20180 1408
rect 32812 1364 32852 1492
rect 35596 1448 35636 1492
rect 46278 1448 46368 1468
rect 34147 1408 34156 1448
rect 34196 1408 35636 1448
rect 45283 1408 45292 1448
rect 45332 1408 46368 1448
rect 46278 1388 46368 1408
rect 20140 1324 20428 1364
rect 20468 1324 20477 1364
rect 27523 1324 27532 1364
rect 27572 1324 32852 1364
rect 34243 1324 34252 1364
rect 34292 1324 41452 1364
rect 41492 1324 41501 1364
rect 14860 1240 18892 1280
rect 18932 1240 18941 1280
rect 0 1112 90 1132
rect 46278 1112 46368 1132
rect 0 1072 1420 1112
rect 1460 1072 1469 1112
rect 44611 1072 44620 1112
rect 44660 1072 46368 1112
rect 0 1052 90 1072
rect 46278 1052 46368 1072
rect 28099 904 28108 944
rect 28148 904 33484 944
rect 33524 904 33533 944
rect 10147 820 10156 860
rect 10196 820 16204 860
rect 16244 820 16253 860
rect 27715 820 27724 860
rect 27764 820 33196 860
rect 33236 820 33245 860
rect 0 776 90 796
rect 46278 776 46368 796
rect 0 736 1132 776
rect 1172 736 1181 776
rect 45379 736 45388 776
rect 45428 736 46368 776
rect 0 716 90 736
rect 46278 716 46368 736
rect 33859 652 33868 692
rect 33908 652 40108 692
rect 40148 652 40157 692
rect 4387 568 4396 608
rect 4436 568 11788 608
rect 11828 568 11837 608
rect 33091 400 33100 440
rect 33140 400 42604 440
rect 42644 400 42653 440
rect 32899 148 32908 188
rect 32948 148 42892 188
rect 42932 148 42941 188
rect 33475 64 33484 104
rect 33524 64 43660 104
rect 43700 64 43709 104
<< via2 >>
rect 32524 11656 32564 11696
rect 42508 11656 42548 11696
rect 35596 11572 35636 11612
rect 42316 11572 42356 11612
rect 37516 11488 37556 11528
rect 44524 11488 44564 11528
rect 35692 11404 35732 11444
rect 44716 11404 44756 11444
rect 32620 11320 32660 11360
rect 44332 11320 44372 11360
rect 16972 11236 17012 11276
rect 38956 11236 38996 11276
rect 76 11152 116 11192
rect 34924 11152 34964 11192
rect 45004 11152 45044 11192
rect 1996 11068 2036 11108
rect 14476 11068 14516 11108
rect 37804 11068 37844 11108
rect 42124 11068 42164 11108
rect 42316 11068 42356 11108
rect 43564 11068 43604 11108
rect 45100 11068 45140 11108
rect 11500 10984 11540 11024
rect 28012 10984 28052 11024
rect 29260 10984 29300 11024
rect 35020 10984 35060 11024
rect 38764 10984 38804 11024
rect 18412 10900 18452 10940
rect 32908 10900 32948 10940
rect 40300 10900 40340 10940
rect 1324 10816 1364 10856
rect 3052 10816 3092 10856
rect 9676 10816 9716 10856
rect 14572 10816 14612 10856
rect 40588 10816 40628 10856
rect 43852 10816 43892 10856
rect 14764 10732 14804 10772
rect 21484 10732 21524 10772
rect 28108 10732 28148 10772
rect 38380 10732 38420 10772
rect 42988 10732 43028 10772
rect 76 10648 116 10688
rect 1996 10396 2036 10436
rect 8236 10648 8276 10688
rect 19564 10648 19604 10688
rect 27532 10648 27572 10688
rect 29260 10648 29300 10688
rect 29452 10648 29492 10688
rect 37516 10648 37556 10688
rect 44428 10648 44468 10688
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 3052 10396 3092 10436
rect 4684 10396 4724 10436
rect 9676 10480 9716 10520
rect 16396 10480 16436 10520
rect 5836 10396 5876 10436
rect 6892 10396 6932 10436
rect 8140 10396 8180 10436
rect 10444 10396 10484 10436
rect 11596 10396 11636 10436
rect 12748 10396 12788 10436
rect 16204 10396 16244 10436
rect 17356 10396 17396 10436
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 25612 10564 25652 10604
rect 28012 10564 28052 10604
rect 34732 10564 34772 10604
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 39052 10564 39092 10604
rect 20140 10396 20180 10436
rect 20716 10396 20756 10436
rect 7276 10312 7316 10352
rect 9292 10312 9332 10352
rect 6796 10228 6836 10268
rect 7084 10228 7124 10268
rect 7660 10228 7700 10268
rect 1132 10144 1172 10184
rect 3532 10144 3572 10184
rect 6700 10144 6740 10184
rect 6988 10144 7028 10184
rect 8908 10144 8948 10184
rect 10924 10228 10964 10268
rect 11692 10228 11732 10268
rect 11116 10144 11156 10184
rect 11500 10144 11540 10184
rect 14476 10228 14516 10268
rect 14860 10228 14900 10268
rect 16396 10259 16436 10268
rect 16396 10228 16436 10259
rect 14380 10144 14420 10184
rect 2284 10060 2324 10100
rect 5356 10060 5396 10100
rect 5740 10060 5780 10100
rect 6220 10060 6260 10100
rect 7180 10060 7220 10100
rect 8428 10060 8468 10100
rect 12844 10060 12884 10100
rect 20140 10228 20180 10268
rect 21292 10228 21332 10268
rect 21484 10228 21524 10268
rect 21868 10228 21908 10268
rect 34348 10480 34388 10520
rect 43276 10480 43316 10520
rect 24268 10396 24308 10436
rect 26572 10396 26612 10436
rect 27724 10396 27764 10436
rect 28876 10396 28916 10436
rect 30028 10396 30068 10436
rect 34636 10396 34676 10436
rect 26860 10312 26900 10352
rect 31180 10312 31220 10352
rect 33580 10312 33620 10352
rect 34252 10312 34292 10352
rect 24172 10228 24212 10268
rect 25036 10228 25076 10268
rect 25804 10228 25844 10268
rect 16972 10144 17012 10184
rect 19468 10144 19508 10184
rect 28108 10228 28148 10268
rect 29644 10228 29684 10268
rect 30700 10228 30740 10268
rect 33196 10228 33236 10268
rect 34828 10228 34868 10268
rect 35020 10228 35060 10268
rect 29452 10144 29492 10184
rect 31468 10144 31508 10184
rect 31660 10144 31700 10184
rect 32524 10144 32564 10184
rect 32908 10144 32948 10184
rect 35788 10396 35828 10436
rect 36940 10396 36980 10436
rect 38092 10396 38132 10436
rect 39244 10396 39284 10436
rect 40588 10396 40628 10436
rect 41548 10396 41588 10436
rect 42700 10396 42740 10436
rect 38956 10312 38996 10352
rect 40396 10312 40436 10352
rect 43180 10312 43220 10352
rect 43372 10312 43412 10352
rect 35788 10228 35828 10268
rect 37804 10144 37844 10184
rect 38380 10144 38420 10184
rect 39244 10228 39284 10268
rect 42028 10228 42068 10268
rect 42892 10228 42932 10268
rect 39148 10144 39188 10184
rect 43276 10144 43316 10184
rect 43564 10144 43604 10184
rect 43756 10144 43796 10184
rect 44332 10144 44372 10184
rect 44716 10144 44756 10184
rect 45100 10144 45140 10184
rect 45484 10144 45524 10184
rect 14668 10060 14708 10100
rect 15148 10060 15188 10100
rect 17452 10060 17492 10100
rect 19948 10060 19988 10100
rect 25900 10060 25940 10100
rect 27340 10060 27380 10100
rect 27628 10060 27668 10100
rect 36268 10060 36308 10100
rect 38284 10060 38324 10100
rect 41740 10060 41780 10100
rect 44236 10060 44276 10100
rect 2956 9976 2996 10016
rect 10732 9976 10772 10016
rect 13324 9976 13364 10016
rect 13516 9976 13556 10016
rect 14956 9976 14996 10016
rect 17644 9976 17684 10016
rect 17836 9976 17876 10016
rect 18700 9976 18740 10016
rect 19276 9976 19316 10016
rect 20044 9976 20084 10016
rect 23308 9976 23348 10016
rect 27052 9976 27092 10016
rect 29452 9976 29492 10016
rect 29740 9976 29780 10016
rect 31756 9976 31796 10016
rect 34540 9976 34580 10016
rect 36652 9976 36692 10016
rect 41836 9976 41876 10016
rect 2092 9892 2132 9932
rect 8524 9892 8564 9932
rect 25132 9892 25172 9932
rect 26956 9892 26996 9932
rect 33100 9892 33140 9932
rect 34828 9892 34868 9932
rect 40396 9892 40436 9932
rect 42028 9892 42068 9932
rect 42220 9892 42260 9932
rect 43276 9892 43316 9932
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 10540 9808 10580 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 21868 9808 21908 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 34636 9808 34676 9848
rect 41932 9808 41972 9848
rect 44812 9808 44852 9848
rect 2668 9724 2708 9764
rect 5740 9724 5780 9764
rect 20140 9724 20180 9764
rect 6316 9640 6356 9680
rect 7276 9640 7316 9680
rect 8428 9640 8468 9680
rect 12460 9640 12500 9680
rect 13900 9640 13940 9680
rect 15052 9640 15092 9680
rect 18508 9640 18548 9680
rect 18700 9640 18740 9680
rect 1132 9556 1172 9596
rect 1324 9556 1364 9596
rect 1228 9472 1268 9512
rect 7948 9472 7988 9512
rect 8524 9472 8564 9512
rect 5548 9388 5588 9428
rect 7084 9388 7124 9428
rect 2188 9220 2228 9260
rect 5740 9220 5780 9260
rect 7276 9304 7316 9344
rect 20812 9640 20852 9680
rect 34444 9724 34484 9764
rect 39052 9724 39092 9764
rect 42796 9724 42836 9764
rect 25420 9640 25460 9680
rect 11788 9556 11828 9596
rect 21964 9556 22004 9596
rect 22156 9556 22196 9596
rect 24940 9556 24980 9596
rect 9004 9472 9044 9512
rect 11308 9472 11348 9512
rect 14092 9472 14132 9512
rect 14572 9472 14612 9512
rect 15532 9472 15572 9512
rect 16972 9472 17012 9512
rect 17836 9472 17876 9512
rect 21004 9472 21044 9512
rect 22252 9472 22292 9512
rect 9676 9388 9716 9428
rect 10924 9388 10964 9428
rect 7852 9304 7892 9344
rect 6796 9136 6836 9176
rect 7756 9136 7796 9176
rect 8620 9220 8660 9260
rect 9100 9220 9140 9260
rect 10060 9220 10100 9260
rect 11212 9220 11252 9260
rect 11596 9360 11627 9400
rect 11627 9360 11636 9400
rect 12076 9388 12116 9428
rect 12748 9388 12788 9428
rect 13324 9388 13364 9428
rect 14956 9388 14996 9428
rect 15436 9388 15476 9428
rect 15820 9388 15860 9428
rect 16588 9388 16596 9428
rect 16596 9388 16628 9428
rect 17740 9388 17780 9428
rect 18124 9388 18164 9428
rect 18508 9388 18548 9428
rect 18988 9388 19028 9428
rect 20044 9388 20084 9428
rect 20908 9388 20948 9428
rect 21484 9388 21524 9428
rect 23308 9388 23348 9428
rect 11884 9304 11924 9344
rect 12652 9304 12692 9344
rect 14668 9304 14708 9344
rect 15052 9304 15092 9344
rect 21580 9304 21620 9344
rect 21772 9304 21812 9344
rect 22060 9304 22100 9344
rect 22732 9304 22772 9344
rect 24652 9388 24692 9428
rect 26476 9472 26516 9512
rect 26956 9472 26996 9512
rect 27340 9472 27380 9512
rect 25420 9388 25460 9428
rect 25900 9388 25908 9428
rect 25908 9388 25940 9428
rect 32332 9640 32372 9680
rect 33484 9640 33524 9680
rect 40300 9640 40340 9680
rect 44428 9640 44468 9680
rect 27820 9472 27860 9512
rect 29548 9472 29588 9512
rect 31660 9472 31700 9512
rect 28396 9388 28436 9428
rect 38956 9556 38996 9596
rect 39244 9556 39284 9596
rect 41548 9556 41588 9596
rect 41740 9556 41780 9596
rect 34156 9472 34196 9512
rect 34540 9472 34580 9512
rect 34828 9472 34868 9512
rect 36748 9472 36788 9512
rect 39148 9472 39188 9512
rect 39340 9472 39380 9512
rect 42028 9472 42068 9512
rect 42508 9472 42548 9512
rect 42892 9472 42932 9512
rect 43084 9472 43124 9512
rect 43276 9472 43316 9512
rect 43660 9472 43700 9512
rect 44044 9472 44084 9512
rect 31468 9388 31508 9428
rect 32332 9388 32372 9428
rect 24364 9304 24404 9344
rect 27436 9304 27476 9344
rect 27916 9304 27956 9344
rect 29548 9304 29588 9344
rect 31756 9304 31796 9344
rect 11788 9220 11828 9260
rect 14380 9220 14420 9260
rect 16972 9220 17012 9260
rect 18508 9220 18548 9260
rect 19372 9220 19412 9260
rect 25900 9220 25940 9260
rect 29068 9220 29108 9260
rect 14284 9136 14324 9176
rect 18700 9136 18740 9176
rect 21100 9136 21140 9176
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 8332 9052 8372 9092
rect 11308 9052 11348 9092
rect 15916 9052 15956 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 20620 9052 20660 9092
rect 20908 9052 20948 9092
rect 21772 9052 21812 9092
rect 24748 9052 24788 9092
rect 25132 9052 25172 9092
rect 32716 9052 32756 9092
rect 9964 8968 10004 9008
rect 12364 8968 12404 9008
rect 34924 9388 34964 9428
rect 35884 9388 35924 9428
rect 36652 9388 36692 9428
rect 37132 9388 37172 9428
rect 38380 9388 38420 9428
rect 38764 9388 38804 9428
rect 40396 9388 40401 9428
rect 40401 9388 40436 9428
rect 41740 9388 41780 9428
rect 34444 9304 34484 9344
rect 36940 9304 36980 9344
rect 40204 9304 40244 9344
rect 41356 9304 41396 9344
rect 43948 9304 43988 9344
rect 33388 9220 33428 9260
rect 36268 9220 36308 9260
rect 36844 9220 36884 9260
rect 40396 9220 40436 9260
rect 42028 9220 42068 9260
rect 42796 9220 42836 9260
rect 43372 9220 43412 9260
rect 37420 9136 37460 9176
rect 41452 9136 41492 9176
rect 43276 9136 43316 9176
rect 44620 9136 44660 9176
rect 33292 9052 33332 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 37324 9052 37364 9092
rect 43084 9052 43124 9092
rect 16588 8968 16628 9008
rect 21196 8968 21236 9008
rect 21484 8968 21524 9008
rect 27916 8968 27956 9008
rect 32524 8968 32564 9008
rect 33196 8968 33236 9008
rect 34828 8968 34868 9008
rect 41740 8968 41780 9008
rect 41932 8968 41972 9008
rect 43372 8968 43412 9008
rect 11020 8884 11060 8924
rect 12460 8884 12500 8924
rect 18124 8884 18164 8924
rect 19468 8884 19508 8924
rect 19660 8884 19700 8924
rect 1228 8800 1268 8840
rect 21964 8884 22004 8924
rect 23980 8884 24020 8924
rect 24364 8884 24404 8924
rect 24940 8884 24980 8924
rect 27820 8884 27860 8924
rect 32812 8884 32852 8924
rect 34924 8884 34964 8924
rect 38476 8884 38516 8924
rect 39724 8884 39764 8924
rect 42028 8884 42068 8924
rect 44044 8884 44084 8924
rect 44524 8884 44564 8924
rect 6988 8800 7028 8840
rect 9100 8800 9140 8840
rect 10540 8800 10580 8840
rect 10732 8800 10772 8840
rect 11212 8800 11252 8840
rect 5548 8747 5588 8756
rect 5548 8716 5588 8747
rect 5932 8716 5972 8756
rect 7084 8716 7124 8756
rect 7948 8716 7979 8756
rect 7979 8716 7988 8756
rect 8428 8716 8468 8756
rect 8812 8716 8852 8756
rect 10060 8716 10100 8756
rect 10828 8716 10868 8756
rect 11308 8716 11348 8756
rect 11884 8716 11924 8756
rect 21868 8800 21908 8840
rect 25804 8800 25844 8840
rect 25996 8800 26036 8840
rect 29644 8800 29684 8840
rect 33196 8800 33236 8840
rect 35980 8800 36020 8840
rect 12844 8716 12876 8756
rect 12876 8716 12884 8756
rect 14284 8716 14324 8756
rect 14860 8716 14900 8756
rect 15916 8716 15956 8756
rect 17452 8716 17492 8756
rect 17740 8716 17780 8756
rect 18124 8716 18164 8756
rect 18508 8716 18548 8756
rect 19276 8716 19316 8756
rect 19948 8716 19988 8756
rect 20812 8716 20852 8756
rect 21676 8716 21716 8756
rect 24076 8747 24116 8756
rect 24076 8716 24116 8747
rect 24652 8716 24692 8756
rect 24940 8716 24980 8756
rect 25708 8716 25748 8756
rect 27052 8716 27092 8756
rect 28012 8716 28052 8756
rect 28300 8747 28340 8756
rect 28300 8716 28340 8747
rect 29740 8716 29780 8756
rect 30220 8716 30260 8756
rect 30508 8716 30548 8756
rect 31084 8747 31124 8756
rect 31084 8716 31124 8747
rect 31564 8747 31604 8756
rect 31564 8716 31604 8747
rect 31852 8716 31892 8756
rect 1228 8632 1268 8672
rect 1996 8632 2036 8672
rect 2572 8632 2612 8672
rect 2764 8632 2804 8672
rect 4300 8632 4340 8672
rect 10636 8632 10676 8672
rect 11404 8632 11444 8672
rect 13036 8632 13076 8672
rect 13996 8632 14036 8672
rect 14188 8632 14228 8672
rect 17548 8632 17588 8672
rect 18604 8632 18644 8672
rect 21388 8632 21428 8672
rect 22060 8632 22100 8672
rect 29068 8632 29108 8672
rect 30892 8632 30932 8672
rect 32140 8632 32180 8672
rect 33004 8632 33044 8672
rect 6604 8548 6644 8588
rect 7372 8548 7412 8588
rect 11884 8548 11924 8588
rect 15820 8548 15860 8588
rect 29452 8548 29492 8588
rect 6796 8464 6836 8504
rect 7468 8464 7508 8504
rect 30412 8548 30452 8588
rect 34540 8716 34580 8756
rect 34828 8716 34868 8756
rect 33196 8632 33236 8672
rect 36268 8716 36308 8756
rect 36748 8716 36788 8756
rect 37036 8716 37076 8756
rect 38380 8716 38420 8756
rect 40492 8716 40532 8756
rect 40780 8716 40820 8756
rect 41356 8747 41396 8756
rect 41356 8716 41396 8747
rect 41644 8716 41684 8756
rect 34444 8632 34484 8672
rect 34924 8632 34964 8672
rect 38572 8632 38612 8672
rect 40396 8632 40436 8672
rect 42796 8632 42836 8672
rect 42988 8632 43028 8672
rect 43372 8632 43412 8672
rect 43756 8632 43796 8672
rect 44716 8632 44756 8672
rect 44908 8632 44948 8672
rect 46252 8632 46292 8672
rect 34540 8548 34580 8588
rect 41452 8548 41492 8588
rect 9292 8464 9332 8504
rect 13420 8464 13460 8504
rect 13804 8464 13844 8504
rect 24364 8464 24404 8504
rect 26668 8464 26708 8504
rect 28492 8464 28532 8504
rect 29260 8464 29300 8504
rect 29836 8464 29876 8504
rect 30028 8464 30068 8504
rect 38188 8464 38228 8504
rect 5452 8380 5492 8420
rect 9676 8380 9716 8420
rect 11308 8380 11348 8420
rect 14188 8380 14228 8420
rect 22540 8380 22580 8420
rect 23404 8380 23444 8420
rect 35884 8380 35924 8420
rect 39820 8464 39860 8504
rect 41548 8464 41588 8504
rect 41644 8380 41684 8420
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 7660 8296 7700 8336
rect 8524 8296 8564 8336
rect 11500 8296 11540 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 25420 8296 25460 8336
rect 28300 8296 28340 8336
rect 28588 8296 28628 8336
rect 31660 8296 31700 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 9868 8212 9908 8252
rect 11884 8212 11924 8252
rect 1228 8128 1268 8168
rect 6988 8128 7028 8168
rect 7372 8128 7412 8168
rect 10252 8128 10292 8168
rect 11020 8128 11060 8168
rect 11500 8128 11540 8168
rect 13612 8128 13652 8168
rect 13804 8128 13844 8168
rect 1228 7960 1268 8000
rect 6508 7960 6548 8000
rect 2572 7876 2612 7916
rect 3436 7876 3476 7916
rect 4300 7876 4340 7916
rect 5932 7876 5972 7916
rect 6604 7876 6644 7916
rect 7468 8044 7508 8084
rect 7660 8044 7700 8084
rect 38092 8212 38132 8252
rect 45004 8296 45044 8336
rect 45484 8212 45524 8252
rect 15244 8128 15284 8168
rect 17740 8128 17780 8168
rect 17932 8128 17972 8168
rect 23116 8128 23156 8168
rect 8044 8044 8084 8084
rect 8140 7960 8171 8000
rect 8171 7960 8180 8000
rect 7372 7876 7412 7916
rect 7660 7876 7700 7916
rect 6988 7792 7028 7832
rect 7276 7792 7316 7832
rect 1708 7708 1748 7748
rect 4972 7708 5012 7748
rect 7084 7708 7124 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 7276 7624 7316 7664
rect 7852 7624 7892 7664
rect 8716 7960 8756 8000
rect 13708 8044 13748 8084
rect 22924 8044 22964 8084
rect 23500 8044 23540 8084
rect 26188 8044 26228 8084
rect 12460 7960 12500 8000
rect 13132 7960 13172 8000
rect 13516 7960 13556 8000
rect 14188 7960 14228 8000
rect 15628 7960 15668 8000
rect 17260 7960 17300 8000
rect 18316 7960 18356 8000
rect 19084 7960 19124 8000
rect 19756 7960 19796 8000
rect 21772 7960 21812 8000
rect 23404 7960 23444 8000
rect 23788 7960 23828 8000
rect 27436 7960 27476 8000
rect 28588 7960 28628 8000
rect 29452 7960 29492 8000
rect 8524 7876 8564 7916
rect 9292 7876 9332 7916
rect 9484 7876 9524 7916
rect 10060 7876 10100 7916
rect 10348 7876 10379 7916
rect 10379 7876 10388 7916
rect 11788 7876 11828 7916
rect 13900 7876 13940 7916
rect 14764 7876 14804 7916
rect 8908 7792 8948 7832
rect 13804 7792 13844 7832
rect 14956 7792 14996 7832
rect 15628 7792 15668 7832
rect 9580 7708 9620 7748
rect 31660 8128 31700 8168
rect 34156 8128 34196 8168
rect 34444 8128 34484 8168
rect 36268 8128 36308 8168
rect 36652 8128 36692 8168
rect 37132 8128 37172 8168
rect 43948 8128 43988 8168
rect 46252 8128 46292 8168
rect 30508 8044 30548 8084
rect 31468 8044 31508 8084
rect 40780 8044 40820 8084
rect 41836 8044 41876 8084
rect 32812 7960 32852 8000
rect 36652 7960 36692 8000
rect 36844 7960 36884 8000
rect 38188 7960 38228 8000
rect 42316 7960 42356 8000
rect 42700 7960 42740 8000
rect 43084 7960 43124 8000
rect 43372 7960 43412 8000
rect 44524 7960 44564 8000
rect 44908 7960 44948 8000
rect 16684 7876 16724 7916
rect 18220 7876 18260 7916
rect 18412 7876 18452 7916
rect 19660 7876 19700 7916
rect 21004 7876 21044 7916
rect 21964 7876 22004 7916
rect 23116 7876 23156 7916
rect 24172 7876 24212 7916
rect 25420 7876 25460 7916
rect 26092 7876 26132 7916
rect 26284 7876 26315 7916
rect 26315 7876 26324 7916
rect 26668 7876 26708 7916
rect 28492 7876 28500 7916
rect 28500 7876 28532 7916
rect 30412 7876 30452 7916
rect 30892 7876 30932 7916
rect 31084 7876 31124 7916
rect 31660 7876 31700 7916
rect 31948 7876 31988 7916
rect 34252 7876 34292 7916
rect 34924 7876 34964 7916
rect 35788 7876 35828 7916
rect 38092 7876 38132 7916
rect 38476 7876 38509 7916
rect 38509 7876 38516 7916
rect 39820 7876 39860 7916
rect 16780 7792 16820 7832
rect 24652 7792 24692 7832
rect 26476 7792 26516 7832
rect 27148 7792 27188 7832
rect 30028 7792 30068 7832
rect 30316 7792 30356 7832
rect 31756 7792 31796 7832
rect 32428 7792 32468 7832
rect 10828 7708 10868 7748
rect 13132 7708 13172 7748
rect 14188 7708 14228 7748
rect 15340 7708 15380 7748
rect 16012 7708 16052 7748
rect 16300 7708 16340 7748
rect 16972 7708 17012 7748
rect 19372 7708 19412 7748
rect 19948 7708 19988 7748
rect 21580 7708 21620 7748
rect 22156 7708 22196 7748
rect 25900 7708 25940 7748
rect 26284 7708 26324 7748
rect 28204 7708 28244 7748
rect 29068 7708 29108 7748
rect 29452 7708 29492 7748
rect 32044 7708 32084 7748
rect 33772 7708 33812 7748
rect 10348 7624 10388 7664
rect 11020 7624 11060 7664
rect 39628 7792 39668 7832
rect 40204 7792 40244 7832
rect 41644 7876 41684 7916
rect 42124 7792 42164 7832
rect 41836 7708 41876 7748
rect 18988 7624 19028 7664
rect 20716 7624 20756 7664
rect 28300 7624 28340 7664
rect 33964 7624 34004 7664
rect 34156 7624 34196 7664
rect 39052 7624 39092 7664
rect 46252 7624 46292 7664
rect 10252 7540 10292 7580
rect 18124 7540 18164 7580
rect 1228 7456 1268 7496
rect 6988 7456 7028 7496
rect 8044 7456 8084 7496
rect 9772 7456 9812 7496
rect 10540 7456 10580 7496
rect 6028 7372 6068 7412
rect 7660 7372 7700 7412
rect 8716 7372 8756 7412
rect 2668 7288 2708 7328
rect 8140 7288 8180 7328
rect 9196 7372 9236 7412
rect 19180 7540 19220 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 21772 7540 21812 7580
rect 29932 7540 29972 7580
rect 30220 7540 30260 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 21196 7456 21236 7496
rect 13420 7372 13460 7412
rect 17644 7372 17684 7412
rect 19756 7372 19796 7412
rect 20236 7372 20276 7412
rect 21772 7372 21812 7412
rect 9580 7288 9620 7328
rect 9964 7288 10004 7328
rect 3436 7235 3476 7244
rect 3436 7204 3476 7235
rect 4396 7204 4436 7244
rect 5548 7204 5588 7244
rect 6796 7204 6836 7244
rect 7180 7204 7220 7244
rect 7468 7204 7508 7244
rect 7660 7204 7691 7244
rect 7691 7204 7700 7244
rect 8812 7204 8852 7244
rect 6412 7120 6452 7160
rect 7276 7120 7299 7160
rect 7299 7120 7316 7160
rect 8044 7120 8084 7160
rect 8428 7120 8468 7160
rect 4300 7036 4340 7076
rect 5836 7036 5876 7076
rect 7180 7036 7220 7076
rect 7756 7036 7796 7076
rect 1612 6952 1652 6992
rect 4780 6952 4820 6992
rect 6124 6952 6164 6992
rect 7948 6952 7988 6992
rect 9868 7204 9908 7244
rect 14284 7288 14324 7328
rect 11212 7204 11252 7244
rect 11692 7204 11732 7244
rect 11884 7204 11924 7244
rect 13420 7204 13460 7244
rect 14572 7204 14612 7244
rect 14956 7235 14996 7244
rect 14956 7204 14996 7235
rect 16396 7204 16436 7244
rect 9196 7120 9236 7160
rect 9484 7120 9524 7160
rect 9676 7120 9716 7160
rect 10156 7120 10196 7160
rect 10732 7120 10772 7160
rect 17644 7204 17684 7244
rect 18508 7204 18548 7244
rect 18700 7204 18740 7244
rect 21292 7288 21332 7328
rect 25804 7456 25844 7496
rect 34252 7456 34292 7496
rect 43372 7456 43412 7496
rect 46252 7456 46292 7496
rect 22348 7372 22388 7412
rect 23788 7372 23828 7412
rect 24460 7372 24500 7412
rect 28204 7372 28244 7412
rect 30316 7372 30356 7412
rect 31948 7372 31988 7412
rect 33772 7372 33812 7412
rect 22636 7288 22676 7328
rect 32908 7288 32948 7328
rect 20236 7204 20276 7244
rect 11020 7120 11060 7160
rect 11308 7120 11348 7160
rect 14860 7120 14900 7160
rect 18412 7120 18452 7160
rect 12844 7036 12884 7076
rect 15148 7036 15188 7076
rect 9676 6952 9716 6992
rect 11692 6952 11732 6992
rect 13036 6952 13076 6992
rect 14380 6952 14420 6992
rect 16204 6952 16244 6992
rect 17452 6952 17492 6992
rect 7276 6868 7316 6908
rect 9484 6868 9524 6908
rect 10732 6868 10772 6908
rect 11500 6868 11540 6908
rect 21484 7204 21524 7244
rect 22060 7204 22100 7244
rect 22444 7204 22484 7244
rect 22732 7204 22772 7244
rect 23500 7235 23540 7244
rect 23500 7204 23540 7235
rect 24556 7204 24596 7244
rect 27340 7235 27380 7244
rect 27340 7204 27380 7235
rect 28780 7204 28820 7244
rect 30028 7235 30068 7244
rect 30028 7204 30068 7235
rect 30508 7204 30548 7244
rect 37132 7372 37172 7412
rect 44812 7372 44852 7412
rect 33580 7288 33620 7328
rect 39052 7288 39092 7328
rect 33868 7204 33908 7244
rect 34924 7204 34964 7244
rect 36940 7204 36980 7244
rect 37516 7204 37556 7244
rect 38380 7204 38420 7244
rect 40492 7204 40532 7244
rect 41356 7235 41396 7244
rect 41356 7204 41396 7235
rect 41836 7235 41876 7244
rect 41836 7204 41876 7235
rect 20140 7120 20180 7160
rect 22252 7120 22292 7160
rect 23404 7120 23444 7160
rect 25708 7120 25748 7160
rect 26188 7120 26228 7160
rect 28684 7120 28724 7160
rect 32236 7120 32276 7160
rect 34540 7120 34580 7160
rect 37132 7120 37172 7160
rect 39148 7120 39188 7160
rect 40396 7120 40436 7160
rect 40588 7120 40628 7160
rect 43372 7120 43412 7160
rect 43756 7120 43796 7160
rect 44044 7120 44084 7160
rect 44908 7120 44948 7160
rect 21484 7036 21524 7076
rect 23212 7036 23252 7076
rect 30796 7036 30836 7076
rect 32428 7036 32468 7076
rect 32812 7036 32852 7076
rect 33772 7036 33812 7076
rect 39820 7036 39860 7076
rect 43852 7036 43892 7076
rect 44428 7036 44468 7076
rect 17836 6952 17876 6992
rect 19660 6952 19700 6992
rect 26860 6952 26900 6992
rect 30412 6952 30452 6992
rect 30604 6952 30644 6992
rect 36748 6952 36788 6992
rect 37132 6952 37172 6992
rect 38092 6952 38132 6992
rect 39244 6952 39284 6992
rect 32236 6868 32276 6908
rect 34924 6868 34964 6908
rect 35692 6868 35732 6908
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4684 6784 4724 6824
rect 9868 6784 9908 6824
rect 18508 6784 18548 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 19756 6784 19796 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 3436 6700 3476 6740
rect 7756 6700 7796 6740
rect 12844 6700 12884 6740
rect 14860 6700 14900 6740
rect 22924 6700 22964 6740
rect 27436 6700 27476 6740
rect 31948 6700 31988 6740
rect 6124 6616 6164 6656
rect 8812 6616 8852 6656
rect 10252 6616 10292 6656
rect 10732 6616 10772 6656
rect 3724 6532 3764 6572
rect 4684 6532 4724 6572
rect 9196 6532 9236 6572
rect 4492 6448 4532 6488
rect 5548 6448 5588 6488
rect 6988 6448 7028 6488
rect 7948 6448 7988 6488
rect 2572 6364 2612 6404
rect 4300 6364 4340 6404
rect 4876 6364 4916 6404
rect 5452 6364 5492 6404
rect 6028 6364 6068 6404
rect 6412 6364 6452 6404
rect 7084 6364 7115 6404
rect 7115 6364 7124 6404
rect 9292 6448 9332 6488
rect 9676 6532 9716 6572
rect 10348 6448 10388 6488
rect 11020 6448 11060 6488
rect 8236 6364 8273 6404
rect 8273 6364 8276 6404
rect 8716 6364 8756 6404
rect 9964 6364 10004 6404
rect 5740 6280 5780 6320
rect 7180 6280 7220 6320
rect 8044 6280 8084 6320
rect 9484 6280 9524 6320
rect 11404 6364 11444 6404
rect 10348 6280 10388 6320
rect 4204 6196 4244 6236
rect 5356 6196 5396 6236
rect 6028 6196 6068 6236
rect 8620 6196 8660 6236
rect 10060 6196 10100 6236
rect 10252 6196 10292 6236
rect 11212 6196 11252 6236
rect 46252 6952 46292 6992
rect 37228 6868 37268 6908
rect 40300 6784 40340 6824
rect 43468 6784 43508 6824
rect 46252 6784 46292 6824
rect 43564 6700 43604 6740
rect 18700 6616 18740 6656
rect 23308 6616 23348 6656
rect 23500 6616 23540 6656
rect 25804 6616 25844 6656
rect 28012 6616 28052 6656
rect 30028 6616 30068 6656
rect 31372 6616 31412 6656
rect 32428 6616 32468 6656
rect 34348 6616 34388 6656
rect 37132 6616 37172 6656
rect 40396 6616 40436 6656
rect 44236 6616 44276 6656
rect 14476 6532 14516 6572
rect 20908 6532 20948 6572
rect 21388 6532 21428 6572
rect 40012 6532 40052 6572
rect 40684 6532 40724 6572
rect 16588 6448 16628 6488
rect 17068 6448 17108 6488
rect 17452 6448 17492 6488
rect 17836 6448 17876 6488
rect 18124 6448 18164 6488
rect 18508 6448 18548 6488
rect 20716 6448 20756 6488
rect 22060 6448 22100 6488
rect 22348 6448 22388 6488
rect 25708 6448 25748 6488
rect 28780 6448 28820 6488
rect 29644 6448 29684 6488
rect 30508 6448 30548 6488
rect 33196 6448 33236 6488
rect 34540 6448 34580 6488
rect 38380 6448 38420 6488
rect 44140 6448 44180 6488
rect 44332 6448 44372 6488
rect 44716 6448 44756 6488
rect 11884 6364 11924 6404
rect 13420 6364 13460 6404
rect 14572 6364 14612 6404
rect 16396 6364 16436 6404
rect 18604 6364 18644 6404
rect 19276 6364 19316 6404
rect 19660 6364 19700 6404
rect 19852 6364 19892 6404
rect 22924 6364 22964 6404
rect 26380 6364 26420 6404
rect 27340 6364 27380 6404
rect 28204 6364 28244 6404
rect 15820 6280 15860 6320
rect 17740 6280 17780 6320
rect 29740 6364 29780 6404
rect 30028 6364 30068 6404
rect 31948 6364 31988 6404
rect 33484 6364 33524 6404
rect 34828 6364 34868 6404
rect 35404 6364 35444 6404
rect 36844 6364 36884 6404
rect 20044 6280 20084 6320
rect 21196 6280 21236 6320
rect 21484 6280 21524 6320
rect 21964 6280 22004 6320
rect 25036 6280 25076 6320
rect 26860 6280 26900 6320
rect 28300 6280 28340 6320
rect 30316 6280 30356 6320
rect 11596 6196 11636 6236
rect 14860 6196 14900 6236
rect 20524 6196 20564 6236
rect 26284 6196 26324 6236
rect 28492 6196 28532 6236
rect 30124 6196 30164 6236
rect 4396 6112 4436 6152
rect 6124 6112 6164 6152
rect 12844 6112 12884 6152
rect 18508 6112 18548 6152
rect 24364 6112 24404 6152
rect 30700 6196 30740 6236
rect 32140 6196 32180 6236
rect 33004 6196 33044 6236
rect 35596 6196 35636 6236
rect 36076 6196 36116 6236
rect 38956 6364 38996 6404
rect 40204 6364 40244 6404
rect 37612 6280 37652 6320
rect 41068 6196 41108 6236
rect 32908 6112 32948 6152
rect 40300 6112 40340 6152
rect 43948 6112 43988 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 7276 6028 7316 6068
rect 8236 6028 8276 6068
rect 8620 6028 8660 6068
rect 14092 6028 14132 6068
rect 18412 6028 18452 6068
rect 19756 6028 19796 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 22060 6028 22100 6068
rect 24172 6028 24212 6068
rect 27436 6028 27476 6068
rect 27724 6028 27764 6068
rect 28780 6028 28820 6068
rect 30124 6028 30164 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 17932 5944 17972 5984
rect 32812 5944 32852 5984
rect 33772 5944 33812 5984
rect 34732 5944 34772 5984
rect 38764 5944 38804 5984
rect 2092 5860 2132 5900
rect 4492 5860 4532 5900
rect 5836 5860 5876 5900
rect 6028 5860 6068 5900
rect 9292 5860 9332 5900
rect 17068 5860 17108 5900
rect 1612 5776 1652 5816
rect 5932 5776 5972 5816
rect 17644 5860 17684 5900
rect 23212 5860 23252 5900
rect 31948 5860 31988 5900
rect 33004 5860 33044 5900
rect 34540 5860 34580 5900
rect 35692 5860 35732 5900
rect 7084 5776 7124 5816
rect 10348 5776 10388 5816
rect 11308 5776 11348 5816
rect 13228 5776 13268 5816
rect 20236 5776 20276 5816
rect 20428 5776 20468 5816
rect 23884 5776 23924 5816
rect 24172 5776 24212 5816
rect 25804 5776 25844 5816
rect 29740 5776 29780 5816
rect 30700 5776 30740 5816
rect 32140 5776 32180 5816
rect 36172 5776 36212 5816
rect 36460 5776 36500 5816
rect 36652 5776 36692 5816
rect 2284 5692 2324 5732
rect 3532 5723 3572 5732
rect 3532 5692 3572 5723
rect 4108 5692 4148 5732
rect 4396 5692 4436 5732
rect 76 5608 116 5648
rect 5644 5692 5684 5732
rect 7180 5692 7211 5732
rect 7211 5692 7220 5732
rect 7468 5692 7508 5732
rect 2188 5524 2228 5564
rect 4300 5524 4340 5564
rect 76 5440 116 5480
rect 5836 5608 5876 5648
rect 6220 5608 6260 5648
rect 2380 5440 2420 5480
rect 2572 5440 2612 5480
rect 5452 5440 5492 5480
rect 7852 5692 7892 5732
rect 8428 5692 8468 5732
rect 8721 5692 8761 5732
rect 9196 5692 9236 5732
rect 10444 5692 10484 5732
rect 11596 5692 11636 5732
rect 11884 5723 11924 5732
rect 11884 5692 11924 5723
rect 12940 5692 12980 5732
rect 13612 5692 13652 5732
rect 6604 5608 6644 5648
rect 8812 5608 8852 5648
rect 9676 5608 9716 5648
rect 10348 5608 10388 5648
rect 11020 5608 11060 5648
rect 14092 5608 14132 5648
rect 7660 5524 7700 5564
rect 9580 5524 9620 5564
rect 9772 5524 9812 5564
rect 14860 5692 14900 5732
rect 15820 5692 15860 5732
rect 15148 5608 15188 5648
rect 16492 5692 16532 5732
rect 17164 5692 17204 5732
rect 17548 5692 17588 5732
rect 15436 5608 15476 5648
rect 18508 5692 18548 5732
rect 18892 5692 18932 5732
rect 20812 5692 20852 5732
rect 22156 5723 22196 5732
rect 22156 5692 22196 5723
rect 23212 5692 23252 5732
rect 24076 5692 24116 5732
rect 24364 5692 24404 5732
rect 20908 5608 20948 5648
rect 21196 5608 21236 5648
rect 25516 5692 25556 5732
rect 25996 5692 26036 5732
rect 22252 5608 22292 5648
rect 20140 5524 20180 5564
rect 20332 5524 20372 5564
rect 26764 5692 26804 5732
rect 25132 5608 25172 5648
rect 25708 5608 25748 5648
rect 30316 5692 30356 5732
rect 30892 5692 30932 5732
rect 31756 5692 31796 5732
rect 34060 5692 34100 5732
rect 34348 5692 34388 5732
rect 34636 5692 34676 5732
rect 27148 5608 27188 5648
rect 27724 5608 27764 5648
rect 28108 5608 28148 5648
rect 29260 5608 29300 5648
rect 30508 5608 30548 5648
rect 31276 5608 31316 5648
rect 33100 5608 33140 5648
rect 24460 5524 24500 5564
rect 25420 5524 25460 5564
rect 29548 5524 29588 5564
rect 7180 5440 7220 5480
rect 8620 5440 8660 5480
rect 9004 5440 9044 5480
rect 9388 5440 9428 5480
rect 10252 5440 10292 5480
rect 11116 5440 11156 5480
rect 11404 5440 11444 5480
rect 14572 5440 14612 5480
rect 18604 5440 18644 5480
rect 20428 5440 20468 5480
rect 23788 5440 23828 5480
rect 28396 5440 28436 5480
rect 29740 5440 29780 5480
rect 5644 5356 5684 5396
rect 18508 5356 18548 5396
rect 20140 5356 20180 5396
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 6892 5272 6932 5312
rect 13420 5272 13460 5312
rect 14284 5272 14324 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 19372 5272 19412 5312
rect 3244 5104 3284 5144
rect 5644 5104 5684 5144
rect 6604 5104 6644 5144
rect 7372 5188 7412 5228
rect 16396 5188 16436 5228
rect 20812 5188 20852 5228
rect 8524 5104 8564 5144
rect 11596 5104 11636 5144
rect 2380 5020 2420 5060
rect 3916 5020 3956 5060
rect 4108 5020 4148 5060
rect 7180 5020 7220 5060
rect 8044 5020 8084 5060
rect 8236 5020 8276 5060
rect 76 4936 116 4976
rect 2188 4936 2228 4976
rect 6028 4936 6068 4976
rect 2284 4852 2324 4892
rect 3724 4852 3764 4892
rect 76 4768 116 4808
rect 4204 4768 4244 4808
rect 5452 4852 5492 4892
rect 5740 4852 5780 4892
rect 6124 4852 6164 4892
rect 6220 4768 6260 4808
rect 2860 4684 2900 4724
rect 5740 4684 5780 4724
rect 6892 4852 6932 4892
rect 7276 4852 7316 4892
rect 7756 4852 7787 4892
rect 7787 4852 7796 4892
rect 9292 4936 9332 4976
rect 10636 5020 10676 5060
rect 11020 5020 11060 5060
rect 12460 5104 12500 5144
rect 17164 5104 17204 5144
rect 13036 5020 13076 5060
rect 18220 5020 18260 5060
rect 8524 4852 8564 4892
rect 9196 4852 9236 4892
rect 10252 4852 10292 4892
rect 10444 4852 10484 4892
rect 11116 4852 11156 4892
rect 11500 4852 11540 4892
rect 8716 4768 8756 4808
rect 9388 4768 9428 4808
rect 10636 4768 10676 4808
rect 12460 4936 12500 4976
rect 13324 4936 13364 4976
rect 12748 4852 12788 4892
rect 13036 4852 13076 4892
rect 13708 4852 13748 4892
rect 12652 4768 12692 4808
rect 15052 4936 15092 4976
rect 15820 4936 15860 4976
rect 16492 4936 16532 4976
rect 14284 4852 14324 4892
rect 14668 4852 14708 4892
rect 15436 4852 15476 4892
rect 16300 4852 16340 4892
rect 16684 4852 16724 4892
rect 18604 5104 18644 5144
rect 18796 5104 18836 5144
rect 21004 5104 21044 5144
rect 21772 5356 21812 5396
rect 22252 5356 22292 5396
rect 27052 5356 27092 5396
rect 27820 5356 27860 5396
rect 27916 5272 27956 5312
rect 21964 5188 22004 5228
rect 28876 5188 28916 5228
rect 26188 5104 26228 5144
rect 27148 5104 27188 5144
rect 30988 5524 31028 5564
rect 32716 5524 32756 5564
rect 33196 5524 33236 5564
rect 33676 5524 33716 5564
rect 30508 5440 30548 5480
rect 33004 5440 33044 5480
rect 35596 5692 35636 5732
rect 36076 5692 36116 5732
rect 36364 5692 36395 5732
rect 36395 5692 36404 5732
rect 36940 5692 36980 5732
rect 38188 5723 38228 5732
rect 38188 5692 38228 5723
rect 40300 5692 40340 5732
rect 41356 5692 41396 5732
rect 33868 5608 33908 5648
rect 38956 5608 38996 5648
rect 40684 5608 40724 5648
rect 44524 5608 44564 5648
rect 44908 5608 44948 5648
rect 36364 5524 36404 5564
rect 34060 5440 34100 5480
rect 37516 5440 37556 5480
rect 38380 5440 38420 5480
rect 38572 5440 38612 5480
rect 43084 5356 43124 5396
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 30316 5104 30356 5144
rect 31372 5104 31412 5144
rect 31564 5104 31604 5144
rect 32236 5104 32276 5144
rect 32716 5104 32756 5144
rect 33580 5104 33620 5144
rect 36460 5104 36500 5144
rect 38380 5104 38420 5144
rect 39148 5104 39188 5144
rect 20524 5020 20564 5060
rect 21964 5020 22004 5060
rect 22444 5020 22484 5060
rect 23980 5020 24020 5060
rect 26380 5020 26420 5060
rect 28588 5020 28628 5060
rect 33388 5020 33428 5060
rect 18700 4936 18740 4976
rect 24556 4936 24596 4976
rect 27340 4936 27380 4976
rect 27532 4936 27572 4976
rect 28876 4936 28916 4976
rect 32044 4936 32084 4976
rect 32428 4936 32468 4976
rect 33004 4936 33044 4976
rect 34828 4936 34868 4976
rect 35692 4936 35732 4976
rect 36940 4936 36980 4976
rect 37900 4936 37940 4976
rect 43948 5020 43988 5060
rect 40972 4936 41012 4976
rect 43564 4936 43604 4976
rect 18796 4852 18836 4892
rect 19564 4852 19604 4892
rect 20332 4852 20372 4892
rect 21676 4852 21716 4892
rect 21964 4852 22004 4892
rect 22636 4852 22676 4892
rect 23980 4852 24020 4892
rect 25132 4852 25172 4892
rect 27628 4852 27668 4892
rect 28108 4852 28148 4892
rect 28684 4852 28724 4892
rect 29356 4852 29396 4892
rect 30028 4852 30068 4892
rect 31564 4852 31604 4892
rect 31756 4852 31796 4892
rect 34252 4852 34292 4892
rect 35596 4852 35604 4892
rect 35604 4852 35636 4892
rect 35788 4852 35828 4892
rect 35980 4852 36020 4892
rect 36460 4852 36500 4892
rect 37516 4852 37556 4892
rect 37996 4852 38036 4892
rect 40300 4852 40331 4892
rect 40331 4852 40340 4892
rect 19948 4768 19988 4808
rect 20428 4768 20468 4808
rect 20908 4768 20948 4808
rect 22732 4768 22772 4808
rect 7180 4684 7220 4724
rect 14284 4684 14324 4724
rect 16108 4684 16148 4724
rect 16588 4684 16628 4724
rect 20044 4684 20084 4724
rect 25420 4684 25460 4724
rect 25996 4684 26036 4724
rect 4012 4600 4052 4640
rect 6988 4600 7028 4640
rect 18604 4600 18644 4640
rect 21292 4600 21332 4640
rect 21868 4600 21908 4640
rect 26188 4600 26228 4640
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 10732 4516 10772 4556
rect 13420 4516 13460 4556
rect 17452 4516 17492 4556
rect 19660 4516 19700 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 20524 4516 20564 4556
rect 25516 4516 25556 4556
rect 26092 4516 26132 4556
rect 27340 4516 27380 4556
rect 32332 4768 32372 4808
rect 35692 4768 35732 4808
rect 37900 4768 37940 4808
rect 39916 4768 39947 4808
rect 39947 4768 39956 4808
rect 28876 4684 28916 4724
rect 30220 4684 30260 4724
rect 29260 4600 29300 4640
rect 32428 4600 32468 4640
rect 34348 4600 34388 4640
rect 29548 4516 29588 4556
rect 33964 4516 34004 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 35884 4516 35924 4556
rect 44620 4516 44660 4556
rect 7756 4432 7796 4472
rect 9196 4432 9236 4472
rect 9580 4432 9620 4472
rect 13324 4432 13364 4472
rect 16684 4432 16724 4472
rect 28684 4432 28724 4472
rect 31180 4432 31220 4472
rect 40300 4432 40340 4472
rect 5548 4348 5588 4388
rect 5836 4348 5867 4388
rect 5867 4348 5876 4388
rect 6988 4348 7028 4388
rect 7276 4348 7316 4388
rect 7660 4348 7700 4388
rect 10732 4348 10772 4388
rect 11308 4348 11348 4388
rect 13228 4348 13268 4388
rect 14668 4348 14708 4388
rect 16300 4348 16340 4388
rect 18220 4348 18260 4388
rect 22156 4348 22196 4388
rect 23212 4348 23252 4388
rect 25708 4348 25748 4388
rect 26380 4348 26420 4388
rect 27052 4348 27092 4388
rect 28108 4348 28148 4388
rect 28780 4348 28820 4388
rect 29740 4348 29780 4388
rect 30028 4348 30068 4388
rect 31852 4348 31892 4388
rect 32428 4348 32468 4388
rect 33580 4348 33620 4388
rect 36076 4348 36116 4388
rect 37900 4348 37940 4388
rect 38092 4348 38132 4388
rect 2476 4264 2516 4304
rect 5740 4264 5780 4304
rect 5932 4264 5972 4304
rect 6604 4264 6644 4304
rect 12940 4264 12980 4304
rect 14284 4264 14324 4304
rect 15148 4264 15188 4304
rect 16588 4264 16628 4304
rect 3052 4180 3092 4220
rect 3532 4180 3572 4220
rect 4108 4180 4148 4220
rect 4492 4180 4532 4220
rect 5356 4180 5396 4220
rect 5836 4180 5876 4220
rect 6028 4180 6057 4220
rect 6057 4180 6068 4220
rect 7180 4180 7220 4220
rect 7756 4180 7796 4220
rect 8044 4180 8084 4220
rect 8428 4180 8468 4220
rect 2668 4096 2708 4136
rect 6796 4096 6836 4136
rect 6988 4096 7028 4136
rect 2380 3928 2420 3968
rect 4300 3928 4340 3968
rect 9100 4211 9140 4220
rect 9100 4180 9140 4211
rect 9484 4180 9524 4220
rect 9772 4180 9812 4220
rect 10636 4211 10676 4220
rect 10636 4180 10676 4211
rect 11116 4211 11156 4220
rect 11116 4180 11156 4211
rect 12844 4180 12884 4220
rect 13324 4180 13364 4220
rect 7660 4096 7700 4136
rect 8236 4096 8276 4136
rect 14860 4180 14900 4220
rect 16492 4180 16532 4220
rect 17548 4180 17588 4220
rect 18700 4180 18740 4220
rect 19276 4180 19316 4220
rect 19756 4180 19796 4220
rect 19948 4180 19988 4220
rect 8044 4012 8084 4052
rect 8812 4012 8852 4052
rect 10252 4096 10292 4136
rect 11692 4096 11732 4136
rect 11980 4096 12020 4136
rect 14764 4096 14804 4136
rect 19468 4096 19508 4136
rect 12364 4012 12404 4052
rect 5740 3928 5780 3968
rect 7564 3928 7604 3968
rect 8428 3928 8468 3968
rect 10252 3928 10292 3968
rect 12172 3928 12212 3968
rect 20332 4264 20372 4304
rect 21004 4264 21044 4304
rect 27340 4264 27380 4304
rect 29644 4264 29684 4304
rect 31276 4264 31316 4304
rect 37708 4264 37748 4304
rect 40012 4264 40052 4304
rect 20620 4180 20660 4220
rect 21196 4180 21236 4220
rect 21868 4211 21908 4220
rect 21868 4180 21908 4211
rect 22444 4180 22484 4220
rect 23404 4180 23444 4220
rect 23884 4180 23924 4220
rect 26284 4180 26324 4220
rect 26668 4180 26708 4220
rect 22348 4096 22388 4136
rect 24268 4096 24308 4136
rect 24844 4096 24884 4136
rect 25036 4096 25076 4136
rect 25612 4096 25652 4136
rect 25900 4096 25940 4136
rect 27052 4096 27092 4136
rect 12940 4012 12980 4052
rect 20332 4012 20372 4052
rect 21964 4012 22004 4052
rect 13036 3928 13076 3968
rect 15052 3928 15092 3968
rect 19468 3928 19508 3968
rect 20236 3928 20276 3968
rect 21196 3928 21236 3968
rect 22828 3928 22868 3968
rect 23020 3928 23060 3968
rect 23500 3928 23540 3968
rect 23884 3928 23924 3968
rect 24460 3928 24500 3968
rect 27244 4180 27284 4220
rect 28588 4180 28628 4220
rect 29932 4180 29972 4220
rect 32044 4180 32084 4220
rect 30508 4096 30548 4136
rect 31276 4096 31316 4136
rect 32428 4180 32468 4220
rect 33868 4180 33908 4220
rect 34252 4180 34292 4220
rect 34636 4180 34676 4220
rect 31852 4096 31892 4136
rect 25228 4012 25268 4052
rect 26572 4012 26612 4052
rect 4492 3844 4532 3884
rect 5644 3844 5684 3884
rect 5836 3844 5876 3884
rect 7372 3844 7412 3884
rect 9196 3844 9236 3884
rect 12268 3844 12308 3884
rect 13708 3844 13748 3884
rect 15820 3844 15860 3884
rect 25036 3844 25076 3884
rect 27148 3928 27188 3968
rect 31564 3928 31604 3968
rect 32332 3844 32372 3884
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 11212 3760 11252 3800
rect 14956 3760 14996 3800
rect 16876 3760 16916 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 21004 3760 21044 3800
rect 25228 3760 25268 3800
rect 28684 3760 28724 3800
rect 30220 3760 30260 3800
rect 5164 3676 5204 3716
rect 14860 3676 14900 3716
rect 21196 3676 21236 3716
rect 26092 3676 26132 3716
rect 26476 3676 26516 3716
rect 27052 3676 27092 3716
rect 29836 3676 29876 3716
rect 30508 3676 30548 3716
rect 32332 3676 32372 3716
rect 35692 4180 35732 4220
rect 36460 4180 36500 4220
rect 37612 4180 37652 4220
rect 43276 4180 43316 4220
rect 33004 4096 33044 4136
rect 33580 4096 33620 4136
rect 34348 4096 34388 4136
rect 38668 4096 38708 4136
rect 38860 4096 38900 4136
rect 39628 4096 39668 4136
rect 32908 4012 32948 4052
rect 34540 4012 34580 4052
rect 40972 4012 41012 4052
rect 34444 3928 34484 3968
rect 35788 3928 35828 3968
rect 41644 3928 41684 3968
rect 35116 3844 35156 3884
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 32908 3676 32948 3716
rect 34540 3676 34580 3716
rect 40492 3676 40532 3716
rect 3148 3592 3188 3632
rect 7276 3592 7316 3632
rect 8620 3592 8660 3632
rect 9196 3592 9236 3632
rect 16588 3592 16628 3632
rect 18892 3592 18932 3632
rect 19180 3592 19220 3632
rect 19564 3592 19604 3632
rect 26572 3592 26612 3632
rect 26956 3592 26996 3632
rect 28204 3592 28244 3632
rect 33580 3592 33620 3632
rect 36556 3592 36596 3632
rect 37420 3592 37460 3632
rect 41068 3592 41108 3632
rect 1132 3508 1172 3548
rect 6316 3508 6356 3548
rect 7372 3508 7412 3548
rect 14668 3508 14708 3548
rect 18220 3508 18260 3548
rect 20236 3508 20276 3548
rect 24364 3508 24404 3548
rect 24556 3508 24596 3548
rect 30124 3508 30164 3548
rect 1420 3424 1460 3464
rect 1996 3424 2036 3464
rect 2956 3424 2996 3464
rect 4204 3424 4244 3464
rect 6220 3424 6260 3464
rect 7468 3424 7508 3464
rect 10732 3424 10772 3464
rect 11020 3424 11060 3464
rect 3052 3340 3092 3380
rect 4300 3340 4340 3380
rect 5548 3340 5588 3380
rect 6316 3340 6356 3380
rect 6796 3340 6836 3380
rect 2092 3256 2132 3296
rect 4396 3256 4436 3296
rect 5740 3256 5780 3296
rect 6124 3256 6164 3296
rect 7180 3340 7220 3380
rect 7564 3340 7604 3380
rect 7852 3340 7892 3380
rect 8812 3340 8852 3380
rect 8620 3256 8660 3296
rect 2572 3172 2612 3212
rect 6508 3172 6548 3212
rect 8812 3172 8852 3212
rect 6796 3088 6836 3128
rect 12076 3424 12116 3464
rect 13900 3424 13940 3464
rect 14476 3424 14516 3464
rect 14764 3424 14804 3464
rect 15052 3424 15092 3464
rect 16108 3424 16148 3464
rect 17356 3424 17396 3464
rect 17932 3424 17972 3464
rect 18508 3424 18548 3464
rect 18892 3424 18932 3464
rect 20140 3424 20180 3464
rect 10252 3340 10292 3380
rect 10636 3340 10676 3380
rect 10828 3340 10868 3380
rect 11500 3340 11540 3380
rect 9676 3256 9707 3296
rect 9707 3256 9716 3296
rect 35116 3508 35156 3548
rect 23692 3424 23732 3464
rect 24748 3424 24788 3464
rect 26668 3424 26708 3464
rect 27244 3424 27284 3464
rect 29164 3424 29204 3464
rect 30316 3424 30356 3464
rect 34540 3424 34580 3464
rect 35596 3424 35636 3464
rect 36076 3424 36116 3464
rect 36268 3424 36308 3464
rect 40300 3424 40340 3464
rect 12556 3340 12596 3380
rect 12844 3340 12884 3380
rect 13708 3340 13748 3380
rect 16588 3340 16628 3380
rect 17836 3340 17876 3380
rect 18988 3340 19028 3380
rect 20524 3340 20564 3380
rect 21964 3340 22004 3380
rect 23212 3340 23252 3380
rect 24844 3340 24884 3380
rect 25612 3340 25652 3380
rect 27052 3340 27092 3380
rect 28204 3340 28244 3380
rect 28780 3340 28820 3380
rect 29260 3340 29300 3380
rect 30700 3340 30740 3380
rect 32332 3340 32372 3380
rect 35692 3340 35732 3380
rect 37900 3340 37940 3380
rect 38956 3340 38996 3380
rect 39244 3340 39284 3380
rect 40492 3340 40532 3380
rect 40780 3340 40820 3380
rect 40972 3340 41012 3380
rect 41740 3340 41780 3380
rect 12076 3256 12116 3296
rect 14476 3256 14516 3296
rect 19948 3256 19988 3296
rect 21484 3256 21524 3296
rect 22828 3256 22868 3296
rect 24460 3256 24500 3296
rect 36268 3256 36308 3296
rect 36460 3256 36500 3296
rect 36940 3256 36980 3296
rect 39916 3256 39956 3296
rect 9388 3172 9428 3212
rect 9964 3172 10004 3212
rect 13516 3172 13556 3212
rect 13900 3172 13940 3212
rect 14572 3172 14612 3212
rect 11308 3088 11348 3128
rect 14860 3088 14900 3128
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 7756 3004 7796 3044
rect 17164 3172 17204 3212
rect 17548 3172 17588 3212
rect 17836 3172 17876 3212
rect 18508 3172 18548 3212
rect 18796 3172 18836 3212
rect 21868 3172 21908 3212
rect 22156 3172 22196 3212
rect 24268 3172 24308 3212
rect 25708 3172 25748 3212
rect 26284 3172 26324 3212
rect 26476 3172 26516 3212
rect 27436 3172 27476 3212
rect 30508 3172 30548 3212
rect 30988 3172 31028 3212
rect 34348 3172 34388 3212
rect 35116 3172 35156 3212
rect 35884 3172 35924 3212
rect 18700 3088 18740 3128
rect 22540 3088 22580 3128
rect 25900 3088 25940 3128
rect 31276 3088 31316 3128
rect 18412 3004 18452 3044
rect 19756 3004 19796 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 22156 3004 22196 3044
rect 24364 3004 24404 3044
rect 29356 3004 29396 3044
rect 30892 3004 30932 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 35596 3004 35636 3044
rect 35884 3004 35924 3044
rect 2668 2920 2708 2960
rect 5452 2920 5492 2960
rect 5932 2920 5972 2960
rect 11692 2920 11732 2960
rect 16492 2920 16532 2960
rect 17548 2920 17588 2960
rect 18604 2920 18644 2960
rect 18892 2920 18932 2960
rect 21964 2920 22004 2960
rect 26476 2920 26516 2960
rect 29260 2920 29300 2960
rect 30028 2920 30068 2960
rect 31660 2920 31700 2960
rect 33004 2920 33044 2960
rect 34924 2920 34964 2960
rect 35692 2920 35732 2960
rect 38668 2920 38708 2960
rect 2380 2836 2420 2876
rect 1996 2752 2036 2792
rect 2860 2752 2900 2792
rect 1516 2500 1556 2540
rect 3436 2836 3476 2876
rect 4204 2836 4244 2876
rect 6220 2836 6260 2876
rect 6700 2836 6731 2876
rect 6731 2836 6740 2876
rect 10252 2836 10292 2876
rect 12652 2836 12692 2876
rect 13708 2836 13748 2876
rect 15436 2836 15476 2876
rect 3340 2752 3380 2792
rect 4108 2752 4148 2792
rect 7276 2752 7316 2792
rect 9484 2752 9524 2792
rect 11500 2752 11540 2792
rect 12556 2752 12596 2792
rect 13420 2752 13460 2792
rect 14284 2752 14324 2792
rect 3436 2668 3476 2708
rect 4972 2668 5012 2708
rect 5452 2668 5492 2708
rect 6124 2668 6164 2708
rect 6796 2668 6836 2708
rect 7084 2668 7124 2708
rect 7372 2668 7412 2708
rect 9004 2668 9044 2708
rect 10924 2668 10964 2708
rect 12268 2668 12296 2687
rect 12296 2668 12308 2687
rect 2476 2584 2516 2624
rect 3244 2584 3284 2624
rect 4204 2584 4244 2624
rect 4396 2584 4436 2624
rect 6508 2584 6539 2624
rect 6539 2584 6548 2624
rect 6700 2584 6740 2624
rect 9676 2584 9716 2624
rect 12268 2647 12308 2668
rect 12748 2668 12788 2708
rect 15148 2699 15188 2708
rect 15148 2668 15188 2699
rect 15820 2668 15860 2708
rect 11884 2584 11924 2624
rect 2956 2500 2996 2540
rect 3148 2416 3188 2456
rect 5644 2500 5684 2540
rect 6028 2500 6068 2540
rect 7852 2500 7892 2540
rect 8140 2500 8180 2540
rect 12556 2500 12596 2540
rect 13804 2500 13844 2540
rect 15148 2500 15188 2540
rect 17836 2836 17876 2876
rect 18988 2836 19028 2876
rect 21868 2836 21908 2876
rect 22732 2836 22772 2876
rect 23692 2836 23732 2876
rect 26668 2836 26708 2876
rect 29644 2836 29684 2876
rect 33964 2836 34004 2876
rect 34348 2836 34388 2876
rect 37516 2836 37556 2876
rect 39532 2836 39572 2876
rect 41740 2836 41780 2876
rect 17452 2752 17492 2792
rect 18316 2752 18356 2792
rect 18508 2752 18548 2792
rect 17164 2699 17204 2708
rect 17164 2668 17204 2699
rect 17356 2668 17396 2708
rect 17644 2668 17684 2708
rect 17836 2668 17876 2708
rect 17548 2584 17588 2624
rect 18412 2584 18452 2624
rect 19180 2668 19220 2708
rect 22444 2752 22484 2792
rect 20236 2668 20276 2708
rect 21100 2668 21140 2708
rect 21676 2668 21716 2708
rect 21964 2668 22004 2708
rect 22924 2668 22964 2708
rect 23116 2668 23156 2708
rect 24556 2668 24596 2708
rect 24844 2668 24884 2708
rect 19276 2584 19316 2624
rect 21292 2584 21332 2624
rect 23308 2584 23348 2624
rect 25324 2668 25364 2708
rect 25612 2699 25652 2708
rect 25612 2668 25652 2699
rect 25900 2668 25940 2708
rect 28588 2752 28628 2792
rect 27628 2699 27668 2708
rect 27628 2668 27668 2699
rect 28396 2668 28436 2708
rect 29164 2699 29204 2708
rect 29164 2668 29204 2699
rect 29356 2668 29396 2708
rect 30508 2752 30548 2792
rect 31084 2752 31124 2792
rect 31660 2752 31700 2792
rect 32428 2752 32468 2792
rect 32620 2752 32660 2792
rect 37804 2752 37844 2792
rect 40780 2752 40820 2792
rect 30700 2668 30740 2708
rect 31276 2626 31316 2666
rect 32044 2668 32084 2708
rect 32908 2668 32948 2708
rect 33868 2668 33908 2708
rect 34156 2668 34196 2708
rect 34732 2668 34772 2708
rect 35116 2699 35156 2708
rect 35116 2668 35156 2699
rect 35596 2699 35636 2708
rect 35596 2668 35636 2699
rect 36268 2668 36308 2708
rect 37900 2668 37940 2708
rect 38668 2668 38708 2708
rect 38956 2668 38996 2708
rect 24748 2584 24788 2624
rect 28588 2584 28628 2624
rect 30508 2584 30548 2624
rect 33964 2584 34004 2624
rect 34348 2584 34388 2624
rect 34540 2584 34580 2624
rect 36748 2584 36788 2624
rect 40684 2584 40724 2624
rect 43084 2584 43124 2624
rect 17740 2500 17780 2540
rect 18796 2500 18836 2540
rect 22732 2500 22772 2540
rect 23116 2500 23156 2540
rect 25708 2500 25748 2540
rect 30220 2500 30260 2540
rect 5740 2416 5780 2456
rect 12268 2416 12308 2456
rect 12460 2416 12500 2456
rect 15436 2416 15476 2456
rect 18220 2416 18260 2456
rect 19276 2416 19316 2456
rect 20524 2416 20564 2456
rect 22924 2416 22964 2456
rect 24460 2416 24500 2456
rect 28780 2416 28820 2456
rect 29164 2416 29204 2456
rect 32332 2416 32372 2456
rect 34540 2416 34580 2456
rect 36076 2416 36116 2456
rect 37420 2416 37460 2456
rect 38188 2416 38228 2456
rect 3340 2332 3380 2372
rect 4396 2332 4436 2372
rect 7660 2332 7700 2372
rect 12556 2332 12596 2372
rect 13420 2332 13460 2372
rect 16204 2332 16244 2372
rect 16876 2332 16916 2372
rect 21388 2332 21428 2372
rect 21580 2332 21620 2372
rect 24076 2332 24116 2372
rect 24652 2332 24692 2372
rect 31660 2332 31700 2372
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 8812 2248 8852 2288
rect 12940 2248 12980 2288
rect 14380 2248 14420 2288
rect 17356 2248 17396 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 20908 2248 20948 2288
rect 30028 2248 30068 2288
rect 30220 2248 30260 2288
rect 31276 2248 31316 2288
rect 32908 2248 32948 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 35116 2248 35156 2288
rect 39916 2248 39956 2288
rect 3532 2164 3572 2204
rect 2284 2080 2324 2120
rect 4012 2080 4052 2120
rect 3532 1996 3572 2036
rect 11980 2164 12020 2204
rect 14476 2164 14516 2204
rect 18508 2164 18548 2204
rect 21676 2164 21716 2204
rect 23020 2164 23060 2204
rect 23212 2164 23252 2204
rect 29164 2164 29204 2204
rect 4492 2080 4532 2120
rect 6028 2080 6068 2120
rect 6412 2080 6452 2120
rect 6892 2080 6932 2120
rect 8428 2080 8468 2120
rect 8620 2080 8660 2120
rect 11788 2080 11828 2120
rect 12076 2080 12116 2120
rect 12748 2080 12788 2120
rect 14188 2080 14228 2120
rect 15148 2080 15188 2120
rect 15532 2080 15572 2120
rect 15916 2080 15956 2120
rect 16684 2080 16724 2120
rect 18604 2080 18644 2120
rect 20236 2080 20276 2120
rect 24748 2080 24788 2120
rect 25708 2080 25748 2120
rect 27244 2080 27284 2120
rect 29356 2080 29396 2120
rect 4300 1996 4340 2036
rect 6988 1996 7028 2036
rect 9772 1996 9812 2036
rect 1420 1912 1460 1952
rect 2764 1912 2804 1952
rect 3436 1912 3476 1952
rect 652 1828 692 1868
rect 4780 1912 4820 1952
rect 7180 1912 7220 1952
rect 7372 1912 7412 1952
rect 8140 1912 8180 1952
rect 12460 1912 12500 1952
rect 12844 1912 12884 1952
rect 4300 1744 4340 1784
rect 4972 1828 5012 1868
rect 4492 1660 4532 1700
rect 4204 1576 4244 1616
rect 4588 1492 4628 1532
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 8236 1828 8276 1868
rect 8620 1828 8660 1868
rect 9676 1828 9716 1868
rect 10060 1744 10100 1784
rect 10540 1828 10580 1868
rect 11884 1828 11924 1868
rect 14476 1912 14516 1952
rect 15916 1912 15956 1952
rect 17068 1912 17108 1952
rect 13804 1828 13844 1868
rect 15340 1828 15380 1868
rect 15724 1828 15764 1868
rect 16972 1828 17012 1868
rect 18220 1828 18260 1868
rect 18604 1828 18644 1868
rect 19372 1828 19412 1868
rect 21004 1996 21044 2036
rect 22348 1996 22388 2036
rect 23116 1996 23156 2036
rect 24556 1996 24596 2036
rect 25420 1996 25460 2036
rect 43468 2500 43508 2540
rect 45292 2416 45332 2456
rect 29836 2164 29876 2204
rect 37996 2164 38036 2204
rect 29932 2080 29972 2120
rect 31564 2080 31604 2120
rect 32044 2080 32084 2120
rect 29164 1996 29204 2036
rect 38764 2080 38804 2120
rect 33964 1996 34004 2036
rect 22060 1912 22100 1952
rect 24940 1912 24980 1952
rect 26956 1912 26996 1952
rect 27436 1912 27476 1952
rect 27628 1912 27668 1952
rect 29740 1912 29780 1952
rect 33004 1912 33044 1952
rect 21580 1828 21620 1868
rect 22828 1828 22868 1868
rect 23308 1828 23348 1868
rect 25708 1828 25748 1868
rect 26284 1828 26324 1868
rect 27532 1828 27572 1868
rect 27724 1828 27764 1868
rect 29932 1828 29972 1868
rect 30412 1828 30452 1868
rect 31564 1828 31604 1868
rect 32044 1828 32084 1868
rect 32428 1828 32468 1868
rect 33484 1912 33524 1952
rect 33772 1912 33812 1952
rect 34732 1996 34772 2036
rect 34540 1912 34580 1952
rect 34924 1912 34964 1952
rect 37900 1996 37940 2036
rect 41644 1996 41684 2036
rect 44620 1996 44660 2036
rect 35884 1912 35924 1952
rect 37420 1828 37460 1868
rect 38284 1912 38324 1952
rect 44140 1912 44180 1952
rect 38956 1828 38996 1868
rect 18028 1744 18068 1784
rect 20044 1744 20084 1784
rect 21484 1744 21524 1784
rect 24940 1744 24980 1784
rect 25324 1744 25364 1784
rect 29260 1744 29300 1784
rect 31276 1744 31316 1784
rect 8620 1660 8660 1700
rect 10156 1660 10196 1700
rect 12940 1660 12980 1700
rect 14572 1660 14612 1700
rect 23692 1660 23732 1700
rect 31660 1660 31700 1700
rect 32428 1660 32468 1700
rect 33196 1660 33236 1700
rect 33484 1660 33524 1700
rect 36172 1660 36212 1700
rect 39724 1660 39764 1700
rect 13036 1492 13076 1532
rect 13708 1576 13748 1616
rect 20716 1576 20756 1616
rect 21196 1576 21236 1616
rect 23308 1576 23348 1616
rect 24652 1576 24692 1616
rect 29548 1576 29588 1616
rect 32908 1576 32948 1616
rect 44620 1744 44660 1784
rect 45388 1660 45428 1700
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 24556 1492 24596 1532
rect 24844 1492 24884 1532
rect 34924 1492 34964 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 39820 1492 39860 1532
rect 652 1408 692 1448
rect 12172 1408 12212 1448
rect 14284 1408 14324 1448
rect 15916 1408 15956 1448
rect 21484 1408 21524 1448
rect 25612 1408 25652 1448
rect 27340 1408 27380 1448
rect 34156 1408 34196 1448
rect 45292 1408 45332 1448
rect 20428 1324 20468 1364
rect 27532 1324 27572 1364
rect 34252 1324 34292 1364
rect 41452 1324 41492 1364
rect 18892 1240 18932 1280
rect 1420 1072 1460 1112
rect 44620 1072 44660 1112
rect 28108 904 28148 944
rect 33484 904 33524 944
rect 10156 820 10196 860
rect 16204 820 16244 860
rect 27724 820 27764 860
rect 33196 820 33236 860
rect 1132 736 1172 776
rect 45388 736 45428 776
rect 33868 652 33908 692
rect 40108 652 40148 692
rect 4396 568 4436 608
rect 11788 568 11828 608
rect 33100 400 33140 440
rect 42604 400 42644 440
rect 32908 148 32948 188
rect 42892 148 42932 188
rect 33484 64 33524 104
rect 43660 64 43700 104
<< metal3 >>
rect 3512 12100 3592 12180
rect 4664 12100 4744 12180
rect 5816 12100 5896 12180
rect 6968 12100 7048 12180
rect 8120 12100 8200 12180
rect 9272 12100 9352 12180
rect 10424 12100 10504 12180
rect 11576 12100 11656 12180
rect 12728 12100 12808 12180
rect 13880 12100 13960 12180
rect 15032 12100 15112 12180
rect 16184 12100 16264 12180
rect 17336 12100 17416 12180
rect 18488 12100 18568 12180
rect 19640 12100 19720 12180
rect 20792 12100 20872 12180
rect 21944 12100 22024 12180
rect 23096 12100 23176 12180
rect 24248 12100 24328 12180
rect 25400 12100 25480 12180
rect 26552 12100 26632 12180
rect 27704 12100 27784 12180
rect 28856 12100 28936 12180
rect 30008 12100 30088 12180
rect 31160 12100 31240 12180
rect 32312 12100 32392 12180
rect 33464 12100 33544 12180
rect 34616 12100 34696 12180
rect 35768 12100 35848 12180
rect 36920 12100 37000 12180
rect 38072 12100 38152 12180
rect 39224 12100 39304 12180
rect 40376 12100 40456 12180
rect 41528 12100 41608 12180
rect 42680 12100 42760 12180
rect 76 11192 116 11201
rect 76 10688 116 11152
rect 1996 11108 2036 11117
rect 76 10639 116 10648
rect 1324 10856 1364 10865
rect 1132 10184 1172 10193
rect 1132 9596 1172 10144
rect 1132 9547 1172 9556
rect 1324 9596 1364 10816
rect 1324 9547 1364 9556
rect 1996 10436 2036 11068
rect 1228 9512 1268 9521
rect 1228 8840 1268 9472
rect 1228 8791 1268 8800
rect 1228 8672 1268 8681
rect 1228 8168 1268 8632
rect 1996 8672 2036 10396
rect 3052 10856 3092 10865
rect 3052 10436 3092 10816
rect 2284 10100 2324 10109
rect 1996 8623 2036 8632
rect 2092 9932 2132 9941
rect 1228 8119 1268 8128
rect 1228 8000 1268 8009
rect 1228 7496 1268 7960
rect 1228 7447 1268 7456
rect 1708 7748 1748 7757
rect 1612 6992 1652 7001
rect 1612 6236 1652 6952
rect 1612 6187 1652 6196
rect 1612 5816 1652 5825
rect 1612 5681 1652 5776
rect 76 5648 116 5657
rect 76 5480 116 5608
rect 76 5431 116 5440
rect 76 4976 116 4985
rect 76 4808 116 4936
rect 76 4759 116 4768
rect 1420 4136 1460 4145
rect 1132 3548 1172 3557
rect 652 1868 692 1877
rect 652 1448 692 1828
rect 652 1399 692 1408
rect 1132 776 1172 3508
rect 1420 3464 1460 4096
rect 1420 3415 1460 3424
rect 1708 2792 1748 7708
rect 2092 6068 2132 9892
rect 1996 6028 2132 6068
rect 2188 9260 2228 9269
rect 1996 3716 2036 6028
rect 1996 3667 2036 3676
rect 2092 5900 2132 5909
rect 1708 2743 1748 2752
rect 1996 3464 2036 3473
rect 1996 2792 2036 3424
rect 2092 3296 2132 5860
rect 2188 5564 2228 9220
rect 2188 4976 2228 5524
rect 2188 4927 2228 4936
rect 2284 5732 2324 10060
rect 2956 10016 2996 10025
rect 2668 9764 2708 9773
rect 2572 8672 2612 8681
rect 2284 4892 2324 5692
rect 2476 7916 2516 7925
rect 2380 5480 2420 5489
rect 2380 5060 2420 5440
rect 2380 5011 2420 5020
rect 2284 4843 2324 4852
rect 2476 4304 2516 7876
rect 2572 7916 2612 8632
rect 2572 6404 2612 7876
rect 2668 7328 2708 9724
rect 2764 8672 2804 8681
rect 2764 8168 2804 8632
rect 2764 8119 2804 8128
rect 2668 7279 2708 7288
rect 2764 7496 2804 7505
rect 2572 6355 2612 6364
rect 2476 4255 2516 4264
rect 2572 5480 2612 5489
rect 2380 3968 2420 3977
rect 2380 3884 2420 3928
rect 2380 3833 2420 3844
rect 2380 3716 2420 3725
rect 2092 3247 2132 3256
rect 2284 3632 2324 3641
rect 1996 2743 2036 2752
rect 1516 2540 1556 2549
rect 1516 2405 1556 2500
rect 2284 2120 2324 3592
rect 2380 2876 2420 3676
rect 2572 3212 2612 5440
rect 2572 3163 2612 3172
rect 2668 4136 2708 4145
rect 2668 2960 2708 4096
rect 2668 2911 2708 2920
rect 2764 2900 2804 7456
rect 2860 4724 2900 4733
rect 2860 4589 2900 4684
rect 2956 3464 2996 9976
rect 2956 3415 2996 3424
rect 3052 4220 3092 10396
rect 3532 10184 3572 12100
rect 4684 10436 4724 12100
rect 4928 10604 5296 10613
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 4928 10555 5296 10564
rect 4684 10387 4724 10396
rect 5836 10436 5876 12100
rect 5836 10387 5876 10396
rect 6892 10436 6932 10445
rect 6796 10268 6836 10277
rect 3532 10135 3572 10144
rect 6700 10184 6740 10193
rect 5356 10100 5396 10109
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 4300 8672 4340 8681
rect 4300 8537 4340 8632
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 4972 8336 5012 8345
rect 3436 7916 3476 7925
rect 3244 7832 3284 7841
rect 3052 3380 3092 4180
rect 3148 6488 3188 6497
rect 3148 3632 3188 6448
rect 3244 5144 3284 7792
rect 3436 7244 3476 7876
rect 4300 7916 4340 7925
rect 3476 7204 3572 7244
rect 3436 7195 3476 7204
rect 3244 5095 3284 5104
rect 3436 6740 3476 6749
rect 3148 3583 3188 3592
rect 3052 3331 3092 3340
rect 2956 3128 2996 3137
rect 2764 2860 2900 2900
rect 2380 2827 2420 2836
rect 2476 2792 2516 2801
rect 2476 2624 2516 2752
rect 2860 2792 2900 2860
rect 2860 2743 2900 2752
rect 2476 2575 2516 2584
rect 2956 2540 2996 3088
rect 3436 2876 3476 6700
rect 3532 5732 3572 7204
rect 4300 7076 4340 7876
rect 4972 7748 5012 8296
rect 4972 7699 5012 7708
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 4876 7328 4916 7337
rect 4300 7027 4340 7036
rect 4396 7244 4436 7253
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 3724 6572 3764 6581
rect 3724 6404 3764 6532
rect 3724 6355 3764 6364
rect 4300 6404 4340 6413
rect 4204 6236 4244 6245
rect 3532 4220 3572 5692
rect 4108 5732 4148 5741
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 3916 5060 3956 5069
rect 4108 5060 4148 5692
rect 3956 5020 4052 5060
rect 3916 5011 3956 5020
rect 3724 4892 3764 4901
rect 3724 4757 3764 4852
rect 4012 4640 4052 5020
rect 4108 5011 4148 5020
rect 4204 4976 4244 6196
rect 4300 5564 4340 6364
rect 4300 5515 4340 5524
rect 4396 6152 4436 7204
rect 4780 6992 4820 7001
rect 4684 6824 4724 6833
rect 4684 6572 4724 6784
rect 4684 6523 4724 6532
rect 4396 5732 4436 6112
rect 4204 4808 4244 4936
rect 4204 4759 4244 4768
rect 4012 4591 4052 4600
rect 3532 4171 3572 4180
rect 4108 4220 4148 4229
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 3436 2827 3476 2836
rect 3532 3716 3572 3725
rect 3340 2792 3380 2801
rect 2956 2491 2996 2500
rect 3244 2624 3284 2633
rect 3244 2489 3284 2584
rect 3148 2456 3188 2465
rect 3148 2372 3188 2416
rect 3148 2321 3188 2332
rect 3340 2372 3380 2752
rect 3340 2323 3380 2332
rect 3436 2708 3476 2717
rect 2284 2071 2324 2080
rect 1420 1952 1460 1961
rect 1420 1112 1460 1912
rect 1420 1063 1460 1072
rect 2764 1952 2804 1961
rect 1132 727 1172 736
rect 2764 104 2804 1912
rect 3436 1952 3476 2668
rect 3532 2204 3572 3676
rect 4108 2792 4148 4180
rect 4300 3968 4340 3977
rect 4396 3968 4436 5692
rect 4492 6488 4532 6497
rect 4492 5900 4532 6448
rect 4780 6152 4820 6952
rect 4876 6404 4916 7288
rect 5356 6992 5396 10060
rect 5740 10100 5780 10109
rect 5740 9764 5780 10060
rect 5548 9428 5588 9437
rect 5548 8756 5588 9388
rect 5740 9260 5780 9724
rect 6220 10100 6260 10109
rect 5740 9211 5780 9220
rect 5932 9512 5972 9521
rect 5356 6943 5396 6952
rect 5452 8420 5492 8429
rect 4876 6355 4916 6364
rect 5452 6404 5492 8380
rect 5548 7244 5588 8716
rect 5932 8756 5972 9472
rect 5932 8707 5972 8716
rect 5548 7195 5588 7204
rect 5932 7916 5972 7925
rect 5836 7076 5876 7085
rect 5548 6488 5588 6497
rect 5836 6488 5876 7036
rect 5588 6448 5876 6488
rect 5548 6439 5588 6448
rect 4780 6103 4820 6112
rect 5356 6236 5396 6245
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 4492 4220 4532 5860
rect 4684 5648 4724 5657
rect 4492 4171 4532 4180
rect 4588 5144 4628 5153
rect 4340 3928 4436 3968
rect 4204 3464 4244 3473
rect 4204 2876 4244 3424
rect 4300 3380 4340 3928
rect 4300 3331 4340 3340
rect 4492 3884 4532 3893
rect 4204 2827 4244 2836
rect 4396 3296 4436 3305
rect 3688 2288 4056 2297
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 3688 2239 4056 2248
rect 3532 2155 3572 2164
rect 4012 2120 4052 2129
rect 3436 1903 3476 1912
rect 3532 2036 3572 2045
rect 3532 1901 3572 1996
rect 4012 1985 4052 2080
rect 4108 1952 4148 2752
rect 4396 2708 4436 3256
rect 4108 1903 4148 1912
rect 4204 2624 4244 2633
rect 4204 1616 4244 2584
rect 4396 2624 4436 2668
rect 4396 2573 4436 2584
rect 4396 2372 4436 2381
rect 4300 2204 4340 2213
rect 4300 2036 4340 2164
rect 4300 1987 4340 1996
rect 4300 1868 4340 1879
rect 4300 1784 4340 1828
rect 4300 1735 4340 1744
rect 4204 1567 4244 1576
rect 4396 608 4436 2332
rect 4492 2120 4532 3844
rect 4492 2071 4532 2080
rect 4492 1700 4532 1709
rect 4492 1565 4532 1660
rect 4588 1532 4628 5104
rect 4684 4892 4724 5608
rect 4684 4843 4724 4852
rect 4780 4808 4820 4817
rect 4780 2120 4820 4768
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 5356 4220 5396 6196
rect 5452 5648 5492 6364
rect 5740 6320 5780 6329
rect 5452 5599 5492 5608
rect 5644 5732 5684 5741
rect 5452 5480 5492 5489
rect 5452 5345 5492 5440
rect 5644 5396 5684 5692
rect 5548 5228 5588 5237
rect 5356 4171 5396 4180
rect 5452 4892 5492 4901
rect 5164 3800 5204 3809
rect 5164 3716 5204 3760
rect 5164 3665 5204 3676
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 5452 2960 5492 4852
rect 5548 4388 5588 5188
rect 5644 5144 5684 5356
rect 5644 5095 5684 5104
rect 5740 5732 5780 6280
rect 5932 5984 5972 7876
rect 6028 7412 6068 7421
rect 6028 7277 6068 7372
rect 6124 6992 6164 7001
rect 6028 6656 6068 6665
rect 6028 6404 6068 6616
rect 6124 6656 6164 6952
rect 6124 6607 6164 6616
rect 6028 6355 6068 6364
rect 5932 5935 5972 5944
rect 6028 6236 6068 6245
rect 5836 5900 5876 5909
rect 5836 5765 5876 5860
rect 6028 5900 6068 6196
rect 6124 6236 6164 6245
rect 6124 6152 6164 6196
rect 6124 6101 6164 6112
rect 6028 5851 6068 5860
rect 6124 5984 6164 5993
rect 5932 5816 5972 5825
rect 5740 4892 5780 5692
rect 5740 4843 5780 4852
rect 5836 5648 5876 5657
rect 5548 4339 5588 4348
rect 5740 4724 5780 4733
rect 5644 4304 5684 4313
rect 5644 3884 5684 4264
rect 5740 4304 5780 4684
rect 5836 4388 5876 5608
rect 5836 4339 5876 4348
rect 5740 4255 5780 4264
rect 5932 4304 5972 5776
rect 6124 5312 6164 5944
rect 6220 5648 6260 10060
rect 6220 5599 6260 5608
rect 6316 9680 6356 9689
rect 6220 5312 6260 5321
rect 6124 5272 6220 5312
rect 5932 4255 5972 4264
rect 6028 4976 6068 4985
rect 5836 4220 5876 4229
rect 5644 3835 5684 3844
rect 5740 3968 5780 3977
rect 5740 3833 5780 3928
rect 5836 3884 5876 4180
rect 6028 4220 6068 4936
rect 6124 4976 6164 4985
rect 6124 4892 6164 4936
rect 6124 4841 6164 4852
rect 6028 4171 6068 4180
rect 6220 4808 6260 5272
rect 5836 3835 5876 3844
rect 6220 3464 6260 4768
rect 5548 3380 5588 3389
rect 5548 3245 5588 3340
rect 6028 3380 6068 3389
rect 5740 3296 5780 3305
rect 4780 2071 4820 2080
rect 4972 2708 5012 2717
rect 4780 1952 4820 1961
rect 4780 1817 4820 1912
rect 4972 1868 5012 2668
rect 5452 2708 5492 2920
rect 5740 2960 5780 3256
rect 5740 2911 5780 2920
rect 5932 2960 5972 2969
rect 5932 2708 5972 2920
rect 5452 2659 5492 2668
rect 5644 2668 5972 2708
rect 5644 2540 5684 2668
rect 5644 2491 5684 2500
rect 6028 2540 6068 3340
rect 6124 3296 6164 3305
rect 6124 2708 6164 3256
rect 6220 3044 6260 3424
rect 6316 4052 6356 9640
rect 6604 8588 6644 8597
rect 6508 8000 6548 8009
rect 6412 7160 6452 7169
rect 6508 7160 6548 7960
rect 6452 7120 6548 7160
rect 6412 7111 6452 7120
rect 6316 3548 6356 4012
rect 6316 3380 6356 3508
rect 6316 3331 6356 3340
rect 6412 6404 6452 6413
rect 6220 2995 6260 3004
rect 6220 2876 6260 2885
rect 6220 2741 6260 2836
rect 6124 2659 6164 2668
rect 6028 2491 6068 2500
rect 5740 2456 5780 2465
rect 5740 2321 5780 2416
rect 6028 2120 6068 2129
rect 6028 1985 6068 2080
rect 6412 2120 6452 6364
rect 6508 6068 6548 7120
rect 6604 7916 6644 8548
rect 6700 8084 6740 10144
rect 6700 8035 6740 8044
rect 6796 9176 6836 10228
rect 6796 8504 6836 9136
rect 6604 6908 6644 7876
rect 6796 7244 6836 8464
rect 6796 7195 6836 7204
rect 6604 6859 6644 6868
rect 6892 6236 6932 10396
rect 6988 10184 7028 12100
rect 8140 10436 8180 12100
rect 8140 10387 8180 10396
rect 8236 10688 8276 10697
rect 7276 10352 7316 10361
rect 6988 10135 7028 10144
rect 7084 10268 7124 10277
rect 7084 10016 7124 10228
rect 6988 9976 7124 10016
rect 7180 10100 7220 10109
rect 6988 8840 7028 9976
rect 6988 8791 7028 8800
rect 7084 9428 7124 9437
rect 7084 8756 7124 9388
rect 7084 8707 7124 8716
rect 7084 8588 7124 8597
rect 6988 8252 7028 8261
rect 6988 8168 7028 8212
rect 6988 8117 7028 8128
rect 6988 7832 7028 7841
rect 6988 7496 7028 7792
rect 6988 7447 7028 7456
rect 7084 7748 7124 8548
rect 6508 6019 6548 6028
rect 6700 6196 6932 6236
rect 6988 7160 7028 7169
rect 6988 6488 7028 7120
rect 6988 6236 7028 6448
rect 7084 6404 7124 7708
rect 7180 7244 7220 10060
rect 7276 9680 7316 10312
rect 7276 9631 7316 9640
rect 7660 10268 7700 10277
rect 7276 9344 7316 9353
rect 7276 7832 7316 9304
rect 7372 8588 7412 8597
rect 7372 8168 7412 8548
rect 7372 7916 7412 8128
rect 7468 8504 7508 8513
rect 7468 8084 7508 8464
rect 7660 8336 7700 10228
rect 7948 9512 7988 9521
rect 7852 9344 7892 9353
rect 7660 8287 7700 8296
rect 7756 9176 7796 9185
rect 7468 8035 7508 8044
rect 7660 8084 7700 8093
rect 7756 8084 7796 9136
rect 7852 8588 7892 9304
rect 7852 8539 7892 8548
rect 7948 8756 7988 9472
rect 7700 8044 7796 8084
rect 7660 8035 7700 8044
rect 7372 7867 7412 7876
rect 7660 7916 7700 7925
rect 7276 7783 7316 7792
rect 7180 7195 7220 7204
rect 7276 7664 7316 7673
rect 7276 7160 7316 7624
rect 7660 7412 7700 7876
rect 7660 7363 7700 7372
rect 7852 7664 7892 7673
rect 7276 7111 7316 7120
rect 7468 7244 7508 7253
rect 7468 7109 7508 7204
rect 7660 7244 7700 7255
rect 7660 7160 7700 7204
rect 7660 7111 7700 7120
rect 7084 6355 7124 6364
rect 7180 7076 7220 7085
rect 6508 5900 6548 5909
rect 6508 3548 6548 5860
rect 6604 5648 6644 5657
rect 6604 5144 6644 5608
rect 6604 5095 6644 5104
rect 6604 4976 6644 4985
rect 6604 4304 6644 4936
rect 6604 4255 6644 4264
rect 6508 3499 6548 3508
rect 6508 3212 6548 3221
rect 6508 2624 6548 3172
rect 6700 2876 6740 6196
rect 6796 6068 6836 6077
rect 6796 4220 6836 6028
rect 6892 5312 6932 5321
rect 6892 4892 6932 5272
rect 6988 4976 7028 6196
rect 7180 6320 7220 7036
rect 7756 7076 7796 7085
rect 7180 6185 7220 6280
rect 7276 6908 7316 6917
rect 7084 6152 7124 6161
rect 7084 5816 7124 6112
rect 7276 6068 7316 6868
rect 7756 6908 7796 7036
rect 7756 6859 7796 6868
rect 7756 6740 7796 6749
rect 7756 6572 7796 6700
rect 7756 6523 7796 6532
rect 7084 5767 7124 5776
rect 7180 5732 7220 5827
rect 7180 5683 7220 5692
rect 6988 4927 7028 4936
rect 7084 5648 7124 5657
rect 6892 4843 6932 4852
rect 6988 4640 7028 4649
rect 6988 4388 7028 4600
rect 6988 4339 7028 4348
rect 6796 4136 6836 4180
rect 7084 4220 7124 5608
rect 7180 5480 7220 5489
rect 7180 5345 7220 5440
rect 7180 5144 7220 5153
rect 7180 5060 7220 5104
rect 7180 5009 7220 5020
rect 7276 4892 7316 6028
rect 7468 5732 7508 5741
rect 7372 5228 7412 5237
rect 7372 5093 7412 5188
rect 7316 4852 7412 4892
rect 7276 4843 7316 4852
rect 7180 4724 7220 4733
rect 7180 4472 7220 4684
rect 7180 4423 7220 4432
rect 7276 4388 7316 4397
rect 7180 4220 7220 4229
rect 7084 4180 7180 4220
rect 6796 3380 6836 4096
rect 6988 4136 7028 4147
rect 6988 4052 7028 4096
rect 6988 4003 7028 4012
rect 6796 3331 6836 3340
rect 6700 2827 6740 2836
rect 6796 3128 6836 3137
rect 7084 3128 7124 4180
rect 7180 4171 7220 4180
rect 7276 3632 7316 4348
rect 7372 3884 7412 4852
rect 7372 3835 7412 3844
rect 7276 3583 7316 3592
rect 7372 3548 7412 3557
rect 7372 3413 7412 3508
rect 7468 3464 7508 5692
rect 7756 5732 7796 5741
rect 7660 5564 7700 5573
rect 7660 4388 7700 5524
rect 7756 4892 7796 5692
rect 7852 5732 7892 7624
rect 7948 7244 7988 8716
rect 8044 8084 8084 8093
rect 8044 7949 8084 8044
rect 8140 8000 8180 8009
rect 7948 7195 7988 7204
rect 8044 7496 8084 7505
rect 8044 7160 8084 7456
rect 8140 7328 8180 7960
rect 8140 7279 8180 7288
rect 8236 7160 8276 10648
rect 9292 10352 9332 12100
rect 9292 10303 9332 10312
rect 9676 10856 9716 10865
rect 9676 10520 9716 10816
rect 8908 10184 8948 10193
rect 8428 10100 8468 10109
rect 8428 9680 8468 10060
rect 8084 7120 8180 7160
rect 8044 7111 8084 7120
rect 7948 6992 7988 7001
rect 7948 6488 7988 6952
rect 7948 6439 7988 6448
rect 7852 5683 7892 5692
rect 8044 6320 8084 6329
rect 8044 5732 8084 6280
rect 8044 5683 8084 5692
rect 8044 5060 8084 5069
rect 8044 4925 8084 5020
rect 7756 4843 7796 4852
rect 7660 4304 7700 4348
rect 7660 4253 7700 4264
rect 7756 4472 7796 4481
rect 7756 4220 7796 4432
rect 7660 4136 7700 4145
rect 6796 2708 6836 3088
rect 6988 3088 7124 3128
rect 7180 3380 7220 3389
rect 6796 2659 6836 2668
rect 6892 3044 6932 3053
rect 6508 2575 6548 2584
rect 6700 2624 6740 2633
rect 6700 2372 6740 2584
rect 6700 2323 6740 2332
rect 6412 2071 6452 2080
rect 6892 2120 6932 3004
rect 6892 2071 6932 2080
rect 6988 2036 7028 3088
rect 7084 2960 7124 2969
rect 7084 2708 7124 2920
rect 7084 2659 7124 2668
rect 7180 2120 7220 3340
rect 7468 3212 7508 3424
rect 7564 3968 7604 3977
rect 7564 3380 7604 3928
rect 7564 3331 7604 3340
rect 7468 3163 7508 3172
rect 7276 2792 7316 2801
rect 7276 2204 7316 2752
rect 7372 2792 7412 2801
rect 7372 2708 7412 2752
rect 7372 2288 7412 2668
rect 7660 2372 7700 4096
rect 7756 3044 7796 4180
rect 8044 4220 8084 4229
rect 8044 4052 8084 4180
rect 7756 2995 7796 3004
rect 7852 3380 7892 3389
rect 7852 2540 7892 3340
rect 7852 2491 7892 2500
rect 7660 2323 7700 2332
rect 7372 2239 7412 2248
rect 7276 2155 7316 2164
rect 7180 2071 7220 2080
rect 6988 1987 7028 1996
rect 4972 1819 5012 1828
rect 7180 1952 7220 1961
rect 4588 1483 4628 1492
rect 4928 1532 5296 1541
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 4928 1483 5296 1492
rect 4396 559 4436 568
rect 7180 272 7220 1912
rect 7372 1952 7412 1961
rect 7372 1028 7412 1912
rect 8044 1700 8084 4012
rect 8140 2708 8180 7120
rect 8236 7111 8276 7120
rect 8332 9092 8372 9101
rect 8236 6404 8276 6413
rect 8236 6068 8276 6364
rect 8236 6019 8276 6028
rect 8236 5060 8276 5069
rect 8236 4136 8276 5020
rect 8236 4087 8276 4096
rect 8332 2900 8372 9052
rect 8428 8756 8468 9640
rect 8524 9932 8564 9941
rect 8524 9512 8564 9892
rect 8524 9463 8564 9472
rect 8908 9344 8948 10144
rect 9004 9512 9044 9521
rect 9004 9377 9044 9472
rect 9676 9428 9716 10480
rect 10444 10436 10484 12100
rect 10444 10387 10484 10396
rect 11500 11024 11540 11033
rect 10924 10268 10964 10277
rect 10732 10016 10772 10025
rect 9676 9379 9716 9388
rect 10540 9848 10580 9857
rect 8908 9295 8948 9304
rect 8428 8707 8468 8716
rect 8620 9260 8660 9269
rect 8524 8336 8564 8345
rect 8524 7916 8564 8296
rect 8428 7496 8468 7505
rect 8428 7160 8468 7456
rect 8524 7328 8564 7876
rect 8524 7279 8564 7288
rect 8428 7111 8468 7120
rect 8620 7076 8660 9220
rect 9100 9260 9140 9269
rect 9100 9176 9140 9220
rect 9100 9125 9140 9136
rect 10060 9260 10100 9269
rect 10060 9125 10100 9220
rect 9964 9008 10004 9017
rect 9100 8840 9140 8849
rect 8812 8756 8852 8765
rect 8716 8336 8756 8345
rect 8716 8000 8756 8296
rect 8812 8252 8852 8716
rect 8812 8203 8852 8212
rect 8716 7951 8756 7960
rect 9004 8084 9044 8093
rect 8908 7832 8948 7841
rect 8812 7748 8852 7757
rect 8812 7496 8852 7708
rect 8812 7447 8852 7456
rect 8620 7027 8660 7036
rect 8716 7412 8756 7421
rect 8428 6656 8468 6665
rect 8428 5900 8468 6616
rect 8716 6404 8756 7372
rect 8812 7244 8852 7253
rect 8812 6656 8852 7204
rect 8812 6607 8852 6616
rect 8716 6355 8756 6364
rect 8620 6236 8660 6331
rect 8660 6196 8756 6236
rect 8620 6187 8660 6196
rect 8620 6068 8660 6077
rect 8428 5860 8564 5900
rect 8428 5732 8468 5741
rect 8428 4220 8468 5692
rect 8524 5312 8564 5860
rect 8620 5480 8660 6028
rect 8620 5431 8660 5440
rect 8716 5741 8756 6196
rect 8716 5732 8761 5741
rect 8716 5692 8721 5732
rect 8716 5683 8761 5692
rect 8524 5272 8660 5312
rect 8524 5144 8564 5153
rect 8524 4892 8564 5104
rect 8524 4808 8564 4852
rect 8524 4759 8564 4768
rect 8428 3968 8468 4180
rect 8428 3919 8468 3928
rect 8620 3632 8660 5272
rect 8716 4808 8756 5683
rect 8716 4759 8756 4768
rect 8812 5648 8852 5657
rect 8812 4052 8852 5608
rect 8908 4976 8948 7792
rect 8908 4927 8948 4936
rect 9004 6908 9044 8044
rect 9004 5480 9044 6868
rect 8812 4003 8852 4012
rect 8620 3583 8660 3592
rect 8812 3380 8852 3475
rect 8812 3331 8852 3340
rect 8620 3296 8660 3305
rect 8620 3161 8660 3256
rect 8812 3212 8852 3221
rect 9004 3212 9044 5440
rect 9100 4220 9140 8800
rect 9868 8588 9908 8597
rect 9292 8504 9332 8513
rect 9292 7916 9332 8464
rect 9676 8420 9716 8429
rect 9196 7412 9236 7421
rect 9196 7328 9236 7372
rect 9196 7277 9236 7288
rect 9196 7160 9236 7169
rect 9196 6572 9236 7120
rect 9292 6656 9332 7876
rect 9484 7916 9524 7925
rect 9292 6607 9332 6616
rect 9388 7328 9428 7337
rect 9196 6523 9236 6532
rect 9292 6488 9332 6497
rect 9292 5900 9332 6448
rect 9196 5816 9236 5825
rect 9196 5732 9236 5776
rect 9196 5681 9236 5692
rect 9292 4976 9332 5860
rect 9388 6320 9428 7288
rect 9388 5480 9428 6280
rect 9388 5431 9428 5440
rect 9484 7160 9524 7876
rect 9580 7748 9620 7757
rect 9580 7328 9620 7708
rect 9676 7412 9716 8380
rect 9868 8252 9908 8548
rect 9676 7363 9716 7372
rect 9772 7496 9812 7505
rect 9580 7279 9620 7288
rect 9484 6908 9524 7120
rect 9676 7244 9716 7253
rect 9676 7160 9716 7204
rect 9676 7109 9716 7120
rect 9484 6320 9524 6868
rect 9676 6992 9716 7001
rect 9676 6572 9716 6952
rect 9676 6523 9716 6532
rect 9292 4927 9332 4936
rect 9196 4892 9236 4901
rect 9196 4808 9236 4852
rect 9388 4808 9428 4817
rect 9196 4768 9388 4808
rect 9196 4472 9236 4768
rect 9388 4759 9428 4768
rect 9196 4423 9236 4432
rect 9100 4171 9140 4180
rect 9484 4220 9524 6280
rect 9676 5648 9716 5657
rect 9580 5564 9620 5573
rect 9580 4472 9620 5524
rect 9580 4423 9620 4432
rect 9484 4171 9524 4180
rect 9196 3884 9236 3893
rect 9196 3632 9236 3844
rect 9196 3583 9236 3592
rect 9676 3296 9716 5608
rect 9772 5564 9812 7456
rect 9868 7244 9908 8212
rect 9868 7195 9908 7204
rect 9964 7328 10004 8968
rect 10540 8840 10580 9808
rect 10540 8791 10580 8800
rect 10732 8840 10772 9976
rect 10924 10016 10964 10228
rect 10924 9428 10964 9976
rect 10924 9379 10964 9388
rect 11116 10184 11156 10193
rect 10732 8791 10772 8800
rect 11020 8924 11060 8933
rect 11020 8789 11060 8884
rect 10060 8756 10100 8765
rect 10060 8336 10100 8716
rect 10828 8756 10868 8765
rect 10636 8672 10676 8681
rect 10060 8296 10292 8336
rect 10252 8168 10292 8296
rect 10252 8119 10292 8128
rect 10348 8084 10388 8093
rect 9964 7193 10004 7288
rect 10060 7916 10100 7925
rect 9772 5515 9812 5524
rect 9868 6824 9908 6833
rect 9772 4892 9812 4901
rect 9772 4220 9812 4852
rect 9772 4171 9812 4180
rect 9676 3247 9716 3256
rect 8852 3172 9044 3212
rect 9388 3212 9428 3221
rect 8332 2860 8468 2900
rect 8140 2668 8276 2708
rect 8140 2540 8180 2549
rect 8140 1952 8180 2500
rect 8140 1903 8180 1912
rect 8236 1868 8276 2668
rect 8428 2120 8468 2860
rect 8812 2288 8852 3172
rect 9388 3077 9428 3172
rect 9484 2792 9524 2801
rect 8812 2239 8852 2248
rect 9004 2708 9044 2717
rect 8428 2071 8468 2080
rect 8620 2120 8660 2129
rect 8236 1819 8276 1828
rect 8620 1868 8660 2080
rect 9004 2036 9044 2668
rect 9484 2657 9524 2752
rect 9004 1987 9044 1996
rect 9676 2624 9716 2633
rect 8620 1819 8660 1828
rect 9676 1868 9716 2584
rect 9772 2036 9812 2045
rect 9868 2036 9908 6784
rect 9964 6404 10004 6415
rect 9964 6320 10004 6364
rect 9964 5312 10004 6280
rect 10060 6236 10100 7876
rect 10348 7916 10388 8044
rect 10636 8084 10676 8632
rect 10636 8035 10676 8044
rect 10828 7916 10868 8716
rect 11020 8168 11060 8177
rect 10348 7867 10388 7876
rect 10636 7876 10868 7916
rect 10924 8084 10964 8093
rect 10348 7664 10388 7673
rect 10252 7580 10292 7589
rect 10060 6187 10100 6196
rect 10156 7160 10196 7169
rect 9964 5263 10004 5272
rect 10060 6068 10100 6077
rect 9812 1996 9908 2036
rect 9964 3212 10004 3221
rect 9964 2036 10004 3172
rect 9772 1987 9812 1996
rect 9964 1987 10004 1996
rect 9676 1819 9716 1828
rect 10060 1784 10100 6028
rect 10156 5648 10196 7120
rect 10252 6656 10292 7540
rect 10252 6607 10292 6616
rect 10348 6488 10388 7624
rect 10540 7580 10580 7589
rect 10540 7496 10580 7540
rect 10540 7445 10580 7456
rect 10348 6439 10388 6448
rect 10540 6404 10580 6413
rect 10348 6320 10388 6329
rect 10156 2792 10196 5608
rect 10252 6236 10292 6245
rect 10252 5480 10292 6196
rect 10348 6068 10388 6280
rect 10348 6019 10388 6028
rect 10348 5816 10388 5911
rect 10348 5767 10388 5776
rect 10444 5732 10484 5741
rect 10252 5431 10292 5440
rect 10348 5648 10388 5657
rect 10252 4892 10292 4903
rect 10252 4808 10292 4852
rect 10252 4759 10292 4768
rect 10252 4304 10292 4313
rect 10252 4136 10292 4264
rect 10252 4087 10292 4096
rect 10252 3968 10292 3977
rect 10252 3800 10292 3928
rect 10252 3751 10292 3760
rect 10252 3380 10292 3389
rect 10252 2876 10292 3340
rect 10252 2827 10292 2836
rect 10156 2743 10196 2752
rect 10060 1735 10100 1744
rect 8044 1651 8084 1660
rect 8620 1700 8660 1709
rect 8620 1565 8660 1660
rect 10156 1700 10196 1709
rect 7372 979 7412 988
rect 10156 860 10196 1660
rect 10348 1616 10388 5608
rect 10444 5597 10484 5692
rect 10444 5060 10484 5069
rect 10444 4892 10484 5020
rect 10444 3548 10484 4852
rect 10444 3499 10484 3508
rect 10540 3464 10580 6364
rect 10636 5060 10676 7876
rect 10828 7748 10868 7757
rect 10732 7160 10772 7169
rect 10732 6908 10772 7120
rect 10732 6656 10772 6868
rect 10732 6607 10772 6616
rect 10636 5011 10676 5020
rect 10732 5396 10772 5405
rect 10636 4808 10676 4817
rect 10636 4640 10676 4768
rect 10636 4591 10676 4600
rect 10732 4556 10772 5356
rect 10732 4507 10772 4516
rect 10732 4388 10772 4397
rect 10540 1868 10580 3424
rect 10636 4220 10676 4229
rect 10636 3380 10676 4180
rect 10732 4200 10772 4348
rect 10828 4304 10868 7708
rect 10828 4255 10868 4264
rect 10732 4160 10868 4200
rect 10828 3800 10868 4160
rect 10732 3548 10772 3557
rect 10732 3464 10772 3508
rect 10732 3413 10772 3424
rect 10636 3331 10676 3340
rect 10828 3380 10868 3760
rect 10828 3331 10868 3340
rect 10924 2900 10964 8044
rect 11020 7664 11060 8128
rect 11020 7615 11060 7624
rect 11020 7160 11060 7169
rect 11020 6488 11060 7120
rect 11116 6740 11156 10144
rect 11500 10184 11540 10984
rect 11596 10436 11636 12100
rect 11596 10387 11636 10396
rect 12748 10436 12788 12100
rect 12748 10387 12788 10396
rect 11500 10135 11540 10144
rect 11692 10268 11732 10277
rect 11308 9512 11348 9521
rect 11212 9260 11252 9269
rect 11212 8840 11252 9220
rect 11212 8791 11252 8800
rect 11308 9092 11348 9472
rect 11500 9400 11636 9428
rect 11500 9388 11596 9400
rect 11308 8756 11348 9052
rect 11308 8707 11348 8716
rect 11404 9092 11444 9101
rect 11404 8672 11444 9052
rect 11404 8623 11444 8632
rect 11308 8504 11348 8513
rect 11308 8420 11348 8464
rect 11308 8369 11348 8380
rect 11500 8336 11540 9388
rect 11596 9351 11636 9360
rect 11500 8168 11540 8296
rect 11500 8119 11540 8128
rect 11692 7412 11732 10228
rect 12844 10100 12884 10109
rect 12364 9764 12404 9773
rect 11788 9596 11828 9605
rect 11788 9260 11828 9556
rect 12268 9512 12308 9521
rect 12076 9428 12116 9437
rect 11788 9211 11828 9220
rect 11884 9344 11924 9353
rect 11884 8756 11924 9304
rect 12076 9092 12116 9388
rect 12076 9043 12116 9052
rect 11884 8707 11924 8716
rect 11884 8588 11924 8597
rect 11884 8252 11924 8548
rect 11788 7916 11828 7925
rect 11884 7916 11924 8212
rect 11828 7876 11924 7916
rect 11788 7867 11828 7876
rect 11116 6691 11156 6700
rect 11212 7244 11252 7253
rect 11020 6439 11060 6448
rect 11212 6236 11252 7204
rect 11692 7244 11732 7372
rect 11308 7160 11348 7169
rect 11308 7025 11348 7120
rect 11596 7160 11636 7169
rect 11596 6992 11636 7120
rect 11596 6943 11636 6952
rect 11692 6992 11732 7204
rect 11692 6943 11732 6952
rect 11884 7244 11924 7253
rect 11500 6908 11540 6917
rect 11212 6187 11252 6196
rect 11404 6404 11444 6413
rect 11308 5816 11348 5825
rect 11020 5648 11060 5657
rect 11020 5513 11060 5608
rect 11116 5480 11156 5489
rect 11156 5440 11252 5480
rect 11116 5431 11156 5440
rect 11020 5060 11060 5069
rect 11020 3464 11060 5020
rect 11116 4892 11156 4901
rect 11116 4220 11156 4852
rect 11116 4171 11156 4180
rect 11212 4220 11252 5440
rect 11308 4388 11348 5776
rect 11404 5480 11444 6364
rect 11404 5431 11444 5440
rect 11500 6236 11540 6868
rect 11884 6404 11924 7204
rect 11596 6236 11636 6245
rect 11500 6196 11596 6236
rect 11500 4892 11540 6196
rect 11596 6187 11636 6196
rect 11596 5732 11636 5741
rect 11596 5144 11636 5692
rect 11596 5095 11636 5104
rect 11884 5732 11924 6364
rect 11500 4843 11540 4852
rect 11308 4339 11348 4348
rect 11212 4171 11252 4180
rect 11692 4136 11732 4145
rect 11020 3415 11060 3424
rect 11212 3800 11252 3809
rect 10924 2860 11060 2900
rect 10924 2708 10964 2717
rect 10924 2573 10964 2668
rect 10540 1819 10580 1828
rect 10348 1567 10388 1576
rect 10156 811 10196 820
rect 7180 223 7220 232
rect 2860 104 2900 113
rect 2764 64 2860 104
rect 11020 80 11060 2860
rect 11212 80 11252 3760
rect 11500 3380 11540 3389
rect 11308 3128 11348 3137
rect 11308 1952 11348 3088
rect 11500 2792 11540 3340
rect 11692 2960 11732 4096
rect 11692 2911 11732 2920
rect 11500 2743 11540 2752
rect 11308 1903 11348 1912
rect 11404 2624 11444 2633
rect 11404 80 11444 2584
rect 11884 2624 11924 5692
rect 12172 7244 12212 7253
rect 12076 5228 12116 5237
rect 11788 2120 11828 2129
rect 11788 1532 11828 2080
rect 11884 1868 11924 2584
rect 11980 4136 12020 4145
rect 11980 2624 12020 4096
rect 12076 3800 12116 5188
rect 12172 3968 12212 7204
rect 12172 3919 12212 3928
rect 12268 3884 12308 9472
rect 12364 9008 12404 9724
rect 12460 9680 12500 9689
rect 12748 9680 12788 9689
rect 12500 9640 12692 9680
rect 12460 9631 12500 9640
rect 12652 9344 12692 9640
rect 12748 9428 12788 9640
rect 12748 9379 12788 9388
rect 12652 9295 12692 9304
rect 12364 8959 12404 8968
rect 12460 8924 12500 8933
rect 12460 8000 12500 8884
rect 12844 8756 12884 10060
rect 13324 10016 13364 10025
rect 13324 9428 13364 9976
rect 13516 10016 13556 10025
rect 13516 9881 13556 9976
rect 13900 9680 13940 12100
rect 14476 11108 14516 11117
rect 14476 10268 14516 11068
rect 13900 9631 13940 9640
rect 14380 10184 14420 10193
rect 13324 9379 13364 9388
rect 13996 9596 14036 9605
rect 12844 8707 12884 8716
rect 13036 8672 13076 8681
rect 12460 7951 12500 7960
rect 12556 8000 12596 8009
rect 12364 6908 12404 6917
rect 12364 4052 12404 6868
rect 12460 6656 12500 6665
rect 12460 5144 12500 6616
rect 12460 5095 12500 5104
rect 12460 4976 12500 4985
rect 12460 4556 12500 4936
rect 12460 4507 12500 4516
rect 12364 4003 12404 4012
rect 12268 3835 12308 3844
rect 12076 3464 12116 3760
rect 12076 3415 12116 3424
rect 12556 3548 12596 7960
rect 13036 7328 13076 8632
rect 13996 8672 14036 9556
rect 13996 8623 14036 8632
rect 14092 9512 14132 9521
rect 13132 8588 13172 8597
rect 13132 8000 13172 8548
rect 13420 8504 13460 8513
rect 13172 7960 13268 8000
rect 13132 7951 13172 7960
rect 13132 7748 13172 7757
rect 13132 7496 13172 7708
rect 13132 7447 13172 7456
rect 13036 7288 13172 7328
rect 12844 7076 12884 7085
rect 12844 6740 12884 7036
rect 12844 6691 12884 6700
rect 13036 6992 13076 7001
rect 12844 6152 12884 6161
rect 12844 5060 12884 6112
rect 12940 5816 12980 5825
rect 12940 5732 12980 5776
rect 12940 5681 12980 5692
rect 13036 5060 13076 6952
rect 12844 5020 12980 5060
rect 12748 4892 12788 4901
rect 12844 4892 12884 4920
rect 12788 4852 12844 4892
rect 12652 4808 12692 4817
rect 12652 4673 12692 4768
rect 12748 4640 12788 4852
rect 12844 4843 12884 4852
rect 12748 4591 12788 4600
rect 12940 4472 12980 5020
rect 13036 5011 13076 5020
rect 13036 4892 13076 4901
rect 13036 4808 13076 4852
rect 13036 4757 13076 4768
rect 13132 4640 13172 7288
rect 13228 5816 13268 7960
rect 13420 7412 13460 8464
rect 13804 8504 13844 8513
rect 13612 8168 13652 8177
rect 13420 7363 13460 7372
rect 13516 8000 13556 8009
rect 13324 7328 13364 7337
rect 13324 6572 13364 7288
rect 13324 6523 13364 6532
rect 13420 7244 13460 7253
rect 13228 5732 13268 5776
rect 13228 5652 13268 5692
rect 13420 6404 13460 7204
rect 13420 5312 13460 6364
rect 13420 5263 13460 5272
rect 13324 4976 13364 4985
rect 13364 4936 13460 4976
rect 13324 4927 13364 4936
rect 12268 3380 12308 3389
rect 11980 2575 12020 2584
rect 12076 3296 12116 3305
rect 11884 1819 11924 1828
rect 11980 2204 12020 2213
rect 11788 1483 11828 1492
rect 11788 608 11828 617
rect 11596 104 11636 113
rect 2860 36 2900 64
rect 11000 0 11080 80
rect 11192 0 11272 80
rect 11384 0 11464 80
rect 11576 64 11596 80
rect 11788 80 11828 568
rect 11980 80 12020 2164
rect 12076 2120 12116 3256
rect 12268 2708 12308 3340
rect 12556 3380 12596 3508
rect 12556 3331 12596 3340
rect 12844 4432 12980 4472
rect 13036 4600 13172 4640
rect 12844 4220 12884 4432
rect 12940 4304 12980 4313
rect 13036 4304 13076 4600
rect 13420 4556 13460 4936
rect 13420 4507 13460 4516
rect 13324 4472 13364 4481
rect 12980 4264 13076 4304
rect 13228 4388 13268 4397
rect 12940 4236 12980 4264
rect 12844 3380 12884 4180
rect 12940 4052 12980 4061
rect 12940 3917 12980 4012
rect 13036 3968 13076 3977
rect 12844 3331 12884 3340
rect 13036 3128 13076 3928
rect 12844 3088 13076 3128
rect 13132 3548 13172 3557
rect 12844 2900 12884 3088
rect 13132 3044 13172 3508
rect 13036 3004 13172 3044
rect 12652 2876 12692 2885
rect 12268 2638 12308 2647
rect 12556 2792 12596 2801
rect 12556 2540 12596 2752
rect 12556 2491 12596 2500
rect 12268 2456 12308 2465
rect 12460 2456 12500 2465
rect 12308 2416 12404 2456
rect 12268 2407 12308 2416
rect 12076 2071 12116 2080
rect 12172 1448 12212 1457
rect 12172 80 12212 1408
rect 12364 80 12404 2416
rect 12460 1952 12500 2416
rect 12460 1903 12500 1912
rect 12556 2372 12596 2381
rect 12556 80 12596 2332
rect 12652 1532 12692 2836
rect 12748 2876 12788 2885
rect 12844 2876 12980 2900
rect 12844 2860 12940 2876
rect 12748 2708 12788 2836
rect 12940 2827 12980 2836
rect 12748 2659 12788 2668
rect 12940 2288 12980 2297
rect 12940 2153 12980 2248
rect 13036 2204 13076 3004
rect 13228 2900 13268 4348
rect 13324 4220 13364 4432
rect 13324 4171 13364 4180
rect 13516 3212 13556 7960
rect 13612 5732 13652 8128
rect 13804 8168 13844 8464
rect 13804 8119 13844 8128
rect 13612 5683 13652 5692
rect 13708 8084 13748 8093
rect 13708 5564 13748 8044
rect 13900 7916 13940 7925
rect 13612 5524 13748 5564
rect 13804 7832 13844 7841
rect 13612 3548 13652 5524
rect 13708 4892 13748 4901
rect 13708 4304 13748 4852
rect 13708 3884 13748 4264
rect 13708 3835 13748 3844
rect 13612 3499 13652 3508
rect 13516 3163 13556 3172
rect 13612 3380 13652 3389
rect 13036 2155 13076 2164
rect 13132 2860 13268 2900
rect 13516 3044 13556 3053
rect 12748 2120 12788 2129
rect 12748 2036 12788 2080
rect 12748 1985 12788 1996
rect 12844 2120 12884 2129
rect 12844 1952 12884 2080
rect 12844 1903 12884 1912
rect 12940 1700 12980 1709
rect 12652 1492 12788 1532
rect 12748 80 12788 1492
rect 12940 1364 12980 1660
rect 12940 1315 12980 1324
rect 13036 1532 13076 1541
rect 12940 440 12980 449
rect 12940 80 12980 400
rect 13036 272 13076 1492
rect 13132 1280 13172 2860
rect 13420 2792 13460 2801
rect 13420 2657 13460 2752
rect 13420 2372 13460 2381
rect 13132 1231 13172 1240
rect 13228 2204 13268 2213
rect 13228 440 13268 2164
rect 13420 2036 13460 2332
rect 13420 1987 13460 1996
rect 13228 391 13268 400
rect 13324 1280 13364 1289
rect 13036 232 13172 272
rect 13132 80 13172 232
rect 13324 80 13364 1240
rect 13516 80 13556 3004
rect 13612 1448 13652 3340
rect 13708 3380 13748 3389
rect 13708 2876 13748 3340
rect 13804 3044 13844 7792
rect 13900 7244 13940 7876
rect 13900 7204 14036 7244
rect 13900 3464 13940 3473
rect 13900 3329 13940 3424
rect 13996 3380 14036 7204
rect 14092 6572 14132 9472
rect 14380 9428 14420 10144
rect 14380 9379 14420 9388
rect 14380 9260 14420 9269
rect 14284 9176 14324 9185
rect 14284 8756 14324 9136
rect 14380 9008 14420 9220
rect 14380 8959 14420 8968
rect 14188 8672 14228 8683
rect 14188 8588 14228 8632
rect 14188 8539 14228 8548
rect 14188 8420 14228 8429
rect 14188 8000 14228 8380
rect 14188 7951 14228 7960
rect 14092 6523 14132 6532
rect 14188 7748 14228 7757
rect 14092 6068 14132 6077
rect 14092 5933 14132 6028
rect 13996 3331 14036 3340
rect 14092 5648 14132 5657
rect 13804 2995 13844 3004
rect 13900 3212 13940 3221
rect 13900 2960 13940 3172
rect 13900 2911 13940 2920
rect 13708 2827 13748 2836
rect 13804 2540 13844 2549
rect 13708 2288 13748 2297
rect 13708 1616 13748 2248
rect 13804 1868 13844 2500
rect 13804 1819 13844 1828
rect 13708 1567 13748 1576
rect 13900 1616 13940 1625
rect 13612 1408 13748 1448
rect 13708 80 13748 1408
rect 13900 80 13940 1576
rect 14092 80 14132 5608
rect 14188 5648 14228 7708
rect 14284 7328 14324 8716
rect 14284 7279 14324 7288
rect 14380 6992 14420 7001
rect 14380 6857 14420 6952
rect 14476 6572 14516 10228
rect 14572 10856 14612 10865
rect 14572 9512 14612 10816
rect 14764 10772 14804 10781
rect 14572 9463 14612 9472
rect 14668 10100 14708 10109
rect 14668 9344 14708 10060
rect 14668 9295 14708 9304
rect 14764 9176 14804 10732
rect 14668 9136 14804 9176
rect 14860 10268 14900 10277
rect 14572 8252 14612 8261
rect 14572 7244 14612 8212
rect 14572 7195 14612 7204
rect 14476 6523 14516 6532
rect 14572 6824 14612 6833
rect 14380 6404 14420 6413
rect 14572 6404 14612 6784
rect 14188 5599 14228 5608
rect 14284 6320 14324 6329
rect 14284 5480 14324 6280
rect 14188 5440 14324 5480
rect 14188 2120 14228 5440
rect 14284 5312 14324 5321
rect 14284 4892 14324 5272
rect 14284 4843 14324 4852
rect 14284 4724 14324 4733
rect 14284 4556 14324 4684
rect 14284 4507 14324 4516
rect 14284 4304 14324 4313
rect 14284 2792 14324 4264
rect 14380 4200 14420 6364
rect 14476 6364 14572 6404
rect 14476 4304 14516 6364
rect 14572 6355 14612 6364
rect 14572 5480 14612 5489
rect 14668 5480 14708 9136
rect 14860 8756 14900 10228
rect 14956 10016 14996 10025
rect 14956 9428 14996 9976
rect 15052 9680 15092 12100
rect 16204 10436 16244 12100
rect 16972 11276 17012 11285
rect 16204 10387 16244 10396
rect 16396 10520 16436 10529
rect 16396 10268 16436 10480
rect 15052 9631 15092 9640
rect 15148 10100 15188 10109
rect 14956 9379 14996 9388
rect 14612 5440 14708 5480
rect 14764 7916 14804 7925
rect 14572 5431 14612 5440
rect 14668 4892 14708 4901
rect 14476 4255 14516 4264
rect 14572 4640 14612 4649
rect 14380 4160 14516 4200
rect 14380 4052 14420 4061
rect 14380 3800 14420 4012
rect 14380 3751 14420 3760
rect 14476 3632 14516 4160
rect 14284 2743 14324 2752
rect 14380 3592 14516 3632
rect 14380 2288 14420 3592
rect 14476 3464 14516 3473
rect 14476 3296 14516 3424
rect 14476 3247 14516 3256
rect 14572 3212 14612 4600
rect 14668 4388 14708 4852
rect 14764 4892 14804 7876
rect 14860 7664 14900 8716
rect 15052 9344 15092 9353
rect 15052 8000 15092 9304
rect 15052 7951 15092 7960
rect 14956 7832 14996 7841
rect 14996 7792 15092 7832
rect 14956 7783 14996 7792
rect 14860 7624 14996 7664
rect 14956 7244 14996 7624
rect 14860 7160 14900 7169
rect 14860 6740 14900 7120
rect 14860 6691 14900 6700
rect 14860 6236 14900 6245
rect 14860 5732 14900 6196
rect 14860 5683 14900 5692
rect 14956 5564 14996 7204
rect 14764 4843 14804 4852
rect 14860 5524 14996 5564
rect 14860 4724 14900 5524
rect 14668 4339 14708 4348
rect 14764 4684 14900 4724
rect 14956 5312 14996 5321
rect 14764 4136 14804 4684
rect 14764 4087 14804 4096
rect 14860 4304 14900 4344
rect 14860 4220 14900 4264
rect 14860 3716 14900 4180
rect 14956 4052 14996 5272
rect 15052 4976 15092 7792
rect 15148 7076 15188 10060
rect 15532 9512 15572 9521
rect 15436 9428 15476 9437
rect 15436 8756 15476 9388
rect 15532 9377 15572 9472
rect 15820 9428 15860 9437
rect 15820 9260 15860 9388
rect 15148 7027 15188 7036
rect 15244 8168 15284 8177
rect 15052 4927 15092 4936
rect 15148 5648 15188 5657
rect 15148 5480 15188 5608
rect 15148 4304 15188 5440
rect 15148 4255 15188 4264
rect 14956 4003 14996 4012
rect 15052 3968 15092 3977
rect 14860 3667 14900 3676
rect 14956 3800 14996 3809
rect 14572 3163 14612 3172
rect 14668 3548 14708 3557
rect 14572 3044 14612 3053
rect 14572 2900 14612 3004
rect 14380 2239 14420 2248
rect 14476 2860 14612 2900
rect 14476 2204 14516 2860
rect 14476 2155 14516 2164
rect 14188 2071 14228 2080
rect 14476 1952 14516 1961
rect 14284 1448 14324 1457
rect 14284 80 14324 1408
rect 14476 1112 14516 1912
rect 14572 1700 14612 1709
rect 14572 1280 14612 1660
rect 14572 1231 14612 1240
rect 14476 1063 14516 1072
rect 14476 272 14516 281
rect 14476 80 14516 232
rect 14668 80 14708 3508
rect 14764 3464 14804 3473
rect 14764 608 14804 3424
rect 14860 3128 14900 3137
rect 14860 1616 14900 3088
rect 14956 1784 14996 3760
rect 15052 3464 15092 3928
rect 15052 3415 15092 3424
rect 15148 3212 15188 3221
rect 15148 2708 15188 3172
rect 15148 2659 15188 2668
rect 15148 2540 15188 2549
rect 15148 2120 15188 2500
rect 15148 2071 15188 2080
rect 14956 1735 14996 1744
rect 14860 1567 14900 1576
rect 14764 559 14804 568
rect 14860 1448 14900 1457
rect 14860 80 14900 1408
rect 15052 1028 15092 1037
rect 15052 80 15092 988
rect 15244 80 15284 8128
rect 15340 7748 15380 7757
rect 15340 1868 15380 7708
rect 15436 6404 15476 8716
rect 15436 6355 15476 6364
rect 15532 9220 15860 9260
rect 15436 5648 15476 5657
rect 15436 4892 15476 5608
rect 15436 2876 15476 4852
rect 15436 2456 15476 2836
rect 15436 2407 15476 2416
rect 15532 2120 15572 9220
rect 15916 9092 15956 9101
rect 15916 8756 15956 9052
rect 15820 8588 15860 8597
rect 15820 8504 15860 8548
rect 15820 8453 15860 8464
rect 15724 8420 15764 8429
rect 15628 8000 15668 8095
rect 15628 7951 15668 7960
rect 15532 2071 15572 2080
rect 15628 7832 15668 7841
rect 15340 1819 15380 1828
rect 15436 1616 15476 1625
rect 15436 80 15476 1576
rect 15628 80 15668 7792
rect 15724 5312 15764 8380
rect 15916 7244 15956 8716
rect 16108 8924 16148 8933
rect 15916 7195 15956 7204
rect 16012 7748 16052 7757
rect 15820 6320 15860 6331
rect 15820 6236 15860 6280
rect 15820 6187 15860 6196
rect 15724 5263 15764 5272
rect 15820 5900 15860 5909
rect 15820 5732 15860 5860
rect 15820 4976 15860 5692
rect 15724 4936 15820 4976
rect 15724 2900 15764 4936
rect 15820 4927 15860 4936
rect 15916 5144 15956 5153
rect 15820 4220 15860 4229
rect 15820 3884 15860 4180
rect 15820 3835 15860 3844
rect 15724 2860 15860 2900
rect 15820 2708 15860 2860
rect 15820 2659 15860 2668
rect 15916 2120 15956 5104
rect 15916 2071 15956 2080
rect 15820 1952 15860 1961
rect 15724 1868 15764 1877
rect 15724 1028 15764 1828
rect 15724 979 15764 988
rect 15820 80 15860 1912
rect 15916 1952 15956 1961
rect 15916 1448 15956 1912
rect 15916 1399 15956 1408
rect 16012 80 16052 7708
rect 16108 5732 16148 8884
rect 16300 7748 16340 7757
rect 16108 5683 16148 5692
rect 16204 6992 16244 7001
rect 16108 4724 16148 4733
rect 16108 4388 16148 4684
rect 16108 4339 16148 4348
rect 16108 3800 16148 3809
rect 16108 3464 16148 3760
rect 16108 3415 16148 3424
rect 16204 2372 16244 6952
rect 16300 5816 16340 7708
rect 16396 7244 16436 10228
rect 16972 10184 17012 11236
rect 17356 10436 17396 12100
rect 17356 10387 17396 10396
rect 18412 10940 18452 10949
rect 16972 10135 17012 10144
rect 17452 10100 17492 10109
rect 16972 9512 17012 9521
rect 16588 9428 16628 9437
rect 16588 9008 16628 9388
rect 16972 9260 17012 9472
rect 16972 9211 17012 9220
rect 16588 8959 16628 8968
rect 17452 8756 17492 10060
rect 17644 10016 17684 10025
rect 17836 10016 17876 10025
rect 17684 9976 17836 10016
rect 17644 9967 17684 9976
rect 17836 9967 17876 9976
rect 17452 8707 17492 8716
rect 17740 9512 17780 9521
rect 17740 9428 17780 9472
rect 17740 8756 17780 9388
rect 17740 8707 17780 8716
rect 17836 9512 17876 9521
rect 17548 8672 17588 8681
rect 17260 8000 17300 8009
rect 16396 6404 16436 7204
rect 16684 7916 16724 7925
rect 16396 6355 16436 6364
rect 16588 6488 16628 6497
rect 16300 5767 16340 5776
rect 16492 5732 16532 5741
rect 16396 5228 16436 5237
rect 16300 4892 16340 4901
rect 16300 4388 16340 4852
rect 16300 4339 16340 4348
rect 16204 2323 16244 2332
rect 16204 860 16244 869
rect 16204 80 16244 820
rect 16396 80 16436 5188
rect 16492 4976 16532 5692
rect 16492 4927 16532 4936
rect 16588 4724 16628 6448
rect 16684 5984 16724 7876
rect 16684 5935 16724 5944
rect 16780 7832 16820 7841
rect 16588 4675 16628 4684
rect 16684 4892 16724 4901
rect 16588 4556 16628 4565
rect 16492 4304 16532 4313
rect 16492 4220 16532 4264
rect 16588 4304 16628 4516
rect 16684 4472 16724 4852
rect 16684 4423 16724 4432
rect 16588 4255 16628 4264
rect 16684 4304 16724 4313
rect 16492 4169 16532 4180
rect 16588 3632 16628 3641
rect 16588 3380 16628 3592
rect 16588 3331 16628 3340
rect 16492 2960 16532 2969
rect 16492 1448 16532 2920
rect 16492 1399 16532 1408
rect 16588 2792 16628 2801
rect 16588 80 16628 2752
rect 16684 2120 16724 4264
rect 16684 2071 16724 2080
rect 16780 80 16820 7792
rect 16972 7748 17012 7757
rect 16972 5060 17012 7708
rect 17068 6488 17108 6497
rect 17068 5900 17108 6448
rect 17068 5851 17108 5860
rect 17164 5732 17204 5741
rect 17164 5564 17204 5692
rect 16972 5011 17012 5020
rect 17068 5312 17108 5321
rect 16876 3800 16916 3809
rect 16876 2372 16916 3760
rect 16972 3380 17012 3389
rect 16972 2960 17012 3340
rect 16972 2911 17012 2920
rect 16876 2323 16916 2332
rect 16972 2372 17012 2381
rect 16972 2036 17012 2332
rect 16972 1868 17012 1996
rect 17068 1952 17108 5272
rect 17164 5144 17204 5524
rect 17164 5095 17204 5104
rect 17164 3212 17204 3221
rect 17164 2708 17204 3172
rect 17164 2659 17204 2668
rect 17068 1903 17108 1912
rect 16972 1819 17012 1828
rect 16972 1448 17012 1457
rect 17260 1448 17300 7960
rect 17452 7244 17492 7253
rect 17452 6992 17492 7204
rect 17452 6943 17492 6952
rect 17452 6488 17492 6497
rect 17452 6404 17492 6448
rect 17452 5984 17492 6364
rect 17452 5935 17492 5944
rect 17548 5732 17588 8632
rect 17740 8168 17780 8179
rect 17740 8084 17780 8128
rect 17740 8035 17780 8044
rect 17644 7412 17684 7452
rect 17644 7328 17684 7372
rect 17644 7244 17684 7288
rect 17644 7193 17684 7204
rect 17836 7160 17876 9472
rect 18412 9512 18452 10900
rect 18508 9680 18548 12100
rect 19564 10688 19604 10697
rect 19468 10184 19508 10193
rect 18700 10016 18740 10025
rect 18508 9631 18548 9640
rect 18604 9764 18644 9773
rect 18604 9512 18644 9724
rect 18700 9680 18740 9976
rect 19276 10016 19316 10025
rect 18808 9848 19176 9857
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 18808 9799 19176 9808
rect 18700 9631 18740 9640
rect 18124 9428 18164 9437
rect 18124 8924 18164 9388
rect 18124 8875 18164 8884
rect 18124 8756 18164 8765
rect 18412 8756 18452 9472
rect 18508 9472 18644 9512
rect 18508 9428 18548 9472
rect 18508 9379 18548 9388
rect 18988 9428 19028 9437
rect 18508 9260 18548 9269
rect 18508 9176 18548 9220
rect 18700 9176 18740 9185
rect 18508 9136 18700 9176
rect 18700 9127 18740 9136
rect 18508 8756 18548 8765
rect 18412 8716 18508 8756
rect 18124 8621 18164 8716
rect 17932 8168 17972 8177
rect 17932 7580 17972 8128
rect 17932 7531 17972 7540
rect 18028 8000 18068 8009
rect 17836 7120 17972 7160
rect 17836 6992 17876 7001
rect 17836 6488 17876 6952
rect 17836 6439 17876 6448
rect 17740 6320 17780 6329
rect 17452 4556 17492 4565
rect 17356 3464 17396 3473
rect 17356 3044 17396 3424
rect 17356 2995 17396 3004
rect 17452 2792 17492 4516
rect 17548 4220 17588 5692
rect 17644 5900 17684 5909
rect 17644 5396 17684 5860
rect 17644 5347 17684 5356
rect 17548 4171 17588 4180
rect 17644 4892 17684 4901
rect 17548 3212 17588 3221
rect 17548 2960 17588 3172
rect 17548 2911 17588 2920
rect 17452 2743 17492 2752
rect 17548 2792 17588 2801
rect 17356 2708 17396 2717
rect 17356 2288 17396 2668
rect 17356 2239 17396 2248
rect 17452 2624 17492 2633
rect 17452 2120 17492 2584
rect 17548 2624 17588 2752
rect 17644 2708 17684 4852
rect 17740 2876 17780 6280
rect 17932 5984 17972 7120
rect 17932 5935 17972 5944
rect 17932 4052 17972 4061
rect 17932 3464 17972 4012
rect 17932 3415 17972 3424
rect 17836 3380 17876 3389
rect 17836 3212 17876 3340
rect 17836 3163 17876 3172
rect 18028 2900 18068 7960
rect 18316 8000 18356 8009
rect 18220 7916 18260 7925
rect 18124 7580 18164 7589
rect 18124 6488 18164 7540
rect 18220 7580 18260 7876
rect 18220 7531 18260 7540
rect 18124 6439 18164 6448
rect 18220 7328 18260 7337
rect 18220 5480 18260 7288
rect 17740 2827 17780 2836
rect 17836 2876 17876 2885
rect 17644 2659 17684 2668
rect 17836 2708 17876 2836
rect 17836 2659 17876 2668
rect 17932 2860 18068 2900
rect 18124 5440 18260 5480
rect 17548 2575 17588 2584
rect 17740 2624 17780 2635
rect 17740 2540 17780 2584
rect 17740 2491 17780 2500
rect 16972 80 17012 1408
rect 17164 1408 17300 1448
rect 17356 2080 17492 2120
rect 17164 80 17204 1408
rect 17356 80 17396 2080
rect 17548 1784 17588 1793
rect 17548 80 17588 1744
rect 17740 1364 17780 1373
rect 17740 80 17780 1324
rect 17932 80 17972 2860
rect 18028 2708 18068 2717
rect 18028 2204 18068 2668
rect 18028 2155 18068 2164
rect 18028 1784 18068 1793
rect 18028 1649 18068 1744
rect 18124 80 18164 5440
rect 18220 5060 18260 5069
rect 18220 4388 18260 5020
rect 18220 4339 18260 4348
rect 18220 3548 18260 3557
rect 18220 2960 18260 3508
rect 18220 2911 18260 2920
rect 18316 2792 18356 7960
rect 18412 7916 18452 7925
rect 18412 7328 18452 7876
rect 18412 7279 18452 7288
rect 18508 7244 18548 8716
rect 18988 8756 19028 9388
rect 18988 8707 19028 8716
rect 19276 8756 19316 9976
rect 19276 8707 19316 8716
rect 19372 9260 19412 9269
rect 19372 9092 19412 9220
rect 18604 8672 18644 8681
rect 18604 8504 18644 8632
rect 18604 8455 18644 8464
rect 19276 8504 19316 8513
rect 18808 8336 19176 8345
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 18808 8287 19176 8296
rect 19084 8000 19124 8009
rect 19084 7865 19124 7960
rect 18988 7664 19028 7673
rect 19028 7624 19220 7664
rect 18988 7615 19028 7624
rect 19180 7580 19220 7624
rect 19180 7531 19220 7540
rect 18508 7195 18548 7204
rect 18700 7244 18740 7253
rect 18412 7160 18452 7169
rect 18412 6320 18452 7120
rect 18508 6824 18548 6833
rect 18508 6488 18548 6784
rect 18700 6656 18740 7204
rect 18808 6824 19176 6833
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 18808 6775 19176 6784
rect 18700 6607 18740 6616
rect 18508 6439 18548 6448
rect 18412 6271 18452 6280
rect 18604 6404 18644 6415
rect 18604 6320 18644 6364
rect 18604 6271 18644 6280
rect 19276 6404 19316 8464
rect 19372 7748 19412 9052
rect 19468 8924 19508 10144
rect 19468 8875 19508 8884
rect 19372 7699 19412 7708
rect 19468 8084 19508 8093
rect 18508 6152 18548 6161
rect 18412 6068 18452 6077
rect 18412 3212 18452 6028
rect 18508 6068 18548 6112
rect 18508 6017 18548 6028
rect 18700 5816 18740 5825
rect 18508 5732 18548 5741
rect 18508 5396 18548 5692
rect 18508 5347 18548 5356
rect 18604 5480 18644 5489
rect 18604 5144 18644 5440
rect 18700 5144 18740 5776
rect 18892 5732 18932 5741
rect 18892 5597 18932 5692
rect 18808 5312 19176 5321
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 18808 5263 19176 5272
rect 18796 5144 18836 5153
rect 19276 5144 19316 6364
rect 19372 7580 19412 7589
rect 19372 5312 19412 7540
rect 19372 5177 19412 5272
rect 18700 5104 18796 5144
rect 18604 5095 18644 5104
rect 18700 4976 18740 4985
rect 18604 4936 18700 4976
rect 18604 4640 18644 4936
rect 18700 4927 18740 4936
rect 18796 4892 18836 5104
rect 18796 4843 18836 4852
rect 19180 5104 19316 5144
rect 18508 3464 18548 3473
rect 18508 3329 18548 3424
rect 18412 3163 18452 3172
rect 18508 3212 18548 3221
rect 18412 3044 18452 3053
rect 18412 2792 18452 3004
rect 18508 2960 18548 3172
rect 18508 2911 18548 2920
rect 18604 2960 18644 4600
rect 19180 4304 19220 5104
rect 19180 4255 19220 4264
rect 19372 4472 19412 4481
rect 18700 4220 18740 4229
rect 18700 4085 18740 4180
rect 19276 4220 19316 4229
rect 18700 3800 18740 3809
rect 18700 3632 18740 3760
rect 18808 3800 19176 3809
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 18808 3751 19176 3760
rect 18892 3632 18932 3641
rect 18700 3592 18836 3632
rect 18796 3212 18836 3592
rect 18796 3163 18836 3172
rect 18892 3464 18932 3592
rect 18604 2911 18644 2920
rect 18700 3128 18740 3137
rect 18508 2792 18548 2801
rect 18412 2752 18508 2792
rect 18316 2743 18356 2752
rect 18508 2743 18548 2752
rect 18412 2624 18452 2633
rect 18452 2584 18644 2624
rect 18412 2575 18452 2584
rect 18220 2456 18260 2465
rect 18220 2372 18260 2416
rect 18220 2332 18548 2372
rect 18508 2204 18548 2332
rect 18508 2155 18548 2164
rect 18412 2120 18452 2129
rect 18220 1952 18260 1961
rect 18220 1868 18260 1912
rect 18220 1817 18260 1828
rect 18316 1280 18356 1289
rect 18316 80 18356 1240
rect 18412 1112 18452 2080
rect 18604 2120 18644 2584
rect 18604 2071 18644 2080
rect 18604 1868 18644 1877
rect 18604 1532 18644 1828
rect 18604 1483 18644 1492
rect 18412 1072 18548 1112
rect 18508 80 18548 1072
rect 18700 80 18740 3088
rect 18892 2960 18932 3424
rect 19180 3632 19220 3641
rect 18892 2911 18932 2920
rect 18988 3380 19028 3389
rect 18796 2876 18836 2885
rect 18796 2540 18836 2836
rect 18988 2876 19028 3340
rect 18988 2827 19028 2836
rect 19084 3212 19124 3221
rect 19084 2876 19124 3172
rect 19084 2827 19124 2836
rect 19180 2708 19220 3592
rect 19180 2659 19220 2668
rect 19276 2624 19316 4180
rect 19372 3212 19412 4432
rect 19468 4136 19508 8044
rect 19564 4892 19604 10648
rect 19660 8924 19700 12100
rect 20048 10604 20416 10613
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20048 10555 20416 10564
rect 20140 10436 20180 10445
rect 20140 10268 20180 10396
rect 20140 10219 20180 10228
rect 20716 10436 20756 10445
rect 19660 8875 19700 8884
rect 19948 10100 19988 10109
rect 19948 8756 19988 10060
rect 20044 10016 20084 10025
rect 20044 9428 20084 9976
rect 20140 9764 20180 9773
rect 20140 9629 20180 9724
rect 20620 9680 20660 9689
rect 20044 9379 20084 9388
rect 20048 9092 20416 9101
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20048 9043 20416 9052
rect 20620 9092 20660 9640
rect 20716 9512 20756 10396
rect 20812 9680 20852 12100
rect 21484 10772 21524 10781
rect 21292 10268 21332 10277
rect 21196 9848 21236 9857
rect 20812 9631 20852 9640
rect 20908 9764 20948 9773
rect 20716 9472 20852 9512
rect 20620 9043 20660 9052
rect 19948 8707 19988 8716
rect 20812 8756 20852 9472
rect 20908 9428 20948 9724
rect 20908 9379 20948 9388
rect 21004 9512 21044 9521
rect 19756 8000 19796 8009
rect 19660 7916 19700 7925
rect 19660 7412 19700 7876
rect 19660 7363 19700 7372
rect 19756 7412 19796 7960
rect 19756 7363 19796 7372
rect 19948 7748 19988 7757
rect 19660 6992 19700 7001
rect 19660 6404 19700 6952
rect 19756 6824 19796 6833
rect 19756 6656 19796 6784
rect 19756 6607 19796 6616
rect 19660 6355 19700 6364
rect 19852 6404 19892 6413
rect 19756 6320 19796 6329
rect 19756 6068 19796 6280
rect 19756 6019 19796 6028
rect 19852 5711 19892 6364
rect 19948 5816 19988 7708
rect 20716 7664 20756 7673
rect 20048 7580 20416 7589
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20048 7531 20416 7540
rect 20620 7496 20660 7505
rect 20236 7412 20276 7452
rect 20236 7328 20276 7372
rect 20044 7288 20276 7328
rect 20044 6320 20084 7288
rect 20236 7244 20276 7288
rect 20236 7195 20276 7204
rect 20140 7160 20180 7169
rect 20140 6824 20180 7120
rect 20140 6775 20180 6784
rect 20044 6271 20084 6280
rect 20524 6236 20564 6245
rect 20048 6068 20416 6077
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20048 6019 20416 6028
rect 19948 5767 19988 5776
rect 20236 5816 20276 5825
rect 20428 5816 20468 5825
rect 20276 5776 20428 5816
rect 20236 5767 20276 5776
rect 20428 5767 20468 5776
rect 19756 5671 19892 5711
rect 19604 4852 19700 4892
rect 19564 4843 19604 4852
rect 19660 4556 19700 4852
rect 19756 4556 19796 5671
rect 20140 5564 20180 5573
rect 20332 5564 20372 5573
rect 20180 5524 20332 5564
rect 20140 5515 20180 5524
rect 20332 5515 20372 5524
rect 20428 5480 20468 5489
rect 20140 5396 20180 5405
rect 20236 5396 20276 5405
rect 20180 5356 20236 5396
rect 20140 5328 20180 5356
rect 20236 5347 20276 5356
rect 20044 5312 20084 5321
rect 19948 4808 19988 4817
rect 19948 4556 19988 4768
rect 20044 4724 20084 5272
rect 20428 4976 20468 5440
rect 20524 5060 20564 6196
rect 20524 5011 20564 5020
rect 20332 4936 20468 4976
rect 20332 4892 20372 4936
rect 20332 4843 20372 4852
rect 20428 4808 20468 4817
rect 20468 4768 20564 4808
rect 20428 4759 20468 4768
rect 20044 4675 20084 4684
rect 19756 4516 19892 4556
rect 19660 4472 19700 4516
rect 19660 4432 19796 4472
rect 19660 4421 19700 4432
rect 19660 4304 19700 4313
rect 19564 4220 19604 4260
rect 19564 4136 19604 4180
rect 19508 4096 19604 4136
rect 19468 4087 19508 4096
rect 19372 3163 19412 3172
rect 19468 3968 19508 3977
rect 19276 2575 19316 2584
rect 18796 2491 18836 2500
rect 19276 2456 19316 2465
rect 18808 2288 19176 2297
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 18808 2239 19176 2248
rect 19276 2036 19316 2416
rect 19276 1987 19316 1996
rect 19372 1952 19412 1961
rect 19372 1868 19412 1912
rect 19372 1817 19412 1828
rect 18892 1280 18932 1289
rect 18892 80 18932 1240
rect 19276 1112 19316 1121
rect 19084 608 19124 617
rect 19084 80 19124 568
rect 19276 80 19316 1072
rect 19468 80 19508 3928
rect 19564 3632 19604 4096
rect 19564 3583 19604 3592
rect 19660 80 19700 4264
rect 19756 4220 19796 4432
rect 19756 4171 19796 4180
rect 19756 3044 19796 3053
rect 19756 2960 19796 3004
rect 19756 2909 19796 2920
rect 19852 80 19892 4516
rect 19948 4507 19988 4516
rect 20048 4556 20416 4565
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20048 4507 20416 4516
rect 20524 4556 20564 4768
rect 20524 4507 20564 4516
rect 20620 4472 20660 7456
rect 20716 6824 20756 7624
rect 20716 6775 20756 6784
rect 20716 6488 20756 6497
rect 20716 4640 20756 6448
rect 20716 4591 20756 4600
rect 20812 5732 20852 8716
rect 20908 9092 20948 9101
rect 20908 6572 20948 9052
rect 21004 8084 21044 9472
rect 21004 8035 21044 8044
rect 21100 9176 21140 9185
rect 20908 6523 20948 6532
rect 21004 7916 21044 7925
rect 21004 6404 21044 7876
rect 21004 5816 21044 6364
rect 21004 5767 21044 5776
rect 20812 5228 20852 5692
rect 20620 4432 20756 4472
rect 20140 4304 20180 4313
rect 20332 4304 20372 4313
rect 20180 4264 20332 4304
rect 20140 4255 20180 4264
rect 20332 4255 20372 4264
rect 20620 4304 20660 4315
rect 19948 4220 19988 4229
rect 19948 3296 19988 4180
rect 20620 4220 20660 4264
rect 20620 4171 20660 4180
rect 20332 4052 20372 4061
rect 20236 3968 20276 3977
rect 20236 3548 20276 3928
rect 20236 3499 20276 3508
rect 20140 3464 20180 3473
rect 20140 3380 20180 3424
rect 20332 3380 20372 4012
rect 20620 4052 20660 4061
rect 20140 3340 20372 3380
rect 20524 3380 20564 3389
rect 19948 3247 19988 3256
rect 19948 3044 19988 3053
rect 19948 1364 19988 3004
rect 20048 3044 20416 3053
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20048 2995 20416 3004
rect 20044 2876 20084 2885
rect 20044 1784 20084 2836
rect 20236 2708 20276 2717
rect 20236 2120 20276 2668
rect 20524 2456 20564 3340
rect 20524 2288 20564 2416
rect 20524 2239 20564 2248
rect 20236 2071 20276 2080
rect 20044 1735 20084 1744
rect 20048 1532 20416 1541
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20048 1483 20416 1492
rect 20428 1364 20468 1373
rect 19948 1324 20276 1364
rect 20044 1028 20084 1037
rect 20044 80 20084 988
rect 20236 80 20276 1324
rect 20428 80 20468 1324
rect 20620 80 20660 4012
rect 20716 3632 20756 4432
rect 20812 4052 20852 5188
rect 20908 5648 20948 5657
rect 20908 4808 20948 5608
rect 21004 5312 21044 5321
rect 21004 5144 21044 5272
rect 21004 5095 21044 5104
rect 20908 4759 20948 4768
rect 20812 4003 20852 4012
rect 21004 4304 21044 4313
rect 21004 3800 21044 4264
rect 21004 3751 21044 3760
rect 20716 3592 21044 3632
rect 20908 3212 20948 3221
rect 20908 2288 20948 3172
rect 20908 2239 20948 2248
rect 21004 2036 21044 3592
rect 21100 2708 21140 9136
rect 21196 9008 21236 9808
rect 21292 9092 21332 10228
rect 21484 10268 21524 10732
rect 21484 10219 21524 10228
rect 21868 10268 21908 10277
rect 21868 9848 21908 10228
rect 21772 9596 21812 9605
rect 21292 9043 21332 9052
rect 21484 9428 21524 9437
rect 21196 8959 21236 8968
rect 21484 9008 21524 9388
rect 21580 9344 21620 9353
rect 21580 9092 21620 9304
rect 21772 9344 21812 9556
rect 21772 9295 21812 9304
rect 21772 9092 21812 9101
rect 21580 9052 21772 9092
rect 21772 9043 21812 9052
rect 21484 8959 21524 8968
rect 21868 8840 21908 9808
rect 21964 9596 22004 12100
rect 21964 9547 22004 9556
rect 22156 9596 22196 9605
rect 22060 9512 22100 9521
rect 22060 9344 22100 9472
rect 22156 9461 22196 9556
rect 22252 9512 22292 9521
rect 22060 9295 22100 9304
rect 22060 9092 22100 9101
rect 21868 8791 21908 8800
rect 21964 8924 22004 8933
rect 21676 8756 21716 8765
rect 21388 8672 21428 8681
rect 21196 7496 21236 7505
rect 21196 6656 21236 7456
rect 21292 7496 21332 7505
rect 21292 7328 21332 7456
rect 21292 7279 21332 7288
rect 21196 6607 21236 6616
rect 21388 6572 21428 8632
rect 21676 8588 21716 8716
rect 21580 7748 21620 7757
rect 21484 7328 21524 7337
rect 21484 7244 21524 7288
rect 21484 7193 21524 7204
rect 21388 6523 21428 6532
rect 21484 7076 21524 7085
rect 21196 6320 21236 6329
rect 21196 5648 21236 6280
rect 21484 6320 21524 7036
rect 21484 6271 21524 6280
rect 21580 5732 21620 7708
rect 21580 5683 21620 5692
rect 21196 5599 21236 5608
rect 21676 4892 21716 8548
rect 21964 8084 22004 8884
rect 21868 8044 22004 8084
rect 22060 8672 22100 9052
rect 21772 8000 21812 8009
rect 21772 7865 21812 7960
rect 21772 7580 21812 7675
rect 21772 7531 21812 7540
rect 21772 7412 21812 7421
rect 21772 7277 21812 7372
rect 21868 6236 21908 8044
rect 21964 7916 22004 7925
rect 21964 6320 22004 7876
rect 22060 7412 22100 8632
rect 22156 7748 22196 7757
rect 22156 7580 22196 7708
rect 22156 7531 22196 7540
rect 22252 7412 22292 9472
rect 22732 9344 22772 9353
rect 22540 8420 22580 8429
rect 22060 7372 22196 7412
rect 22060 7244 22100 7253
rect 22060 6824 22100 7204
rect 22156 6992 22196 7372
rect 22252 7160 22292 7372
rect 22348 7412 22388 7421
rect 22348 7328 22388 7372
rect 22348 7277 22388 7288
rect 22252 7111 22292 7120
rect 22444 7244 22484 7253
rect 22444 7109 22484 7204
rect 22156 6952 22388 6992
rect 22060 6775 22100 6784
rect 21964 6271 22004 6280
rect 22060 6488 22100 6497
rect 21868 6187 21908 6196
rect 22060 6068 22100 6448
rect 22060 6019 22100 6028
rect 22348 6488 22388 6952
rect 22252 5816 22292 5825
rect 22156 5732 22196 5741
rect 21676 4843 21716 4852
rect 21772 5396 21812 5405
rect 21388 4808 21428 4817
rect 21292 4640 21332 4649
rect 21196 4220 21236 4229
rect 21196 4085 21236 4180
rect 21196 3968 21236 3977
rect 21196 3716 21236 3928
rect 21196 3667 21236 3676
rect 21100 2659 21140 2668
rect 21292 2624 21332 4600
rect 21388 4052 21428 4768
rect 21388 4012 21620 4052
rect 21484 3296 21524 3305
rect 21484 3212 21524 3256
rect 21484 3161 21524 3172
rect 21292 2575 21332 2584
rect 21004 1987 21044 1996
rect 21388 2372 21428 2381
rect 20812 1784 20852 1793
rect 20716 1616 20756 1625
rect 20716 1481 20756 1576
rect 20812 80 20852 1744
rect 21196 1616 21236 1625
rect 21196 80 21236 1576
rect 21388 80 21428 2332
rect 21580 2372 21620 4012
rect 21676 3800 21716 3809
rect 21676 2960 21716 3760
rect 21676 2911 21716 2920
rect 21580 2323 21620 2332
rect 21676 2708 21716 2717
rect 21676 2372 21716 2668
rect 21676 2323 21716 2332
rect 21676 2204 21716 2213
rect 21580 1868 21620 1877
rect 21484 1784 21524 1793
rect 21484 1448 21524 1744
rect 21580 1733 21620 1828
rect 21484 1399 21524 1408
rect 21580 1364 21620 1373
rect 21580 80 21620 1324
rect 21676 1280 21716 2164
rect 21772 1448 21812 5356
rect 21964 5228 22004 5237
rect 21964 5060 22004 5188
rect 21964 4892 22004 5020
rect 21964 4843 22004 4852
rect 21868 4640 21908 4649
rect 21868 4220 21908 4600
rect 21868 4171 21908 4180
rect 21964 4556 22004 4565
rect 21964 4052 22004 4516
rect 22156 4388 22196 5692
rect 22252 5648 22292 5776
rect 22252 5599 22292 5608
rect 22156 4339 22196 4348
rect 22252 5396 22292 5405
rect 21964 4003 22004 4012
rect 22156 4220 22196 4229
rect 22060 3632 22100 3641
rect 21964 3380 22004 3389
rect 21868 3212 21908 3221
rect 21868 2876 21908 3172
rect 21964 2960 22004 3340
rect 21964 2911 22004 2920
rect 21868 2827 21908 2836
rect 21964 2792 22004 2803
rect 21964 2708 22004 2752
rect 21964 2659 22004 2668
rect 22060 1952 22100 3592
rect 22156 3212 22196 4180
rect 22156 3163 22196 3172
rect 22060 1903 22100 1912
rect 22156 3044 22196 3053
rect 21772 1408 22004 1448
rect 21676 1240 21812 1280
rect 21772 80 21812 1240
rect 21964 80 22004 1408
rect 22156 80 22196 3004
rect 22252 1448 22292 5356
rect 22348 5396 22388 6448
rect 22540 5816 22580 8380
rect 22636 7496 22676 7505
rect 22636 7328 22676 7456
rect 22636 7279 22676 7288
rect 22540 5767 22580 5776
rect 22732 7244 22772 9304
rect 23116 8168 23156 12100
rect 24268 10436 24308 12100
rect 24268 10387 24308 10396
rect 24172 10268 24212 10277
rect 23308 10016 23348 10025
rect 23308 9428 23348 9976
rect 23308 9379 23348 9388
rect 23980 8924 24020 8933
rect 23116 8119 23156 8128
rect 23404 8420 23444 8429
rect 22924 8084 22964 8093
rect 22924 7496 22964 8044
rect 23116 8000 23156 8011
rect 23116 7916 23156 7960
rect 23404 8000 23444 8380
rect 23500 8420 23540 8429
rect 23500 8084 23540 8380
rect 23500 8035 23540 8044
rect 23404 7951 23444 7960
rect 23788 8000 23828 8009
rect 23116 7867 23156 7876
rect 22924 7447 22964 7456
rect 22348 4136 22388 5356
rect 22444 5060 22484 5069
rect 22444 4220 22484 5020
rect 22444 4171 22484 4180
rect 22636 4892 22676 4901
rect 22348 4087 22388 4096
rect 22540 3128 22580 3137
rect 22348 2792 22388 2801
rect 22348 2036 22388 2752
rect 22444 2792 22484 2801
rect 22444 2288 22484 2752
rect 22444 2239 22484 2248
rect 22348 1987 22388 1996
rect 22252 1408 22388 1448
rect 22348 80 22388 1408
rect 22540 80 22580 3088
rect 22636 2372 22676 4852
rect 22732 4808 22772 7204
rect 22732 4759 22772 4768
rect 22828 7412 22868 7421
rect 22828 3968 22868 7372
rect 23788 7412 23828 7960
rect 23788 7363 23828 7372
rect 23500 7244 23540 7253
rect 23404 7160 23444 7169
rect 23212 7076 23252 7085
rect 22924 6740 22964 6749
rect 22924 6404 22964 6700
rect 22924 6320 22964 6364
rect 23212 6404 23252 7036
rect 23212 6355 23252 6364
rect 23308 6656 23348 6665
rect 22924 6271 22964 6280
rect 23212 5900 23252 5909
rect 23212 5732 23252 5860
rect 23212 5683 23252 5692
rect 23212 4388 23252 4397
rect 22828 3919 22868 3928
rect 23020 3968 23060 3977
rect 23020 3632 23060 3928
rect 23020 3583 23060 3592
rect 23212 3380 23252 4348
rect 23212 3331 23252 3340
rect 22828 3296 22868 3305
rect 22732 2876 22772 2885
rect 22732 2792 22772 2836
rect 22732 2741 22772 2752
rect 22636 2323 22676 2332
rect 22732 2540 22772 2549
rect 22732 80 22772 2500
rect 22828 1868 22868 3256
rect 22924 3212 22964 3221
rect 22924 2792 22964 3172
rect 23116 3044 23156 3053
rect 23116 2876 23156 3004
rect 23116 2827 23156 2836
rect 22924 2708 22964 2752
rect 23212 2792 23252 2801
rect 22924 2657 22964 2668
rect 23020 2708 23060 2717
rect 23116 2708 23156 2717
rect 23060 2668 23116 2708
rect 23020 2659 23060 2668
rect 23116 2659 23156 2668
rect 23116 2540 23156 2549
rect 22828 1819 22868 1828
rect 22924 2456 22964 2465
rect 22924 80 22964 2416
rect 23020 2204 23060 2213
rect 23116 2204 23156 2500
rect 23060 2164 23156 2204
rect 23212 2204 23252 2752
rect 23308 2624 23348 6616
rect 23404 4220 23444 7120
rect 23500 6656 23540 7204
rect 23500 6607 23540 6616
rect 23884 6236 23924 6245
rect 23884 5816 23924 6196
rect 23884 5767 23924 5776
rect 23788 5480 23828 5489
rect 23788 5345 23828 5440
rect 23980 5060 24020 8884
rect 24076 8756 24116 8765
rect 24076 5732 24116 8716
rect 24172 7916 24212 10228
rect 25036 10268 25076 10277
rect 24940 9596 24980 9605
rect 24652 9428 24692 9437
rect 24364 9344 24404 9353
rect 24364 8924 24404 9304
rect 24364 8875 24404 8884
rect 24652 8756 24692 9388
rect 24652 8707 24692 8716
rect 24748 9092 24788 9101
rect 24172 7867 24212 7876
rect 24364 8504 24404 8513
rect 24268 7580 24308 7589
rect 24172 6068 24212 6077
rect 24172 5816 24212 6028
rect 24172 5767 24212 5776
rect 24076 5683 24116 5692
rect 23980 4892 24020 5020
rect 23980 4843 24020 4852
rect 24172 5312 24212 5321
rect 23404 4171 23444 4180
rect 23884 4472 23924 4481
rect 23884 4220 23924 4432
rect 23884 4171 23924 4180
rect 23308 2575 23348 2584
rect 23500 3968 23540 3977
rect 23020 2155 23060 2164
rect 23212 2155 23252 2164
rect 23308 2120 23348 2129
rect 23116 2036 23156 2045
rect 23116 80 23156 1996
rect 23308 1868 23348 2080
rect 23308 1819 23348 1828
rect 23308 1616 23348 1625
rect 23308 80 23348 1576
rect 23500 80 23540 3928
rect 23884 3968 23924 3977
rect 23692 3464 23732 3473
rect 23692 2876 23732 3424
rect 23692 2827 23732 2836
rect 23692 1700 23732 1709
rect 23692 80 23732 1660
rect 23884 80 23924 3928
rect 24172 2792 24212 5272
rect 24268 4136 24308 7540
rect 24364 6152 24404 8464
rect 24652 7832 24692 7841
rect 24364 6103 24404 6112
rect 24460 7412 24500 7421
rect 24268 4087 24308 4096
rect 24364 5732 24404 5741
rect 24364 3968 24404 5692
rect 24460 5564 24500 7372
rect 24460 5515 24500 5524
rect 24556 7244 24596 7253
rect 24556 6320 24596 7204
rect 24556 4976 24596 6280
rect 24556 4927 24596 4936
rect 24556 4304 24596 4313
rect 24460 3968 24500 3977
rect 24364 3928 24460 3968
rect 24460 3632 24500 3928
rect 24460 3583 24500 3592
rect 24364 3548 24404 3557
rect 24172 2743 24212 2752
rect 24268 3212 24308 3221
rect 24076 2372 24116 2381
rect 24076 80 24116 2332
rect 24268 80 24308 3172
rect 24364 3044 24404 3508
rect 24556 3548 24596 4264
rect 24556 3499 24596 3508
rect 24460 3296 24500 3305
rect 24460 3212 24500 3256
rect 24460 3161 24500 3172
rect 24364 2995 24404 3004
rect 24556 2708 24596 2717
rect 24460 2456 24500 2465
rect 24460 80 24500 2416
rect 24556 2036 24596 2668
rect 24652 2624 24692 7792
rect 24748 3464 24788 9052
rect 24940 8924 24980 9556
rect 24940 8875 24980 8884
rect 24940 8756 24980 8765
rect 24940 8000 24980 8716
rect 25036 8756 25076 10228
rect 25132 9932 25172 9941
rect 25132 9092 25172 9892
rect 25420 9680 25460 12100
rect 25420 9631 25460 9640
rect 25612 10604 25652 10613
rect 25420 9428 25460 9437
rect 25420 9293 25460 9388
rect 25132 9043 25172 9052
rect 25036 8707 25076 8716
rect 24940 5144 24980 7960
rect 25420 8336 25460 8345
rect 25420 7916 25460 8296
rect 25420 7867 25460 7876
rect 25132 7496 25172 7505
rect 24940 5095 24980 5104
rect 25036 6320 25076 6329
rect 24844 4304 24884 4313
rect 24844 4136 24884 4264
rect 25036 4136 25076 6280
rect 25132 5648 25172 7456
rect 25132 5599 25172 5608
rect 25516 5816 25556 5825
rect 25516 5732 25556 5776
rect 25420 5564 25460 5573
rect 24844 4087 24884 4096
rect 24940 4096 25036 4136
rect 24748 3415 24788 3424
rect 24844 3548 24884 3557
rect 24844 3380 24884 3508
rect 24844 3331 24884 3340
rect 24844 2708 24884 2717
rect 24748 2624 24788 2633
rect 24652 2584 24748 2624
rect 24556 1987 24596 1996
rect 24652 2372 24692 2381
rect 24652 1784 24692 2332
rect 24748 2120 24788 2584
rect 24844 2624 24884 2668
rect 24844 2573 24884 2584
rect 24748 2071 24788 2080
rect 24940 1952 24980 4096
rect 25036 4087 25076 4096
rect 25132 5312 25172 5321
rect 25132 4892 25172 5272
rect 24940 1903 24980 1912
rect 25036 3884 25076 3893
rect 24556 1744 24692 1784
rect 24940 1784 24980 1793
rect 24556 1532 24596 1744
rect 24556 1483 24596 1492
rect 24652 1616 24692 1625
rect 24652 80 24692 1576
rect 24940 1616 24980 1744
rect 24940 1567 24980 1576
rect 24844 1532 24884 1541
rect 24844 80 24884 1492
rect 25036 80 25076 3844
rect 25132 2540 25172 4852
rect 25420 4724 25460 5524
rect 25516 5396 25556 5692
rect 25516 5347 25556 5356
rect 25420 4675 25460 4684
rect 25516 4556 25556 4565
rect 25516 4472 25556 4516
rect 25516 4421 25556 4432
rect 25612 4388 25652 10564
rect 26572 10436 26612 12100
rect 26572 10387 26612 10396
rect 27532 10688 27572 10697
rect 26860 10352 26900 10361
rect 25804 10268 25844 10277
rect 25804 8840 25844 10228
rect 25900 10100 25940 10109
rect 26860 10100 26900 10312
rect 25900 9428 25940 10060
rect 26764 10060 26900 10100
rect 27340 10100 27380 10109
rect 26476 9596 26516 9607
rect 26476 9512 26516 9556
rect 26476 9463 26516 9472
rect 25900 9379 25940 9388
rect 26284 9428 26324 9437
rect 25900 9260 25940 9269
rect 25940 9220 26036 9260
rect 25900 9211 25940 9220
rect 25804 8791 25844 8800
rect 25996 8840 26036 9220
rect 25996 8791 26036 8800
rect 25708 8756 25748 8765
rect 25708 7160 25748 8716
rect 26188 8084 26228 8093
rect 26092 7916 26132 7925
rect 25900 7748 25940 7757
rect 25708 6488 25748 7120
rect 25804 7496 25844 7505
rect 25804 6656 25844 7456
rect 25804 6607 25844 6616
rect 25708 6404 25748 6448
rect 25708 6355 25748 6364
rect 25804 5816 25844 5825
rect 25708 5648 25748 5657
rect 25708 4892 25748 5608
rect 25708 4843 25748 4852
rect 25708 4388 25748 4397
rect 25612 4348 25708 4388
rect 25228 4052 25268 4147
rect 25228 4003 25268 4012
rect 25612 4136 25652 4145
rect 25132 2491 25172 2500
rect 25228 3800 25268 3809
rect 25228 80 25268 3760
rect 25612 3380 25652 4096
rect 25612 3331 25652 3340
rect 25612 3212 25652 3221
rect 25324 2708 25364 2717
rect 25324 1784 25364 2668
rect 25612 2708 25652 3172
rect 25708 3212 25748 4348
rect 25804 3800 25844 5776
rect 25900 4136 25940 7708
rect 26092 6824 26132 7876
rect 26188 7160 26228 8044
rect 26284 7916 26324 9388
rect 26284 7867 26324 7876
rect 26572 9008 26612 9017
rect 26476 7832 26516 7841
rect 26284 7748 26324 7757
rect 26284 7580 26324 7708
rect 26284 7531 26324 7540
rect 26188 7111 26228 7120
rect 26092 6775 26132 6784
rect 26380 6404 26420 6413
rect 26284 6236 26324 6245
rect 25996 5900 26036 5909
rect 25996 5732 26036 5860
rect 25996 5683 26036 5692
rect 26188 5144 26228 5153
rect 26188 5009 26228 5104
rect 25900 4087 25940 4096
rect 25996 4724 26036 4733
rect 25804 3751 25844 3760
rect 25708 3163 25748 3172
rect 25612 2659 25652 2668
rect 25900 3128 25940 3137
rect 25900 2708 25940 3088
rect 25900 2659 25940 2668
rect 25708 2540 25748 2549
rect 25708 2120 25748 2500
rect 25324 1735 25364 1744
rect 25420 2036 25460 2045
rect 25420 80 25460 1996
rect 25708 1868 25748 2080
rect 25708 1819 25748 1828
rect 25804 1616 25844 1625
rect 25612 1448 25652 1457
rect 25612 80 25652 1408
rect 25804 80 25844 1576
rect 25996 80 26036 4684
rect 26188 4640 26228 4649
rect 26092 4556 26132 4565
rect 26092 3716 26132 4516
rect 26092 3667 26132 3676
rect 26188 80 26228 4600
rect 26284 4220 26324 6196
rect 26380 5060 26420 6364
rect 26476 5228 26516 7792
rect 26572 6152 26612 8968
rect 26668 8504 26708 8513
rect 26668 7916 26708 8464
rect 26668 7867 26708 7876
rect 26764 6656 26804 10060
rect 27052 10016 27092 10025
rect 26956 9932 26996 9941
rect 26956 9512 26996 9892
rect 26956 9463 26996 9472
rect 27052 8756 27092 9976
rect 27340 9512 27380 10060
rect 27340 9463 27380 9472
rect 27052 8707 27092 8716
rect 27436 9344 27476 9353
rect 27148 8000 27188 8009
rect 27148 7832 27188 7960
rect 27148 7783 27188 7792
rect 27436 8000 27476 9304
rect 27436 7412 27476 7960
rect 27436 7363 27476 7372
rect 27340 7244 27380 7253
rect 26572 6103 26612 6112
rect 26668 6616 26804 6656
rect 26860 6992 26900 7001
rect 26476 5179 26516 5188
rect 26668 5984 26708 6616
rect 26860 6320 26900 6952
rect 27340 6404 27380 7204
rect 27340 6355 27380 6364
rect 27436 6740 27476 6749
rect 26860 6271 26900 6280
rect 26420 5020 26516 5060
rect 26380 5011 26420 5020
rect 26284 4171 26324 4180
rect 26380 4388 26420 4397
rect 26284 3212 26324 3221
rect 26284 1868 26324 3172
rect 26284 1819 26324 1828
rect 26380 80 26420 4348
rect 26476 3716 26516 5020
rect 26668 4220 26708 5944
rect 26860 6152 26900 6161
rect 26764 5900 26804 5909
rect 26764 5732 26804 5860
rect 26764 5683 26804 5692
rect 26668 4171 26708 4180
rect 26764 5480 26804 5489
rect 26476 3667 26516 3676
rect 26572 4052 26612 4061
rect 26572 3632 26612 4012
rect 26572 3583 26612 3592
rect 26668 3464 26708 3473
rect 26476 3212 26516 3221
rect 26476 2960 26516 3172
rect 26476 2911 26516 2920
rect 26668 2876 26708 3424
rect 26668 2827 26708 2836
rect 26572 692 26612 701
rect 26572 80 26612 652
rect 26764 80 26804 5440
rect 26860 2900 26900 6112
rect 27436 6068 27476 6700
rect 27436 6019 27476 6028
rect 27148 5648 27188 5657
rect 27052 5396 27092 5405
rect 26956 5228 26996 5237
rect 26956 4640 26996 5188
rect 26956 4591 26996 4600
rect 27052 4388 27092 5356
rect 27148 5144 27188 5608
rect 27148 5095 27188 5104
rect 27340 4976 27380 4985
rect 27340 4556 27380 4936
rect 27532 4976 27572 10648
rect 27724 10436 27764 12100
rect 28012 11024 28052 11033
rect 28012 10604 28052 10984
rect 28012 10555 28052 10564
rect 28108 10772 28148 10781
rect 27724 10387 27764 10396
rect 28108 10268 28148 10732
rect 28876 10436 28916 12100
rect 28876 10387 28916 10396
rect 29260 11024 29300 11033
rect 29260 10688 29300 10984
rect 28108 10219 28148 10228
rect 27628 10100 27668 10109
rect 27628 10016 27668 10060
rect 27628 9965 27668 9976
rect 27820 9512 27860 9521
rect 27820 8924 27860 9472
rect 28396 9428 28436 9437
rect 27916 9344 27956 9353
rect 27916 9008 27956 9304
rect 28396 9293 28436 9388
rect 27916 8959 27956 8968
rect 29068 9260 29108 9269
rect 27820 8875 27860 8884
rect 28012 8756 28052 8765
rect 28012 8621 28052 8716
rect 28300 8756 28340 8765
rect 28300 8336 28340 8716
rect 28972 8756 29012 8765
rect 28012 8084 28052 8093
rect 28012 6656 28052 8044
rect 28204 7748 28244 7757
rect 28204 7412 28244 7708
rect 28300 7664 28340 8296
rect 28492 8504 28532 8513
rect 28492 7916 28532 8464
rect 28588 8336 28628 8345
rect 28588 8000 28628 8296
rect 28588 7951 28628 7960
rect 28780 8252 28820 8261
rect 28492 7867 28532 7876
rect 28300 7615 28340 7624
rect 28204 7363 28244 7372
rect 28780 7244 28820 8212
rect 28780 7195 28820 7204
rect 28684 7160 28724 7169
rect 28012 6607 28052 6616
rect 28108 6656 28148 6665
rect 27724 6068 27764 6077
rect 27724 5648 27764 6028
rect 27724 5599 27764 5608
rect 28108 5648 28148 6616
rect 28108 5599 28148 5608
rect 28204 6404 28244 6413
rect 27532 4927 27572 4936
rect 27820 5396 27860 5405
rect 27340 4507 27380 4516
rect 27628 4892 27668 4901
rect 27052 4339 27092 4348
rect 27340 4304 27380 4313
rect 27244 4220 27284 4229
rect 27052 4180 27244 4220
rect 27052 4136 27092 4180
rect 27244 4171 27284 4180
rect 27340 4169 27380 4264
rect 27052 4087 27092 4096
rect 27148 3968 27188 3977
rect 26956 3716 26996 3725
rect 26956 3632 26996 3676
rect 26956 3581 26996 3592
rect 27052 3716 27092 3725
rect 27052 3380 27092 3676
rect 27052 3331 27092 3340
rect 26860 2860 26996 2900
rect 26956 1952 26996 2860
rect 26956 1903 26996 1912
rect 26956 860 26996 869
rect 26956 80 26996 820
rect 27148 80 27188 3928
rect 27244 3464 27284 3473
rect 27244 2120 27284 3424
rect 27244 2071 27284 2080
rect 27436 3212 27476 3221
rect 27436 1952 27476 3172
rect 27436 1903 27476 1912
rect 27628 2708 27668 4852
rect 27628 1952 27668 2668
rect 27628 1903 27668 1912
rect 27532 1868 27572 1877
rect 27340 1448 27380 1457
rect 27340 80 27380 1408
rect 27532 1364 27572 1828
rect 27724 1868 27764 1877
rect 27724 1733 27764 1828
rect 27532 1315 27572 1324
rect 27820 1028 27860 5356
rect 27532 988 27860 1028
rect 27916 5312 27956 5321
rect 27532 80 27572 988
rect 27724 860 27764 869
rect 27724 80 27764 820
rect 27916 80 27956 5272
rect 28108 4892 28148 4901
rect 28108 4388 28148 4852
rect 28108 4339 28148 4348
rect 28204 3632 28244 6364
rect 28204 3583 28244 3592
rect 28300 6320 28340 6329
rect 28204 3380 28244 3389
rect 28204 3128 28244 3340
rect 28204 3079 28244 3088
rect 28108 944 28148 953
rect 28108 80 28148 904
rect 28300 80 28340 6280
rect 28492 6236 28532 6245
rect 28396 5480 28436 5489
rect 28396 5345 28436 5440
rect 28396 4388 28436 4397
rect 28396 2708 28436 4348
rect 28396 2659 28436 2668
rect 28492 80 28532 6196
rect 28588 5564 28628 5573
rect 28588 5060 28628 5524
rect 28684 5228 28724 7120
rect 28780 6488 28820 6497
rect 28780 6068 28820 6448
rect 28780 6019 28820 6028
rect 28684 5179 28724 5188
rect 28876 5480 28916 5489
rect 28876 5228 28916 5440
rect 28876 5179 28916 5188
rect 28588 4220 28628 5020
rect 28780 5144 28820 5153
rect 28684 4892 28724 4901
rect 28684 4472 28724 4852
rect 28684 4337 28724 4432
rect 28780 4388 28820 5104
rect 28876 4976 28916 4987
rect 28876 4892 28916 4936
rect 28876 4843 28916 4852
rect 28780 4339 28820 4348
rect 28876 4724 28916 4733
rect 28588 4171 28628 4180
rect 28780 4220 28820 4229
rect 28684 3800 28724 3809
rect 28588 2792 28628 2801
rect 28588 2624 28628 2752
rect 28588 2575 28628 2584
rect 28684 80 28724 3760
rect 28780 3380 28820 4180
rect 28780 3331 28820 3340
rect 28780 2708 28820 2717
rect 28780 2456 28820 2668
rect 28780 2407 28820 2416
rect 28876 80 28916 4684
rect 28972 2036 29012 8716
rect 29068 8672 29108 9220
rect 29068 8623 29108 8632
rect 29260 8504 29300 10648
rect 29452 10688 29492 10697
rect 29452 10184 29492 10648
rect 30028 10436 30068 12100
rect 30028 10387 30068 10396
rect 31180 10352 31220 12100
rect 31180 10303 31220 10312
rect 29452 10135 29492 10144
rect 29644 10268 29684 10277
rect 29452 10016 29492 10025
rect 29452 9512 29492 9976
rect 29644 10016 29684 10228
rect 30700 10268 30740 10277
rect 29548 9512 29588 9521
rect 29452 9472 29548 9512
rect 29548 9463 29588 9472
rect 29548 9344 29588 9353
rect 29644 9344 29684 9976
rect 29588 9304 29684 9344
rect 29740 10016 29780 10025
rect 29260 8455 29300 8464
rect 29452 8588 29492 8597
rect 29452 8000 29492 8548
rect 29452 7951 29492 7960
rect 28972 1987 29012 1996
rect 29068 7748 29108 7757
rect 29068 80 29108 7708
rect 29452 7748 29492 7757
rect 29260 5648 29300 5657
rect 29260 4640 29300 5608
rect 29260 4591 29300 4600
rect 29356 4892 29396 4901
rect 29164 3632 29204 3641
rect 29164 3464 29204 3592
rect 29164 3415 29204 3424
rect 29260 3380 29300 3389
rect 29260 2960 29300 3340
rect 29356 3044 29396 4852
rect 29356 2995 29396 3004
rect 29164 2708 29204 2717
rect 29164 2456 29204 2668
rect 29164 2204 29204 2416
rect 29164 2155 29204 2164
rect 29260 2120 29300 2920
rect 29260 2071 29300 2080
rect 29356 2708 29396 2717
rect 29356 2120 29396 2668
rect 29356 2071 29396 2080
rect 29164 2036 29204 2045
rect 29164 1901 29204 1996
rect 29260 1784 29300 1793
rect 29260 80 29300 1744
rect 29452 80 29492 7708
rect 29548 6320 29588 9304
rect 29644 8840 29684 8849
rect 29644 6488 29684 8800
rect 29740 8756 29780 9976
rect 29740 8707 29780 8716
rect 30220 8756 30260 8765
rect 30508 8756 30548 8765
rect 30260 8716 30452 8756
rect 30220 8707 30260 8716
rect 30412 8588 30452 8716
rect 29644 6439 29684 6448
rect 29836 8504 29876 8513
rect 29740 6404 29780 6413
rect 29548 6280 29684 6320
rect 29548 5564 29588 5573
rect 29548 4556 29588 5524
rect 29548 4507 29588 4516
rect 29644 4304 29684 6280
rect 29740 5816 29780 6364
rect 29740 5767 29780 5776
rect 29740 5480 29780 5489
rect 29740 4556 29780 5440
rect 29740 4507 29780 4516
rect 29644 4255 29684 4264
rect 29740 4388 29780 4397
rect 29644 2876 29684 2885
rect 29644 2792 29684 2836
rect 29644 2741 29684 2752
rect 29740 1952 29780 4348
rect 29836 3716 29876 8464
rect 30028 8504 30068 8513
rect 30028 7832 30068 8464
rect 30412 7916 30452 8548
rect 30508 8084 30548 8716
rect 30508 8035 30548 8044
rect 30028 7783 30068 7792
rect 30316 7832 30356 7841
rect 29932 7580 29972 7589
rect 29932 6404 29972 7540
rect 30220 7580 30260 7589
rect 30220 7445 30260 7540
rect 30316 7412 30356 7792
rect 30316 7363 30356 7372
rect 29932 4220 29972 6364
rect 30028 7244 30068 7253
rect 30028 6656 30068 7204
rect 30412 6992 30452 7876
rect 30412 6943 30452 6952
rect 30508 7412 30548 7421
rect 30508 7244 30548 7372
rect 30220 6656 30260 6665
rect 30028 6404 30068 6616
rect 30028 6355 30068 6364
rect 30124 6616 30220 6656
rect 30124 6404 30164 6616
rect 30220 6588 30260 6616
rect 30508 6488 30548 7204
rect 30508 6439 30548 6448
rect 30604 6992 30644 7001
rect 30124 6355 30164 6364
rect 30316 6320 30356 6329
rect 30124 6236 30164 6245
rect 30316 6236 30356 6280
rect 30164 6196 30356 6236
rect 30124 6187 30164 6196
rect 30124 6068 30164 6077
rect 30164 6028 30260 6068
rect 30124 6019 30164 6028
rect 30220 5144 30260 6028
rect 30316 5732 30356 5741
rect 30316 5564 30356 5692
rect 30508 5648 30548 5657
rect 30316 5515 30356 5524
rect 30412 5608 30508 5648
rect 30412 5396 30452 5608
rect 30508 5599 30548 5608
rect 30412 5347 30452 5356
rect 30508 5480 30548 5489
rect 30508 5345 30548 5440
rect 30316 5144 30356 5153
rect 30220 5104 30316 5144
rect 30316 5095 30356 5104
rect 30028 4892 30068 4901
rect 30028 4388 30068 4852
rect 30028 4339 30068 4348
rect 30220 4724 30260 4733
rect 29932 4171 29972 4180
rect 30220 3800 30260 4684
rect 30508 4472 30548 4481
rect 30508 4136 30548 4432
rect 30508 4087 30548 4096
rect 30220 3751 30260 3760
rect 29836 3667 29876 3676
rect 30508 3716 30548 3725
rect 30316 3632 30356 3641
rect 30124 3548 30164 3557
rect 30028 2960 30068 2969
rect 29836 2876 29876 2885
rect 29836 2204 29876 2836
rect 30028 2288 30068 2920
rect 30028 2239 30068 2248
rect 29836 2155 29876 2164
rect 29740 1903 29780 1912
rect 29932 2120 29972 2129
rect 29932 1868 29972 2080
rect 29932 1819 29972 1828
rect 29548 1616 29588 1625
rect 29548 1481 29588 1576
rect 29836 1280 29876 1289
rect 29644 440 29684 449
rect 29644 80 29684 400
rect 29836 80 29876 1240
rect 30124 692 30164 3508
rect 30316 3464 30356 3592
rect 30508 3581 30548 3676
rect 30316 3415 30356 3424
rect 30412 3548 30452 3557
rect 30220 2540 30260 2549
rect 30220 2405 30260 2500
rect 30220 2288 30260 2297
rect 30220 2153 30260 2248
rect 30412 1868 30452 3508
rect 30508 3212 30548 3221
rect 30508 2792 30548 3172
rect 30508 2743 30548 2752
rect 30508 2624 30548 2633
rect 30508 2489 30548 2584
rect 30412 1819 30452 1828
rect 30604 1616 30644 6952
rect 30700 6656 30740 10228
rect 31468 10184 31508 10193
rect 31660 10184 31700 10193
rect 31508 10144 31660 10184
rect 31468 10135 31508 10144
rect 31660 10135 31700 10144
rect 31756 10016 31796 10025
rect 31660 9512 31700 9521
rect 31468 9428 31508 9437
rect 31084 8756 31124 8765
rect 30892 8672 30932 8681
rect 30892 7916 30932 8632
rect 30892 7867 30932 7876
rect 31084 7916 31124 8716
rect 31084 7867 31124 7876
rect 31468 8084 31508 9388
rect 30700 6404 30740 6616
rect 30700 6355 30740 6364
rect 30796 7076 30836 7085
rect 30700 6236 30740 6245
rect 30700 5816 30740 6196
rect 30700 5767 30740 5776
rect 30700 3884 30740 3893
rect 30700 3380 30740 3844
rect 30700 3044 30740 3340
rect 30700 2995 30740 3004
rect 30700 2708 30740 2717
rect 30700 2573 30740 2668
rect 30028 652 30164 692
rect 30220 1576 30644 1616
rect 30028 80 30068 652
rect 30220 80 30260 1576
rect 30604 1448 30644 1457
rect 30412 944 30452 953
rect 30412 80 30452 904
rect 30604 80 30644 1408
rect 30796 80 30836 7036
rect 31372 6656 31412 6665
rect 31372 6152 31412 6616
rect 31372 6103 31412 6112
rect 30892 5816 30932 5827
rect 30892 5732 30932 5776
rect 30892 5683 30932 5692
rect 31276 5648 31316 5657
rect 30988 5564 31028 5573
rect 30988 3884 31028 5524
rect 31276 4892 31316 5608
rect 31180 4472 31220 4481
rect 30988 3844 31124 3884
rect 30988 3212 31028 3221
rect 30892 3044 30932 3053
rect 30892 1448 30932 3004
rect 30892 1399 30932 1408
rect 30988 80 31028 3172
rect 31084 2792 31124 3844
rect 31084 2743 31124 2752
rect 31180 80 31220 4432
rect 31276 4304 31316 4852
rect 31276 4255 31316 4264
rect 31372 5144 31412 5153
rect 31276 4136 31316 4145
rect 31276 3128 31316 4096
rect 31276 3079 31316 3088
rect 31276 2876 31316 2885
rect 31276 2666 31316 2836
rect 31276 2617 31316 2626
rect 31276 2288 31316 2297
rect 31276 1784 31316 2248
rect 31276 1735 31316 1744
rect 31372 80 31412 5104
rect 31468 1700 31508 8044
rect 31564 8756 31604 8765
rect 31564 5144 31604 8716
rect 31660 8336 31700 9472
rect 31756 9344 31796 9976
rect 32332 9680 32372 12100
rect 32524 11696 32564 11705
rect 32524 10184 32564 11656
rect 32524 10135 32564 10144
rect 32620 11360 32660 11369
rect 32332 9631 32372 9640
rect 32332 9512 32372 9521
rect 32332 9428 32372 9472
rect 32332 9377 32372 9388
rect 32524 9428 32564 9437
rect 31756 9295 31796 9304
rect 32524 9008 32564 9388
rect 32524 8959 32564 8968
rect 32524 8840 32564 8849
rect 31660 8168 31700 8296
rect 31660 8119 31700 8128
rect 31852 8756 31892 8765
rect 31564 5095 31604 5104
rect 31660 7916 31700 7925
rect 31660 5816 31700 7876
rect 31756 7832 31796 7841
rect 31756 6656 31796 7792
rect 31852 6740 31892 8716
rect 32140 8672 32180 8681
rect 31948 7916 31988 7925
rect 31948 7412 31988 7876
rect 31948 7363 31988 7372
rect 32044 7748 32084 7757
rect 31948 6740 31988 6749
rect 31852 6700 31948 6740
rect 31756 6616 31892 6656
rect 31564 4892 31604 4901
rect 31564 3968 31604 4852
rect 31564 2120 31604 3928
rect 31660 3128 31700 5776
rect 31756 5900 31796 5909
rect 31756 5732 31796 5860
rect 31756 5683 31796 5692
rect 31660 3079 31700 3088
rect 31756 4892 31796 4901
rect 31660 2960 31700 2969
rect 31660 2792 31700 2920
rect 31660 2743 31700 2752
rect 31660 2372 31700 2381
rect 31660 2237 31700 2332
rect 31564 1868 31604 2080
rect 31564 1819 31604 1828
rect 31468 1651 31508 1660
rect 31660 1700 31700 1709
rect 31564 1364 31604 1373
rect 31564 80 31604 1324
rect 31660 692 31700 1660
rect 31756 1280 31796 4852
rect 31852 4892 31892 6616
rect 31948 6404 31988 6700
rect 31948 6355 31988 6364
rect 31852 4843 31892 4852
rect 31948 5900 31988 5909
rect 31852 4388 31892 4397
rect 31852 4136 31892 4348
rect 31852 4087 31892 4096
rect 31756 1231 31796 1240
rect 31852 3800 31892 3809
rect 31852 692 31892 3760
rect 31660 643 31700 652
rect 31756 652 31892 692
rect 31756 80 31796 652
rect 31948 80 31988 5860
rect 32044 4976 32084 7708
rect 32140 6404 32180 8632
rect 32428 7832 32468 7841
rect 32332 7412 32372 7421
rect 32236 7244 32276 7255
rect 32236 7160 32276 7204
rect 32236 7111 32276 7120
rect 32236 6908 32276 6917
rect 32236 6656 32276 6868
rect 32236 6607 32276 6616
rect 32140 6364 32276 6404
rect 32140 6236 32180 6245
rect 32140 5816 32180 6196
rect 32140 5767 32180 5776
rect 32236 5648 32276 6364
rect 32044 4927 32084 4936
rect 32140 5608 32276 5648
rect 32044 4220 32084 4229
rect 32044 4085 32084 4180
rect 32044 2708 32084 2717
rect 32044 2120 32084 2668
rect 32044 2071 32084 2080
rect 32044 1868 32084 1877
rect 32044 1733 32084 1828
rect 32140 80 32180 5608
rect 32236 5144 32276 5153
rect 32236 440 32276 5104
rect 32332 4808 32372 7372
rect 32428 7328 32468 7792
rect 32428 7279 32468 7288
rect 32428 7076 32468 7085
rect 32428 6656 32468 7036
rect 32428 6607 32468 6616
rect 32428 4976 32468 4985
rect 32428 4841 32468 4936
rect 32332 4759 32372 4768
rect 32428 4640 32468 4649
rect 32428 4388 32468 4600
rect 32428 4339 32468 4348
rect 32428 4220 32468 4229
rect 32332 3884 32372 3979
rect 32332 3835 32372 3844
rect 32332 3716 32372 3725
rect 32332 3548 32372 3676
rect 32332 3380 32372 3508
rect 32332 3331 32372 3340
rect 32428 2792 32468 4180
rect 32332 2456 32372 2465
rect 32332 2372 32372 2416
rect 32332 2321 32372 2332
rect 32428 1868 32468 2752
rect 32428 1819 32468 1828
rect 32428 1700 32468 1709
rect 32236 391 32276 400
rect 32332 1448 32372 1457
rect 32332 80 32372 1408
rect 32428 860 32468 1660
rect 32428 811 32468 820
rect 32524 80 32564 8800
rect 32620 2900 32660 11320
rect 32908 10940 32948 10949
rect 32908 10184 32948 10900
rect 32908 10135 32948 10144
rect 33196 10268 33236 10277
rect 33004 9932 33044 9941
rect 32716 9092 32756 9101
rect 32716 8924 32756 9052
rect 32908 9008 32948 9017
rect 32716 8875 32756 8884
rect 32812 8924 32852 8933
rect 32812 8000 32852 8884
rect 32812 7951 32852 7960
rect 32908 7664 32948 8968
rect 33004 8672 33044 9892
rect 33004 8623 33044 8632
rect 33100 9932 33140 9941
rect 33100 8420 33140 9892
rect 33196 9764 33236 10228
rect 33196 9715 33236 9724
rect 33484 9680 33524 12100
rect 34348 10520 34388 10529
rect 33484 9631 33524 9640
rect 33580 10352 33620 10361
rect 33388 9260 33428 9269
rect 33292 9092 33332 9101
rect 33196 9008 33236 9017
rect 33196 8840 33236 8968
rect 33292 9008 33332 9052
rect 33292 8957 33332 8968
rect 33196 8791 33236 8800
rect 33196 8672 33236 8683
rect 33196 8588 33236 8632
rect 33196 8539 33236 8548
rect 33100 8380 33332 8420
rect 32716 7624 32948 7664
rect 32716 5816 32756 7624
rect 33100 7540 33236 7580
rect 32908 7496 32948 7505
rect 32908 7328 32948 7456
rect 33100 7496 33140 7540
rect 33100 7447 33140 7456
rect 32908 7279 32948 7288
rect 32812 7076 32852 7085
rect 32812 5984 32852 7036
rect 33196 6488 33236 7540
rect 33196 6439 33236 6448
rect 33196 6320 33236 6329
rect 33004 6236 33044 6245
rect 32812 5935 32852 5944
rect 32908 6152 32948 6161
rect 32716 5776 32852 5816
rect 32716 5564 32756 5573
rect 32716 5144 32756 5524
rect 32716 5095 32756 5104
rect 32716 4892 32756 4901
rect 32716 4304 32756 4852
rect 32716 4255 32756 4264
rect 32716 3884 32756 3893
rect 32716 3212 32756 3844
rect 32716 3163 32756 3172
rect 32620 2860 32756 2900
rect 32620 2792 32660 2801
rect 32620 2657 32660 2752
rect 32716 80 32756 2860
rect 32812 1448 32852 5776
rect 32908 4052 32948 6112
rect 33004 5900 33044 6196
rect 33004 5851 33044 5860
rect 33100 5648 33140 5657
rect 33004 5480 33044 5489
rect 33004 4976 33044 5440
rect 33004 4927 33044 4936
rect 33100 4640 33140 5608
rect 33196 5564 33236 6280
rect 33196 5515 33236 5524
rect 33100 4591 33140 4600
rect 33196 5396 33236 5405
rect 32908 4003 32948 4012
rect 33004 4136 33044 4145
rect 32908 3716 32948 3725
rect 32908 3044 32948 3676
rect 32908 2708 32948 3004
rect 33004 2960 33044 4096
rect 33196 3128 33236 5356
rect 33004 2911 33044 2920
rect 33100 3088 33236 3128
rect 33100 2792 33140 3088
rect 32908 2659 32948 2668
rect 33004 2752 33140 2792
rect 32908 2288 32948 2297
rect 32908 1616 32948 2248
rect 33004 1952 33044 2752
rect 33292 2708 33332 8380
rect 33388 5396 33428 9220
rect 33580 7496 33620 10312
rect 34252 10352 34292 10361
rect 34252 10016 34292 10312
rect 34252 9967 34292 9976
rect 33928 9848 34296 9857
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 33928 9799 34296 9808
rect 34156 9596 34196 9607
rect 34156 9512 34196 9556
rect 34156 9463 34196 9472
rect 33580 7447 33620 7456
rect 33676 8924 33716 8933
rect 33580 7328 33620 7337
rect 33484 6404 33524 6413
rect 33484 6269 33524 6364
rect 33388 5347 33428 5356
rect 33580 5312 33620 7288
rect 33676 5816 33716 8884
rect 33928 8336 34296 8345
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 33928 8287 34296 8296
rect 34156 8168 34196 8177
rect 33964 8000 34004 8009
rect 33772 7748 33812 7757
rect 33772 7580 33812 7708
rect 33964 7664 34004 7960
rect 33964 7615 34004 7624
rect 34156 7664 34196 8128
rect 34156 7615 34196 7624
rect 34252 7916 34292 7925
rect 33772 7412 33812 7540
rect 34252 7496 34292 7876
rect 34252 7447 34292 7456
rect 33772 7363 33812 7372
rect 33868 7412 33908 7421
rect 33868 7244 33908 7372
rect 33868 7195 33908 7204
rect 33772 7076 33812 7085
rect 33772 5984 33812 7036
rect 33928 6824 34296 6833
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 33928 6775 34296 6784
rect 34348 6656 34388 10480
rect 34636 10436 34676 12100
rect 35596 11612 35636 11621
rect 34924 11192 34964 11201
rect 34636 10387 34676 10396
rect 34732 10604 34772 10613
rect 34540 10016 34580 10025
rect 34444 9764 34484 9773
rect 34444 9344 34484 9724
rect 34540 9512 34580 9976
rect 34636 9932 34676 9943
rect 34636 9848 34676 9892
rect 34636 9799 34676 9808
rect 34540 9463 34580 9472
rect 34444 9092 34484 9304
rect 34444 9052 34580 9092
rect 34540 8756 34580 9052
rect 34540 8707 34580 8716
rect 34444 8672 34484 8681
rect 34444 8168 34484 8632
rect 34444 8119 34484 8128
rect 34540 8588 34580 8597
rect 34540 7328 34580 8548
rect 34348 6607 34388 6616
rect 34444 7288 34580 7328
rect 33772 5935 33812 5944
rect 33676 5776 34100 5816
rect 34060 5732 34100 5776
rect 33868 5648 33908 5657
rect 33772 5608 33868 5648
rect 33676 5564 33716 5573
rect 33676 5429 33716 5524
rect 33580 5272 33716 5312
rect 33580 5144 33620 5153
rect 33388 5060 33428 5069
rect 33388 4052 33428 5020
rect 33580 4388 33620 5104
rect 33580 4339 33620 4348
rect 33388 4003 33428 4012
rect 33580 4136 33620 4145
rect 33580 3632 33620 4096
rect 33580 3583 33620 3592
rect 33484 3044 33524 3053
rect 33484 2876 33524 3004
rect 33484 2827 33524 2836
rect 33292 2668 33524 2708
rect 33004 1903 33044 1912
rect 33388 2372 33428 2381
rect 32908 1567 32948 1576
rect 33196 1700 33236 1709
rect 32812 1399 32852 1408
rect 33196 860 33236 1660
rect 33196 811 33236 820
rect 33292 1616 33332 1625
rect 33100 440 33140 449
rect 32908 188 32948 197
rect 32908 80 32948 148
rect 33100 80 33140 400
rect 33292 80 33332 1576
rect 33388 776 33428 2332
rect 33484 1952 33524 2668
rect 33484 1903 33524 1912
rect 33484 1700 33524 1709
rect 33484 944 33524 1660
rect 33676 1448 33716 5272
rect 33772 4220 33812 5608
rect 33868 5599 33908 5608
rect 34060 5480 34100 5692
rect 34060 5431 34100 5440
rect 34348 5732 34388 5741
rect 33928 5312 34296 5321
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 33928 5263 34296 5272
rect 34252 5144 34292 5153
rect 34252 4892 34292 5104
rect 34252 4843 34292 4852
rect 34348 4640 34388 5692
rect 34348 4591 34388 4600
rect 33964 4556 34004 4565
rect 33868 4220 33908 4229
rect 33812 4180 33868 4220
rect 33772 4171 33812 4180
rect 33868 4171 33908 4180
rect 33964 4052 34004 4516
rect 34252 4388 34292 4397
rect 34252 4220 34292 4348
rect 34252 4171 34292 4180
rect 34444 4220 34484 7288
rect 34540 7160 34580 7169
rect 34540 6488 34580 7120
rect 34540 6439 34580 6448
rect 34732 5984 34772 10564
rect 34828 10268 34868 10277
rect 34828 10133 34868 10228
rect 34828 9932 34868 9941
rect 34828 9764 34868 9892
rect 34828 9715 34868 9724
rect 34924 9596 34964 11152
rect 35020 11024 35060 11033
rect 35020 10268 35060 10984
rect 35168 10604 35536 10613
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35168 10555 35536 10564
rect 35020 10219 35060 10228
rect 34924 9556 35060 9596
rect 34828 9512 34868 9521
rect 34828 9008 34868 9472
rect 34828 8756 34868 8968
rect 34828 8707 34868 8716
rect 34924 9428 34964 9437
rect 34924 8924 34964 9388
rect 34924 8672 34964 8884
rect 34924 8623 34964 8632
rect 34924 7916 34964 7925
rect 34732 5935 34772 5944
rect 34828 7496 34868 7505
rect 34828 6404 34868 7456
rect 34924 7244 34964 7876
rect 34924 7195 34964 7204
rect 34444 4171 34484 4180
rect 34540 5900 34580 5909
rect 33772 4012 34004 4052
rect 34348 4136 34388 4145
rect 33772 1952 33812 4012
rect 33928 3800 34296 3809
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 33928 3751 34296 3760
rect 34348 3548 34388 4096
rect 34540 4052 34580 5860
rect 34636 5816 34676 5827
rect 34636 5732 34676 5776
rect 34636 5683 34676 5692
rect 34828 4976 34868 6364
rect 34828 4927 34868 4936
rect 34924 6908 34964 6917
rect 34732 4388 34772 4397
rect 34540 4003 34580 4012
rect 34636 4220 34676 4229
rect 34156 3508 34388 3548
rect 34444 3968 34484 3977
rect 33964 2876 34004 2885
rect 33964 2741 34004 2836
rect 33868 2708 33908 2717
rect 33868 2573 33908 2668
rect 34156 2708 34196 3508
rect 34348 3212 34388 3221
rect 34444 3212 34484 3928
rect 34540 3716 34580 3725
rect 34540 3464 34580 3676
rect 34540 3415 34580 3424
rect 34636 3296 34676 4180
rect 34388 3172 34484 3212
rect 34540 3256 34676 3296
rect 34348 3163 34388 3172
rect 34444 3044 34484 3053
rect 34156 2659 34196 2668
rect 34348 2876 34388 2885
rect 33964 2624 34004 2635
rect 33964 2540 34004 2584
rect 34348 2624 34388 2836
rect 34348 2575 34388 2584
rect 33964 2491 34004 2500
rect 33928 2288 34296 2297
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 33928 2239 34296 2248
rect 33964 2036 34004 2045
rect 34004 1996 34196 2036
rect 33964 1987 34004 1996
rect 33772 1903 33812 1912
rect 34156 1448 34196 1996
rect 33676 1408 34100 1448
rect 33484 895 33524 904
rect 33388 736 33716 776
rect 33484 104 33524 113
rect 11636 64 11656 80
rect 11576 0 11656 64
rect 11768 0 11848 80
rect 11960 0 12040 80
rect 12152 0 12232 80
rect 12344 0 12424 80
rect 12536 0 12616 80
rect 12728 0 12808 80
rect 12920 0 13000 80
rect 13112 0 13192 80
rect 13304 0 13384 80
rect 13496 0 13576 80
rect 13688 0 13768 80
rect 13880 0 13960 80
rect 14072 0 14152 80
rect 14264 0 14344 80
rect 14456 0 14536 80
rect 14648 0 14728 80
rect 14840 0 14920 80
rect 15032 0 15112 80
rect 15224 0 15304 80
rect 15416 0 15496 80
rect 15608 0 15688 80
rect 15800 0 15880 80
rect 15992 0 16072 80
rect 16184 0 16264 80
rect 16376 0 16456 80
rect 16568 0 16648 80
rect 16760 0 16840 80
rect 16952 0 17032 80
rect 17144 0 17224 80
rect 17336 0 17416 80
rect 17528 0 17608 80
rect 17720 0 17800 80
rect 17912 0 17992 80
rect 18104 0 18184 80
rect 18296 0 18376 80
rect 18488 0 18568 80
rect 18680 0 18760 80
rect 18872 0 18952 80
rect 19064 0 19144 80
rect 19256 0 19336 80
rect 19448 0 19528 80
rect 19640 0 19720 80
rect 19832 0 19912 80
rect 20024 0 20104 80
rect 20216 0 20296 80
rect 20408 0 20488 80
rect 20600 0 20680 80
rect 20792 0 20872 80
rect 20984 0 21064 80
rect 21176 0 21256 80
rect 21368 0 21448 80
rect 21560 0 21640 80
rect 21752 0 21832 80
rect 21944 0 22024 80
rect 22136 0 22216 80
rect 22328 0 22408 80
rect 22520 0 22600 80
rect 22712 0 22792 80
rect 22904 0 22984 80
rect 23096 0 23176 80
rect 23288 0 23368 80
rect 23480 0 23560 80
rect 23672 0 23752 80
rect 23864 0 23944 80
rect 24056 0 24136 80
rect 24248 0 24328 80
rect 24440 0 24520 80
rect 24632 0 24712 80
rect 24824 0 24904 80
rect 25016 0 25096 80
rect 25208 0 25288 80
rect 25400 0 25480 80
rect 25592 0 25672 80
rect 25784 0 25864 80
rect 25976 0 26056 80
rect 26168 0 26248 80
rect 26360 0 26440 80
rect 26552 0 26632 80
rect 26744 0 26824 80
rect 26936 0 27016 80
rect 27128 0 27208 80
rect 27320 0 27400 80
rect 27512 0 27592 80
rect 27704 0 27784 80
rect 27896 0 27976 80
rect 28088 0 28168 80
rect 28280 0 28360 80
rect 28472 0 28552 80
rect 28664 0 28744 80
rect 28856 0 28936 80
rect 29048 0 29128 80
rect 29240 0 29320 80
rect 29432 0 29512 80
rect 29624 0 29704 80
rect 29816 0 29896 80
rect 30008 0 30088 80
rect 30200 0 30280 80
rect 30392 0 30472 80
rect 30584 0 30664 80
rect 30776 0 30856 80
rect 30968 0 31048 80
rect 31160 0 31240 80
rect 31352 0 31432 80
rect 31544 0 31624 80
rect 31736 0 31816 80
rect 31928 0 32008 80
rect 32120 0 32200 80
rect 32312 0 32392 80
rect 32504 0 32584 80
rect 32696 0 32776 80
rect 32888 0 32968 80
rect 33080 0 33160 80
rect 33272 0 33352 80
rect 33464 64 33484 80
rect 33676 80 33716 736
rect 33868 692 33908 701
rect 33868 80 33908 652
rect 34060 80 34100 1408
rect 34156 1399 34196 1408
rect 34252 1364 34292 1373
rect 34252 80 34292 1324
rect 34444 80 34484 3004
rect 34540 2624 34580 3256
rect 34540 2575 34580 2584
rect 34636 3044 34676 3053
rect 34540 2456 34580 2465
rect 34540 1952 34580 2416
rect 34540 1903 34580 1912
rect 34636 80 34676 3004
rect 34732 2708 34772 4348
rect 34924 3128 34964 6868
rect 34732 2036 34772 2668
rect 34732 1987 34772 1996
rect 34828 3088 34964 3128
rect 34828 80 34868 3088
rect 34924 2960 34964 2971
rect 34924 2876 34964 2920
rect 34924 2827 34964 2836
rect 34924 1952 34964 1961
rect 34924 1532 34964 1912
rect 34924 1483 34964 1492
rect 35020 80 35060 9556
rect 35168 9092 35536 9101
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35168 9043 35536 9052
rect 35168 7580 35536 7589
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35168 7531 35536 7540
rect 35404 6404 35444 6413
rect 35404 6236 35444 6364
rect 35596 6404 35636 11572
rect 35692 11444 35732 11453
rect 35692 6908 35732 11404
rect 35788 10436 35828 12100
rect 35788 10387 35828 10396
rect 36940 10436 36980 12100
rect 37516 11528 37556 11537
rect 37516 10688 37556 11488
rect 37516 10639 37556 10648
rect 37804 11108 37844 11117
rect 36940 10387 36980 10396
rect 35692 6859 35732 6868
rect 35788 10268 35828 10277
rect 35788 7916 35828 10228
rect 37804 10184 37844 11068
rect 38092 10436 38132 12100
rect 38956 11276 38996 11285
rect 38764 11024 38804 11033
rect 38092 10387 38132 10396
rect 38380 10772 38420 10781
rect 37804 10135 37844 10144
rect 38380 10184 38420 10732
rect 38380 10135 38420 10144
rect 38764 10268 38804 10984
rect 38956 10352 38996 11236
rect 38956 10303 38996 10312
rect 39052 10604 39092 10613
rect 36268 10100 36308 10109
rect 35884 9428 35924 9437
rect 35884 9293 35924 9388
rect 36268 9260 36308 10060
rect 38284 10100 38324 10109
rect 36652 10016 36692 10025
rect 36652 9428 36692 9976
rect 37420 9596 37460 9605
rect 36652 9379 36692 9388
rect 36748 9512 36788 9521
rect 36268 9211 36308 9220
rect 35980 8840 36020 8849
rect 35596 6355 35636 6364
rect 35404 6187 35444 6196
rect 35596 6236 35636 6245
rect 35168 6068 35536 6077
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35168 6019 35536 6028
rect 35596 5732 35636 6196
rect 35596 5683 35636 5692
rect 35692 5900 35732 5909
rect 35692 4976 35732 5860
rect 35692 4927 35732 4936
rect 35596 4892 35636 4901
rect 35168 4556 35536 4565
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35168 4507 35536 4516
rect 35116 3884 35156 3893
rect 35116 3716 35156 3844
rect 35116 3667 35156 3676
rect 35116 3548 35156 3557
rect 35116 3212 35156 3508
rect 35596 3464 35636 4852
rect 35788 4892 35828 7876
rect 35788 4843 35828 4852
rect 35884 8420 35924 8429
rect 35692 4808 35732 4817
rect 35692 4220 35732 4768
rect 35884 4556 35924 8380
rect 35980 5564 36020 8800
rect 36268 8756 36308 8765
rect 36268 8168 36308 8716
rect 36748 8756 36788 9472
rect 37132 9428 37172 9437
rect 36940 9344 36980 9353
rect 36748 8621 36788 8716
rect 36844 9260 36884 9269
rect 36844 8252 36884 9220
rect 36940 9209 36980 9304
rect 36844 8203 36884 8212
rect 37036 8756 37076 8765
rect 36268 8119 36308 8128
rect 36652 8168 36692 8177
rect 36652 8000 36692 8128
rect 36652 7951 36692 7960
rect 36844 8000 36884 8009
rect 36268 7328 36308 7337
rect 36076 6236 36116 6245
rect 36076 5732 36116 6196
rect 36076 5683 36116 5692
rect 36172 5816 36212 5825
rect 35980 5515 36020 5524
rect 36172 5396 36212 5776
rect 36076 5356 36212 5396
rect 35980 4892 36020 4901
rect 35980 4757 36020 4852
rect 36076 4556 36116 5356
rect 35884 4507 35924 4516
rect 35980 4516 36116 4556
rect 35692 4171 35732 4180
rect 35788 3968 35828 3977
rect 35788 3833 35828 3928
rect 35596 3415 35636 3424
rect 35116 3163 35156 3172
rect 35692 3380 35732 3389
rect 35168 3044 35536 3053
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35168 2995 35536 3004
rect 35596 3044 35636 3053
rect 35116 2708 35156 2717
rect 35116 2540 35156 2668
rect 35596 2708 35636 3004
rect 35692 2960 35732 3340
rect 35884 3212 35924 3221
rect 35884 3044 35924 3172
rect 35884 2995 35924 3004
rect 35692 2911 35732 2920
rect 35980 2900 36020 4516
rect 36076 4388 36116 4397
rect 36076 3464 36116 4348
rect 36076 3415 36116 3424
rect 36268 3464 36308 7288
rect 36748 6992 36788 7001
rect 36748 6824 36788 6952
rect 36748 6775 36788 6784
rect 36844 6404 36884 7960
rect 36844 6355 36884 6364
rect 36940 7244 36980 7253
rect 36652 5900 36692 5911
rect 36460 5816 36500 5825
rect 36364 5732 36404 5741
rect 36364 5564 36404 5692
rect 36364 5515 36404 5524
rect 36460 5144 36500 5776
rect 36652 5816 36692 5860
rect 36652 5767 36692 5776
rect 36940 5732 36980 7204
rect 36940 5228 36980 5692
rect 36940 5179 36980 5188
rect 36460 5095 36500 5104
rect 36940 4976 36980 4985
rect 37036 4976 37076 8716
rect 37132 8168 37172 9388
rect 37420 9176 37460 9556
rect 37420 9127 37460 9136
rect 37132 8119 37172 8128
rect 37324 9092 37364 9101
rect 37132 8000 37172 8009
rect 37132 7412 37172 7960
rect 37132 7160 37172 7372
rect 37132 7111 37172 7120
rect 37132 6992 37172 7001
rect 37132 6656 37172 6952
rect 37132 6607 37172 6616
rect 37228 6908 37268 6917
rect 37228 6656 37268 6868
rect 37228 6607 37268 6616
rect 36980 4936 37076 4976
rect 36460 4892 36500 4901
rect 36460 4220 36500 4852
rect 36460 4171 36500 4180
rect 36556 4052 36596 4061
rect 36556 3632 36596 4012
rect 36556 3583 36596 3592
rect 36268 3415 36308 3424
rect 35596 2659 35636 2668
rect 35884 2860 36020 2900
rect 36268 3296 36308 3305
rect 35116 2288 35156 2500
rect 35116 2239 35156 2248
rect 35884 1952 35924 2860
rect 36076 2708 36116 2717
rect 36076 2456 36116 2668
rect 36268 2708 36308 3256
rect 36460 3296 36500 3307
rect 36460 3212 36500 3256
rect 36940 3296 36980 4936
rect 36940 3247 36980 3256
rect 36460 3163 36500 3172
rect 36268 2659 36308 2668
rect 36076 2407 36116 2416
rect 36748 2624 36788 2633
rect 35884 1903 35924 1912
rect 36172 1700 36212 1709
rect 35168 1532 35536 1541
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35168 1483 35536 1492
rect 36172 944 36212 1660
rect 36748 1364 36788 2584
rect 37324 1616 37364 9052
rect 38188 8504 38228 8513
rect 37804 8252 37844 8261
rect 37516 7244 37556 7253
rect 37420 6572 37460 6581
rect 37420 3632 37460 6532
rect 37516 6320 37556 7204
rect 37708 7244 37748 7253
rect 37516 6271 37556 6280
rect 37612 6320 37652 6329
rect 37516 5480 37556 5489
rect 37516 4892 37556 5440
rect 37516 4843 37556 4852
rect 37420 3583 37460 3592
rect 37612 4220 37652 6280
rect 37708 4304 37748 7204
rect 37708 4255 37748 4264
rect 37612 3632 37652 4180
rect 37612 3583 37652 3592
rect 37420 2960 37460 2969
rect 37420 2900 37460 2920
rect 37420 2876 37556 2900
rect 37420 2860 37516 2876
rect 37516 2796 37556 2836
rect 37804 2792 37844 8212
rect 38092 8252 38132 8261
rect 38092 7916 38132 8212
rect 38188 8000 38228 8464
rect 38188 7951 38228 7960
rect 38092 7867 38132 7876
rect 38092 6992 38132 7001
rect 38092 6740 38132 6952
rect 38092 6691 38132 6700
rect 38188 5732 38228 5741
rect 37900 5060 37940 5071
rect 37900 4976 37940 5020
rect 37900 4927 37940 4936
rect 37996 4892 38036 4901
rect 37900 4808 37940 4817
rect 37900 4388 37940 4768
rect 37900 4339 37940 4348
rect 37804 2743 37844 2752
rect 37900 4136 37940 4145
rect 37900 3380 37940 4096
rect 37900 2708 37940 3340
rect 37420 2456 37460 2465
rect 37420 1868 37460 2416
rect 37900 2036 37940 2668
rect 37996 2204 38036 4852
rect 38092 4640 38132 4649
rect 38092 4388 38132 4600
rect 38092 4339 38132 4348
rect 38188 2456 38228 5692
rect 38188 2407 38228 2416
rect 37996 2155 38036 2164
rect 37900 1987 37940 1996
rect 38284 1952 38324 10060
rect 38380 9512 38420 9521
rect 38380 9428 38420 9472
rect 38380 9377 38420 9388
rect 38764 9428 38804 10228
rect 39052 9764 39092 10564
rect 39244 10436 39284 12100
rect 40300 10940 40340 10949
rect 40300 10805 40340 10900
rect 39244 10387 39284 10396
rect 40396 10352 40436 12100
rect 40588 10856 40628 10865
rect 40588 10436 40628 10816
rect 40588 10387 40628 10396
rect 41548 10436 41588 12100
rect 42508 11696 42548 11705
rect 42316 11612 42356 11621
rect 41548 10387 41588 10396
rect 42124 11108 42164 11117
rect 40396 10303 40436 10312
rect 39244 10268 39284 10277
rect 39052 9715 39092 9724
rect 39148 10184 39188 10193
rect 38956 9680 38996 9691
rect 38956 9596 38996 9640
rect 38956 9547 38996 9556
rect 38764 9379 38804 9388
rect 39148 9512 39188 10144
rect 39244 10133 39284 10228
rect 42028 10268 42068 10277
rect 41740 10100 41780 10109
rect 39340 10016 39380 10025
rect 38476 8924 38516 8933
rect 38380 8756 38420 8765
rect 38380 7244 38420 8716
rect 38476 8672 38516 8884
rect 38572 8672 38612 8700
rect 38476 8632 38572 8672
rect 38476 7916 38516 8632
rect 38572 8623 38612 8632
rect 38476 7867 38516 7876
rect 39052 7664 39092 7673
rect 39052 7328 39092 7624
rect 39052 7279 39092 7288
rect 38380 6488 38420 7204
rect 39148 7160 39188 9472
rect 39244 9596 39284 9605
rect 39244 9461 39284 9556
rect 39340 9512 39380 9976
rect 39340 9463 39380 9472
rect 40108 9932 40148 9941
rect 39724 8924 39764 8933
rect 39148 7111 39188 7120
rect 39628 7832 39668 7841
rect 38380 6439 38420 6448
rect 39244 6992 39284 7001
rect 38956 6404 38996 6413
rect 38764 5984 38804 5993
rect 38380 5480 38420 5489
rect 38380 5144 38420 5440
rect 38380 5095 38420 5104
rect 38572 5480 38612 5489
rect 38572 4808 38612 5440
rect 38572 4759 38612 4768
rect 38668 4136 38708 4145
rect 38668 2960 38708 4096
rect 38668 2911 38708 2920
rect 38668 2708 38708 2717
rect 38668 2372 38708 2668
rect 38668 2323 38708 2332
rect 38764 2120 38804 5944
rect 38956 5648 38996 6364
rect 38956 5144 38996 5608
rect 38956 5095 38996 5104
rect 39148 5480 39188 5489
rect 39148 5144 39188 5440
rect 39148 5095 39188 5104
rect 38860 4136 38900 4145
rect 38860 4001 38900 4096
rect 38764 2071 38804 2080
rect 38956 3380 38996 3389
rect 38956 2708 38996 3340
rect 39244 3380 39284 6952
rect 39244 3331 39284 3340
rect 39532 4472 39572 4481
rect 39532 2876 39572 4432
rect 39628 4136 39668 7792
rect 39628 3548 39668 4096
rect 39628 3499 39668 3508
rect 39532 2827 39572 2836
rect 38284 1903 38324 1912
rect 37420 1819 37460 1828
rect 38956 1868 38996 2668
rect 38956 1819 38996 1828
rect 39724 1700 39764 8884
rect 39820 8504 39860 8513
rect 39820 7916 39860 8464
rect 39820 7867 39860 7876
rect 39724 1651 39764 1660
rect 39820 7076 39860 7085
rect 37324 1567 37364 1576
rect 39820 1532 39860 7036
rect 40012 6572 40052 6581
rect 39916 4808 39956 4817
rect 39916 3296 39956 4768
rect 40012 4304 40052 6532
rect 40012 4255 40052 4264
rect 39916 2288 39956 3256
rect 39916 2239 39956 2248
rect 39820 1483 39860 1492
rect 36748 1315 36788 1324
rect 36172 895 36212 904
rect 40108 692 40148 9892
rect 40396 9932 40436 9941
rect 40300 9680 40340 9689
rect 40300 9545 40340 9640
rect 40204 9428 40244 9439
rect 40204 9344 40244 9388
rect 40396 9428 40436 9892
rect 40396 9379 40436 9388
rect 41548 9596 41588 9605
rect 40204 9295 40244 9304
rect 41356 9344 41396 9353
rect 40396 9260 40436 9269
rect 40396 8672 40436 9220
rect 40396 8623 40436 8632
rect 40492 8756 40532 8765
rect 40204 7832 40244 7841
rect 40204 6404 40244 7792
rect 40492 7244 40532 8716
rect 40780 8756 40820 8765
rect 40780 8084 40820 8716
rect 40780 8035 40820 8044
rect 41356 8756 41396 9304
rect 41452 9344 41492 9353
rect 41452 9176 41492 9304
rect 41452 9127 41492 9136
rect 40396 7160 40436 7169
rect 40300 6824 40340 6833
rect 40300 6689 40340 6784
rect 40396 6656 40436 7120
rect 40396 6607 40436 6616
rect 40204 6355 40244 6364
rect 40300 6152 40340 6161
rect 40300 6017 40340 6112
rect 40300 5732 40340 5741
rect 40300 4892 40340 5692
rect 40300 4472 40340 4852
rect 40300 4423 40340 4432
rect 40492 3884 40532 7204
rect 41356 7244 41396 8716
rect 40588 7160 40628 7169
rect 40588 6908 40628 7120
rect 40588 6859 40628 6868
rect 40684 6572 40724 6581
rect 40684 5648 40724 6532
rect 40684 5599 40724 5608
rect 41068 6236 41108 6245
rect 40972 4976 41012 4985
rect 40972 4052 41012 4936
rect 40972 4003 41012 4012
rect 40492 3835 40532 3844
rect 40972 3884 41012 3893
rect 40492 3716 40532 3725
rect 40300 3464 40340 3473
rect 40300 3329 40340 3424
rect 40492 3380 40532 3676
rect 40492 2900 40532 3340
rect 40780 3380 40820 3389
rect 40492 2860 40724 2900
rect 40684 2624 40724 2860
rect 40780 2792 40820 3340
rect 40972 3380 41012 3844
rect 41068 3632 41108 6196
rect 41356 5732 41396 7204
rect 41356 5683 41396 5692
rect 41452 8588 41492 8597
rect 41068 3583 41108 3592
rect 40972 3331 41012 3340
rect 40780 2743 40820 2752
rect 40684 2575 40724 2584
rect 41452 1364 41492 8548
rect 41548 8504 41588 9556
rect 41740 9596 41780 10060
rect 41740 9547 41780 9556
rect 41836 10016 41876 10025
rect 41740 9428 41780 9437
rect 41644 9092 41684 9101
rect 41644 8756 41684 9052
rect 41740 9008 41780 9388
rect 41740 8959 41780 8968
rect 41644 8707 41684 8716
rect 41548 8455 41588 8464
rect 41644 8420 41684 8429
rect 41644 7916 41684 8380
rect 41836 8084 41876 9976
rect 42028 9932 42068 10228
rect 41932 9848 41972 9857
rect 41932 9008 41972 9808
rect 42028 9512 42068 9892
rect 42028 9463 42068 9472
rect 42028 9260 42068 9269
rect 42028 9092 42068 9220
rect 42028 9043 42068 9052
rect 41932 8959 41972 8968
rect 41836 8035 41876 8044
rect 42028 8924 42068 8933
rect 41644 7867 41684 7876
rect 41836 7748 41876 7757
rect 41836 7244 41876 7708
rect 41836 7195 41876 7204
rect 41644 3968 41684 3977
rect 41644 2036 41684 3928
rect 41740 3380 41780 3389
rect 41740 2876 41780 3340
rect 42028 3128 42068 8884
rect 42124 7832 42164 11068
rect 42316 11108 42356 11572
rect 42316 11059 42356 11068
rect 42220 9932 42260 9941
rect 42220 9797 42260 9892
rect 42508 9512 42548 11656
rect 42700 10436 42740 12100
rect 44524 11528 44564 11537
rect 44332 11360 44372 11369
rect 43564 11108 43604 11117
rect 42700 10387 42740 10396
rect 42988 10772 43028 10781
rect 42892 10268 42932 10277
rect 42508 9463 42548 9472
rect 42604 10228 42892 10268
rect 42316 8000 42356 8009
rect 42316 7916 42356 7960
rect 42316 7865 42356 7876
rect 42124 7783 42164 7792
rect 42028 3079 42068 3088
rect 41740 2827 41780 2836
rect 41644 1987 41684 1996
rect 41452 1315 41492 1324
rect 40108 643 40148 652
rect 42604 440 42644 10228
rect 42892 10219 42932 10228
rect 42796 9764 42836 9773
rect 42796 9260 42836 9724
rect 42796 9211 42836 9220
rect 42892 9512 42932 9521
rect 42796 8672 42836 8681
rect 42796 8537 42836 8632
rect 42700 8000 42740 8009
rect 42700 7832 42740 7960
rect 42700 7783 42740 7792
rect 42604 391 42644 400
rect 42892 188 42932 9472
rect 42988 8672 43028 10732
rect 43276 10520 43316 10529
rect 43180 10352 43220 10361
rect 43276 10352 43316 10480
rect 43220 10312 43316 10352
rect 43372 10352 43412 10361
rect 43180 10303 43220 10312
rect 43276 10184 43316 10193
rect 43372 10184 43412 10312
rect 43316 10144 43412 10184
rect 43564 10184 43604 11068
rect 43276 10135 43316 10144
rect 43564 10135 43604 10144
rect 43756 10940 43796 10949
rect 43756 10184 43796 10900
rect 43756 10135 43796 10144
rect 43852 10856 43892 10865
rect 43276 9932 43316 9941
rect 43084 9512 43124 9521
rect 43084 9092 43124 9472
rect 43276 9512 43316 9892
rect 43276 9463 43316 9472
rect 43660 9512 43700 9521
rect 43372 9344 43412 9355
rect 43372 9260 43412 9304
rect 43372 9211 43412 9220
rect 43084 9043 43124 9052
rect 43276 9176 43316 9185
rect 42988 8623 43028 8632
rect 43084 8168 43124 8177
rect 43084 8000 43124 8128
rect 43084 7951 43124 7960
rect 43084 5396 43124 5405
rect 43084 2624 43124 5356
rect 43276 4220 43316 9136
rect 43372 9008 43412 9017
rect 43372 8672 43412 8968
rect 43372 8623 43412 8632
rect 43372 8000 43412 8009
rect 43372 7496 43412 7960
rect 43372 7447 43412 7456
rect 43372 7160 43412 7169
rect 43372 7025 43412 7120
rect 43276 4171 43316 4180
rect 43468 6824 43508 6833
rect 43084 2575 43124 2584
rect 43468 2540 43508 6784
rect 43564 6740 43604 6749
rect 43564 4976 43604 6700
rect 43564 4927 43604 4936
rect 43468 2491 43508 2500
rect 42892 139 42932 148
rect 43660 104 43700 9472
rect 43756 9176 43796 9185
rect 43756 8672 43796 9136
rect 43756 8623 43796 8632
rect 43756 7160 43796 7169
rect 43756 7076 43796 7120
rect 43756 7025 43796 7036
rect 43852 7076 43892 10816
rect 44332 10184 44372 11320
rect 44332 10135 44372 10144
rect 44428 10688 44468 10697
rect 44236 10100 44276 10109
rect 44044 9512 44084 9521
rect 43948 9344 43988 9353
rect 43948 8168 43988 9304
rect 44044 8924 44084 9472
rect 44044 8875 44084 8884
rect 43948 8119 43988 8128
rect 43852 7027 43892 7036
rect 44044 7160 44084 7169
rect 43948 6152 43988 6161
rect 43948 5060 43988 6112
rect 43948 5011 43988 5020
rect 44044 4724 44084 7120
rect 44236 6656 44276 10060
rect 44428 9680 44468 10648
rect 44428 9631 44468 9640
rect 44524 8924 44564 11488
rect 44716 11444 44756 11453
rect 44716 10184 44756 11404
rect 44716 10135 44756 10144
rect 45004 11192 45044 11201
rect 44812 9848 44852 9857
rect 44524 8875 44564 8884
rect 44620 9176 44660 9185
rect 44524 8000 44564 8009
rect 44524 7748 44564 7960
rect 44524 7699 44564 7708
rect 44428 7076 44468 7085
rect 44620 7076 44660 9136
rect 44716 8840 44756 8849
rect 44716 8672 44756 8800
rect 44716 8623 44756 8632
rect 44812 7412 44852 9808
rect 44908 9260 44948 9269
rect 44908 8672 44948 9220
rect 44908 8623 44948 8632
rect 45004 8336 45044 11152
rect 45100 11108 45140 11117
rect 45100 10184 45140 11068
rect 45100 10135 45140 10144
rect 45484 10184 45524 10193
rect 45004 8287 45044 8296
rect 45484 8252 45524 10144
rect 45484 8203 45524 8212
rect 46252 8672 46292 8681
rect 46252 8168 46292 8632
rect 46252 8119 46292 8128
rect 44908 8000 44948 8009
rect 44908 7664 44948 7960
rect 44908 7615 44948 7624
rect 46252 7664 46292 7673
rect 46252 7496 46292 7624
rect 46252 7447 46292 7456
rect 44812 7363 44852 7372
rect 44468 7036 44660 7076
rect 44908 7160 44948 7169
rect 44428 7027 44468 7036
rect 44908 6992 44948 7120
rect 44908 6943 44948 6952
rect 46252 6992 46292 7001
rect 46252 6824 46292 6952
rect 46252 6775 46292 6784
rect 44236 6607 44276 6616
rect 44140 6488 44180 6497
rect 44140 6353 44180 6448
rect 44332 6488 44372 6497
rect 44044 4675 44084 4684
rect 44332 3296 44372 6448
rect 44716 6488 44756 6497
rect 44524 5648 44564 5657
rect 44524 5513 44564 5608
rect 44332 3247 44372 3256
rect 44620 4556 44660 4565
rect 44140 2456 44180 2465
rect 44140 1952 44180 2416
rect 44620 2036 44660 4516
rect 44716 3380 44756 6448
rect 44908 5732 44948 5743
rect 44908 5648 44948 5692
rect 44908 5599 44948 5608
rect 44716 3331 44756 3340
rect 44620 1987 44660 1996
rect 45292 2456 45332 2465
rect 44140 1903 44180 1912
rect 44620 1784 44660 1793
rect 44620 1112 44660 1744
rect 45292 1448 45332 2416
rect 45292 1399 45332 1408
rect 45388 1700 45428 1709
rect 44620 1063 44660 1072
rect 45388 776 45428 1660
rect 45388 727 45428 736
rect 33524 64 33544 80
rect 33464 0 33544 64
rect 33656 0 33736 80
rect 33848 0 33928 80
rect 34040 0 34120 80
rect 34232 0 34312 80
rect 34424 0 34504 80
rect 34616 0 34696 80
rect 34808 0 34888 80
rect 35000 0 35080 80
rect 43660 55 43700 64
<< via3 >>
rect 1612 6196 1652 6236
rect 1612 5776 1652 5816
rect 1420 4096 1460 4136
rect 1996 3676 2036 3716
rect 1708 2752 1748 2792
rect 2476 7876 2516 7916
rect 2764 8128 2804 8168
rect 2764 7456 2804 7496
rect 2380 3844 2420 3884
rect 2380 3676 2420 3716
rect 2284 3592 2324 3632
rect 1516 2500 1556 2540
rect 2860 4684 2900 4724
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 4300 8632 4340 8672
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 4972 8296 5012 8336
rect 3244 7792 3284 7832
rect 3148 6448 3188 6488
rect 2956 3088 2996 3128
rect 2476 2752 2516 2792
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 4876 7288 4916 7328
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 3724 6364 3764 6404
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 3724 4852 3764 4892
rect 4204 4936 4244 4976
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 3532 3676 3572 3716
rect 3244 2584 3284 2624
rect 3148 2332 3188 2372
rect 5932 9472 5972 9512
rect 5356 6952 5396 6992
rect 4780 6112 4820 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 4684 5608 4724 5648
rect 4588 5104 4628 5144
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 4012 2080 4052 2120
rect 3532 1996 3572 2036
rect 4396 2668 4436 2708
rect 4108 1912 4148 1952
rect 4300 2164 4340 2204
rect 4300 1828 4340 1868
rect 4492 1660 4532 1700
rect 4684 4852 4724 4892
rect 4780 4768 4820 4808
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 5452 5608 5492 5648
rect 5452 5440 5492 5480
rect 5548 5188 5588 5228
rect 5164 3760 5204 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 6028 7372 6068 7412
rect 6028 6616 6068 6656
rect 5932 5944 5972 5984
rect 5836 5860 5876 5900
rect 6124 6196 6164 6236
rect 6124 5944 6164 5984
rect 5740 5692 5780 5732
rect 5644 4264 5684 4304
rect 6220 5272 6260 5312
rect 5740 3928 5780 3968
rect 6124 4936 6164 4976
rect 5548 3340 5588 3380
rect 6028 3340 6068 3380
rect 4780 2080 4820 2120
rect 4780 1912 4820 1952
rect 5740 2920 5780 2960
rect 6316 4012 6356 4052
rect 6220 3004 6260 3044
rect 6220 2836 6260 2876
rect 5740 2416 5780 2456
rect 6028 2080 6068 2120
rect 6700 8044 6740 8084
rect 6604 6868 6644 6908
rect 7084 8548 7124 8588
rect 6988 8212 7028 8252
rect 6508 6028 6548 6068
rect 6988 7120 7028 7160
rect 7852 8548 7892 8588
rect 7468 7204 7508 7244
rect 7660 7120 7700 7160
rect 6988 6196 7028 6236
rect 6508 5860 6548 5900
rect 6604 4936 6644 4976
rect 6508 3508 6548 3548
rect 6796 6028 6836 6068
rect 7180 6280 7220 6320
rect 7084 6112 7124 6152
rect 7756 6868 7796 6908
rect 7756 6532 7796 6572
rect 7180 5692 7220 5732
rect 6988 4936 7028 4976
rect 7084 5608 7124 5648
rect 6796 4180 6836 4220
rect 7180 5440 7220 5480
rect 7180 5104 7220 5144
rect 7372 5188 7412 5228
rect 7180 4432 7220 4472
rect 6988 4012 7028 4052
rect 7372 3508 7412 3548
rect 7756 5692 7796 5732
rect 8044 8044 8084 8084
rect 7948 7204 7988 7244
rect 8044 5692 8084 5732
rect 8044 5020 8084 5060
rect 7660 4264 7700 4304
rect 6892 3004 6932 3044
rect 6700 2332 6740 2372
rect 7084 2920 7124 2960
rect 7468 3172 7508 3212
rect 7372 2752 7412 2792
rect 7372 2248 7412 2288
rect 7276 2164 7316 2204
rect 7180 2080 7220 2120
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 8236 7120 8276 7160
rect 9004 9472 9044 9512
rect 8908 9304 8948 9344
rect 8428 7456 8468 7496
rect 8524 7288 8564 7328
rect 9100 9136 9140 9176
rect 10060 9220 10100 9260
rect 8716 8296 8756 8336
rect 8812 8212 8852 8252
rect 9004 8044 9044 8084
rect 8812 7708 8852 7748
rect 8812 7456 8852 7496
rect 8620 7036 8660 7076
rect 8428 6616 8468 6656
rect 8620 6196 8660 6236
rect 8524 4768 8564 4808
rect 8908 4936 8948 4976
rect 9004 6868 9044 6908
rect 8812 3340 8852 3380
rect 8620 3256 8660 3296
rect 9868 8548 9908 8588
rect 9196 7288 9236 7328
rect 9292 6616 9332 6656
rect 9388 7288 9428 7328
rect 9196 5776 9236 5816
rect 9388 6280 9428 6320
rect 9676 7372 9716 7412
rect 9676 7204 9716 7244
rect 10924 9976 10964 10016
rect 11020 8884 11060 8924
rect 10348 8044 10388 8084
rect 9964 7288 10004 7328
rect 9772 4852 9812 4892
rect 9388 3172 9428 3212
rect 9484 2752 9524 2792
rect 9004 1996 9044 2036
rect 9964 6280 10004 6320
rect 10636 8044 10676 8084
rect 10924 8044 10964 8084
rect 9964 5272 10004 5312
rect 10060 6028 10100 6068
rect 9964 1996 10004 2036
rect 10540 7540 10580 7580
rect 10540 6364 10580 6404
rect 10156 5608 10196 5648
rect 10348 6028 10388 6068
rect 10348 5776 10388 5816
rect 10444 5692 10484 5732
rect 10252 4768 10292 4808
rect 10252 4264 10292 4304
rect 10252 3760 10292 3800
rect 10156 2752 10196 2792
rect 8044 1660 8084 1700
rect 8620 1660 8660 1700
rect 7372 988 7412 1028
rect 10444 5020 10484 5060
rect 10444 3508 10484 3548
rect 10732 5356 10772 5396
rect 10636 4600 10676 4640
rect 10540 3424 10580 3464
rect 10828 4264 10868 4304
rect 10828 3760 10868 3800
rect 10732 3508 10772 3548
rect 11404 9052 11444 9092
rect 11308 8464 11348 8504
rect 12364 9724 12404 9764
rect 12268 9472 12308 9512
rect 12076 9052 12116 9092
rect 11692 7372 11732 7412
rect 11116 6700 11156 6740
rect 11308 7120 11348 7160
rect 11596 7120 11636 7160
rect 11596 6952 11636 6992
rect 11020 5608 11060 5648
rect 11212 4180 11252 4220
rect 10924 2668 10964 2708
rect 10348 1576 10388 1616
rect 7180 232 7220 272
rect 2860 64 2900 104
rect 11308 1912 11348 1952
rect 11404 2584 11444 2624
rect 12172 7204 12212 7244
rect 12076 5188 12116 5228
rect 12748 9640 12788 9680
rect 13516 9976 13556 10016
rect 13996 9556 14036 9596
rect 12556 7960 12596 8000
rect 12364 6868 12404 6908
rect 12460 6616 12500 6656
rect 12460 4516 12500 4556
rect 12076 3760 12116 3800
rect 13132 8548 13172 8588
rect 13132 7456 13172 7496
rect 12940 5776 12980 5816
rect 12844 4852 12884 4892
rect 12652 4768 12692 4808
rect 12748 4600 12788 4640
rect 13036 4768 13076 4808
rect 13324 7288 13364 7328
rect 13324 6532 13364 6572
rect 13228 5692 13268 5732
rect 12556 3508 12596 3548
rect 12268 3340 12308 3380
rect 11980 2584 12020 2624
rect 11788 1492 11828 1532
rect 11596 64 11636 104
rect 12940 4012 12980 4052
rect 13132 3508 13172 3548
rect 12268 2687 12308 2708
rect 12268 2668 12308 2687
rect 12748 2836 12788 2876
rect 12940 2836 12980 2876
rect 12940 2248 12980 2288
rect 13708 4264 13748 4304
rect 13612 3508 13652 3548
rect 13612 3340 13652 3380
rect 13036 2164 13076 2204
rect 13516 3004 13556 3044
rect 12748 1996 12788 2036
rect 12844 2080 12884 2120
rect 12940 1324 12980 1364
rect 12940 400 12980 440
rect 13420 2752 13460 2792
rect 13132 1240 13172 1280
rect 13228 2164 13268 2204
rect 13420 1996 13460 2036
rect 13228 400 13268 440
rect 13324 1240 13364 1280
rect 13900 3424 13940 3464
rect 14380 9388 14420 9428
rect 14380 8968 14420 9008
rect 14188 8548 14228 8588
rect 14092 6532 14132 6572
rect 14092 6028 14132 6068
rect 13996 3340 14036 3380
rect 13804 3004 13844 3044
rect 13900 2920 13940 2960
rect 13708 2248 13748 2288
rect 13900 1576 13940 1616
rect 14380 6952 14420 6992
rect 14572 8212 14612 8252
rect 14572 6784 14612 6824
rect 14380 6364 14420 6404
rect 14188 5608 14228 5648
rect 14284 6280 14324 6320
rect 14284 4516 14324 4556
rect 14476 4264 14516 4304
rect 14572 4600 14612 4640
rect 14380 4012 14420 4052
rect 14380 3760 14420 3800
rect 15052 7960 15092 8000
rect 14764 4852 14804 4892
rect 14956 5272 14996 5312
rect 14860 4264 14900 4304
rect 15532 9472 15572 9512
rect 15436 8716 15476 8756
rect 15148 5440 15188 5480
rect 14956 4012 14996 4052
rect 14572 3004 14612 3044
rect 14572 1240 14612 1280
rect 14476 1072 14516 1112
rect 14476 232 14516 272
rect 15148 3172 15188 3212
rect 14956 1744 14996 1784
rect 14860 1576 14900 1616
rect 14764 568 14804 608
rect 14860 1408 14900 1448
rect 15052 988 15092 1028
rect 15436 6364 15476 6404
rect 15820 8464 15860 8504
rect 15724 8380 15764 8420
rect 15628 7960 15668 8000
rect 15436 1576 15476 1616
rect 16108 8884 16148 8924
rect 15916 7204 15956 7244
rect 15820 6196 15860 6236
rect 15724 5272 15764 5312
rect 15820 5860 15860 5900
rect 15916 5104 15956 5144
rect 15820 4180 15860 4220
rect 15820 1912 15860 1952
rect 15724 988 15764 1028
rect 16108 5692 16148 5732
rect 16108 4348 16148 4388
rect 16108 3760 16148 3800
rect 17740 9472 17780 9512
rect 16300 5776 16340 5816
rect 16684 5944 16724 5984
rect 16588 4516 16628 4556
rect 16492 4264 16532 4304
rect 16684 4264 16724 4304
rect 16492 1408 16532 1448
rect 16588 2752 16628 2792
rect 17164 5524 17204 5564
rect 16972 5020 17012 5060
rect 17068 5272 17108 5312
rect 16972 3340 17012 3380
rect 16972 2920 17012 2960
rect 16972 2332 17012 2372
rect 16972 1996 17012 2036
rect 17452 7204 17492 7244
rect 17452 6364 17492 6404
rect 17452 5944 17492 5984
rect 17740 8044 17780 8084
rect 17644 7288 17684 7328
rect 18604 9724 18644 9764
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 18412 9472 18452 9512
rect 18124 8716 18164 8756
rect 17932 7540 17972 7580
rect 18028 7960 18068 8000
rect 17356 3004 17396 3044
rect 17644 5356 17684 5396
rect 17644 4852 17684 4892
rect 17548 2752 17588 2792
rect 17452 2584 17492 2624
rect 17932 4012 17972 4052
rect 18220 7540 18260 7580
rect 18220 7288 18260 7328
rect 17740 2836 17780 2876
rect 17740 2584 17780 2624
rect 16972 1408 17012 1448
rect 17548 1744 17588 1784
rect 17740 1324 17780 1364
rect 18028 2668 18068 2708
rect 18028 2164 18068 2204
rect 18028 1744 18068 1784
rect 18220 2920 18260 2960
rect 18412 7288 18452 7328
rect 18988 8716 19028 8756
rect 19372 9052 19412 9092
rect 18604 8464 18644 8504
rect 19276 8464 19316 8504
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 19084 7960 19124 8000
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 18412 6280 18452 6320
rect 18604 6280 18644 6320
rect 19468 8044 19508 8084
rect 18508 6028 18548 6068
rect 18700 5776 18740 5816
rect 18892 5692 18932 5732
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 19372 7540 19412 7580
rect 19372 5272 19412 5312
rect 18508 3424 18548 3464
rect 18412 3172 18452 3212
rect 18508 2920 18548 2960
rect 19180 4264 19220 4304
rect 19372 4432 19412 4472
rect 18700 4180 18740 4220
rect 18700 3760 18740 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 18412 2080 18452 2120
rect 18220 1912 18260 1952
rect 18316 1240 18356 1280
rect 18604 1492 18644 1532
rect 18796 2836 18836 2876
rect 19084 3172 19124 3212
rect 19084 2836 19124 2876
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 20140 9724 20180 9764
rect 20620 9640 20660 9680
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 21196 9808 21236 9848
rect 20908 9724 20948 9764
rect 19660 7372 19700 7412
rect 19756 6616 19796 6656
rect 19756 6280 19796 6320
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 20620 7456 20660 7496
rect 20140 6784 20180 6824
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 19948 5776 19988 5816
rect 20236 5356 20276 5396
rect 20044 5272 20084 5312
rect 19660 4264 19700 4304
rect 19564 4180 19604 4220
rect 19372 3172 19412 3212
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 19276 1996 19316 2036
rect 19372 1912 19412 1952
rect 19276 1072 19316 1112
rect 19084 568 19124 608
rect 19756 2920 19796 2960
rect 19948 4516 19988 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 20716 6784 20756 6824
rect 20716 4600 20756 4640
rect 21004 8044 21044 8084
rect 21004 6364 21044 6404
rect 21004 5776 21044 5816
rect 20140 4264 20180 4304
rect 20620 4264 20660 4304
rect 20620 4012 20660 4052
rect 19948 3004 19988 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 20044 2836 20084 2876
rect 20524 2248 20564 2288
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 20044 988 20084 1028
rect 21004 5272 21044 5312
rect 20812 4012 20852 4052
rect 20908 3172 20948 3212
rect 21772 9556 21812 9596
rect 21292 9052 21332 9092
rect 22156 9556 22196 9596
rect 22060 9472 22100 9512
rect 22060 9052 22100 9092
rect 21292 7456 21332 7496
rect 21196 6616 21236 6656
rect 21676 8548 21716 8588
rect 21484 7288 21524 7328
rect 21580 5692 21620 5732
rect 21772 7960 21812 8000
rect 21772 7540 21812 7580
rect 21772 7372 21812 7412
rect 22156 7540 22196 7580
rect 22252 7372 22292 7412
rect 22348 7288 22388 7328
rect 22444 7204 22484 7244
rect 22060 6784 22100 6824
rect 21868 6196 21908 6236
rect 22252 5776 22292 5816
rect 21388 4768 21428 4808
rect 21196 4180 21236 4220
rect 21484 3172 21524 3212
rect 20812 1744 20852 1784
rect 20716 1576 20756 1616
rect 21676 3760 21716 3800
rect 21676 2920 21716 2960
rect 21676 2332 21716 2372
rect 21580 1828 21620 1868
rect 21580 1324 21620 1364
rect 21964 4516 22004 4556
rect 22156 4180 22196 4220
rect 22060 3592 22100 3632
rect 21964 2752 22004 2792
rect 22636 7456 22676 7496
rect 22540 5776 22580 5816
rect 23116 7960 23156 8000
rect 23500 8380 23540 8420
rect 22924 7456 22964 7496
rect 22348 5356 22388 5396
rect 22348 2752 22388 2792
rect 22444 2248 22484 2288
rect 22828 7372 22868 7412
rect 23212 6364 23252 6404
rect 22924 6280 22964 6320
rect 23020 3592 23060 3632
rect 22732 2752 22772 2792
rect 22636 2332 22676 2372
rect 22924 3172 22964 3212
rect 23116 3004 23156 3044
rect 23116 2836 23156 2876
rect 22924 2752 22964 2792
rect 23212 2752 23252 2792
rect 23020 2668 23060 2708
rect 23884 6196 23924 6236
rect 23788 5440 23828 5480
rect 24076 8716 24116 8756
rect 24268 7540 24308 7580
rect 24172 5272 24212 5312
rect 23884 4432 23924 4472
rect 23308 2080 23348 2120
rect 24556 6280 24596 6320
rect 24556 4264 24596 4304
rect 24460 3592 24500 3632
rect 24172 2752 24212 2792
rect 24460 3172 24500 3212
rect 24556 2668 24596 2708
rect 25420 9388 25460 9428
rect 25036 8716 25076 8756
rect 24940 7960 24980 8000
rect 25132 7456 25172 7496
rect 24940 5104 24980 5144
rect 24844 4264 24884 4304
rect 25516 5776 25556 5816
rect 24844 3508 24884 3548
rect 24844 2584 24884 2624
rect 25132 5272 25172 5312
rect 24940 1576 24980 1616
rect 25516 5356 25556 5396
rect 25516 4432 25556 4472
rect 26476 9556 26516 9596
rect 26284 9388 26324 9428
rect 25708 6364 25748 6404
rect 25708 4852 25748 4892
rect 25228 4012 25268 4052
rect 25132 2500 25172 2540
rect 25612 3172 25652 3212
rect 26572 8968 26612 9008
rect 26284 7540 26324 7580
rect 26092 6784 26132 6824
rect 25996 5860 26036 5900
rect 26188 5104 26228 5144
rect 25804 3760 25844 3800
rect 25804 1576 25844 1616
rect 27148 7960 27188 8000
rect 27436 7372 27476 7412
rect 26572 6112 26612 6152
rect 26476 5188 26516 5228
rect 26668 5944 26708 5984
rect 26860 6112 26900 6152
rect 26764 5860 26804 5900
rect 26764 5440 26804 5480
rect 26572 652 26612 692
rect 26956 5188 26996 5228
rect 26956 4600 26996 4640
rect 27628 9976 27668 10016
rect 28396 9388 28436 9428
rect 28012 8716 28052 8756
rect 28972 8716 29012 8756
rect 28012 8044 28052 8084
rect 28780 8212 28820 8252
rect 28108 6616 28148 6656
rect 27340 4264 27380 4304
rect 26956 3676 26996 3716
rect 26956 820 26996 860
rect 27724 1828 27764 1868
rect 28204 3088 28244 3128
rect 28396 5440 28436 5480
rect 28396 4348 28436 4388
rect 28588 5524 28628 5564
rect 28684 5188 28724 5228
rect 28876 5440 28916 5480
rect 28780 5104 28820 5144
rect 28684 4432 28724 4472
rect 28876 4852 28916 4892
rect 28780 4180 28820 4220
rect 28588 2752 28628 2792
rect 28780 2668 28820 2708
rect 29644 9976 29684 10016
rect 28972 1996 29012 2036
rect 29164 3592 29204 3632
rect 29260 2080 29300 2120
rect 29164 1996 29204 2036
rect 29740 4516 29780 4556
rect 29644 2752 29684 2792
rect 30220 7540 30260 7580
rect 29932 6364 29972 6404
rect 30508 7372 30548 7412
rect 30220 6616 30260 6656
rect 30124 6364 30164 6404
rect 30316 5524 30356 5564
rect 30412 5356 30452 5396
rect 30508 5440 30548 5480
rect 30508 4432 30548 4472
rect 30508 3676 30548 3716
rect 30316 3592 30356 3632
rect 29836 2836 29876 2876
rect 29548 1576 29588 1616
rect 29836 1240 29876 1280
rect 29644 400 29684 440
rect 30412 3508 30452 3548
rect 30220 2500 30260 2540
rect 30220 2248 30260 2288
rect 30508 2584 30548 2624
rect 30700 6616 30740 6656
rect 30700 6364 30740 6404
rect 30700 3844 30740 3884
rect 30700 3004 30740 3044
rect 30700 2668 30740 2708
rect 30604 1408 30644 1448
rect 30412 904 30452 944
rect 31372 6112 31412 6152
rect 30892 5776 30932 5816
rect 31276 4852 31316 4892
rect 30892 1408 30932 1448
rect 31276 2836 31316 2876
rect 32332 9472 32372 9512
rect 32524 9388 32564 9428
rect 32524 8800 32564 8840
rect 31852 8716 31892 8756
rect 31660 5776 31700 5816
rect 31756 5860 31796 5900
rect 31660 3088 31700 3128
rect 31660 2332 31700 2372
rect 31468 1660 31508 1700
rect 31564 1324 31604 1364
rect 31852 4852 31892 4892
rect 31756 1240 31796 1280
rect 31852 3760 31892 3800
rect 31660 652 31700 692
rect 32332 7372 32372 7412
rect 32236 7204 32276 7244
rect 32236 6616 32276 6656
rect 32044 4180 32084 4220
rect 32044 1828 32084 1868
rect 32428 7288 32468 7328
rect 32428 4936 32468 4976
rect 32332 3844 32372 3884
rect 32332 3508 32372 3548
rect 32332 2332 32372 2372
rect 32236 400 32276 440
rect 32332 1408 32372 1448
rect 32428 820 32468 860
rect 33004 9892 33044 9932
rect 32908 8968 32948 9008
rect 32716 8884 32756 8924
rect 33196 9724 33236 9764
rect 33292 8968 33332 9008
rect 33196 8548 33236 8588
rect 32908 7456 32948 7496
rect 33100 7456 33140 7496
rect 33196 6280 33236 6320
rect 32716 4852 32756 4892
rect 32716 4264 32756 4304
rect 32716 3844 32756 3884
rect 32716 3172 32756 3212
rect 32620 2752 32660 2792
rect 33100 4600 33140 4640
rect 33196 5356 33236 5396
rect 32908 3004 32948 3044
rect 34252 9976 34292 10016
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 34156 9556 34196 9596
rect 33580 7456 33620 7496
rect 33676 8884 33716 8924
rect 33484 6364 33524 6404
rect 33388 5356 33428 5396
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 33964 7960 34004 8000
rect 33772 7540 33812 7580
rect 33868 7372 33908 7412
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 34636 9892 34676 9932
rect 33676 5524 33716 5564
rect 33388 4012 33428 4052
rect 33484 3004 33524 3044
rect 33484 2836 33524 2876
rect 33388 2332 33428 2372
rect 32812 1408 32852 1448
rect 33292 1576 33332 1616
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 34252 5104 34292 5144
rect 33772 4180 33812 4220
rect 34252 4348 34292 4388
rect 34828 10228 34868 10268
rect 34828 9724 34868 9764
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 34924 9388 34964 9428
rect 34828 7456 34868 7496
rect 34444 4180 34484 4220
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 34636 5776 34676 5816
rect 34732 4348 34772 4388
rect 33964 2836 34004 2876
rect 33868 2668 33908 2708
rect 34444 3004 34484 3044
rect 33964 2500 34004 2540
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 34540 2584 34580 2624
rect 34636 3004 34676 3044
rect 34924 2836 34964 2876
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 35788 10228 35828 10268
rect 38764 10228 38804 10268
rect 35884 9388 35924 9428
rect 37420 9556 37460 9596
rect 36748 9472 36788 9512
rect 35596 6364 35636 6404
rect 35404 6196 35444 6236
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 35116 3676 35156 3716
rect 36940 9304 36980 9344
rect 36748 8716 36788 8756
rect 36844 8212 36884 8252
rect 36844 7960 36884 8000
rect 36268 7288 36308 7328
rect 35980 5524 36020 5564
rect 35980 4852 36020 4892
rect 35788 3928 35828 3968
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 36748 6784 36788 6824
rect 36652 5860 36692 5900
rect 36940 5188 36980 5228
rect 37132 7960 37172 8000
rect 37228 6616 37268 6656
rect 36556 4012 36596 4052
rect 35116 2500 35156 2540
rect 36076 2668 36116 2708
rect 36460 3172 36500 3212
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 37804 8212 37844 8252
rect 37420 6532 37460 6572
rect 37708 7204 37748 7244
rect 37516 6280 37556 6320
rect 37612 3592 37652 3632
rect 37420 2920 37460 2960
rect 38092 6700 38132 6740
rect 37900 5020 37940 5060
rect 37900 4096 37940 4136
rect 38092 4600 38132 4640
rect 38380 9472 38420 9512
rect 40300 10900 40340 10940
rect 39244 10228 39284 10268
rect 38956 9640 38996 9680
rect 39340 9976 39380 10016
rect 39244 9556 39284 9596
rect 40108 9892 40148 9932
rect 38572 4768 38612 4808
rect 38668 2332 38708 2372
rect 38956 5104 38996 5144
rect 39148 5440 39188 5480
rect 38860 4096 38900 4136
rect 39532 4432 39572 4472
rect 39628 3508 39668 3548
rect 37324 1576 37364 1616
rect 36748 1324 36788 1364
rect 36172 904 36212 944
rect 40300 9640 40340 9680
rect 40204 9388 40244 9428
rect 41452 9304 41492 9344
rect 40300 6784 40340 6824
rect 40300 6112 40340 6152
rect 40588 6868 40628 6908
rect 40492 3844 40532 3884
rect 40972 3844 41012 3884
rect 40300 3424 40340 3464
rect 41644 9052 41684 9092
rect 42028 9052 42068 9092
rect 42220 9892 42260 9932
rect 42316 7876 42356 7916
rect 42028 3088 42068 3128
rect 42796 8632 42836 8672
rect 42700 7792 42740 7832
rect 43756 10900 43796 10940
rect 43372 9304 43412 9344
rect 43084 8128 43124 8168
rect 43372 7120 43412 7160
rect 43756 9136 43796 9176
rect 43756 7036 43796 7076
rect 44524 7708 44564 7748
rect 44716 8800 44756 8840
rect 44908 9220 44948 9260
rect 44908 7624 44948 7664
rect 44908 6952 44948 6992
rect 44140 6448 44180 6488
rect 44044 4684 44084 4724
rect 44524 5608 44564 5648
rect 44332 3256 44372 3296
rect 44140 2416 44180 2456
rect 44908 5692 44948 5732
rect 44716 3340 44756 3380
<< metal4 >>
rect 40291 10900 40300 10940
rect 40340 10900 43756 10940
rect 43796 10900 43805 10940
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 20039 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20425 10604
rect 35159 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 35545 10604
rect 34819 10228 34828 10268
rect 34868 10228 35788 10268
rect 35828 10228 35837 10268
rect 38755 10228 38764 10268
rect 38804 10228 39244 10268
rect 39284 10228 39293 10268
rect 10915 9976 10924 10016
rect 10964 9976 13516 10016
rect 13556 9976 13565 10016
rect 27619 9976 27628 10016
rect 27668 9976 29644 10016
rect 29684 9976 29693 10016
rect 34243 9976 34252 10016
rect 34292 9976 39340 10016
rect 39380 9976 39389 10016
rect 32995 9892 33004 9932
rect 33044 9892 34636 9932
rect 34676 9892 34685 9932
rect 40099 9892 40108 9932
rect 40148 9892 42220 9932
rect 42260 9892 42269 9932
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 21187 9808 21196 9848
rect 21236 9808 33236 9848
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 33196 9764 33236 9808
rect 12355 9724 12364 9764
rect 12404 9724 18604 9764
rect 18644 9724 18653 9764
rect 20131 9724 20140 9764
rect 20180 9724 20908 9764
rect 20948 9724 20957 9764
rect 33187 9724 33196 9764
rect 33236 9724 34828 9764
rect 34868 9724 34877 9764
rect 12739 9640 12748 9680
rect 12788 9640 20620 9680
rect 20660 9640 20669 9680
rect 30220 9640 37556 9680
rect 38947 9640 38956 9680
rect 38996 9640 40300 9680
rect 40340 9640 40349 9680
rect 30220 9596 30260 9640
rect 37516 9596 37556 9640
rect 13987 9556 13996 9596
rect 14036 9556 21772 9596
rect 21812 9556 22156 9596
rect 22196 9556 22205 9596
rect 26467 9556 26476 9596
rect 26516 9556 30260 9596
rect 34147 9556 34156 9596
rect 34196 9556 37420 9596
rect 37460 9556 37469 9596
rect 37516 9556 39244 9596
rect 39284 9556 39293 9596
rect 5923 9472 5932 9512
rect 5972 9472 9004 9512
rect 9044 9472 9053 9512
rect 12259 9472 12268 9512
rect 12308 9472 15532 9512
rect 15572 9472 17740 9512
rect 17780 9472 17789 9512
rect 18403 9472 18412 9512
rect 18452 9472 22060 9512
rect 22100 9472 22109 9512
rect 32323 9472 32332 9512
rect 32372 9472 35924 9512
rect 36739 9472 36748 9512
rect 36788 9472 38380 9512
rect 38420 9472 38429 9512
rect 35884 9428 35924 9472
rect 14371 9388 14380 9428
rect 14420 9388 14572 9428
rect 14612 9388 14621 9428
rect 25411 9388 25420 9428
rect 25460 9388 26284 9428
rect 26324 9388 28396 9428
rect 28436 9388 28445 9428
rect 32515 9388 32524 9428
rect 32564 9388 34924 9428
rect 34964 9388 34973 9428
rect 35875 9388 35884 9428
rect 35924 9388 40204 9428
rect 40244 9388 40253 9428
rect 8899 9304 8908 9344
rect 8948 9304 36940 9344
rect 36980 9304 36989 9344
rect 41443 9304 41452 9344
rect 41492 9304 43372 9344
rect 43412 9304 43421 9344
rect 10051 9220 10060 9260
rect 10100 9220 44908 9260
rect 44948 9220 44957 9260
rect 9091 9136 9100 9176
rect 9140 9136 43756 9176
rect 43796 9136 43805 9176
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 11395 9052 11404 9092
rect 11444 9052 12076 9092
rect 12116 9052 19372 9092
rect 19412 9052 19421 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 21283 9052 21292 9092
rect 21332 9052 22060 9092
rect 22100 9052 22109 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 41635 9052 41644 9092
rect 41684 9052 42028 9092
rect 42068 9052 42077 9092
rect 14371 8968 14380 9008
rect 14420 8968 26572 9008
rect 26612 8968 26621 9008
rect 32899 8968 32908 9008
rect 32948 8968 33292 9008
rect 33332 8968 33341 9008
rect 11011 8884 11020 8924
rect 11060 8884 16108 8924
rect 16148 8884 16157 8924
rect 32707 8884 32716 8924
rect 32756 8884 33676 8924
rect 33716 8884 33725 8924
rect 32515 8800 32524 8840
rect 32564 8800 44716 8840
rect 44756 8800 44765 8840
rect 15427 8716 15436 8756
rect 15476 8716 18124 8756
rect 18164 8716 18988 8756
rect 19028 8716 19037 8756
rect 24067 8716 24076 8756
rect 24116 8716 25036 8756
rect 25076 8716 25085 8756
rect 28003 8716 28012 8756
rect 28052 8716 28972 8756
rect 29012 8716 29021 8756
rect 31843 8716 31852 8756
rect 31892 8716 36748 8756
rect 36788 8716 36797 8756
rect 4291 8632 4300 8672
rect 4340 8632 42796 8672
rect 42836 8632 42845 8672
rect 7075 8548 7084 8588
rect 7124 8548 7852 8588
rect 7892 8548 9868 8588
rect 9908 8548 9917 8588
rect 13123 8548 13132 8588
rect 13172 8548 14188 8588
rect 14228 8548 21676 8588
rect 21716 8548 21725 8588
rect 33101 8548 33196 8588
rect 33236 8548 33245 8588
rect 11299 8464 11308 8504
rect 11348 8464 15820 8504
rect 15860 8464 15869 8504
rect 18595 8464 18604 8504
rect 18644 8464 19276 8504
rect 19316 8464 19325 8504
rect 15715 8380 15724 8420
rect 15764 8380 23500 8420
rect 23540 8380 23549 8420
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 4963 8296 4972 8336
rect 5012 8296 8716 8336
rect 8756 8296 8765 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 6979 8212 6988 8252
rect 7028 8212 8812 8252
rect 8852 8212 8861 8252
rect 14563 8212 14572 8252
rect 14612 8212 28780 8252
rect 28820 8212 28829 8252
rect 36835 8212 36844 8252
rect 36884 8212 37804 8252
rect 37844 8212 37853 8252
rect 2755 8128 2764 8168
rect 2804 8128 43084 8168
rect 43124 8128 43133 8168
rect 6691 8044 6700 8084
rect 6740 8044 8044 8084
rect 8084 8044 8093 8084
rect 8995 8044 9004 8084
rect 9044 8044 10348 8084
rect 10388 8044 10397 8084
rect 10627 8044 10636 8084
rect 10676 8044 10924 8084
rect 10964 8044 10973 8084
rect 17731 8044 17740 8084
rect 17780 8044 19468 8084
rect 19508 8044 19517 8084
rect 20995 8044 21004 8084
rect 21044 8044 28012 8084
rect 28052 8044 28061 8084
rect 12547 7960 12556 8000
rect 12596 7960 15052 8000
rect 15092 7960 15101 8000
rect 15533 7960 15628 8000
rect 15668 7960 15677 8000
rect 18019 7960 18028 8000
rect 18068 7960 19084 8000
rect 19124 7960 19133 8000
rect 21763 7960 21772 8000
rect 21812 7960 23116 8000
rect 23156 7960 23165 8000
rect 24931 7960 24940 8000
rect 24980 7960 27148 8000
rect 27188 7960 27197 8000
rect 33955 7960 33964 8000
rect 34004 7960 36844 8000
rect 36884 7960 37132 8000
rect 37172 7960 37181 8000
rect 2467 7876 2476 7916
rect 2516 7876 42316 7916
rect 42356 7876 42365 7916
rect 3235 7792 3244 7832
rect 3284 7792 42700 7832
rect 42740 7792 42749 7832
rect 8803 7708 8812 7748
rect 8852 7708 44524 7748
rect 44564 7708 44573 7748
rect 2860 7624 44908 7664
rect 44948 7624 44957 7664
rect 2860 7496 2900 7624
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 10531 7540 10540 7580
rect 10580 7540 17932 7580
rect 17972 7540 17981 7580
rect 18211 7540 18220 7580
rect 18260 7540 19372 7580
rect 19412 7540 19421 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 21763 7540 21772 7580
rect 21812 7540 22156 7580
rect 22196 7540 22205 7580
rect 24259 7540 24268 7580
rect 24308 7540 26284 7580
rect 26324 7540 26333 7580
rect 30211 7540 30220 7580
rect 30260 7540 33772 7580
rect 33812 7540 33821 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 2755 7456 2764 7496
rect 2804 7456 2900 7496
rect 8419 7456 8428 7496
rect 8468 7456 8812 7496
rect 8852 7456 8861 7496
rect 13123 7456 13132 7496
rect 13172 7456 20620 7496
rect 20660 7456 20669 7496
rect 21283 7456 21292 7496
rect 21332 7456 22636 7496
rect 22676 7456 22685 7496
rect 22915 7456 22924 7496
rect 22964 7456 25132 7496
rect 25172 7456 25181 7496
rect 32899 7456 32908 7496
rect 32948 7456 33100 7496
rect 33140 7456 33149 7496
rect 33571 7456 33580 7496
rect 33620 7456 34828 7496
rect 34868 7456 34877 7496
rect 6019 7372 6028 7412
rect 6068 7372 9676 7412
rect 9716 7372 9725 7412
rect 11683 7372 11692 7412
rect 11732 7372 19660 7412
rect 19700 7372 19709 7412
rect 21763 7372 21772 7412
rect 21812 7372 22252 7412
rect 22292 7372 22301 7412
rect 22819 7372 22828 7412
rect 22868 7372 27436 7412
rect 27476 7372 27485 7412
rect 30499 7372 30508 7412
rect 30548 7372 32332 7412
rect 32372 7372 33868 7412
rect 33908 7372 33917 7412
rect 4867 7288 4876 7328
rect 4916 7288 8524 7328
rect 8564 7288 8573 7328
rect 9187 7288 9196 7328
rect 9236 7288 9245 7328
rect 9379 7288 9388 7328
rect 9428 7288 9964 7328
rect 10004 7288 10013 7328
rect 13315 7288 13324 7328
rect 13364 7288 17644 7328
rect 17684 7288 17693 7328
rect 18211 7288 18220 7328
rect 18260 7288 18412 7328
rect 18452 7288 18461 7328
rect 21475 7288 21484 7328
rect 21524 7288 22348 7328
rect 22388 7288 22397 7328
rect 32419 7288 32428 7328
rect 32468 7288 36268 7328
rect 36308 7288 36317 7328
rect 9196 7244 9236 7288
rect 7459 7204 7468 7244
rect 7508 7204 7948 7244
rect 7988 7204 7997 7244
rect 9196 7204 9676 7244
rect 9716 7204 9725 7244
rect 12163 7204 12172 7244
rect 12212 7204 15916 7244
rect 15956 7204 15965 7244
rect 17443 7204 17452 7244
rect 17492 7204 22444 7244
rect 22484 7204 22493 7244
rect 32227 7204 32236 7244
rect 32276 7204 37708 7244
rect 37748 7204 37757 7244
rect 6979 7120 6988 7160
rect 7028 7120 7660 7160
rect 7700 7120 7709 7160
rect 8227 7120 8236 7160
rect 8276 7120 11308 7160
rect 11348 7120 11357 7160
rect 11587 7120 11596 7160
rect 11636 7120 43372 7160
rect 43412 7120 43421 7160
rect 8611 7036 8620 7076
rect 8660 7036 43756 7076
rect 43796 7036 43805 7076
rect 5347 6952 5356 6992
rect 5396 6952 11596 6992
rect 11636 6952 11645 6992
rect 14371 6952 14380 6992
rect 14420 6952 44908 6992
rect 44948 6952 44957 6992
rect 6595 6868 6604 6908
rect 6644 6868 7756 6908
rect 7796 6868 9004 6908
rect 9044 6868 9053 6908
rect 12355 6868 12364 6908
rect 12404 6868 40588 6908
rect 40628 6868 40637 6908
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 14477 6784 14572 6824
rect 14612 6784 14621 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 19555 6784 19564 6824
rect 19604 6784 20140 6824
rect 20180 6784 20189 6824
rect 20707 6784 20716 6824
rect 20756 6784 22060 6824
rect 22100 6784 26092 6824
rect 26132 6784 26141 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 36739 6784 36748 6824
rect 36788 6784 40300 6824
rect 40340 6784 40349 6824
rect 11107 6700 11116 6740
rect 11156 6700 38092 6740
rect 38132 6700 38141 6740
rect 6019 6616 6028 6656
rect 6068 6616 8428 6656
rect 8468 6616 9292 6656
rect 9332 6616 9341 6656
rect 12451 6616 12460 6656
rect 12500 6616 19756 6656
rect 19796 6616 19805 6656
rect 21187 6616 21196 6656
rect 21236 6616 28108 6656
rect 28148 6616 28157 6656
rect 30211 6616 30220 6656
rect 30260 6616 30700 6656
rect 30740 6616 30749 6656
rect 32227 6616 32236 6656
rect 32276 6616 37228 6656
rect 37268 6616 37277 6656
rect 7747 6532 7756 6572
rect 7796 6532 13324 6572
rect 13364 6532 13373 6572
rect 14083 6532 14092 6572
rect 14132 6532 37420 6572
rect 37460 6532 37469 6572
rect 3139 6448 3148 6488
rect 3188 6448 44140 6488
rect 44180 6448 44189 6488
rect 3715 6364 3724 6404
rect 3764 6364 10540 6404
rect 10580 6364 10589 6404
rect 14371 6364 14380 6404
rect 14420 6364 15436 6404
rect 15476 6364 15485 6404
rect 17443 6364 17452 6404
rect 17492 6364 21004 6404
rect 21044 6364 21053 6404
rect 21196 6364 23212 6404
rect 23252 6364 23261 6404
rect 25699 6364 25708 6404
rect 25748 6364 29932 6404
rect 29972 6364 29981 6404
rect 30115 6364 30124 6404
rect 30164 6364 30173 6404
rect 30691 6364 30700 6404
rect 30740 6364 33484 6404
rect 33524 6364 33533 6404
rect 34627 6364 34636 6404
rect 34676 6364 35596 6404
rect 35636 6364 35645 6404
rect 21196 6320 21236 6364
rect 7171 6280 7180 6320
rect 7220 6280 9388 6320
rect 9428 6280 9437 6320
rect 9955 6280 9964 6320
rect 10004 6280 10100 6320
rect 14275 6280 14284 6320
rect 14324 6280 18412 6320
rect 18452 6280 18604 6320
rect 18644 6280 19564 6320
rect 19604 6280 19613 6320
rect 19747 6280 19756 6320
rect 19796 6280 21236 6320
rect 22915 6280 22924 6320
rect 22964 6280 24556 6320
rect 24596 6280 24605 6320
rect 1603 6196 1612 6236
rect 1652 6196 6124 6236
rect 6164 6196 6173 6236
rect 6979 6196 6988 6236
rect 7028 6196 8620 6236
rect 8660 6196 8669 6236
rect 10060 6152 10100 6280
rect 30124 6236 30164 6364
rect 33187 6280 33196 6320
rect 33236 6280 37516 6320
rect 37556 6280 37565 6320
rect 15811 6196 15820 6236
rect 15860 6196 21868 6236
rect 21908 6196 21917 6236
rect 23875 6196 23884 6236
rect 23924 6196 30164 6236
rect 32131 6196 32140 6236
rect 32180 6196 35404 6236
rect 35444 6196 35453 6236
rect 4771 6112 4780 6152
rect 4820 6112 7084 6152
rect 7124 6112 7133 6152
rect 10060 6112 19852 6152
rect 19892 6112 19901 6152
rect 26563 6112 26572 6152
rect 26612 6112 26860 6152
rect 26900 6112 26909 6152
rect 31363 6112 31372 6152
rect 31412 6112 40300 6152
rect 40340 6112 40349 6152
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 6499 6028 6508 6068
rect 6548 6028 6796 6068
rect 6836 6028 6845 6068
rect 10051 6028 10060 6068
rect 10100 6028 10348 6068
rect 10388 6028 10397 6068
rect 14083 6028 14092 6068
rect 14132 6028 18508 6068
rect 18548 6028 18557 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 5923 5944 5932 5984
rect 5972 5944 6124 5984
rect 6164 5944 6173 5984
rect 12940 5944 16684 5984
rect 16724 5944 17452 5984
rect 17492 5944 17501 5984
rect 20803 5944 20812 5984
rect 20852 5944 26668 5984
rect 26708 5944 26717 5984
rect 5827 5860 5836 5900
rect 5876 5860 6508 5900
rect 6548 5860 6557 5900
rect 12940 5816 12980 5944
rect 15811 5860 15820 5900
rect 15860 5860 25996 5900
rect 26036 5860 26045 5900
rect 26755 5860 26764 5900
rect 26804 5860 31756 5900
rect 31796 5860 36652 5900
rect 36692 5860 36701 5900
rect 25996 5816 26036 5860
rect 1603 5776 1612 5816
rect 1652 5776 9196 5816
rect 9236 5776 9245 5816
rect 10339 5776 10348 5816
rect 10388 5776 12940 5816
rect 12980 5776 12989 5816
rect 16291 5776 16300 5816
rect 16340 5776 18700 5816
rect 18740 5776 18749 5816
rect 19747 5776 19756 5816
rect 19796 5776 19948 5816
rect 19988 5776 19997 5816
rect 20140 5776 20812 5816
rect 20852 5776 20861 5816
rect 20995 5776 21004 5816
rect 21044 5776 22252 5816
rect 22292 5776 22301 5816
rect 22531 5776 22540 5816
rect 22580 5776 24556 5816
rect 24596 5776 25516 5816
rect 25556 5776 25565 5816
rect 25996 5776 30892 5816
rect 30932 5776 30941 5816
rect 31651 5776 31660 5816
rect 31700 5776 34636 5816
rect 34676 5776 34685 5816
rect 20140 5732 20180 5776
rect 5731 5692 5740 5732
rect 5780 5692 7180 5732
rect 7220 5692 7756 5732
rect 7796 5692 8044 5732
rect 8084 5692 8093 5732
rect 10435 5692 10444 5732
rect 10484 5692 13228 5732
rect 13268 5692 13277 5732
rect 16099 5692 16108 5732
rect 16148 5692 18892 5732
rect 18932 5692 20180 5732
rect 21571 5692 21580 5732
rect 21620 5692 44908 5732
rect 44948 5692 44957 5732
rect 4675 5608 4684 5648
rect 4724 5608 5452 5648
rect 5492 5608 7084 5648
rect 7124 5608 7133 5648
rect 10147 5608 10156 5648
rect 10196 5608 11020 5648
rect 11060 5608 11069 5648
rect 14179 5608 14188 5648
rect 14228 5608 44524 5648
rect 44564 5608 44573 5648
rect 17155 5524 17164 5564
rect 17204 5524 28588 5564
rect 28628 5524 28637 5564
rect 30307 5524 30316 5564
rect 30356 5524 31028 5564
rect 33667 5524 33676 5564
rect 33716 5524 35980 5564
rect 36020 5524 36029 5564
rect 30988 5480 31028 5524
rect 5443 5440 5452 5480
rect 5492 5440 7180 5480
rect 7220 5440 7229 5480
rect 15139 5440 15148 5480
rect 15188 5440 20180 5480
rect 20803 5440 20812 5480
rect 20852 5440 23788 5480
rect 23828 5440 23837 5480
rect 26755 5440 26764 5480
rect 26804 5440 28396 5480
rect 28436 5440 28445 5480
rect 28867 5440 28876 5480
rect 28916 5440 30508 5480
rect 30548 5440 30557 5480
rect 30988 5440 39148 5480
rect 39188 5440 39197 5480
rect 10723 5356 10732 5396
rect 10772 5356 17644 5396
rect 17684 5356 17693 5396
rect 18700 5356 20084 5396
rect 18700 5312 18740 5356
rect 20044 5312 20084 5356
rect 20140 5312 20180 5440
rect 20227 5356 20236 5396
rect 20276 5356 22348 5396
rect 22388 5356 22397 5396
rect 25507 5356 25516 5396
rect 25556 5356 30412 5396
rect 30452 5356 30461 5396
rect 33187 5356 33196 5396
rect 33236 5356 33388 5396
rect 33428 5356 33437 5396
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 6211 5272 6220 5312
rect 6260 5272 9964 5312
rect 10004 5272 10013 5312
rect 14947 5272 14956 5312
rect 14996 5272 15724 5312
rect 15764 5272 15773 5312
rect 17059 5272 17068 5312
rect 17108 5272 18740 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 19277 5272 19372 5312
rect 19412 5272 19421 5312
rect 20035 5272 20044 5312
rect 20084 5272 20093 5312
rect 20140 5272 20812 5312
rect 20852 5272 20861 5312
rect 20995 5272 21004 5312
rect 21044 5272 24172 5312
rect 24212 5272 24221 5312
rect 25123 5272 25132 5312
rect 25172 5272 33140 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 33100 5228 33140 5272
rect 5539 5188 5548 5228
rect 5588 5188 7372 5228
rect 7412 5188 7421 5228
rect 12067 5188 12076 5228
rect 12116 5188 26476 5228
rect 26516 5188 26525 5228
rect 26947 5188 26956 5228
rect 26996 5188 28684 5228
rect 28724 5188 30260 5228
rect 33100 5188 36940 5228
rect 36980 5188 36989 5228
rect 30220 5144 30260 5188
rect 4579 5104 4588 5144
rect 4628 5104 7180 5144
rect 7220 5104 7229 5144
rect 15907 5104 15916 5144
rect 15956 5104 24940 5144
rect 24980 5104 24989 5144
rect 26179 5104 26188 5144
rect 26228 5104 28780 5144
rect 28820 5104 28829 5144
rect 30220 5104 34252 5144
rect 34292 5104 38956 5144
rect 38996 5104 39005 5144
rect 8035 5020 8044 5060
rect 8084 5020 10444 5060
rect 10484 5020 10493 5060
rect 16963 5020 16972 5060
rect 17012 5020 37900 5060
rect 37940 5020 37949 5060
rect 4195 4936 4204 4976
rect 4244 4936 6124 4976
rect 6164 4936 6604 4976
rect 6644 4936 6988 4976
rect 7028 4936 7037 4976
rect 8899 4936 8908 4976
rect 8948 4936 32428 4976
rect 32468 4936 32477 4976
rect 3715 4852 3724 4892
rect 3764 4852 4684 4892
rect 4724 4852 4733 4892
rect 9763 4852 9772 4892
rect 9812 4852 12788 4892
rect 12835 4852 12844 4892
rect 12884 4852 13268 4892
rect 14755 4852 14764 4892
rect 14804 4852 14860 4892
rect 14900 4852 14909 4892
rect 17635 4852 17644 4892
rect 17684 4852 23060 4892
rect 25699 4852 25708 4892
rect 25748 4852 28876 4892
rect 28916 4852 31276 4892
rect 31316 4852 31325 4892
rect 31843 4852 31852 4892
rect 31892 4852 32716 4892
rect 32756 4852 35980 4892
rect 36020 4852 36029 4892
rect 12748 4808 12788 4852
rect 13228 4808 13268 4852
rect 23020 4808 23060 4852
rect 4771 4768 4780 4808
rect 4820 4768 8524 4808
rect 8564 4768 8573 4808
rect 10243 4768 10252 4808
rect 10292 4768 12652 4808
rect 12692 4768 12701 4808
rect 12748 4768 13036 4808
rect 13076 4768 13085 4808
rect 13228 4768 21388 4808
rect 21428 4768 21437 4808
rect 23020 4768 38572 4808
rect 38612 4768 38621 4808
rect 2851 4684 2860 4724
rect 2900 4684 44044 4724
rect 44084 4684 44093 4724
rect 10627 4600 10636 4640
rect 10676 4600 12748 4640
rect 12788 4600 12797 4640
rect 14563 4600 14572 4640
rect 14612 4600 19604 4640
rect 19651 4600 19660 4640
rect 19700 4600 20716 4640
rect 20756 4600 20765 4640
rect 21859 4600 21868 4640
rect 21908 4600 26956 4640
rect 26996 4600 27005 4640
rect 33091 4600 33100 4640
rect 33140 4600 38092 4640
rect 38132 4600 38141 4640
rect 19564 4556 19604 4600
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 12451 4516 12460 4556
rect 12500 4516 14284 4556
rect 14324 4516 14333 4556
rect 16579 4516 16588 4556
rect 16628 4516 19508 4556
rect 19564 4516 19948 4556
rect 19988 4516 19997 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 21955 4516 21964 4556
rect 22004 4516 29740 4556
rect 29780 4516 29789 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 19468 4472 19508 4516
rect 7171 4432 7180 4472
rect 7220 4432 19372 4472
rect 19412 4432 19421 4472
rect 19468 4432 23884 4472
rect 23924 4432 23933 4472
rect 25507 4432 25516 4472
rect 25556 4432 28684 4472
rect 28724 4432 28733 4472
rect 30499 4432 30508 4472
rect 30548 4432 39532 4472
rect 39572 4432 39581 4472
rect 16099 4348 16108 4388
rect 16148 4348 28396 4388
rect 28436 4348 34252 4388
rect 34292 4348 34732 4388
rect 34772 4348 34781 4388
rect 5635 4264 5644 4304
rect 5684 4264 7660 4304
rect 7700 4264 7709 4304
rect 10243 4264 10252 4304
rect 10292 4264 10828 4304
rect 10868 4264 13708 4304
rect 13748 4264 13757 4304
rect 14467 4264 14476 4304
rect 14516 4264 14611 4304
rect 14851 4264 14860 4304
rect 14900 4264 16492 4304
rect 16532 4264 16541 4304
rect 16675 4264 16684 4304
rect 16724 4264 19180 4304
rect 19220 4264 19229 4304
rect 19565 4264 19660 4304
rect 19700 4264 19709 4304
rect 19843 4264 19852 4304
rect 19892 4264 20140 4304
rect 20180 4264 20189 4304
rect 20611 4264 20620 4304
rect 20660 4264 24556 4304
rect 24596 4264 24605 4304
rect 24835 4264 24844 4304
rect 24884 4264 27340 4304
rect 27380 4264 27389 4304
rect 28780 4264 32716 4304
rect 32756 4264 32765 4304
rect 28780 4220 28820 4264
rect 6787 4180 6796 4220
rect 6836 4180 11212 4220
rect 11252 4180 15820 4220
rect 15860 4180 15869 4220
rect 18595 4180 18604 4220
rect 18644 4180 18700 4220
rect 18740 4180 18749 4220
rect 19555 4180 19564 4220
rect 19604 4180 21196 4220
rect 21236 4180 22156 4220
rect 22196 4180 22205 4220
rect 28771 4180 28780 4220
rect 28820 4180 28829 4220
rect 32035 4180 32044 4220
rect 32084 4180 33772 4220
rect 33812 4180 33821 4220
rect 34349 4180 34444 4220
rect 34484 4180 34493 4220
rect 1411 4096 1420 4136
rect 1460 4096 37900 4136
rect 37940 4096 38860 4136
rect 38900 4096 38909 4136
rect 6307 4012 6316 4052
rect 6356 4012 6988 4052
rect 7028 4012 7037 4052
rect 12931 4012 12940 4052
rect 12980 4012 14380 4052
rect 14420 4012 14429 4052
rect 14861 4012 14956 4052
rect 14996 4012 15005 4052
rect 17923 4012 17932 4052
rect 17972 4012 20620 4052
rect 20660 4012 20669 4052
rect 20803 4012 20812 4052
rect 20852 4012 25228 4052
rect 25268 4012 25277 4052
rect 33379 4012 33388 4052
rect 33428 4012 36556 4052
rect 36596 4012 36605 4052
rect 5731 3928 5740 3968
rect 5780 3928 33140 3968
rect 33283 3928 33292 3968
rect 33332 3928 35788 3968
rect 35828 3928 35837 3968
rect 33100 3884 33140 3928
rect 2371 3844 2380 3884
rect 2420 3844 30700 3884
rect 30740 3844 30749 3884
rect 32323 3844 32332 3884
rect 32372 3844 32716 3884
rect 32756 3844 32765 3884
rect 33100 3844 40492 3884
rect 40532 3844 40972 3884
rect 41012 3844 41021 3884
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 5155 3760 5164 3800
rect 5204 3760 10252 3800
rect 10292 3760 10301 3800
rect 10819 3760 10828 3800
rect 10868 3760 12076 3800
rect 12116 3760 12125 3800
rect 14371 3760 14380 3800
rect 14420 3760 15628 3800
rect 15668 3760 16108 3800
rect 16148 3760 16157 3800
rect 18499 3760 18508 3800
rect 18548 3760 18700 3800
rect 18740 3760 18749 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 19267 3760 19276 3800
rect 19316 3760 21676 3800
rect 21716 3760 21725 3800
rect 25795 3760 25804 3800
rect 25844 3760 31852 3800
rect 31892 3760 31901 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 1987 3676 1996 3716
rect 2036 3676 2380 3716
rect 2420 3676 2429 3716
rect 3523 3676 3532 3716
rect 3572 3676 26956 3716
rect 26996 3676 27005 3716
rect 30499 3676 30508 3716
rect 30548 3676 35116 3716
rect 35156 3676 35165 3716
rect 2275 3592 2284 3632
rect 2324 3592 21868 3632
rect 21908 3592 21917 3632
rect 22051 3592 22060 3632
rect 22100 3592 23020 3632
rect 23060 3592 23069 3632
rect 24451 3592 24460 3632
rect 24500 3592 29164 3632
rect 29204 3592 29213 3632
rect 30307 3592 30316 3632
rect 30356 3592 33196 3632
rect 33236 3592 37612 3632
rect 37652 3592 37661 3632
rect 6499 3508 6508 3548
rect 6548 3508 7372 3548
rect 7412 3508 7421 3548
rect 10435 3508 10444 3548
rect 10484 3508 10732 3548
rect 10772 3508 12556 3548
rect 12596 3508 12605 3548
rect 13123 3508 13132 3548
rect 13172 3508 13612 3548
rect 13652 3508 13661 3548
rect 14380 3508 24844 3548
rect 24884 3508 30412 3548
rect 30452 3508 32140 3548
rect 32180 3508 32189 3548
rect 32323 3508 32332 3548
rect 32372 3508 39628 3548
rect 39668 3508 39677 3548
rect 14380 3464 14420 3508
rect 10531 3424 10540 3464
rect 10580 3424 13900 3464
rect 13940 3424 14420 3464
rect 18499 3424 18508 3464
rect 18548 3424 40300 3464
rect 40340 3424 40349 3464
rect 5539 3340 5548 3380
rect 5588 3340 6028 3380
rect 6068 3340 6077 3380
rect 8803 3340 8812 3380
rect 8852 3340 12268 3380
rect 12308 3340 12317 3380
rect 13603 3340 13612 3380
rect 13652 3340 13996 3380
rect 14036 3340 14045 3380
rect 16963 3340 16972 3380
rect 17012 3340 44716 3380
rect 44756 3340 44765 3380
rect 8611 3256 8620 3296
rect 8660 3256 44332 3296
rect 44372 3256 44381 3296
rect 7459 3172 7468 3212
rect 7508 3172 9388 3212
rect 9428 3172 9437 3212
rect 14467 3172 14476 3212
rect 14516 3172 15148 3212
rect 15188 3172 15197 3212
rect 17539 3172 17548 3212
rect 17588 3172 18412 3212
rect 18452 3172 18461 3212
rect 19075 3172 19084 3212
rect 19124 3172 19372 3212
rect 19412 3172 19421 3212
rect 19747 3172 19756 3212
rect 19796 3172 20908 3212
rect 20948 3172 20957 3212
rect 21475 3172 21484 3212
rect 21524 3172 22924 3212
rect 22964 3172 22973 3212
rect 24451 3172 24460 3212
rect 24500 3172 25612 3212
rect 25652 3172 25661 3212
rect 32707 3172 32716 3212
rect 32756 3172 36460 3212
rect 36500 3172 36509 3212
rect 2947 3088 2956 3128
rect 2996 3088 28204 3128
rect 28244 3088 28253 3128
rect 31267 3088 31276 3128
rect 31316 3088 31660 3128
rect 31700 3088 31709 3128
rect 33484 3088 42028 3128
rect 42068 3088 42077 3128
rect 33484 3044 33524 3088
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 6211 3004 6220 3044
rect 6260 3004 6892 3044
rect 6932 3004 6941 3044
rect 13507 3004 13516 3044
rect 13556 3004 13804 3044
rect 13844 3004 13853 3044
rect 14563 3004 14572 3044
rect 14612 3004 14956 3044
rect 14996 3004 15005 3044
rect 17347 3004 17356 3044
rect 17396 3004 19948 3044
rect 19988 3004 19997 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 21100 3004 23116 3044
rect 23156 3004 23165 3044
rect 30691 3004 30700 3044
rect 30740 3004 32908 3044
rect 32948 3004 32957 3044
rect 33475 3004 33484 3044
rect 33524 3004 33533 3044
rect 34349 3004 34444 3044
rect 34484 3004 34493 3044
rect 34627 3004 34636 3044
rect 34676 3004 34771 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 21100 2960 21140 3004
rect 5731 2920 5740 2960
rect 5780 2920 7084 2960
rect 7124 2920 7133 2960
rect 13891 2920 13900 2960
rect 13940 2920 16972 2960
rect 17012 2920 17021 2960
rect 18125 2920 18220 2960
rect 18260 2920 18269 2960
rect 18499 2920 18508 2960
rect 18548 2920 19276 2960
rect 19316 2920 19325 2960
rect 19747 2920 19756 2960
rect 19796 2920 21140 2960
rect 21667 2920 21676 2960
rect 21716 2920 37420 2960
rect 37460 2920 37469 2960
rect 6211 2836 6220 2876
rect 6260 2836 12748 2876
rect 12788 2836 12797 2876
rect 12931 2836 12940 2876
rect 12980 2836 17684 2876
rect 17731 2836 17740 2876
rect 17780 2836 18796 2876
rect 18836 2836 18845 2876
rect 19075 2836 19084 2876
rect 19124 2836 20044 2876
rect 20084 2836 20093 2876
rect 23107 2836 23116 2876
rect 23156 2836 29836 2876
rect 29876 2836 29885 2876
rect 31181 2836 31276 2876
rect 31316 2836 31325 2876
rect 33389 2836 33484 2876
rect 33524 2836 33533 2876
rect 33955 2836 33964 2876
rect 34004 2836 34924 2876
rect 34964 2836 34973 2876
rect 17644 2792 17684 2836
rect 1699 2752 1708 2792
rect 1748 2752 2476 2792
rect 2516 2752 7372 2792
rect 7412 2752 7421 2792
rect 9475 2752 9484 2792
rect 9524 2752 10156 2792
rect 10196 2752 10205 2792
rect 13411 2752 13420 2792
rect 13460 2752 16588 2792
rect 16628 2752 16637 2792
rect 17453 2752 17548 2792
rect 17588 2752 17597 2792
rect 17644 2752 21964 2792
rect 22004 2752 22013 2792
rect 22339 2752 22348 2792
rect 22388 2752 22732 2792
rect 22772 2752 22781 2792
rect 22915 2752 22924 2792
rect 22964 2752 23212 2792
rect 23252 2752 23261 2792
rect 24163 2752 24172 2792
rect 24212 2752 28588 2792
rect 28628 2752 28637 2792
rect 29635 2752 29644 2792
rect 29684 2752 32620 2792
rect 32660 2752 32669 2792
rect 4387 2668 4396 2708
rect 4436 2668 10924 2708
rect 10964 2668 10973 2708
rect 12259 2668 12268 2708
rect 12308 2668 18028 2708
rect 18068 2668 18077 2708
rect 18124 2668 23020 2708
rect 23060 2668 23069 2708
rect 24461 2668 24556 2708
rect 24596 2668 24605 2708
rect 28771 2668 28780 2708
rect 28820 2668 30700 2708
rect 30740 2668 30749 2708
rect 33187 2668 33196 2708
rect 33236 2668 33868 2708
rect 33908 2668 36076 2708
rect 36116 2668 36125 2708
rect 18124 2624 18164 2668
rect 3235 2584 3244 2624
rect 3284 2584 11404 2624
rect 11444 2584 11453 2624
rect 11971 2584 11980 2624
rect 12020 2584 17452 2624
rect 17492 2584 17501 2624
rect 17731 2584 17740 2624
rect 17780 2584 18164 2624
rect 18211 2584 18220 2624
rect 18260 2584 24844 2624
rect 24884 2584 24893 2624
rect 30499 2584 30508 2624
rect 30548 2584 34540 2624
rect 34580 2584 34589 2624
rect 1507 2500 1516 2540
rect 1556 2500 25132 2540
rect 25172 2500 25181 2540
rect 30211 2500 30220 2540
rect 30260 2500 33292 2540
rect 33332 2500 33341 2540
rect 33955 2500 33964 2540
rect 34004 2500 35116 2540
rect 35156 2500 35165 2540
rect 5731 2416 5740 2456
rect 5780 2416 22828 2456
rect 22868 2416 22877 2456
rect 23011 2416 23020 2456
rect 23060 2416 44140 2456
rect 44180 2416 44189 2456
rect 3139 2332 3148 2372
rect 3188 2332 6700 2372
rect 6740 2332 6749 2372
rect 10060 2332 16972 2372
rect 17012 2332 17021 2372
rect 18595 2332 18604 2372
rect 18644 2332 21676 2372
rect 21716 2332 22636 2372
rect 22676 2332 22685 2372
rect 31651 2332 31660 2372
rect 31700 2332 32332 2372
rect 32372 2332 32381 2372
rect 33379 2332 33388 2372
rect 33428 2332 33484 2372
rect 33524 2332 33533 2372
rect 33580 2332 38668 2372
rect 38708 2332 38717 2372
rect 10060 2288 10100 2332
rect 33580 2288 33620 2332
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 7363 2248 7372 2288
rect 7412 2248 10100 2288
rect 12931 2248 12940 2288
rect 12980 2248 13708 2288
rect 13748 2248 13757 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 20515 2248 20524 2288
rect 20564 2248 22444 2288
rect 22484 2248 22493 2288
rect 30211 2248 30220 2288
rect 30260 2248 33620 2288
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 4291 2164 4300 2204
rect 4340 2164 7276 2204
rect 7316 2164 7325 2204
rect 13027 2164 13036 2204
rect 13076 2164 13228 2204
rect 13268 2164 13277 2204
rect 18019 2164 18028 2204
rect 18068 2164 22964 2204
rect 22924 2120 22964 2164
rect 4003 2080 4012 2120
rect 4052 2080 4780 2120
rect 4820 2080 4829 2120
rect 6019 2080 6028 2120
rect 6068 2080 7180 2120
rect 7220 2080 7229 2120
rect 12835 2080 12844 2120
rect 12884 2080 18412 2120
rect 18452 2080 18461 2120
rect 22924 2080 23308 2120
rect 23348 2080 29260 2120
rect 29300 2080 29309 2120
rect 3523 1996 3532 2036
rect 3572 1996 9004 2036
rect 9044 1996 9964 2036
rect 10004 1996 10013 2036
rect 12739 1996 12748 2036
rect 12788 1996 13420 2036
rect 13460 1996 13469 2036
rect 16963 1996 16972 2036
rect 17012 1996 19276 2036
rect 19316 1996 19325 2036
rect 28963 1996 28972 2036
rect 29012 1996 29164 2036
rect 29204 1996 29213 2036
rect 4099 1912 4108 1952
rect 4148 1912 4780 1952
rect 4820 1912 4829 1952
rect 11299 1912 11308 1952
rect 11348 1912 15820 1952
rect 15860 1912 15869 1952
rect 18211 1912 18220 1952
rect 18260 1912 19372 1952
rect 19412 1912 19421 1952
rect 4291 1828 4300 1868
rect 4340 1828 18604 1868
rect 18644 1828 18653 1868
rect 21571 1828 21580 1868
rect 21620 1828 27724 1868
rect 27764 1828 27773 1868
rect 32035 1828 32044 1868
rect 32084 1828 33196 1868
rect 33236 1828 33245 1868
rect 14947 1744 14956 1784
rect 14996 1744 17548 1784
rect 17588 1744 17597 1784
rect 18019 1744 18028 1784
rect 18068 1744 20812 1784
rect 20852 1744 20861 1784
rect 4483 1660 4492 1700
rect 4532 1660 8044 1700
rect 8084 1660 8093 1700
rect 8611 1660 8620 1700
rect 8660 1660 31468 1700
rect 31508 1660 31517 1700
rect 10339 1576 10348 1616
rect 10388 1576 13900 1616
rect 13940 1576 13949 1616
rect 14851 1576 14860 1616
rect 14900 1576 15436 1616
rect 15476 1576 15485 1616
rect 20707 1576 20716 1616
rect 20756 1576 24940 1616
rect 24980 1576 24989 1616
rect 25795 1576 25804 1616
rect 25844 1576 29548 1616
rect 29588 1576 29597 1616
rect 33283 1576 33292 1616
rect 33332 1576 37324 1616
rect 37364 1576 37373 1616
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 11779 1492 11788 1532
rect 11828 1492 18604 1532
rect 18644 1492 18653 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 14765 1408 14860 1448
rect 14900 1408 14909 1448
rect 16483 1408 16492 1448
rect 16532 1408 16972 1448
rect 17012 1408 17021 1448
rect 30595 1408 30604 1448
rect 30644 1408 30892 1448
rect 30932 1408 30941 1448
rect 32323 1408 32332 1448
rect 32372 1408 32812 1448
rect 32852 1408 32861 1448
rect 12931 1324 12940 1364
rect 12980 1324 17740 1364
rect 17780 1324 17789 1364
rect 18499 1324 18508 1364
rect 18548 1324 21580 1364
rect 21620 1324 21629 1364
rect 31555 1324 31564 1364
rect 31604 1324 36748 1364
rect 36788 1324 36797 1364
rect 13123 1240 13132 1280
rect 13172 1240 13324 1280
rect 13364 1240 13373 1280
rect 14563 1240 14572 1280
rect 14612 1240 18316 1280
rect 18356 1240 18365 1280
rect 29827 1240 29836 1280
rect 29876 1240 31756 1280
rect 31796 1240 31805 1280
rect 14467 1072 14476 1112
rect 14516 1072 19276 1112
rect 19316 1072 19325 1112
rect 7363 988 7372 1028
rect 7412 988 15052 1028
rect 15092 988 15101 1028
rect 15715 988 15724 1028
rect 15764 988 20044 1028
rect 20084 988 20093 1028
rect 30403 904 30412 944
rect 30452 904 36172 944
rect 36212 904 36221 944
rect 26947 820 26956 860
rect 26996 820 32428 860
rect 32468 820 32477 860
rect 26563 652 26572 692
rect 26612 652 31660 692
rect 31700 652 31709 692
rect 14755 568 14764 608
rect 14804 568 19084 608
rect 19124 568 19133 608
rect 12931 400 12940 440
rect 12980 400 13228 440
rect 13268 400 13277 440
rect 29635 400 29644 440
rect 29684 400 32236 440
rect 32276 400 32285 440
rect 7171 232 7180 272
rect 7220 232 14476 272
rect 14516 232 14525 272
rect 2851 64 2860 104
rect 2900 64 11596 104
rect 11636 64 11645 104
<< via4 >>
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 14572 9388 14612 9428
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 33196 8548 33236 8588
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 15628 7960 15668 8000
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 14572 6784 14612 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 19564 6784 19604 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 34636 6364 34676 6404
rect 19564 6280 19604 6320
rect 32140 6196 32180 6236
rect 19852 6112 19892 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 20812 5944 20852 5984
rect 19756 5776 19796 5816
rect 20812 5776 20852 5816
rect 24556 5776 24596 5816
rect 20812 5440 20852 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 19372 5272 19412 5312
rect 20812 5272 20852 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 14860 4852 14900 4892
rect 19660 4600 19700 4640
rect 21868 4600 21908 4640
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 14476 4264 14516 4304
rect 19660 4264 19700 4304
rect 19852 4264 19892 4304
rect 18604 4180 18644 4220
rect 34444 4180 34484 4220
rect 14956 4012 14996 4052
rect 33292 3928 33332 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 15628 3760 15668 3800
rect 18508 3760 18548 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 19276 3760 19316 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 21868 3592 21908 3632
rect 33196 3592 33236 3632
rect 32140 3508 32180 3548
rect 14476 3172 14516 3212
rect 17548 3172 17588 3212
rect 19756 3172 19796 3212
rect 31276 3088 31316 3128
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 14956 3004 14996 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 34444 3004 34484 3044
rect 34636 3004 34676 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 18220 2920 18260 2960
rect 19276 2920 19316 2960
rect 31276 2836 31316 2876
rect 33484 2836 33524 2876
rect 17548 2752 17588 2792
rect 24556 2668 24596 2708
rect 33196 2668 33236 2708
rect 18220 2584 18260 2624
rect 33292 2500 33332 2540
rect 22828 2416 22868 2456
rect 23020 2416 23060 2456
rect 18604 2332 18644 2372
rect 33484 2332 33524 2372
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 19372 1912 19412 1952
rect 18604 1828 18644 1868
rect 33196 1828 33236 1868
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 14860 1408 14900 1448
rect 18508 1324 18548 1364
<< metal5 >>
rect 3652 9848 4092 12180
rect 3652 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4092 9848
rect 3652 8336 4092 9808
rect 3652 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4092 8336
rect 3652 6824 4092 8296
rect 3652 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4092 6824
rect 3652 5312 4092 6784
rect 3652 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4092 5312
rect 3652 3800 4092 5272
rect 3652 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4092 3800
rect 3652 2288 4092 3760
rect 3652 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4092 2288
rect 3652 0 4092 2248
rect 4892 10604 5332 12180
rect 4892 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5332 10604
rect 4892 9092 5332 10564
rect 18772 9848 19212 12180
rect 18772 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19212 9848
rect 4892 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5332 9092
rect 4892 7580 5332 9052
rect 4892 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5332 7580
rect 4892 6068 5332 7540
rect 14572 9428 14612 9437
rect 14572 6824 14612 9388
rect 18772 8336 19212 9808
rect 18772 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19212 8336
rect 14572 6775 14612 6784
rect 15628 8000 15668 8009
rect 4892 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5332 6068
rect 4892 4556 5332 6028
rect 4892 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5332 4556
rect 4892 3044 5332 4516
rect 14860 4892 14900 4901
rect 14476 4304 14516 4313
rect 14476 3212 14516 4264
rect 14476 3163 14516 3172
rect 4892 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5332 3044
rect 4892 1532 5332 3004
rect 4892 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5332 1532
rect 4892 0 5332 1492
rect 14860 1448 14900 4852
rect 14956 4052 14996 4061
rect 14956 3044 14996 4012
rect 15628 3800 15668 7960
rect 18772 6824 19212 8296
rect 20012 10604 20452 12180
rect 20012 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20452 10604
rect 20012 9092 20452 10564
rect 20012 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20452 9092
rect 20012 7580 20452 9052
rect 33892 9848 34332 12180
rect 33892 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34332 9848
rect 20012 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20452 7580
rect 18772 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19212 6824
rect 18772 5312 19212 6784
rect 19564 6824 19604 6833
rect 19564 6320 19604 6784
rect 19564 6271 19604 6280
rect 19852 6152 19892 6161
rect 19756 5816 19796 5825
rect 18772 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19212 5312
rect 18604 4220 18644 4229
rect 15628 3751 15668 3760
rect 18508 3800 18548 3809
rect 14956 2995 14996 3004
rect 17548 3212 17588 3221
rect 17548 2792 17588 3172
rect 17548 2743 17588 2752
rect 18220 2960 18260 2969
rect 18220 2624 18260 2920
rect 18220 2575 18260 2584
rect 14860 1399 14900 1408
rect 18508 1364 18548 3760
rect 18604 2372 18644 4180
rect 18604 1868 18644 2332
rect 18604 1819 18644 1828
rect 18772 3800 19212 5272
rect 19372 5312 19412 5321
rect 18772 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19212 3800
rect 18772 2288 19212 3760
rect 19276 3800 19316 3809
rect 19276 2960 19316 3760
rect 19276 2911 19316 2920
rect 18772 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19212 2288
rect 18508 1315 18548 1324
rect 18772 0 19212 2248
rect 19372 1952 19412 5272
rect 19660 4640 19700 4649
rect 19660 4304 19700 4600
rect 19660 4255 19700 4264
rect 19756 3212 19796 5776
rect 19852 4304 19892 6112
rect 19852 4255 19892 4264
rect 20012 6068 20452 7540
rect 33196 8588 33236 8597
rect 20012 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20452 6068
rect 20012 4556 20452 6028
rect 32140 6236 32180 6245
rect 20812 5984 20852 5993
rect 20812 5816 20852 5944
rect 20812 5767 20852 5776
rect 24556 5816 24596 5825
rect 20812 5480 20852 5489
rect 20812 5312 20852 5440
rect 20812 5263 20852 5272
rect 20012 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20452 4556
rect 19756 3163 19796 3172
rect 19372 1903 19412 1912
rect 20012 3044 20452 4516
rect 21868 4640 21908 4649
rect 21868 3632 21908 4600
rect 21868 3583 21908 3592
rect 20012 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20452 3044
rect 20012 1532 20452 3004
rect 24556 2708 24596 5776
rect 32140 3548 32180 6196
rect 33196 3632 33236 8548
rect 33892 8336 34332 9808
rect 33892 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34332 8336
rect 33892 6824 34332 8296
rect 33892 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34332 6824
rect 33892 5312 34332 6784
rect 35132 10604 35572 12180
rect 35132 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 35572 10604
rect 35132 9092 35572 10564
rect 35132 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35572 9092
rect 35132 7580 35572 9052
rect 35132 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35572 7580
rect 33892 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34332 5312
rect 33196 3583 33236 3592
rect 33292 3968 33332 3977
rect 32140 3499 32180 3508
rect 31276 3128 31316 3137
rect 31276 2876 31316 3088
rect 31276 2827 31316 2836
rect 24556 2659 24596 2668
rect 33196 2708 33236 2717
rect 22828 2552 23060 2592
rect 22828 2456 22868 2552
rect 22828 2407 22868 2416
rect 23020 2456 23060 2552
rect 23020 2407 23060 2416
rect 33196 1868 33236 2668
rect 33292 2540 33332 3928
rect 33892 3800 34332 5272
rect 34636 6404 34676 6413
rect 33892 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34332 3800
rect 33292 2491 33332 2500
rect 33484 2876 33524 2885
rect 33484 2372 33524 2836
rect 33484 2323 33524 2332
rect 33196 1819 33236 1828
rect 33892 2288 34332 3760
rect 34444 4220 34484 4229
rect 34444 3044 34484 4180
rect 34444 2995 34484 3004
rect 34636 3044 34676 6364
rect 34636 2995 34676 3004
rect 35132 6068 35572 7540
rect 35132 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35572 6068
rect 35132 4556 35572 6028
rect 35132 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35572 4556
rect 35132 3044 35572 4516
rect 35132 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35572 3044
rect 33892 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34332 2288
rect 20012 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20452 1532
rect 20012 0 20452 1492
rect 33892 0 34332 2248
rect 35132 1532 35572 3004
rect 35132 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35572 1532
rect 35132 0 35572 1492
use sg13g2_mux4_1  _049_
timestamp 1677257233
transform 1 0 21504 0 1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _050_
timestamp 1677257233
transform 1 0 21312 0 -1 3024
box -48 -56 2064 834
use sg13g2_mux4_1  _051_
timestamp 1677257233
transform 1 0 21792 0 -1 7560
box -48 -56 2064 834
use sg13g2_mux4_1  _052_
timestamp 1677257233
transform 1 0 24768 0 1 1512
box -48 -56 2064 834
use sg13g2_mux4_1  _053_
timestamp 1677257233
transform 1 0 11328 0 1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _054_
timestamp 1677257233
transform 1 0 15072 0 -1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _055_
timestamp 1677257233
transform 1 0 18240 0 1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _056_
timestamp 1677257233
transform 1 0 31104 0 -1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _057_
timestamp 1677257233
transform 1 0 37824 0 1 7560
box -48 -56 2064 834
use sg13g2_mux4_1  _058_
timestamp 1677257233
transform 1 0 20640 0 -1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _059_
timestamp 1677257233
transform 1 0 19392 0 -1 7560
box -48 -56 2064 834
use sg13g2_mux4_1  _060_
timestamp 1677257233
transform 1 0 23904 0 -1 3024
box -48 -56 2064 834
use sg13g2_mux4_1  _061_
timestamp 1677257233
transform 1 0 10560 0 -1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _062_
timestamp 1677257233
transform 1 0 14688 0 1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _063_
timestamp 1677257233
transform 1 0 14880 0 1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _064_
timestamp 1677257233
transform 1 0 28128 0 1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _065_
timestamp 1677257233
transform 1 0 26784 0 1 7560
box -48 -56 2064 834
use sg13g2_mux4_1  _066_
timestamp 1677257233
transform 1 0 18240 0 -1 3024
box -48 -56 2064 834
use sg13g2_mux4_1  _067_
timestamp 1677257233
transform 1 0 17856 0 1 6048
box -48 -56 2064 834
use sg13g2_mux2_1  _068_
timestamp 1677247768
transform 1 0 35904 0 -1 6048
box -48 -56 1008 834
use sg13g2_mux2_1  _069_
timestamp 1677247768
transform 1 0 40608 0 1 3024
box -48 -56 1008 834
use sg13g2_mux2_1  _070_
timestamp 1677247768
transform 1 0 25728 0 1 7560
box -48 -56 1008 834
use sg13g2_mux2_1  _071_
timestamp 1677247768
transform 1 0 22272 0 1 4536
box -48 -56 1008 834
use sg13g2_nand2b_1  _072_
timestamp 1676567195
transform 1 0 6432 0 -1 7560
box -48 -56 528 834
use sg13g2_o21ai_1  _073_
timestamp 1685175443
transform -1 0 7968 0 1 7560
box -48 -56 538 834
use sg13g2_nand3_1  _074_
timestamp 1683988354
transform 1 0 7008 0 -1 10584
box -48 -56 528 834
use sg13g2_o21ai_1  _075_
timestamp 1685175443
transform -1 0 7488 0 -1 7560
box -48 -56 538 834
use sg13g2_nand3b_1  _076_
timestamp 1676573470
transform -1 0 8160 0 -1 9072
box -48 -56 720 834
use sg13g2_o21ai_1  _077_
timestamp 1685175443
transform -1 0 7968 0 1 9072
box -48 -56 538 834
use sg13g2_nand2_1  _078_
timestamp 1676557249
transform 1 0 6048 0 -1 7560
box -48 -56 432 834
use sg13g2_nand4_1  _079_
timestamp 1685201930
transform 1 0 6912 0 1 7560
box -48 -56 624 834
use sg13g2_o21ai_1  _080_
timestamp 1685175443
transform 1 0 7968 0 1 7560
box -48 -56 538 834
use sg13g2_nand2b_1  _081_
timestamp 1676567195
transform 1 0 6912 0 -1 4536
box -48 -56 528 834
use sg13g2_mux4_1  _082_
timestamp 1677257233
transform -1 0 7872 0 1 3024
box -48 -56 2064 834
use sg13g2_o21ai_1  _083_
timestamp 1685175443
transform -1 0 5856 0 1 3024
box -48 -56 538 834
use sg13g2_o21ai_1  _084_
timestamp 1685175443
transform -1 0 5376 0 1 3024
box -48 -56 538 834
use sg13g2_nand2b_1  _085_
timestamp 1676567195
transform 1 0 6816 0 -1 3024
box -48 -56 528 834
use sg13g2_o21ai_1  _086_
timestamp 1685175443
transform 1 0 6336 0 -1 3024
box -48 -56 538 834
use sg13g2_inv_1  _087_
timestamp 1676382929
transform -1 0 9120 0 1 7560
box -48 -56 336 834
use sg13g2_inv_1  _088_
timestamp 1676382929
transform 1 0 6720 0 -1 10584
box -48 -56 336 834
use sg13g2_mux2_1  _089_
timestamp 1677247768
transform 1 0 6624 0 1 6048
box -48 -56 1008 834
use sg13g2_or2_1  _090_
timestamp 1684236171
transform 1 0 7488 0 -1 7560
box -48 -56 528 834
use sg13g2_a21oi_1  _091_
timestamp 1683973020
transform 1 0 8352 0 1 6048
box -48 -56 528 834
use sg13g2_a221oi_1  _092_
timestamp 1685197497
transform -1 0 8352 0 1 6048
box -48 -56 816 834
use sg13g2_nand2_1  _093_
timestamp 1676557249
transform 1 0 3648 0 1 4536
box -48 -56 432 834
use sg13g2_nand2b_1  _094_
timestamp 1676567195
transform -1 0 6912 0 -1 4536
box -48 -56 528 834
use sg13g2_a21oi_1  _095_
timestamp 1683973020
transform 1 0 5952 0 -1 4536
box -48 -56 528 834
use sg13g2_nor2b_1  _096_
timestamp 1685181386
transform 1 0 4992 0 -1 4536
box -54 -56 528 834
use sg13g2_o21ai_1  _097_
timestamp 1685175443
transform -1 0 6144 0 1 4536
box -48 -56 538 834
use sg13g2_o21ai_1  _098_
timestamp 1685175443
transform 1 0 5472 0 -1 4536
box -48 -56 538 834
use sg13g2_o21ai_1  _099_
timestamp 1685175443
transform -1 0 5952 0 -1 6048
box -48 -56 538 834
use sg13g2_mux4_1  _100_
timestamp 1677257233
transform -1 0 8928 0 -1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _101_
timestamp 1677257233
transform -1 0 9504 0 1 4536
box -48 -56 2064 834
use sg13g2_mux2_1  _102_
timestamp 1677247768
transform -1 0 7488 0 1 4536
box -48 -56 1008 834
use sg13g2_nand2b_1  _103_
timestamp 1676567195
transform 1 0 6432 0 -1 6048
box -48 -56 528 834
use sg13g2_o21ai_1  _104_
timestamp 1685175443
transform 1 0 5952 0 -1 6048
box -48 -56 538 834
use sg13g2_mux2_1  _105_
timestamp 1677247768
transform 1 0 9312 0 -1 7560
box -48 -56 1008 834
use sg13g2_or2_1  _106_
timestamp 1684236171
transform 1 0 10176 0 1 7560
box -48 -56 528 834
use sg13g2_a21oi_1  _107_
timestamp 1683973020
transform -1 0 8832 0 -1 7560
box -48 -56 528 834
use sg13g2_a221oi_1  _108_
timestamp 1685197497
transform 1 0 10272 0 -1 7560
box -48 -56 816 834
use sg13g2_nand2_1  _109_
timestamp 1676557249
transform 1 0 10656 0 1 7560
box -48 -56 432 834
use sg13g2_nand2b_1  _110_
timestamp 1676567195
transform -1 0 10368 0 1 6048
box -48 -56 528 834
use sg13g2_a21oi_1  _111_
timestamp 1683973020
transform 1 0 9696 0 1 7560
box -48 -56 528 834
use sg13g2_nor2b_1  _112_
timestamp 1685181386
transform -1 0 9696 0 1 7560
box -54 -56 528 834
use sg13g2_o21ai_1  _113_
timestamp 1685175443
transform -1 0 9888 0 1 6048
box -48 -56 538 834
use sg13g2_o21ai_1  _114_
timestamp 1685175443
transform -1 0 9312 0 -1 7560
box -48 -56 538 834
use sg13g2_o21ai_1  _115_
timestamp 1685175443
transform 1 0 10368 0 1 6048
box -48 -56 538 834
use sg13g2_mux4_1  _116_
timestamp 1677257233
transform 1 0 9504 0 1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _117_
timestamp 1677257233
transform 1 0 9408 0 -1 4536
box -48 -56 2064 834
use sg13g2_mux2_1  _118_
timestamp 1677247768
transform 1 0 10560 0 -1 6048
box -48 -56 1008 834
use sg13g2_nand2b_1  _119_
timestamp 1676567195
transform 1 0 10848 0 1 6048
box -48 -56 528 834
use sg13g2_o21ai_1  _120_
timestamp 1685175443
transform 1 0 11040 0 -1 7560
box -48 -56 538 834
use sg13g2_mux4_1  _121_
timestamp 1677257233
transform 1 0 11616 0 1 3024
box -48 -56 2064 834
use sg13g2_mux4_1  _122_
timestamp 1677257233
transform 1 0 12480 0 1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _123_
timestamp 1677257233
transform 1 0 30144 0 1 7560
box -48 -56 2064 834
use sg13g2_mux4_1  _124_
timestamp 1677257233
transform 1 0 34368 0 1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _125_
timestamp 1677257233
transform 1 0 33888 0 -1 3024
box -48 -56 2064 834
use sg13g2_mux4_1  _126_
timestamp 1677257233
transform 1 0 30432 0 -1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _127_
timestamp 1677257233
transform 1 0 34176 0 -1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _128_
timestamp 1677257233
transform 1 0 33600 0 -1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _129_
timestamp 1677257233
transform -1 0 11616 0 1 3024
box -48 -56 2064 834
use sg13g2_mux4_1  _130_
timestamp 1677257233
transform 1 0 7392 0 -1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _131_
timestamp 1677257233
transform 1 0 4608 0 1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _132_
timestamp 1677257233
transform -1 0 6912 0 1 7560
box -48 -56 2064 834
use sg13g2_mux4_1  _133_
timestamp 1677257233
transform 1 0 29856 0 -1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _134_
timestamp 1677257233
transform 1 0 27168 0 1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _135_
timestamp 1677257233
transform 1 0 27936 0 -1 3024
box -48 -56 2064 834
use sg13g2_mux4_1  _136_
timestamp 1677257233
transform 1 0 25248 0 -1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _137_
timestamp 1677257233
transform 1 0 30048 0 -1 3024
box -48 -56 2064 834
use sg13g2_mux4_1  _138_
timestamp 1677257233
transform 1 0 24192 0 1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _139_
timestamp 1677257233
transform 1 0 33696 0 -1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _140_
timestamp 1677257233
transform 1 0 40128 0 -1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _141_
timestamp 1677257233
transform 1 0 34080 0 1 1512
box -48 -56 2064 834
use sg13g2_mux4_1  _142_
timestamp 1677257233
transform 1 0 31104 0 1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _143_
timestamp 1677257233
transform 1 0 37248 0 1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _144_
timestamp 1677257233
transform 1 0 40128 0 -1 7560
box -48 -56 2064 834
use sg13g2_mux4_1  _145_
timestamp 1677257233
transform 1 0 15456 0 -1 3024
box -48 -56 2064 834
use sg13g2_mux4_1  _146_
timestamp 1677257233
transform 1 0 17472 0 -1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _147_
timestamp 1677257233
transform 1 0 18432 0 -1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _148_
timestamp 1677257233
transform 1 0 17376 0 -1 7560
box -48 -56 2064 834
use sg13g2_mux4_1  _149_
timestamp 1677257233
transform 1 0 18528 0 1 4536
box -48 -56 2064 834
use sg13g2_dlhq_1  _150_
timestamp 1678805552
transform -1 0 38496 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _151_
timestamp 1678805552
transform -1 0 39648 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _152_
timestamp 1678805552
transform -1 0 40320 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _153_
timestamp 1678805552
transform -1 0 40608 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _154_
timestamp 1678805552
transform -1 0 42144 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _155_
timestamp 1678805552
transform -1 0 40512 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _156_
timestamp 1678805552
transform 1 0 13632 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _157_
timestamp 1678805552
transform -1 0 34848 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _158_
timestamp 1678805552
transform 1 0 20640 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _159_
timestamp 1678805552
transform 1 0 24096 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _160_
timestamp 1678805552
transform 1 0 38592 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _161_
timestamp 1678805552
transform 1 0 35520 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _162_
timestamp 1678805552
transform 1 0 16608 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _163_
timestamp 1678805552
transform -1 0 25632 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _164_
timestamp 1678805552
transform 1 0 16896 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _165_
timestamp 1678805552
transform 1 0 18528 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _166_
timestamp 1678805552
transform 1 0 25152 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _167_
timestamp 1678805552
transform 1 0 26976 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _168_
timestamp 1678805552
transform 1 0 26592 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _169_
timestamp 1678805552
transform 1 0 28512 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _170_
timestamp 1678805552
transform 1 0 13440 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _171_
timestamp 1678805552
transform 1 0 14208 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _172_
timestamp 1678805552
transform 1 0 13152 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _173_
timestamp 1678805552
transform 1 0 14784 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _174_
timestamp 1678805552
transform 1 0 9216 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _175_
timestamp 1678805552
transform 1 0 9600 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _176_
timestamp 1678805552
transform 1 0 13824 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _177_
timestamp 1678805552
transform 1 0 21984 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _178_
timestamp 1678805552
transform -1 0 28704 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _179_
timestamp 1678805552
transform -1 0 28320 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _180_
timestamp 1678805552
transform -1 0 28512 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _181_
timestamp 1678805552
transform -1 0 25344 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _182_
timestamp 1678805552
transform 1 0 36672 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _183_
timestamp 1678805552
transform 1 0 38304 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _184_
timestamp 1678805552
transform -1 0 38688 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _185_
timestamp 1678805552
transform 1 0 30624 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _186_
timestamp 1678805552
transform 1 0 15840 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _187_
timestamp 1678805552
transform -1 0 21600 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _188_
timestamp 1678805552
transform 1 0 13344 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _189_
timestamp 1678805552
transform -1 0 23520 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _190_
timestamp 1678805552
transform -1 0 14208 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _191_
timestamp 1678805552
transform 1 0 11808 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _192_
timestamp 1678805552
transform 1 0 23136 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _193_
timestamp 1678805552
transform 1 0 24768 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _194_
timestamp 1678805552
transform 1 0 20640 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _195_
timestamp 1678805552
transform 1 0 22176 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _196_
timestamp 1678805552
transform 1 0 20352 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _197_
timestamp 1678805552
transform 1 0 21504 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _198_
timestamp 1678805552
transform 1 0 21792 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _199_
timestamp 1678805552
transform 1 0 20160 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _200_
timestamp 1678805552
transform 1 0 18816 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _201_
timestamp 1678805552
transform 1 0 17088 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _202_
timestamp 1678805552
transform 1 0 14976 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _203_
timestamp 1678805552
transform 1 0 15456 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _204_
timestamp 1678805552
transform 1 0 16896 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _205_
timestamp 1678805552
transform 1 0 16512 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _206_
timestamp 1678805552
transform 1 0 15072 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _207_
timestamp 1678805552
transform 1 0 17472 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _208_
timestamp 1678805552
transform 1 0 13728 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _209_
timestamp 1678805552
transform 1 0 15360 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _210_
timestamp 1678805552
transform 1 0 38880 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _211_
timestamp 1678805552
transform 1 0 40032 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _212_
timestamp 1678805552
transform 1 0 36384 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _213_
timestamp 1678805552
transform 1 0 36864 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _214_
timestamp 1678805552
transform 1 0 31872 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _215_
timestamp 1678805552
transform 1 0 30240 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _216_
timestamp 1678805552
transform -1 0 38016 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _217_
timestamp 1678805552
transform 1 0 32256 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _218_
timestamp 1678805552
transform 1 0 40320 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _219_
timestamp 1678805552
transform 1 0 38688 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _220_
timestamp 1678805552
transform 1 0 33888 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _221_
timestamp 1678805552
transform 1 0 32544 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _222_
timestamp 1678805552
transform 1 0 22752 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _223_
timestamp 1678805552
transform 1 0 24096 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _224_
timestamp 1678805552
transform 1 0 28992 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _225_
timestamp 1678805552
transform 1 0 30528 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _226_
timestamp 1678805552
transform 1 0 23520 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _227_
timestamp 1678805552
transform 1 0 25440 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _228_
timestamp 1678805552
transform 1 0 26304 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _229_
timestamp 1678805552
transform 1 0 27648 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _230_
timestamp 1678805552
transform 1 0 25728 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _231_
timestamp 1678805552
transform -1 0 30816 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _232_
timestamp 1678805552
transform 1 0 28224 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _233_
timestamp 1678805552
transform 1 0 30144 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _234_
timestamp 1678805552
transform 1 0 2688 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _235_
timestamp 1678805552
transform 1 0 2112 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _236_
timestamp 1678805552
transform 1 0 2208 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _237_
timestamp 1678805552
transform 1 0 4896 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _238_
timestamp 1678805552
transform 1 0 8160 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _239_
timestamp 1678805552
transform 1 0 2976 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _240_
timestamp 1678805552
transform -1 0 12192 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _241_
timestamp 1678805552
transform 1 0 8928 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _242_
timestamp 1678805552
transform 1 0 34272 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _243_
timestamp 1678805552
transform 1 0 32256 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _244_
timestamp 1678805552
transform 1 0 32928 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _245_
timestamp 1678805552
transform 1 0 34752 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _246_
timestamp 1678805552
transform -1 0 32256 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _247_
timestamp 1678805552
transform -1 0 33888 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _248_
timestamp 1678805552
transform -1 0 38016 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _249_
timestamp 1678805552
transform 1 0 34176 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _250_
timestamp 1678805552
transform 1 0 33024 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _251_
timestamp 1678805552
transform 1 0 35136 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _252_
timestamp 1678805552
transform 1 0 28704 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _253_
timestamp 1678805552
transform 1 0 30432 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _254_
timestamp 1678805552
transform 1 0 13248 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _255_
timestamp 1678805552
transform 1 0 11520 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _256_
timestamp 1678805552
transform 1 0 12192 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _257_
timestamp 1678805552
transform 1 0 10560 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _258_
timestamp 1678805552
transform -1 0 13248 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _259_
timestamp 1678805552
transform -1 0 13152 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _260_
timestamp 1678805552
transform 1 0 7296 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _261_
timestamp 1678805552
transform 1 0 8448 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _262_
timestamp 1678805552
transform 1 0 5856 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _263_
timestamp 1678805552
transform 1 0 5856 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _264_
timestamp 1678805552
transform 1 0 4224 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _265_
timestamp 1678805552
transform 1 0 3840 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _266_
timestamp 1678805552
transform 1 0 2592 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _267_
timestamp 1678805552
transform 1 0 3744 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _268_
timestamp 1678805552
transform 1 0 4032 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _269_
timestamp 1678805552
transform 1 0 4704 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _270_
timestamp 1678805552
transform 1 0 4224 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _271_
timestamp 1678805552
transform 1 0 3168 0 1 3024
box -50 -56 1692 834
use sg13g2_tiehi  _272__205
timestamp 1680000651
transform -1 0 40992 0 1 6048
box -48 -56 432 834
use sg13g2_dfrbp_1  _272_
timestamp 1678705109
transform 1 0 39648 0 -1 6048
box -60 -56 2556 834
use sg13g2_dfrbp_1  _273_
timestamp 1678705109
transform 1 0 39840 0 1 4536
box -60 -56 2556 834
use sg13g2_tiehi  _273__206
timestamp 1680000651
transform -1 0 41280 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _276_
timestamp 1676381911
transform 1 0 4320 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _277_
timestamp 1676381911
transform 1 0 18816 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _278_
timestamp 1676381911
transform 1 0 38880 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _279_
timestamp 1676381911
transform 1 0 39648 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _280_
timestamp 1676381911
transform 1 0 36288 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _281_
timestamp 1676381911
transform 1 0 36384 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _282_
timestamp 1676381911
transform 1 0 36480 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _283_
timestamp 1676381911
transform 1 0 38304 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _284_
timestamp 1676381911
transform 1 0 38784 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _285_
timestamp 1676381911
transform 1 0 40608 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _286_
timestamp 1676381911
transform 1 0 41952 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _287_
timestamp 1676381911
transform 1 0 29472 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _288_
timestamp 1676381911
transform 1 0 34848 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _289_
timestamp 1676381911
transform 1 0 30048 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _290_
timestamp 1676381911
transform 1 0 12960 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _291_
timestamp 1676381911
transform 1 0 20256 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _292_
timestamp 1676381911
transform 1 0 8064 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _293_
timestamp 1676381911
transform 1 0 13824 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _294_
timestamp 1676381911
transform 1 0 17472 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _295_
timestamp 1676381911
transform 1 0 13248 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _296_
timestamp 1676381911
transform 1 0 2400 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _297_
timestamp 1676381911
transform 1 0 7968 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _298_
timestamp 1676381911
transform 1 0 8928 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _299_
timestamp 1676381911
transform 1 0 8448 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _300_
timestamp 1676381911
transform 1 0 3840 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _301_
timestamp 1676381911
transform 1 0 2496 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _302_
timestamp 1676381911
transform 1 0 2496 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _303_
timestamp 1676381911
transform 1 0 8064 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _304_
timestamp 1676381911
transform 1 0 2880 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _305_
timestamp 1676381911
transform 1 0 2784 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _306_
timestamp 1676381911
transform 1 0 4896 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  _307_
timestamp 1676381911
transform 1 0 2208 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _308_
timestamp 1676381911
transform -1 0 28704 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _309_
timestamp 1676381911
transform 1 0 2016 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _310_
timestamp 1676381911
transform -1 0 37056 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _311_
timestamp 1676381911
transform -1 0 37536 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _312_
timestamp 1676381911
transform -1 0 43488 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _313_
timestamp 1676381911
transform -1 0 44928 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _314_
timestamp 1676381911
transform -1 0 44832 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _315_
timestamp 1676381911
transform -1 0 44448 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  _316_
timestamp 1676381911
transform -1 0 43008 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _317_
timestamp 1676381911
transform -1 0 44064 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  _318_
timestamp 1676381911
transform -1 0 44544 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _319_
timestamp 1676381911
transform -1 0 43776 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _320_
timestamp 1676381911
transform -1 0 44160 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _321_
timestamp 1676381911
transform -1 0 43392 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _322_
timestamp 1676381911
transform -1 0 43776 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _323_
timestamp 1676381911
transform -1 0 44448 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _324_
timestamp 1676381911
transform -1 0 44448 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _325_
timestamp 1676381911
transform -1 0 43680 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  _326_
timestamp 1676381911
transform -1 0 44832 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  _327_
timestamp 1676381911
transform -1 0 45216 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  _328_
timestamp 1676381911
transform -1 0 23616 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _329_
timestamp 1676381911
transform -1 0 26304 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _330_
timestamp 1676381911
transform -1 0 41952 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _331_
timestamp 1676381911
transform -1 0 38880 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _332_
timestamp 1676381911
transform 1 0 19872 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _333_
timestamp 1676381911
transform 1 0 18048 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _334_
timestamp 1676381911
transform -1 0 29184 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _335_
timestamp 1676381911
transform -1 0 30336 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _336_
timestamp 1676381911
transform 1 0 16896 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _337_
timestamp 1676381911
transform 1 0 16608 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _338_
timestamp 1676381911
transform 1 0 12384 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _339_
timestamp 1676381911
transform -1 0 26784 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _340_
timestamp 1676381911
transform 1 0 21408 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _341_
timestamp 1676381911
transform -1 0 23424 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _342_
timestamp 1676381911
transform -1 0 42048 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _343_
timestamp 1676381911
transform -1 0 36384 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _344_
timestamp 1676381911
transform 1 0 20256 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _345_
timestamp 1676381911
transform 1 0 16992 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _346_
timestamp 1676381911
transform 1 0 13344 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _347_
timestamp 1676381911
transform -1 0 28896 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _348_
timestamp 1676381911
transform 1 0 23712 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _349_
timestamp 1676381911
transform 1 0 23616 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _350_
timestamp 1676381911
transform 1 0 23520 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _351_
timestamp 1676381911
transform 1 0 20448 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _352_
timestamp 1676381911
transform 1 0 19680 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _353_
timestamp 1676381911
transform 1 0 19584 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _354_
timestamp 1676381911
transform 1 0 19392 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  _355_
timestamp 1676381911
transform 1 0 18240 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _356_
timestamp 1676381911
transform -1 0 42528 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _357_
timestamp 1676381911
transform -1 0 39648 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _358_
timestamp 1676381911
transform -1 0 33888 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _359_
timestamp 1676381911
transform -1 0 40608 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _360_
timestamp 1676381911
transform -1 0 42528 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _361_
timestamp 1676381911
transform -1 0 36288 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _362_
timestamp 1676381911
transform 1 0 26592 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _363_
timestamp 1676381911
transform -1 0 36960 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _364_
timestamp 1676381911
transform 1 0 27840 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _365_
timestamp 1676381911
transform -1 0 33504 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _366_
timestamp 1676381911
transform 1 0 29088 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _367_
timestamp 1676381911
transform -1 0 32928 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _368_
timestamp 1676381911
transform 1 0 8448 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _369_
timestamp 1676381911
transform 1 0 5664 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _370_
timestamp 1676381911
transform 1 0 6144 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _371_
timestamp 1676381911
transform 1 0 9408 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _372_
timestamp 1676381911
transform -1 0 38400 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _373_
timestamp 1676381911
transform -1 0 36576 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _374_
timestamp 1676381911
transform 1 0 32448 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _375_
timestamp 1676381911
transform -1 0 38784 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _376_
timestamp 1676381911
transform 1 0 37152 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  _377_
timestamp 1676381911
transform 1 0 32160 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _378_
timestamp 1676381911
transform 1 0 12096 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _379_
timestamp 1676381911
transform 1 0 13440 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _380_
timestamp 1676381911
transform -1 0 40512 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  fanout69
timestamp 1676381911
transform -1 0 4608 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  fanout70
timestamp 1676381911
transform -1 0 9408 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  fanout71
timestamp 1676381911
transform -1 0 40128 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  fanout72
timestamp 1676381911
transform 1 0 25632 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  fanout73
timestamp 1676381911
transform -1 0 36768 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  fanout74
timestamp 1676381911
transform 1 0 36768 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  fanout75
timestamp 1676381911
transform 1 0 36768 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  fanout76
timestamp 1676381911
transform 1 0 21792 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  fanout77
timestamp 1676381911
transform 1 0 22656 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  fanout78
timestamp 1676381911
transform -1 0 21792 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  fanout79
timestamp 1676381911
transform 1 0 24960 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  fanout80
timestamp 1676381911
transform 1 0 25344 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  fanout81
timestamp 1676381911
transform 1 0 21792 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  fanout82
timestamp 1676381911
transform -1 0 15840 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  fanout83
timestamp 1676381911
transform -1 0 24960 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  fanout84
timestamp 1676381911
transform 1 0 31872 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  fanout85
timestamp 1676381911
transform -1 0 30912 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  fanout86
timestamp 1676381911
transform 1 0 12768 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  fanout87
timestamp 1676381911
transform 1 0 2592 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  fanout88
timestamp 1676381911
transform 1 0 2784 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  fanout89
timestamp 1676381911
transform -1 0 27840 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  fanout90
timestamp 1676381911
transform 1 0 32832 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  fanout91
timestamp 1676381911
transform 1 0 28704 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_12
timestamp 1677580104
transform 1 0 2304 0 1 1512
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_14
timestamp 1677579658
transform 1 0 2496 0 1 1512
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_93
timestamp 1677579658
transform 1 0 10080 0 1 1512
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_198
timestamp 1677580104
transform 1 0 20160 0 1 1512
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_275
timestamp 1677579658
transform 1 0 27552 0 1 1512
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_305
timestamp 1677579658
transform 1 0 30432 0 1 1512
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_364
timestamp 1677580104
transform 1 0 36096 0 1 1512
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_366
timestamp 1677579658
transform 1 0 36288 0 1 1512
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_388
timestamp 1677580104
transform 1 0 38400 0 1 1512
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_390
timestamp 1677579658
transform 1 0 38592 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_408
timestamp 1679581782
transform 1 0 40320 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_415
timestamp 1679581782
transform 1 0 40992 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_422
timestamp 1679581782
transform 1 0 41664 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_429
timestamp 1679581782
transform 1 0 42336 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_436
timestamp 1679581782
transform 1 0 43008 0 1 1512
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_8
timestamp 1677579658
transform 1 0 1920 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_199
timestamp 1677580104
transform 1 0 20256 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_201
timestamp 1677579658
transform 1 0 20448 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_231
timestamp 1677580104
transform 1 0 23328 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_300
timestamp 1677579658
transform 1 0 29952 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_322
timestamp 1677580104
transform 1 0 32064 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_366
timestamp 1677579658
transform 1 0 36288 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_388
timestamp 1677580104
transform 1 0 38400 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_415
timestamp 1679581782
transform 1 0 40992 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_422
timestamp 1679581782
transform 1 0 41664 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_429
timestamp 1679581782
transform 1 0 42336 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_436
timestamp 1679581782
transform 1 0 43008 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_443
timestamp 1679577901
transform 1 0 43680 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_16
timestamp 1677579658
transform 1 0 2688 0 1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_38
timestamp 1677579658
transform 1 0 4800 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_70
timestamp 1677580104
transform 1 0 7872 0 1 3024
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_130
timestamp 1677580104
transform 1 0 13632 0 1 3024
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_165
timestamp 1677580104
transform 1 0 16992 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_167
timestamp 1677579658
transform 1 0 17184 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_238
timestamp 1677580104
transform 1 0 24000 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_240
timestamp 1677579658
transform 1 0 24192 0 1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_245
timestamp 1677579658
transform 1 0 24672 0 1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_267
timestamp 1677579658
transform 1 0 26784 0 1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_289
timestamp 1677579658
transform 1 0 28896 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_341
timestamp 1677580104
transform 1 0 33888 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_343
timestamp 1677579658
transform 1 0 34080 0 1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_373
timestamp 1677579658
transform 1 0 36960 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_391
timestamp 1677580104
transform 1 0 38688 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_393
timestamp 1677579658
transform 1 0 38880 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_425
timestamp 1679581782
transform 1 0 41952 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_432
timestamp 1679581782
transform 1 0 42624 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_439
timestamp 1679581782
transform 1 0 43296 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_446
timestamp 1679577901
transform 1 0 43968 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_450
timestamp 1677579658
transform 1 0 44352 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_8
timestamp 1677580104
transform 1 0 1920 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_10
timestamp 1677579658
transform 1 0 2112 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_107
timestamp 1677580104
transform 1 0 11424 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_159
timestamp 1677579658
transform 1 0 16416 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_177
timestamp 1677580104
transform 1 0 18144 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_179
timestamp 1677579658
transform 1 0 18336 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_201
timestamp 1677580104
transform 1 0 20448 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_232
timestamp 1677579658
transform 1 0 23424 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_241
timestamp 1677580104
transform 1 0 24288 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_243
timestamp 1677579658
transform 1 0 24480 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_264
timestamp 1677579658
transform 1 0 26496 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_282
timestamp 1677580104
transform 1 0 28224 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_284
timestamp 1677579658
transform 1 0 28416 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_310
timestamp 1677580104
transform 1 0 30912 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_337
timestamp 1677579658
transform 1 0 33504 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_396
timestamp 1679577901
transform 1 0 39168 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_400
timestamp 1677579658
transform 1 0 39552 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_405
timestamp 1677579658
transform 1 0 40032 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_410
timestamp 1679577901
transform 1 0 40512 0 -1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_418
timestamp 1679581782
transform 1 0 41280 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_425
timestamp 1679581782
transform 1 0 41952 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_432
timestamp 1679581782
transform 1 0 42624 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_439
timestamp 1679581782
transform 1 0 43296 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_446
timestamp 1677579658
transform 1 0 43968 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_8
timestamp 1679577901
transform 1 0 1920 0 1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_12
timestamp 1677580104
transform 1 0 2304 0 1 4536
box -48 -56 240 834
use sg13g2_decap_4  FILLER_4_22
timestamp 1679577901
transform 1 0 3264 0 1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_108
timestamp 1677580104
transform 1 0 11520 0 1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_139
timestamp 1677580104
transform 1 0 14496 0 1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_162
timestamp 1677580104
transform 1 0 16704 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_202
timestamp 1677579658
transform 1 0 20544 0 1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_234
timestamp 1677579658
transform 1 0 23616 0 1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_252
timestamp 1677579658
transform 1 0 25344 0 1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_278
timestamp 1677580104
transform 1 0 27840 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_280
timestamp 1677579658
transform 1 0 28032 0 1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_344
timestamp 1677579658
transform 1 0 34176 0 1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_374
timestamp 1677580104
transform 1 0 37056 0 1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_401
timestamp 1677580104
transform 1 0 39648 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_429
timestamp 1679581782
transform 1 0 42336 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_436
timestamp 1679581782
transform 1 0 43008 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_443
timestamp 1679581782
transform 1 0 43680 0 1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_450
timestamp 1677579658
transform 1 0 44352 0 1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_8
timestamp 1677580104
transform 1 0 1920 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_10
timestamp 1677579658
transform 1 0 2112 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_81
timestamp 1677579658
transform 1 0 8928 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_108
timestamp 1677579658
transform 1 0 11520 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_143
timestamp 1677580104
transform 1 0 14880 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_183
timestamp 1677579658
transform 1 0 18720 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_205
timestamp 1677580104
transform 1 0 20832 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_207
timestamp 1677579658
transform 1 0 21024 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_250
timestamp 1677579658
transform 1 0 25152 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_272
timestamp 1677580104
transform 1 0 27264 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_298
timestamp 1677580104
transform 1 0 29760 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_304
timestamp 1677579658
transform 1 0 30336 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_338
timestamp 1677579658
transform 1 0 33600 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_360
timestamp 1677580104
transform 1 0 35712 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_4  FILLER_5_397
timestamp 1679577901
transform 1 0 39264 0 -1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_427
timestamp 1679581782
transform 1 0 42144 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_434
timestamp 1679581782
transform 1 0 42816 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_441
timestamp 1679581782
transform 1 0 43488 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_448
timestamp 1677580104
transform 1 0 44160 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_450
timestamp 1677579658
transform 1 0 44352 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_12
timestamp 1677580104
transform 1 0 2304 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_14
timestamp 1677579658
transform 1 0 2496 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_80
timestamp 1677580104
transform 1 0 8832 0 1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_106
timestamp 1677580104
transform 1 0 11328 0 1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_125
timestamp 1677580104
transform 1 0 13152 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_169
timestamp 1677579658
transform 1 0 17376 0 1 6048
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_207
timestamp 1679577901
transform 1 0 21024 0 1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_236
timestamp 1679581782
transform 1 0 23808 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_243
timestamp 1679581782
transform 1 0 24480 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_250
timestamp 1679577901
transform 1 0 25152 0 1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_254
timestamp 1677579658
transform 1 0 25536 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_259
timestamp 1679581782
transform 1 0 26016 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_299
timestamp 1677580104
transform 1 0 29856 0 1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_305
timestamp 1677580104
transform 1 0 30432 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_375
timestamp 1679581782
transform 1 0 37152 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_382
timestamp 1679577901
transform 1 0 37824 0 1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_386
timestamp 1677579658
transform 1 0 38208 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_391
timestamp 1677580104
transform 1 0 38688 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_410
timestamp 1677579658
transform 1 0 40512 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_415
timestamp 1679581782
transform 1 0 40992 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_422
timestamp 1679581782
transform 1 0 41664 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_429
timestamp 1679581782
transform 1 0 42336 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_436
timestamp 1679581782
transform 1 0 43008 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_443
timestamp 1679577901
transform 1 0 43680 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_8
timestamp 1677580104
transform 1 0 1920 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_44
timestamp 1677580104
transform 1 0 5376 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_46
timestamp 1677579658
transform 1 0 5568 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_60
timestamp 1677579658
transform 1 0 6912 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_125
timestamp 1677579658
transform 1 0 13152 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_147
timestamp 1677580104
transform 1 0 15264 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_166
timestamp 1677580104
transform 1 0 17088 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_168
timestamp 1677579658
transform 1 0 17280 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_236
timestamp 1677580104
transform 1 0 23808 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_255
timestamp 1677580104
transform 1 0 25632 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_257
timestamp 1677579658
transform 1 0 25824 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_262
timestamp 1679581782
transform 1 0 26304 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_269
timestamp 1677579658
transform 1 0 26976 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_304
timestamp 1677579658
transform 1 0 30336 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_355
timestamp 1679581782
transform 1 0 35232 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_362
timestamp 1679577901
transform 1 0 35904 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_366
timestamp 1677579658
transform 1 0 36288 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_379
timestamp 1679577901
transform 1 0 37536 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_383
timestamp 1677579658
transform 1 0 37920 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_401
timestamp 1677579658
transform 1 0 39648 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_431
timestamp 1679581782
transform 1 0 42528 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_438
timestamp 1677579658
transform 1 0 43200 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_8
timestamp 1679581782
transform 1 0 1920 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_15
timestamp 1677579658
transform 1 0 2592 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_33
timestamp 1679577901
transform 1 0 4320 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_37
timestamp 1677580104
transform 1 0 4704 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_83
timestamp 1677579658
transform 1 0 9120 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_103
timestamp 1677580104
transform 1 0 11040 0 1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_121
timestamp 1677580104
transform 1 0 12768 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_127
timestamp 1677579658
transform 1 0 13344 0 1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_132
timestamp 1677579658
transform 1 0 13824 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_190
timestamp 1677580104
transform 1 0 19392 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_192
timestamp 1677579658
transform 1 0 19584 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_197
timestamp 1677580104
transform 1 0 20064 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_220
timestamp 1679581782
transform 1 0 22272 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_227
timestamp 1677580104
transform 1 0 22944 0 1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_233
timestamp 1677580104
transform 1 0 23520 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_266
timestamp 1677579658
transform 1 0 26688 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_300
timestamp 1677580104
transform 1 0 29952 0 1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_348
timestamp 1677580104
transform 1 0 34560 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_375
timestamp 1679581782
transform 1 0 37152 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_403
timestamp 1677580104
transform 1 0 39840 0 1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_426
timestamp 1677580104
transform 1 0 42048 0 1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_444
timestamp 1677580104
transform 1 0 43776 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_446
timestamp 1677579658
transform 1 0 43968 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_8
timestamp 1679577901
transform 1 0 1920 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_12
timestamp 1677580104
transform 1 0 2304 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_18
timestamp 1679581782
transform 1 0 2880 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_25
timestamp 1677580104
transform 1 0 3552 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_27
timestamp 1677579658
transform 1 0 3744 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_90
timestamp 1679577901
transform 1 0 9792 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_191
timestamp 1677580104
transform 1 0 19488 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_197
timestamp 1677579658
transform 1 0 20064 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_219
timestamp 1679577901
transform 1 0 22176 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_223
timestamp 1677580104
transform 1 0 22560 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_242
timestamp 1679581782
transform 1 0 24384 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_249
timestamp 1677579658
transform 1 0 25056 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_267
timestamp 1677580104
transform 1 0 26784 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_9_286
timestamp 1679577901
transform 1 0 28608 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_290
timestamp 1677579658
transform 1 0 28992 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_337
timestamp 1679581782
transform 1 0 33504 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_369
timestamp 1677579658
transform 1 0 36576 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_404
timestamp 1677580104
transform 1 0 39936 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_431
timestamp 1677580104
transform 1 0 42528 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_441
timestamp 1677580104
transform 1 0 43488 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_12
timestamp 1679581782
transform 1 0 2304 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_19
timestamp 1679581782
transform 1 0 2976 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_26
timestamp 1679577901
transform 1 0 3648 0 1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_30
timestamp 1677580104
transform 1 0 4032 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_71
timestamp 1677579658
transform 1 0 7968 0 1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_80
timestamp 1677579658
transform 1 0 8832 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_85
timestamp 1677580104
transform 1 0 9312 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_87
timestamp 1677579658
transform 1 0 9504 0 1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_105
timestamp 1677579658
transform 1 0 11232 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_131
timestamp 1677580104
transform 1 0 13728 0 1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_137
timestamp 1677580104
transform 1 0 14304 0 1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_168
timestamp 1679577901
transform 1 0 17280 0 1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_172
timestamp 1677580104
transform 1 0 17664 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_203
timestamp 1677579658
transform 1 0 20640 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_237
timestamp 1677580104
transform 1 0 23904 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_239
timestamp 1677579658
transform 1 0 24096 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_269
timestamp 1677580104
transform 1 0 26976 0 1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_309
timestamp 1677580104
transform 1 0 30816 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_311
timestamp 1677579658
transform 1 0 31008 0 1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_345
timestamp 1677579658
transform 1 0 34272 0 1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_367
timestamp 1677579658
transform 1 0 36384 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_389
timestamp 1677580104
transform 1 0 38496 0 1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_429
timestamp 1677580104
transform 1 0 42336 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_431
timestamp 1677579658
transform 1 0 42528 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_456
timestamp 1677580104
transform 1 0 44928 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_458
timestamp 1677579658
transform 1 0 45120 0 1 9072
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_20
timestamp 1679577901
transform 1 0 3072 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_24
timestamp 1677579658
transform 1 0 3456 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_29
timestamp 1679581782
transform 1 0 3936 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_36
timestamp 1677580104
transform 1 0 4608 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_38
timestamp 1677579658
transform 1 0 4800 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_47
timestamp 1677580104
transform 1 0 5664 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_53
timestamp 1679577901
transform 1 0 6240 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_57
timestamp 1677579658
transform 1 0 6624 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_70
timestamp 1677580104
transform 1 0 7872 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_101
timestamp 1677580104
transform 1 0 10848 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_187
timestamp 1677580104
transform 1 0 19104 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_189
timestamp 1677579658
transform 1 0 19296 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_194
timestamp 1677580104
transform 1 0 19776 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_213
timestamp 1677580104
transform 1 0 21600 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_232
timestamp 1677580104
transform 1 0 23424 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_234
timestamp 1677579658
transform 1 0 23616 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_281
timestamp 1677579658
transform 1 0 28128 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_353
timestamp 1677579658
transform 1 0 35040 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_383
timestamp 1677580104
transform 1 0 37920 0 -1 10584
box -48 -56 240 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform 1 0 3552 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1676381911
transform 1 0 7488 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  input3
timestamp 1676381911
transform 1 0 2304 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input4
timestamp 1676381911
transform 1 0 1152 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  input5
timestamp 1676381911
transform 1 0 1536 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  input6
timestamp 1676381911
transform 1 0 1152 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  input7
timestamp 1676381911
transform 1 0 1536 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input8
timestamp 1676381911
transform 1 0 1152 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input9
timestamp 1676381911
transform 1 0 1920 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  input10
timestamp 1676381911
transform 1 0 1536 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  input11
timestamp 1676381911
transform 1 0 1152 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  input12
timestamp 1676381911
transform 1 0 1536 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input13
timestamp 1676381911
transform 1 0 1152 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input14
timestamp 1676381911
transform 1 0 1536 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input15
timestamp 1676381911
transform 1 0 1152 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input16
timestamp 1676381911
transform 1 0 1536 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input17
timestamp 1676381911
transform 1 0 1152 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input18
timestamp 1676381911
transform 1 0 1536 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input19
timestamp 1676381911
transform 1 0 1152 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input20
timestamp 1676381911
transform 1 0 1536 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input21
timestamp 1676381911
transform 1 0 1152 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  input22
timestamp 1676381911
transform 1 0 1536 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  input23
timestamp 1676381911
transform 1 0 1920 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  input24
timestamp 1676381911
transform 1 0 2304 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  input25
timestamp 1676381911
transform 1 0 1920 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input26
timestamp 1676381911
transform 1 0 1920 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input27
timestamp 1676381911
transform 1 0 2688 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  input28
timestamp 1676381911
transform 1 0 1152 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input29
timestamp 1676381911
transform 1 0 1536 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input30
timestamp 1676381911
transform 1 0 1152 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input31
timestamp 1676381911
transform 1 0 1920 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input32
timestamp 1676381911
transform 1 0 1536 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input33
timestamp 1676381911
transform 1 0 1152 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input34
timestamp 1676381911
transform 1 0 1536 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  input35
timestamp 1676381911
transform -1 0 38400 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input36
timestamp 1676381911
transform 1 0 10176 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input37
timestamp 1676381911
transform 1 0 4608 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  input38
timestamp 1676381911
transform 1 0 3168 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input39
timestamp 1676381911
transform 1 0 2592 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input40
timestamp 1676381911
transform -1 0 9408 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input41
timestamp 1676381911
transform -1 0 12000 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input42
timestamp 1676381911
transform -1 0 12384 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input43
timestamp 1676381911
transform -1 0 10176 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input44
timestamp 1676381911
transform -1 0 10560 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input45
timestamp 1676381911
transform -1 0 6912 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input46
timestamp 1676381911
transform -1 0 7296 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input47
timestamp 1676381911
transform -1 0 8832 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input48
timestamp 1676381911
transform 1 0 3552 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input49
timestamp 1676381911
transform 1 0 2976 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input50
timestamp 1676381911
transform 1 0 3936 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input51
timestamp 1676381911
transform 1 0 3360 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input52
timestamp 1676381911
transform 1 0 3744 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input53
timestamp 1676381911
transform 1 0 4128 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input54
timestamp 1676381911
transform -1 0 11616 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input55
timestamp 1676381911
transform 1 0 4512 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input56
timestamp 1676381911
transform 1 0 13920 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input57
timestamp 1676381911
transform 1 0 15840 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input58
timestamp 1676381911
transform 1 0 11616 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  input59
timestamp 1676381911
transform 1 0 16224 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input60
timestamp 1676381911
transform 1 0 12000 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  input61
timestamp 1676381911
transform 1 0 12384 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  input62
timestamp 1676381911
transform 1 0 10176 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input63
timestamp 1676381911
transform 1 0 7296 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input64
timestamp 1676381911
transform 1 0 14304 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input65
timestamp 1676381911
transform 1 0 8832 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input66
timestamp 1676381911
transform 1 0 14688 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input67
timestamp 1676381911
transform 1 0 9216 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input68
timestamp 1676381911
transform 1 0 15072 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input69
timestamp 1676381911
transform 1 0 7680 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input70
timestamp 1676381911
transform 1 0 11712 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  input71
timestamp 1676381911
transform 1 0 8064 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input72
timestamp 1676381911
transform 1 0 19008 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input73
timestamp 1676381911
transform -1 0 20640 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  input74
timestamp 1676381911
transform 1 0 15360 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input75
timestamp 1676381911
transform 1 0 17280 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input76
timestamp 1676381911
transform 1 0 15744 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input77
timestamp 1676381911
transform -1 0 18048 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input78
timestamp 1676381911
transform 1 0 16128 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input79
timestamp 1676381911
transform 1 0 18624 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input80
timestamp 1676381911
transform 1 0 12192 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input81
timestamp 1676381911
transform 1 0 12576 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input82
timestamp 1676381911
transform 1 0 14208 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input83
timestamp 1676381911
transform 1 0 12960 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input84
timestamp 1676381911
transform 1 0 14592 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input85
timestamp 1676381911
transform 1 0 13344 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input86
timestamp 1676381911
transform 1 0 14976 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input87
timestamp 1676381911
transform 1 0 20640 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output88
timestamp 1676381911
transform -1 0 5664 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output89
timestamp 1676381911
transform -1 0 6240 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output90
timestamp 1676381911
transform 1 0 8832 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output91
timestamp 1676381911
transform 1 0 11040 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output92
timestamp 1676381911
transform 1 0 11424 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output93
timestamp 1676381911
transform -1 0 14304 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output94
timestamp 1676381911
transform -1 0 8448 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output95
timestamp 1676381911
transform 1 0 8448 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output96
timestamp 1676381911
transform 1 0 14496 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output97
timestamp 1676381911
transform -1 0 17088 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output98
timestamp 1676381911
transform 1 0 17088 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output99
timestamp 1676381911
transform 1 0 17856 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output100
timestamp 1676381911
transform 1 0 44064 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output101
timestamp 1676381911
transform 1 0 44448 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output102
timestamp 1676381911
transform 1 0 44832 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output103
timestamp 1676381911
transform 1 0 44448 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output104
timestamp 1676381911
transform 1 0 44832 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output105
timestamp 1676381911
transform 1 0 44448 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output106
timestamp 1676381911
transform 1 0 44832 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output107
timestamp 1676381911
transform 1 0 44448 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output108
timestamp 1676381911
transform 1 0 44832 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output109
timestamp 1676381911
transform 1 0 44448 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output110
timestamp 1676381911
transform 1 0 44832 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output111
timestamp 1676381911
transform 1 0 43680 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output112
timestamp 1676381911
transform 1 0 44832 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output113
timestamp 1676381911
transform 1 0 44448 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output114
timestamp 1676381911
transform 1 0 44832 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output115
timestamp 1676381911
transform 1 0 43680 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output116
timestamp 1676381911
transform 1 0 42720 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output117
timestamp 1676381911
transform 1 0 44064 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output118
timestamp 1676381911
transform 1 0 43008 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output119
timestamp 1676381911
transform 1 0 43680 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output120
timestamp 1676381911
transform 1 0 42624 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output121
timestamp 1676381911
transform 1 0 44064 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output122
timestamp 1676381911
transform 1 0 44064 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output123
timestamp 1676381911
transform 1 0 43296 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output124
timestamp 1676381911
transform 1 0 42240 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output125
timestamp 1676381911
transform 1 0 44448 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output126
timestamp 1676381911
transform 1 0 44832 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output127
timestamp 1676381911
transform 1 0 44448 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output128
timestamp 1676381911
transform 1 0 44832 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output129
timestamp 1676381911
transform 1 0 44448 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output130
timestamp 1676381911
transform 1 0 44064 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output131
timestamp 1676381911
transform 1 0 44832 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output132
timestamp 1676381911
transform -1 0 21120 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output133
timestamp 1676381911
transform -1 0 33504 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output134
timestamp 1676381911
transform -1 0 34272 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output135
timestamp 1676381911
transform -1 0 35040 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output136
timestamp 1676381911
transform -1 0 37152 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output137
timestamp 1676381911
transform -1 0 37920 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output138
timestamp 1676381911
transform -1 0 38496 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output139
timestamp 1676381911
transform 1 0 38496 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output140
timestamp 1676381911
transform -1 0 42528 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output141
timestamp 1676381911
transform -1 0 42912 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output142
timestamp 1676381911
transform -1 0 43296 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output143
timestamp 1676381911
transform 1 0 21120 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output144
timestamp 1676381911
transform -1 0 23520 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output145
timestamp 1676381911
transform 1 0 23712 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output146
timestamp 1676381911
transform -1 0 26592 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output147
timestamp 1676381911
transform -1 0 27744 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output148
timestamp 1676381911
transform -1 0 28128 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output149
timestamp 1676381911
transform -1 0 30240 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output150
timestamp 1676381911
transform -1 0 32640 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output151
timestamp 1676381911
transform -1 0 33024 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output152
timestamp 1676381911
transform 1 0 16512 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output153
timestamp 1676381911
transform 1 0 17472 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output154
timestamp 1676381911
transform 1 0 18432 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output155
timestamp 1676381911
transform 1 0 17856 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output156
timestamp 1676381911
transform 1 0 21120 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output157
timestamp 1676381911
transform 1 0 19200 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output158
timestamp 1676381911
transform 1 0 21504 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output159
timestamp 1676381911
transform 1 0 19968 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output160
timestamp 1676381911
transform 1 0 20544 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output161
timestamp 1676381911
transform 1 0 20928 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output162
timestamp 1676381911
transform 1 0 20352 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output163
timestamp 1676381911
transform 1 0 20736 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output164
timestamp 1676381911
transform -1 0 23904 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output165
timestamp 1676381911
transform 1 0 21120 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output166
timestamp 1676381911
transform -1 0 24288 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output167
timestamp 1676381911
transform -1 0 26304 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output168
timestamp 1676381911
transform -1 0 24672 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output169
timestamp 1676381911
transform 1 0 23520 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output170
timestamp 1676381911
transform -1 0 27168 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output171
timestamp 1676381911
transform -1 0 27552 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output172
timestamp 1676381911
transform -1 0 26112 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output173
timestamp 1676381911
transform -1 0 32928 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output174
timestamp 1676381911
transform -1 0 30528 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output175
timestamp 1676381911
transform -1 0 33312 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output176
timestamp 1676381911
transform -1 0 29376 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output177
timestamp 1676381911
transform -1 0 33696 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output178
timestamp 1676381911
transform -1 0 29760 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output179
timestamp 1676381911
transform -1 0 26496 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output180
timestamp 1676381911
transform -1 0 29664 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output181
timestamp 1676381911
transform -1 0 30048 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output182
timestamp 1676381911
transform -1 0 30432 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output183
timestamp 1676381911
transform -1 0 27456 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output184
timestamp 1676381911
transform -1 0 27840 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output185
timestamp 1676381911
transform -1 0 28608 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output186
timestamp 1676381911
transform -1 0 32544 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output187
timestamp 1676381911
transform -1 0 28992 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output188
timestamp 1676381911
transform -1 0 34080 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output189
timestamp 1676381911
transform -1 0 36192 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output190
timestamp 1676381911
transform -1 0 32448 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output191
timestamp 1676381911
transform -1 0 38400 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output192
timestamp 1676381911
transform -1 0 36576 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output193
timestamp 1676381911
transform -1 0 32832 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output194
timestamp 1676381911
transform -1 0 36000 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output195
timestamp 1676381911
transform -1 0 29472 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output196
timestamp 1676381911
transform -1 0 29856 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output197
timestamp 1676381911
transform -1 0 32160 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output198
timestamp 1676381911
transform -1 0 32544 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output199
timestamp 1676381911
transform -1 0 29568 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output200
timestamp 1676381911
transform -1 0 36288 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output201
timestamp 1676381911
transform -1 0 29952 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output202
timestamp 1676381911
transform -1 0 33216 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output203
timestamp 1676381911
transform -1 0 33600 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output204
timestamp 1676381911
transform -1 0 20064 0 -1 9072
box -48 -56 432 834
<< labels >>
flabel metal3 s 4664 12100 4744 12180 0 FreeSans 320 0 0 0 A_I_top
port 0 nsew signal output
flabel metal3 s 3512 12100 3592 12180 0 FreeSans 320 0 0 0 A_O_top
port 1 nsew signal input
flabel metal3 s 5816 12100 5896 12180 0 FreeSans 320 0 0 0 A_T_top
port 2 nsew signal output
flabel metal3 s 10424 12100 10504 12180 0 FreeSans 320 0 0 0 A_config_C_bit0
port 3 nsew signal output
flabel metal3 s 11576 12100 11656 12180 0 FreeSans 320 0 0 0 A_config_C_bit1
port 4 nsew signal output
flabel metal3 s 12728 12100 12808 12180 0 FreeSans 320 0 0 0 A_config_C_bit2
port 5 nsew signal output
flabel metal3 s 13880 12100 13960 12180 0 FreeSans 320 0 0 0 A_config_C_bit3
port 6 nsew signal output
flabel metal3 s 8120 12100 8200 12180 0 FreeSans 320 0 0 0 B_I_top
port 7 nsew signal output
flabel metal3 s 6968 12100 7048 12180 0 FreeSans 320 0 0 0 B_O_top
port 8 nsew signal input
flabel metal3 s 9272 12100 9352 12180 0 FreeSans 320 0 0 0 B_T_top
port 9 nsew signal output
flabel metal3 s 15032 12100 15112 12180 0 FreeSans 320 0 0 0 B_config_C_bit0
port 10 nsew signal output
flabel metal3 s 16184 12100 16264 12180 0 FreeSans 320 0 0 0 B_config_C_bit1
port 11 nsew signal output
flabel metal3 s 17336 12100 17416 12180 0 FreeSans 320 0 0 0 B_config_C_bit2
port 12 nsew signal output
flabel metal3 s 18488 12100 18568 12180 0 FreeSans 320 0 0 0 B_config_C_bit3
port 13 nsew signal output
flabel metal3 s 20984 0 21064 80 0 FreeSans 320 0 0 0 Ci
port 14 nsew signal input
flabel metal2 s 0 716 90 796 0 FreeSans 320 0 0 0 FrameData[0]
port 15 nsew signal input
flabel metal2 s 0 4076 90 4156 0 FreeSans 320 0 0 0 FrameData[10]
port 16 nsew signal input
flabel metal2 s 0 4412 90 4492 0 FreeSans 320 0 0 0 FrameData[11]
port 17 nsew signal input
flabel metal2 s 0 4748 90 4828 0 FreeSans 320 0 0 0 FrameData[12]
port 18 nsew signal input
flabel metal2 s 0 5084 90 5164 0 FreeSans 320 0 0 0 FrameData[13]
port 19 nsew signal input
flabel metal2 s 0 5420 90 5500 0 FreeSans 320 0 0 0 FrameData[14]
port 20 nsew signal input
flabel metal2 s 0 5756 90 5836 0 FreeSans 320 0 0 0 FrameData[15]
port 21 nsew signal input
flabel metal2 s 0 6092 90 6172 0 FreeSans 320 0 0 0 FrameData[16]
port 22 nsew signal input
flabel metal2 s 0 6428 90 6508 0 FreeSans 320 0 0 0 FrameData[17]
port 23 nsew signal input
flabel metal2 s 0 6764 90 6844 0 FreeSans 320 0 0 0 FrameData[18]
port 24 nsew signal input
flabel metal2 s 0 7100 90 7180 0 FreeSans 320 0 0 0 FrameData[19]
port 25 nsew signal input
flabel metal2 s 0 1052 90 1132 0 FreeSans 320 0 0 0 FrameData[1]
port 26 nsew signal input
flabel metal2 s 0 7436 90 7516 0 FreeSans 320 0 0 0 FrameData[20]
port 27 nsew signal input
flabel metal2 s 0 7772 90 7852 0 FreeSans 320 0 0 0 FrameData[21]
port 28 nsew signal input
flabel metal2 s 0 8108 90 8188 0 FreeSans 320 0 0 0 FrameData[22]
port 29 nsew signal input
flabel metal2 s 0 8444 90 8524 0 FreeSans 320 0 0 0 FrameData[23]
port 30 nsew signal input
flabel metal2 s 0 8780 90 8860 0 FreeSans 320 0 0 0 FrameData[24]
port 31 nsew signal input
flabel metal2 s 0 9116 90 9196 0 FreeSans 320 0 0 0 FrameData[25]
port 32 nsew signal input
flabel metal2 s 0 9452 90 9532 0 FreeSans 320 0 0 0 FrameData[26]
port 33 nsew signal input
flabel metal2 s 0 9788 90 9868 0 FreeSans 320 0 0 0 FrameData[27]
port 34 nsew signal input
flabel metal2 s 0 10124 90 10204 0 FreeSans 320 0 0 0 FrameData[28]
port 35 nsew signal input
flabel metal2 s 0 10460 90 10540 0 FreeSans 320 0 0 0 FrameData[29]
port 36 nsew signal input
flabel metal2 s 0 1388 90 1468 0 FreeSans 320 0 0 0 FrameData[2]
port 37 nsew signal input
flabel metal2 s 0 10796 90 10876 0 FreeSans 320 0 0 0 FrameData[30]
port 38 nsew signal input
flabel metal2 s 0 11132 90 11212 0 FreeSans 320 0 0 0 FrameData[31]
port 39 nsew signal input
flabel metal2 s 0 1724 90 1804 0 FreeSans 320 0 0 0 FrameData[3]
port 40 nsew signal input
flabel metal2 s 0 2060 90 2140 0 FreeSans 320 0 0 0 FrameData[4]
port 41 nsew signal input
flabel metal2 s 0 2396 90 2476 0 FreeSans 320 0 0 0 FrameData[5]
port 42 nsew signal input
flabel metal2 s 0 2732 90 2812 0 FreeSans 320 0 0 0 FrameData[6]
port 43 nsew signal input
flabel metal2 s 0 3068 90 3148 0 FreeSans 320 0 0 0 FrameData[7]
port 44 nsew signal input
flabel metal2 s 0 3404 90 3484 0 FreeSans 320 0 0 0 FrameData[8]
port 45 nsew signal input
flabel metal2 s 0 3740 90 3820 0 FreeSans 320 0 0 0 FrameData[9]
port 46 nsew signal input
flabel metal2 s 46278 716 46368 796 0 FreeSans 320 0 0 0 FrameData_O[0]
port 47 nsew signal output
flabel metal2 s 46278 4076 46368 4156 0 FreeSans 320 0 0 0 FrameData_O[10]
port 48 nsew signal output
flabel metal2 s 46278 4412 46368 4492 0 FreeSans 320 0 0 0 FrameData_O[11]
port 49 nsew signal output
flabel metal2 s 46278 4748 46368 4828 0 FreeSans 320 0 0 0 FrameData_O[12]
port 50 nsew signal output
flabel metal2 s 46278 5084 46368 5164 0 FreeSans 320 0 0 0 FrameData_O[13]
port 51 nsew signal output
flabel metal2 s 46278 5420 46368 5500 0 FreeSans 320 0 0 0 FrameData_O[14]
port 52 nsew signal output
flabel metal2 s 46278 5756 46368 5836 0 FreeSans 320 0 0 0 FrameData_O[15]
port 53 nsew signal output
flabel metal2 s 46278 6092 46368 6172 0 FreeSans 320 0 0 0 FrameData_O[16]
port 54 nsew signal output
flabel metal2 s 46278 6428 46368 6508 0 FreeSans 320 0 0 0 FrameData_O[17]
port 55 nsew signal output
flabel metal2 s 46278 6764 46368 6844 0 FreeSans 320 0 0 0 FrameData_O[18]
port 56 nsew signal output
flabel metal2 s 46278 7100 46368 7180 0 FreeSans 320 0 0 0 FrameData_O[19]
port 57 nsew signal output
flabel metal2 s 46278 1052 46368 1132 0 FreeSans 320 0 0 0 FrameData_O[1]
port 58 nsew signal output
flabel metal2 s 46278 7436 46368 7516 0 FreeSans 320 0 0 0 FrameData_O[20]
port 59 nsew signal output
flabel metal2 s 46278 7772 46368 7852 0 FreeSans 320 0 0 0 FrameData_O[21]
port 60 nsew signal output
flabel metal2 s 46278 8108 46368 8188 0 FreeSans 320 0 0 0 FrameData_O[22]
port 61 nsew signal output
flabel metal2 s 46278 8444 46368 8524 0 FreeSans 320 0 0 0 FrameData_O[23]
port 62 nsew signal output
flabel metal2 s 46278 8780 46368 8860 0 FreeSans 320 0 0 0 FrameData_O[24]
port 63 nsew signal output
flabel metal2 s 46278 9116 46368 9196 0 FreeSans 320 0 0 0 FrameData_O[25]
port 64 nsew signal output
flabel metal2 s 46278 9452 46368 9532 0 FreeSans 320 0 0 0 FrameData_O[26]
port 65 nsew signal output
flabel metal2 s 46278 9788 46368 9868 0 FreeSans 320 0 0 0 FrameData_O[27]
port 66 nsew signal output
flabel metal2 s 46278 10124 46368 10204 0 FreeSans 320 0 0 0 FrameData_O[28]
port 67 nsew signal output
flabel metal2 s 46278 10460 46368 10540 0 FreeSans 320 0 0 0 FrameData_O[29]
port 68 nsew signal output
flabel metal2 s 46278 1388 46368 1468 0 FreeSans 320 0 0 0 FrameData_O[2]
port 69 nsew signal output
flabel metal2 s 46278 10796 46368 10876 0 FreeSans 320 0 0 0 FrameData_O[30]
port 70 nsew signal output
flabel metal2 s 46278 11132 46368 11212 0 FreeSans 320 0 0 0 FrameData_O[31]
port 71 nsew signal output
flabel metal2 s 46278 1724 46368 1804 0 FreeSans 320 0 0 0 FrameData_O[3]
port 72 nsew signal output
flabel metal2 s 46278 2060 46368 2140 0 FreeSans 320 0 0 0 FrameData_O[4]
port 73 nsew signal output
flabel metal2 s 46278 2396 46368 2476 0 FreeSans 320 0 0 0 FrameData_O[5]
port 74 nsew signal output
flabel metal2 s 46278 2732 46368 2812 0 FreeSans 320 0 0 0 FrameData_O[6]
port 75 nsew signal output
flabel metal2 s 46278 3068 46368 3148 0 FreeSans 320 0 0 0 FrameData_O[7]
port 76 nsew signal output
flabel metal2 s 46278 3404 46368 3484 0 FreeSans 320 0 0 0 FrameData_O[8]
port 77 nsew signal output
flabel metal2 s 46278 3740 46368 3820 0 FreeSans 320 0 0 0 FrameData_O[9]
port 78 nsew signal output
flabel metal3 s 31352 0 31432 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 79 nsew signal input
flabel metal3 s 33272 0 33352 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 80 nsew signal input
flabel metal3 s 33464 0 33544 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 81 nsew signal input
flabel metal3 s 33656 0 33736 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 82 nsew signal input
flabel metal3 s 33848 0 33928 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 83 nsew signal input
flabel metal3 s 34040 0 34120 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 84 nsew signal input
flabel metal3 s 34232 0 34312 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 85 nsew signal input
flabel metal3 s 34424 0 34504 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 86 nsew signal input
flabel metal3 s 34616 0 34696 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 87 nsew signal input
flabel metal3 s 34808 0 34888 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 88 nsew signal input
flabel metal3 s 35000 0 35080 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 89 nsew signal input
flabel metal3 s 31544 0 31624 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 90 nsew signal input
flabel metal3 s 31736 0 31816 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 91 nsew signal input
flabel metal3 s 31928 0 32008 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 92 nsew signal input
flabel metal3 s 32120 0 32200 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 93 nsew signal input
flabel metal3 s 32312 0 32392 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 94 nsew signal input
flabel metal3 s 32504 0 32584 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 95 nsew signal input
flabel metal3 s 32696 0 32776 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 96 nsew signal input
flabel metal3 s 32888 0 32968 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 97 nsew signal input
flabel metal3 s 33080 0 33160 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 98 nsew signal input
flabel metal3 s 20792 12100 20872 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 99 nsew signal output
flabel metal3 s 32312 12100 32392 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 100 nsew signal output
flabel metal3 s 33464 12100 33544 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 101 nsew signal output
flabel metal3 s 34616 12100 34696 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 102 nsew signal output
flabel metal3 s 35768 12100 35848 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 103 nsew signal output
flabel metal3 s 36920 12100 37000 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 104 nsew signal output
flabel metal3 s 38072 12100 38152 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 105 nsew signal output
flabel metal3 s 39224 12100 39304 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 106 nsew signal output
flabel metal3 s 40376 12100 40456 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 107 nsew signal output
flabel metal3 s 41528 12100 41608 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 108 nsew signal output
flabel metal3 s 42680 12100 42760 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 109 nsew signal output
flabel metal3 s 21944 12100 22024 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 110 nsew signal output
flabel metal3 s 23096 12100 23176 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 111 nsew signal output
flabel metal3 s 24248 12100 24328 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 112 nsew signal output
flabel metal3 s 25400 12100 25480 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 113 nsew signal output
flabel metal3 s 26552 12100 26632 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 114 nsew signal output
flabel metal3 s 27704 12100 27784 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 115 nsew signal output
flabel metal3 s 28856 12100 28936 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 116 nsew signal output
flabel metal3 s 30008 12100 30088 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 117 nsew signal output
flabel metal3 s 31160 12100 31240 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 118 nsew signal output
flabel metal3 s 11000 0 11080 80 0 FreeSans 320 0 0 0 N1END[0]
port 119 nsew signal input
flabel metal3 s 11192 0 11272 80 0 FreeSans 320 0 0 0 N1END[1]
port 120 nsew signal input
flabel metal3 s 11384 0 11464 80 0 FreeSans 320 0 0 0 N1END[2]
port 121 nsew signal input
flabel metal3 s 11576 0 11656 80 0 FreeSans 320 0 0 0 N1END[3]
port 122 nsew signal input
flabel metal3 s 13304 0 13384 80 0 FreeSans 320 0 0 0 N2END[0]
port 123 nsew signal input
flabel metal3 s 13496 0 13576 80 0 FreeSans 320 0 0 0 N2END[1]
port 124 nsew signal input
flabel metal3 s 13688 0 13768 80 0 FreeSans 320 0 0 0 N2END[2]
port 125 nsew signal input
flabel metal3 s 13880 0 13960 80 0 FreeSans 320 0 0 0 N2END[3]
port 126 nsew signal input
flabel metal3 s 14072 0 14152 80 0 FreeSans 320 0 0 0 N2END[4]
port 127 nsew signal input
flabel metal3 s 14264 0 14344 80 0 FreeSans 320 0 0 0 N2END[5]
port 128 nsew signal input
flabel metal3 s 14456 0 14536 80 0 FreeSans 320 0 0 0 N2END[6]
port 129 nsew signal input
flabel metal3 s 14648 0 14728 80 0 FreeSans 320 0 0 0 N2END[7]
port 130 nsew signal input
flabel metal3 s 11768 0 11848 80 0 FreeSans 320 0 0 0 N2MID[0]
port 131 nsew signal input
flabel metal3 s 11960 0 12040 80 0 FreeSans 320 0 0 0 N2MID[1]
port 132 nsew signal input
flabel metal3 s 12152 0 12232 80 0 FreeSans 320 0 0 0 N2MID[2]
port 133 nsew signal input
flabel metal3 s 12344 0 12424 80 0 FreeSans 320 0 0 0 N2MID[3]
port 134 nsew signal input
flabel metal3 s 12536 0 12616 80 0 FreeSans 320 0 0 0 N2MID[4]
port 135 nsew signal input
flabel metal3 s 12728 0 12808 80 0 FreeSans 320 0 0 0 N2MID[5]
port 136 nsew signal input
flabel metal3 s 12920 0 13000 80 0 FreeSans 320 0 0 0 N2MID[6]
port 137 nsew signal input
flabel metal3 s 13112 0 13192 80 0 FreeSans 320 0 0 0 N2MID[7]
port 138 nsew signal input
flabel metal3 s 14840 0 14920 80 0 FreeSans 320 0 0 0 N4END[0]
port 139 nsew signal input
flabel metal3 s 16760 0 16840 80 0 FreeSans 320 0 0 0 N4END[10]
port 140 nsew signal input
flabel metal3 s 16952 0 17032 80 0 FreeSans 320 0 0 0 N4END[11]
port 141 nsew signal input
flabel metal3 s 17144 0 17224 80 0 FreeSans 320 0 0 0 N4END[12]
port 142 nsew signal input
flabel metal3 s 17336 0 17416 80 0 FreeSans 320 0 0 0 N4END[13]
port 143 nsew signal input
flabel metal3 s 17528 0 17608 80 0 FreeSans 320 0 0 0 N4END[14]
port 144 nsew signal input
flabel metal3 s 17720 0 17800 80 0 FreeSans 320 0 0 0 N4END[15]
port 145 nsew signal input
flabel metal3 s 15032 0 15112 80 0 FreeSans 320 0 0 0 N4END[1]
port 146 nsew signal input
flabel metal3 s 15224 0 15304 80 0 FreeSans 320 0 0 0 N4END[2]
port 147 nsew signal input
flabel metal3 s 15416 0 15496 80 0 FreeSans 320 0 0 0 N4END[3]
port 148 nsew signal input
flabel metal3 s 15608 0 15688 80 0 FreeSans 320 0 0 0 N4END[4]
port 149 nsew signal input
flabel metal3 s 15800 0 15880 80 0 FreeSans 320 0 0 0 N4END[5]
port 150 nsew signal input
flabel metal3 s 15992 0 16072 80 0 FreeSans 320 0 0 0 N4END[6]
port 151 nsew signal input
flabel metal3 s 16184 0 16264 80 0 FreeSans 320 0 0 0 N4END[7]
port 152 nsew signal input
flabel metal3 s 16376 0 16456 80 0 FreeSans 320 0 0 0 N4END[8]
port 153 nsew signal input
flabel metal3 s 16568 0 16648 80 0 FreeSans 320 0 0 0 N4END[9]
port 154 nsew signal input
flabel metal3 s 17912 0 17992 80 0 FreeSans 320 0 0 0 NN4END[0]
port 155 nsew signal input
flabel metal3 s 19832 0 19912 80 0 FreeSans 320 0 0 0 NN4END[10]
port 156 nsew signal input
flabel metal3 s 20024 0 20104 80 0 FreeSans 320 0 0 0 NN4END[11]
port 157 nsew signal input
flabel metal3 s 20216 0 20296 80 0 FreeSans 320 0 0 0 NN4END[12]
port 158 nsew signal input
flabel metal3 s 20408 0 20488 80 0 FreeSans 320 0 0 0 NN4END[13]
port 159 nsew signal input
flabel metal3 s 20600 0 20680 80 0 FreeSans 320 0 0 0 NN4END[14]
port 160 nsew signal input
flabel metal3 s 20792 0 20872 80 0 FreeSans 320 0 0 0 NN4END[15]
port 161 nsew signal input
flabel metal3 s 18104 0 18184 80 0 FreeSans 320 0 0 0 NN4END[1]
port 162 nsew signal input
flabel metal3 s 18296 0 18376 80 0 FreeSans 320 0 0 0 NN4END[2]
port 163 nsew signal input
flabel metal3 s 18488 0 18568 80 0 FreeSans 320 0 0 0 NN4END[3]
port 164 nsew signal input
flabel metal3 s 18680 0 18760 80 0 FreeSans 320 0 0 0 NN4END[4]
port 165 nsew signal input
flabel metal3 s 18872 0 18952 80 0 FreeSans 320 0 0 0 NN4END[5]
port 166 nsew signal input
flabel metal3 s 19064 0 19144 80 0 FreeSans 320 0 0 0 NN4END[6]
port 167 nsew signal input
flabel metal3 s 19256 0 19336 80 0 FreeSans 320 0 0 0 NN4END[7]
port 168 nsew signal input
flabel metal3 s 19448 0 19528 80 0 FreeSans 320 0 0 0 NN4END[8]
port 169 nsew signal input
flabel metal3 s 19640 0 19720 80 0 FreeSans 320 0 0 0 NN4END[9]
port 170 nsew signal input
flabel metal3 s 21176 0 21256 80 0 FreeSans 320 0 0 0 S1BEG[0]
port 171 nsew signal output
flabel metal3 s 21368 0 21448 80 0 FreeSans 320 0 0 0 S1BEG[1]
port 172 nsew signal output
flabel metal3 s 21560 0 21640 80 0 FreeSans 320 0 0 0 S1BEG[2]
port 173 nsew signal output
flabel metal3 s 21752 0 21832 80 0 FreeSans 320 0 0 0 S1BEG[3]
port 174 nsew signal output
flabel metal3 s 21944 0 22024 80 0 FreeSans 320 0 0 0 S2BEG[0]
port 175 nsew signal output
flabel metal3 s 22136 0 22216 80 0 FreeSans 320 0 0 0 S2BEG[1]
port 176 nsew signal output
flabel metal3 s 22328 0 22408 80 0 FreeSans 320 0 0 0 S2BEG[2]
port 177 nsew signal output
flabel metal3 s 22520 0 22600 80 0 FreeSans 320 0 0 0 S2BEG[3]
port 178 nsew signal output
flabel metal3 s 22712 0 22792 80 0 FreeSans 320 0 0 0 S2BEG[4]
port 179 nsew signal output
flabel metal3 s 22904 0 22984 80 0 FreeSans 320 0 0 0 S2BEG[5]
port 180 nsew signal output
flabel metal3 s 23096 0 23176 80 0 FreeSans 320 0 0 0 S2BEG[6]
port 181 nsew signal output
flabel metal3 s 23288 0 23368 80 0 FreeSans 320 0 0 0 S2BEG[7]
port 182 nsew signal output
flabel metal3 s 23480 0 23560 80 0 FreeSans 320 0 0 0 S2BEGb[0]
port 183 nsew signal output
flabel metal3 s 23672 0 23752 80 0 FreeSans 320 0 0 0 S2BEGb[1]
port 184 nsew signal output
flabel metal3 s 23864 0 23944 80 0 FreeSans 320 0 0 0 S2BEGb[2]
port 185 nsew signal output
flabel metal3 s 24056 0 24136 80 0 FreeSans 320 0 0 0 S2BEGb[3]
port 186 nsew signal output
flabel metal3 s 24248 0 24328 80 0 FreeSans 320 0 0 0 S2BEGb[4]
port 187 nsew signal output
flabel metal3 s 24440 0 24520 80 0 FreeSans 320 0 0 0 S2BEGb[5]
port 188 nsew signal output
flabel metal3 s 24632 0 24712 80 0 FreeSans 320 0 0 0 S2BEGb[6]
port 189 nsew signal output
flabel metal3 s 24824 0 24904 80 0 FreeSans 320 0 0 0 S2BEGb[7]
port 190 nsew signal output
flabel metal3 s 25016 0 25096 80 0 FreeSans 320 0 0 0 S4BEG[0]
port 191 nsew signal output
flabel metal3 s 26936 0 27016 80 0 FreeSans 320 0 0 0 S4BEG[10]
port 192 nsew signal output
flabel metal3 s 27128 0 27208 80 0 FreeSans 320 0 0 0 S4BEG[11]
port 193 nsew signal output
flabel metal3 s 27320 0 27400 80 0 FreeSans 320 0 0 0 S4BEG[12]
port 194 nsew signal output
flabel metal3 s 27512 0 27592 80 0 FreeSans 320 0 0 0 S4BEG[13]
port 195 nsew signal output
flabel metal3 s 27704 0 27784 80 0 FreeSans 320 0 0 0 S4BEG[14]
port 196 nsew signal output
flabel metal3 s 27896 0 27976 80 0 FreeSans 320 0 0 0 S4BEG[15]
port 197 nsew signal output
flabel metal3 s 25208 0 25288 80 0 FreeSans 320 0 0 0 S4BEG[1]
port 198 nsew signal output
flabel metal3 s 25400 0 25480 80 0 FreeSans 320 0 0 0 S4BEG[2]
port 199 nsew signal output
flabel metal3 s 25592 0 25672 80 0 FreeSans 320 0 0 0 S4BEG[3]
port 200 nsew signal output
flabel metal3 s 25784 0 25864 80 0 FreeSans 320 0 0 0 S4BEG[4]
port 201 nsew signal output
flabel metal3 s 25976 0 26056 80 0 FreeSans 320 0 0 0 S4BEG[5]
port 202 nsew signal output
flabel metal3 s 26168 0 26248 80 0 FreeSans 320 0 0 0 S4BEG[6]
port 203 nsew signal output
flabel metal3 s 26360 0 26440 80 0 FreeSans 320 0 0 0 S4BEG[7]
port 204 nsew signal output
flabel metal3 s 26552 0 26632 80 0 FreeSans 320 0 0 0 S4BEG[8]
port 205 nsew signal output
flabel metal3 s 26744 0 26824 80 0 FreeSans 320 0 0 0 S4BEG[9]
port 206 nsew signal output
flabel metal3 s 28088 0 28168 80 0 FreeSans 320 0 0 0 SS4BEG[0]
port 207 nsew signal output
flabel metal3 s 30008 0 30088 80 0 FreeSans 320 0 0 0 SS4BEG[10]
port 208 nsew signal output
flabel metal3 s 30200 0 30280 80 0 FreeSans 320 0 0 0 SS4BEG[11]
port 209 nsew signal output
flabel metal3 s 30392 0 30472 80 0 FreeSans 320 0 0 0 SS4BEG[12]
port 210 nsew signal output
flabel metal3 s 30584 0 30664 80 0 FreeSans 320 0 0 0 SS4BEG[13]
port 211 nsew signal output
flabel metal3 s 30776 0 30856 80 0 FreeSans 320 0 0 0 SS4BEG[14]
port 212 nsew signal output
flabel metal3 s 30968 0 31048 80 0 FreeSans 320 0 0 0 SS4BEG[15]
port 213 nsew signal output
flabel metal3 s 28280 0 28360 80 0 FreeSans 320 0 0 0 SS4BEG[1]
port 214 nsew signal output
flabel metal3 s 28472 0 28552 80 0 FreeSans 320 0 0 0 SS4BEG[2]
port 215 nsew signal output
flabel metal3 s 28664 0 28744 80 0 FreeSans 320 0 0 0 SS4BEG[3]
port 216 nsew signal output
flabel metal3 s 28856 0 28936 80 0 FreeSans 320 0 0 0 SS4BEG[4]
port 217 nsew signal output
flabel metal3 s 29048 0 29128 80 0 FreeSans 320 0 0 0 SS4BEG[5]
port 218 nsew signal output
flabel metal3 s 29240 0 29320 80 0 FreeSans 320 0 0 0 SS4BEG[6]
port 219 nsew signal output
flabel metal3 s 29432 0 29512 80 0 FreeSans 320 0 0 0 SS4BEG[7]
port 220 nsew signal output
flabel metal3 s 29624 0 29704 80 0 FreeSans 320 0 0 0 SS4BEG[8]
port 221 nsew signal output
flabel metal3 s 29816 0 29896 80 0 FreeSans 320 0 0 0 SS4BEG[9]
port 222 nsew signal output
flabel metal3 s 31160 0 31240 80 0 FreeSans 320 0 0 0 UserCLK
port 223 nsew signal input
flabel metal3 s 19640 12100 19720 12180 0 FreeSans 320 0 0 0 UserCLKo
port 224 nsew signal output
flabel metal5 s 4892 0 5332 12180 0 FreeSans 2560 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal5 s 4892 0 5332 40 0 FreeSans 320 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal5 s 4892 12140 5332 12180 0 FreeSans 320 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal5 s 20012 0 20452 12180 0 FreeSans 2560 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal5 s 20012 0 20452 40 0 FreeSans 320 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal5 s 20012 12140 20452 12180 0 FreeSans 320 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal5 s 35132 0 35572 12180 0 FreeSans 2560 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal5 s 35132 0 35572 40 0 FreeSans 320 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal5 s 35132 12140 35572 12180 0 FreeSans 320 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal5 s 3652 0 4092 12180 0 FreeSans 2560 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal5 s 3652 0 4092 40 0 FreeSans 320 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal5 s 3652 12140 4092 12180 0 FreeSans 320 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal5 s 18772 0 19212 12180 0 FreeSans 2560 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal5 s 18772 0 19212 40 0 FreeSans 320 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal5 s 18772 12140 19212 12180 0 FreeSans 320 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal5 s 33892 0 34332 12180 0 FreeSans 2560 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal5 s 33892 0 34332 40 0 FreeSans 320 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal5 s 33892 12140 34332 12180 0 FreeSans 320 0 0 0 VPWR
port 226 nsew power bidirectional
rlabel metal1 23184 10584 23184 10584 0 VGND
rlabel metal1 23184 9828 23184 9828 0 VPWR
rlabel metal2 5016 10416 5016 10416 0 A_I_top
rlabel metal3 3552 11142 3552 11142 0 A_O_top
rlabel metal2 5880 10416 5880 10416 0 A_T_top
rlabel metal2 9816 10416 9816 10416 0 A_config_C_bit0
rlabel metal2 11496 10416 11496 10416 0 A_config_C_bit1
rlabel metal2 12264 10416 12264 10416 0 A_config_C_bit2
rlabel metal2 13944 9660 13944 9660 0 A_config_C_bit3
rlabel metal2 8136 10416 8136 10416 0 B_I_top
rlabel metal3 7008 11142 7008 11142 0 B_O_top
rlabel metal2 9048 10332 9048 10332 0 B_T_top
rlabel metal2 14952 9660 14952 9660 0 B_config_C_bit0
rlabel metal2 16488 10416 16488 10416 0 B_config_C_bit1
rlabel metal2 17400 10416 17400 10416 0 B_config_C_bit2
rlabel metal2 18360 9660 18360 9660 0 B_config_C_bit3
rlabel metal2 608 756 608 756 0 FrameData[0]
rlabel metal2 656 4116 656 4116 0 FrameData[10]
rlabel metal2 128 4452 128 4452 0 FrameData[11]
rlabel via2 80 4788 80 4788 0 FrameData[12]
rlabel metal2 464 5124 464 5124 0 FrameData[13]
rlabel via2 80 5460 80 5460 0 FrameData[14]
rlabel metal2 128 5796 128 5796 0 FrameData[15]
rlabel metal2 80 6132 80 6132 0 FrameData[16]
rlabel metal2 656 6468 656 6468 0 FrameData[17]
rlabel metal2 128 6804 128 6804 0 FrameData[18]
rlabel metal2 656 7140 656 7140 0 FrameData[19]
rlabel metal2 752 1092 752 1092 0 FrameData[1]
rlabel metal2 656 7476 656 7476 0 FrameData[20]
rlabel metal2 848 7812 848 7812 0 FrameData[21]
rlabel metal2 656 8148 656 8148 0 FrameData[22]
rlabel metal2 464 8484 464 8484 0 FrameData[23]
rlabel metal2 656 8820 656 8820 0 FrameData[24]
rlabel metal2 128 9156 128 9156 0 FrameData[25]
rlabel metal2 368 9492 368 9492 0 FrameData[26]
rlabel metal2 848 9828 848 9828 0 FrameData[27]
rlabel metal2 560 10164 560 10164 0 FrameData[28]
rlabel metal2 1232 10500 1232 10500 0 FrameData[29]
rlabel metal2 368 1428 368 1428 0 FrameData[2]
rlabel metal2 704 10836 704 10836 0 FrameData[30]
rlabel via2 80 11172 80 11172 0 FrameData[31]
rlabel metal2 320 1764 320 1764 0 FrameData[3]
rlabel metal2 128 2100 128 2100 0 FrameData[4]
rlabel metal2 656 2436 656 2436 0 FrameData[5]
rlabel metal2 1040 2772 1040 2772 0 FrameData[6]
rlabel metal2 896 3108 896 3108 0 FrameData[7]
rlabel metal2 656 3444 656 3444 0 FrameData[8]
rlabel metal2 128 3780 128 3780 0 FrameData[9]
rlabel metal2 45855 756 45855 756 0 FrameData_O[0]
rlabel metal2 45999 4116 45999 4116 0 FrameData_O[10]
rlabel metal2 45168 4368 45168 4368 0 FrameData_O[11]
rlabel metal2 45543 4788 45543 4788 0 FrameData_O[12]
rlabel metal2 45735 5124 45735 5124 0 FrameData_O[13]
rlabel metal2 45951 5460 45951 5460 0 FrameData_O[14]
rlabel metal2 45735 5796 45735 5796 0 FrameData_O[15]
rlabel metal2 45543 6132 45543 6132 0 FrameData_O[16]
rlabel metal2 45735 6468 45735 6468 0 FrameData_O[17]
rlabel via2 46287 6804 46287 6804 0 FrameData_O[18]
rlabel metal2 45735 7140 45735 7140 0 FrameData_O[19]
rlabel metal2 45471 1092 45471 1092 0 FrameData_O[1]
rlabel via2 46287 7476 46287 7476 0 FrameData_O[20]
rlabel metal2 45543 7812 45543 7812 0 FrameData_O[21]
rlabel via2 46287 8148 46287 8148 0 FrameData_O[22]
rlabel metal2 45807 8484 45807 8484 0 FrameData_O[23]
rlabel metal2 44679 8820 44679 8820 0 FrameData_O[24]
rlabel metal2 44424 7056 44424 7056 0 FrameData_O[25]
rlabel metal2 43656 8148 43656 8148 0 FrameData_O[26]
rlabel metal2 44424 7392 44424 7392 0 FrameData_O[27]
rlabel metal2 43080 8148 43080 8148 0 FrameData_O[28]
rlabel metal2 44328 6636 44328 6636 0 FrameData_O[29]
rlabel metal2 45807 1428 45807 1428 0 FrameData_O[2]
rlabel metal2 43752 7056 43752 7056 0 FrameData_O[30]
rlabel metal2 42600 8148 42600 8148 0 FrameData_O[31]
rlabel metal2 45543 1764 45543 1764 0 FrameData_O[3]
rlabel metal2 45735 2100 45735 2100 0 FrameData_O[4]
rlabel metal2 46047 2436 46047 2436 0 FrameData_O[5]
rlabel metal2 45735 2772 45735 2772 0 FrameData_O[6]
rlabel metal2 45543 3108 45543 3108 0 FrameData_O[7]
rlabel metal2 45855 3444 45855 3444 0 FrameData_O[8]
rlabel metal2 45168 3696 45168 3696 0 FrameData_O[9]
rlabel metal3 28800 6258 28800 6258 0 FrameStrobe[0]
rlabel metal3 43104 9282 43104 9282 0 FrameStrobe[10]
rlabel via2 33504 72 33504 72 0 FrameStrobe[11]
rlabel metal3 33696 408 33696 408 0 FrameStrobe[12]
rlabel metal3 33888 366 33888 366 0 FrameStrobe[13]
rlabel metal3 34080 744 34080 744 0 FrameStrobe[14]
rlabel metal3 34272 702 34272 702 0 FrameStrobe[15]
rlabel metal5 34464 3612 34464 3612 0 FrameStrobe[16]
rlabel metal2 38976 11592 38976 11592 0 FrameStrobe[17]
rlabel metal3 44736 10794 44736 10794 0 FrameStrobe[18]
rlabel metal3 34992 9576 34992 9576 0 FrameStrobe[19]
rlabel metal3 36768 1974 36768 1974 0 FrameStrobe[1]
rlabel metal2 21984 6468 21984 6468 0 FrameStrobe[2]
rlabel metal3 33792 6510 33792 6510 0 FrameStrobe[3]
rlabel metal3 34656 9870 34656 9870 0 FrameStrobe[4]
rlabel metal3 33312 9030 33312 9030 0 FrameStrobe[5]
rlabel metal3 32544 4440 32544 4440 0 FrameStrobe[6]
rlabel metal2 39072 11298 39072 11298 0 FrameStrobe[7]
rlabel metal3 42912 4830 42912 4830 0 FrameStrobe[8]
rlabel metal3 42768 10248 42768 10248 0 FrameStrobe[9]
rlabel metal2 20808 9660 20808 9660 0 FrameStrobe_O[0]
rlabel metal3 32352 10890 32352 10890 0 FrameStrobe_O[10]
rlabel metal2 33720 9660 33720 9660 0 FrameStrobe_O[11]
rlabel metal2 34680 10416 34680 10416 0 FrameStrobe_O[12]
rlabel metal2 36312 10416 36312 10416 0 FrameStrobe_O[13]
rlabel metal2 37272 10416 37272 10416 0 FrameStrobe_O[14]
rlabel metal2 38136 10416 38136 10416 0 FrameStrobe_O[15]
rlabel metal2 39048 10416 39048 10416 0 FrameStrobe_O[16]
rlabel metal2 41304 10332 41304 10332 0 FrameStrobe_O[17]
rlabel metal2 42072 10416 42072 10416 0 FrameStrobe_O[18]
rlabel metal2 42840 10416 42840 10416 0 FrameStrobe_O[19]
rlabel metal2 21720 9576 21720 9576 0 FrameStrobe_O[1]
rlabel metal2 23160 8148 23160 8148 0 FrameStrobe_O[2]
rlabel metal2 24168 10416 24168 10416 0 FrameStrobe_O[3]
rlabel metal2 25848 9660 25848 9660 0 FrameStrobe_O[4]
rlabel metal2 27000 10416 27000 10416 0 FrameStrobe_O[5]
rlabel metal2 27768 10416 27768 10416 0 FrameStrobe_O[6]
rlabel metal2 29400 10416 29400 10416 0 FrameStrobe_O[7]
rlabel metal2 31176 10416 31176 10416 0 FrameStrobe_O[8]
rlabel metal2 31944 10332 31944 10332 0 FrameStrobe_O[9]
rlabel metal3 41376 9030 41376 9030 0 Inst_A_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 35616 1932 35616 1932 0 Inst_B_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 10464 2856 10464 2856 0 Inst_N_IO_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 10992 2772 10992 2772 0 Inst_N_IO_ConfigMem.Inst_frame0_bit1.Q
rlabel via1 34558 9408 34558 9408 0 Inst_N_IO_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 36408 9408 36408 9408 0 Inst_N_IO_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 30288 7392 30288 7392 0 Inst_N_IO_ConfigMem.Inst_frame0_bit12.Q
rlabel metal3 31968 7644 31968 7644 0 Inst_N_IO_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 14280 4872 14280 4872 0 Inst_N_IO_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 13056 4998 13056 4998 0 Inst_N_IO_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 13560 3360 13560 3360 0 Inst_N_IO_ConfigMem.Inst_frame0_bit16.Q
rlabel metal3 12096 2688 12096 2688 0 Inst_N_IO_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 9696 4914 9696 4914 0 Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 11192 4872 11192 4872 0 Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 35520 4200 35520 4200 0 Inst_N_IO_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 9168 2772 9168 2772 0 Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 10032 1764 10032 1764 0 Inst_N_IO_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 8016 7938 8016 7938 0 Inst_N_IO_ConfigMem.Inst_frame0_bit22.Q
rlabel via1 7217 10248 7217 10248 0 Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q
rlabel via1 7787 9408 7787 9408 0 Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 4944 5880 4944 5880 0 Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 5808 4872 5808 4872 0 Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q
rlabel metal3 7296 5880 7296 5880 0 Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q
rlabel metal3 5664 5418 5664 5418 0 Inst_N_IO_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 7056 2520 7056 2520 0 Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 33696 3612 33696 3612 0 Inst_N_IO_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 6240 3360 6240 3360 0 Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 6261 2688 6261 2688 0 Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q
rlabel metal3 34464 8400 34464 8400 0 Inst_N_IO_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 36096 8736 36096 8736 0 Inst_N_IO_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 30624 5754 30624 5754 0 Inst_N_IO_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 32160 5754 32160 5754 0 Inst_N_IO_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 34080 2646 34080 2646 0 Inst_N_IO_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 35760 3024 35760 3024 0 Inst_N_IO_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 15216 2100 15216 2100 0 Inst_N_IO_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 17040 3192 17040 3192 0 Inst_N_IO_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 41760 8736 41760 8736 0 Inst_N_IO_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 40320 8694 40320 8694 0 Inst_N_IO_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 35520 5712 35520 5712 0 Inst_N_IO_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 33934 5124 33934 5124 0 Inst_N_IO_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 24336 8904 24336 8904 0 Inst_N_IO_ConfigMem.Inst_frame1_bit14.Q
rlabel via2 25928 9408 25928 9408 0 Inst_N_IO_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 30384 2772 30384 2772 0 Inst_N_IO_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 31920 2688 31920 2688 0 Inst_N_IO_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 25248 5712 25248 5712 0 Inst_N_IO_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 27072 5124 27072 5124 0 Inst_N_IO_ConfigMem.Inst_frame1_bit19.Q
rlabel metal3 40416 6888 40416 6888 0 Inst_N_IO_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 28128 2730 28128 2730 0 Inst_N_IO_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 29280 2100 29280 2100 0 Inst_N_IO_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 27360 9450 27360 9450 0 Inst_N_IO_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 29112 9408 29112 9408 0 Inst_N_IO_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 29904 8736 29904 8736 0 Inst_N_IO_ConfigMem.Inst_frame1_bit24.Q
rlabel metal3 31584 6930 31584 6930 0 Inst_N_IO_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 6776 7876 6776 7876 0 Inst_N_IO_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 3984 7056 3984 7056 0 Inst_N_IO_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 4032 5544 4032 5544 0 Inst_N_IO_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 6408 6384 6408 6384 0 Inst_N_IO_ConfigMem.Inst_frame1_bit29.Q
rlabel metal3 41856 7476 41856 7476 0 Inst_N_IO_ConfigMem.Inst_frame1_bit3.Q
rlabel metal3 9120 6510 9120 6510 0 Inst_N_IO_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 7584 4116 7584 4116 0 Inst_N_IO_ConfigMem.Inst_frame1_bit31.Q
rlabel metal3 37920 4578 37920 4578 0 Inst_N_IO_ConfigMem.Inst_frame1_bit4.Q
rlabel via1 38984 4872 38984 4872 0 Inst_N_IO_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 33264 8904 33264 8904 0 Inst_N_IO_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 31296 9366 31296 9366 0 Inst_N_IO_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 36168 1848 36168 1848 0 Inst_N_IO_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 34272 1890 34272 1890 0 Inst_N_IO_ConfigMem.Inst_frame1_bit9.Q
rlabel metal4 18144 2646 18144 2646 0 Inst_N_IO_ConfigMem.Inst_frame2_bit0.Q
rlabel metal4 25056 3192 25056 3192 0 Inst_N_IO_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 17760 8904 17760 8904 0 Inst_N_IO_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 20040 9408 20040 9408 0 Inst_N_IO_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 15072 5712 15072 5712 0 Inst_N_IO_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 20856 5544 20856 5544 0 Inst_N_IO_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 12672 8988 12672 8988 0 Inst_N_IO_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 13224 9408 13224 9408 0 Inst_N_IO_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 24816 1848 24816 1848 0 Inst_N_IO_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 26408 1848 26408 1848 0 Inst_N_IO_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 21984 7371 21984 7371 0 Inst_N_IO_ConfigMem.Inst_frame2_bit18.Q
rlabel metal3 23520 6930 23520 6930 0 Inst_N_IO_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 19584 7266 19584 7266 0 Inst_N_IO_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 21696 2856 21696 2856 0 Inst_N_IO_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 23040 2142 23040 2142 0 Inst_N_IO_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 23304 9408 23304 9408 0 Inst_N_IO_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 21696 8946 21696 8946 0 Inst_N_IO_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 20328 4872 20328 4872 0 Inst_N_IO_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 18672 4872 18672 4872 0 Inst_N_IO_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 17616 6636 17616 6636 0 Inst_N_IO_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 17568 7182 17568 7182 0 Inst_N_IO_ConfigMem.Inst_frame2_bit27.Q
rlabel metal3 18240 4704 18240 4704 0 Inst_N_IO_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 18624 4242 18624 4242 0 Inst_N_IO_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 21312 7224 21312 7224 0 Inst_N_IO_ConfigMem.Inst_frame2_bit3.Q
rlabel metal2 17568 8736 17568 8736 0 Inst_N_IO_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 19248 8736 19248 8736 0 Inst_N_IO_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 25776 3528 25776 3528 0 Inst_N_IO_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 22440 4200 22440 4200 0 Inst_N_IO_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 38016 7938 38016 7938 0 Inst_N_IO_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 39720 7896 39720 7896 0 Inst_N_IO_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 34560 3150 34560 3150 0 Inst_N_IO_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 32496 3612 32496 3612 0 Inst_N_IO_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 22320 4872 22320 4872 0 Inst_N_IO_ConfigMem.Inst_frame3_bit14.Q
rlabel metal2 25776 7896 25776 7896 0 Inst_N_IO_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 40464 2772 40464 2772 0 Inst_N_IO_ConfigMem.Inst_frame3_bit16.Q
rlabel metal3 36096 5964 36096 5964 0 Inst_N_IO_ConfigMem.Inst_frame3_bit17.Q
rlabel metal2 18048 6426 18048 6426 0 Inst_N_IO_ConfigMem.Inst_frame3_bit18.Q
rlabel metal3 19680 6678 19680 6678 0 Inst_N_IO_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 18528 2100 18528 2100 0 Inst_N_IO_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 20112 2688 20112 2688 0 Inst_N_IO_ConfigMem.Inst_frame3_bit21.Q
rlabel metal2 26832 7896 26832 7896 0 Inst_N_IO_ConfigMem.Inst_frame3_bit22.Q
rlabel via2 28520 7896 28520 7896 0 Inst_N_IO_ConfigMem.Inst_frame3_bit23.Q
rlabel metal3 28128 4620 28128 4620 0 Inst_N_IO_ConfigMem.Inst_frame3_bit24.Q
rlabel metal3 30048 4620 30048 4620 0 Inst_N_IO_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 15009 9408 15009 9408 0 Inst_N_IO_ConfigMem.Inst_frame3_bit26.Q
rlabel via2 16616 9408 16616 9408 0 Inst_N_IO_ConfigMem.Inst_frame3_bit27.Q
rlabel metal3 14688 4620 14688 4620 0 Inst_N_IO_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 16376 4872 16376 4872 0 Inst_N_IO_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 10752 8778 10752 8778 0 Inst_N_IO_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 12288 8778 12288 8778 0 Inst_N_IO_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 23328 4956 23328 4956 0 Inst_N_IO_switch_matrix.S1BEG0
rlabel metal3 26208 7602 26208 7602 0 Inst_N_IO_switch_matrix.S1BEG1
rlabel metal2 41856 3486 41856 3486 0 Inst_N_IO_switch_matrix.S1BEG2
rlabel metal2 38784 5586 38784 5586 0 Inst_N_IO_switch_matrix.S1BEG3
rlabel metal2 19896 6468 19896 6468 0 Inst_N_IO_switch_matrix.S2BEG0
rlabel metal2 19584 2856 19584 2856 0 Inst_N_IO_switch_matrix.S2BEG1
rlabel metal2 28920 7980 28920 7980 0 Inst_N_IO_switch_matrix.S2BEG2
rlabel metal2 30168 5124 30168 5124 0 Inst_N_IO_switch_matrix.S2BEG3
rlabel metal3 16992 9366 16992 9366 0 Inst_N_IO_switch_matrix.S2BEG4
rlabel metal3 16608 5586 16608 5586 0 Inst_N_IO_switch_matrix.S2BEG5
rlabel metal3 12480 8442 12480 8442 0 Inst_N_IO_switch_matrix.S2BEG6
rlabel metal2 26256 2856 26256 2856 0 Inst_N_IO_switch_matrix.S2BEG7
rlabel metal2 21432 7140 21432 7140 0 Inst_N_IO_switch_matrix.S2BEGb0
rlabel metal2 23328 4158 23328 4158 0 Inst_N_IO_switch_matrix.S2BEGb1
rlabel metal2 41712 7980 41712 7980 0 Inst_N_IO_switch_matrix.S2BEGb2
rlabel metal2 36288 4200 36288 4200 0 Inst_N_IO_switch_matrix.S2BEGb3
rlabel metal2 20280 9492 20280 9492 0 Inst_N_IO_switch_matrix.S2BEGb4
rlabel metal3 17088 6174 17088 6174 0 Inst_N_IO_switch_matrix.S2BEGb5
rlabel metal2 13368 9492 13368 9492 0 Inst_N_IO_switch_matrix.S2BEGb6
rlabel metal2 27000 2100 27000 2100 0 Inst_N_IO_switch_matrix.S2BEGb7
rlabel metal3 23808 7686 23808 7686 0 Inst_N_IO_switch_matrix.S4BEG0
rlabel metal2 23472 2856 23472 2856 0 Inst_N_IO_switch_matrix.S4BEG1
rlabel metal2 33792 9408 33792 9408 0 Inst_N_IO_switch_matrix.S4BEG10
rlabel metal2 37128 2100 37128 2100 0 Inst_N_IO_switch_matrix.S4BEG11
rlabel metal2 42264 8652 42264 8652 0 Inst_N_IO_switch_matrix.S4BEG12
rlabel metal2 35664 5880 35664 5880 0 Inst_N_IO_switch_matrix.S4BEG13
rlabel metal2 26736 9408 26736 9408 0 Inst_N_IO_switch_matrix.S4BEG14
rlabel metal4 34464 2856 34464 2856 0 Inst_N_IO_switch_matrix.S4BEG15
rlabel metal2 23544 9492 23544 9492 0 Inst_N_IO_switch_matrix.S4BEG2
rlabel metal2 20520 4872 20520 4872 0 Inst_N_IO_switch_matrix.S4BEG3
rlabel metal3 19776 7686 19776 7686 0 Inst_N_IO_switch_matrix.S4BEG4
rlabel metal2 20328 3948 20328 3948 0 Inst_N_IO_switch_matrix.S4BEG5
rlabel metal3 19488 9534 19488 9534 0 Inst_N_IO_switch_matrix.S4BEG6
rlabel metal2 18288 2772 18288 2772 0 Inst_N_IO_switch_matrix.S4BEG7
rlabel metal2 42264 7140 42264 7140 0 Inst_N_IO_switch_matrix.S4BEG8
rlabel metal2 39384 4956 39384 4956 0 Inst_N_IO_switch_matrix.S4BEG9
rlabel metal2 27936 5586 27936 5586 0 Inst_N_IO_switch_matrix.SS4BEG0
rlabel metal2 30864 2856 30864 2856 0 Inst_N_IO_switch_matrix.SS4BEG1
rlabel metal2 32544 5586 32544 5586 0 Inst_N_IO_switch_matrix.SS4BEG10
rlabel metal2 36624 2856 36624 2856 0 Inst_N_IO_switch_matrix.SS4BEG11
rlabel metal3 36288 9660 36288 9660 0 Inst_N_IO_switch_matrix.SS4BEG12
rlabel metal2 32184 7980 32184 7980 0 Inst_N_IO_switch_matrix.SS4BEG13
rlabel metal2 12336 4956 12336 4956 0 Inst_N_IO_switch_matrix.SS4BEG14
rlabel metal3 13536 5586 13536 5586 0 Inst_N_IO_switch_matrix.SS4BEG15
rlabel metal2 29112 8652 29112 8652 0 Inst_N_IO_switch_matrix.SS4BEG2
rlabel metal2 32304 8904 32304 8904 0 Inst_N_IO_switch_matrix.SS4BEG3
rlabel metal2 8640 7980 8640 7980 0 Inst_N_IO_switch_matrix.SS4BEG4
rlabel metal2 6360 6636 6360 6636 0 Inst_N_IO_switch_matrix.SS4BEG5
rlabel metal2 6288 4956 6288 4956 0 Inst_N_IO_switch_matrix.SS4BEG6
rlabel metal3 9696 4452 9696 4452 0 Inst_N_IO_switch_matrix.SS4BEG7
rlabel metal2 38304 4074 38304 4074 0 Inst_N_IO_switch_matrix.SS4BEG8
rlabel metal2 36312 8652 36312 8652 0 Inst_N_IO_switch_matrix.SS4BEG9
rlabel metal3 11040 1470 11040 1470 0 N1END[0]
rlabel metal2 7824 3780 7824 3780 0 N1END[1]
rlabel metal3 11424 1332 11424 1332 0 N1END[2]
rlabel metal3 2784 1008 2784 1008 0 N1END[3]
rlabel metal3 13344 660 13344 660 0 N2END[0]
rlabel metal3 13824 5418 13824 5418 0 N2END[1]
rlabel metal3 13728 744 13728 744 0 N2END[2]
rlabel metal2 10224 5628 10224 5628 0 N2END[3]
rlabel metal2 13440 5586 13440 5586 0 N2END[4]
rlabel metal3 14304 744 14304 744 0 N2END[5]
rlabel metal3 14496 156 14496 156 0 N2END[6]
rlabel metal3 14688 1794 14688 1794 0 N2END[7]
rlabel metal3 11808 324 11808 324 0 N2MID[0]
rlabel metal3 12000 1122 12000 1122 0 N2MID[1]
rlabel metal3 12192 744 12192 744 0 N2MID[2]
rlabel metal3 12384 1248 12384 1248 0 N2MID[3]
rlabel metal3 12576 1206 12576 1206 0 N2MID[4]
rlabel metal2 9360 2856 9360 2856 0 N2MID[5]
rlabel metal3 13248 1302 13248 1302 0 N2MID[6]
rlabel metal3 13152 156 13152 156 0 N2MID[7]
rlabel metal3 14880 744 14880 744 0 N4END[0]
rlabel metal2 16368 7812 16368 7812 0 N4END[10]
rlabel metal3 16992 744 16992 744 0 N4END[11]
rlabel metal3 17184 744 17184 744 0 N4END[12]
rlabel metal3 17376 1080 17376 1080 0 N4END[13]
rlabel metal3 17568 912 17568 912 0 N4END[14]
rlabel metal3 17760 702 17760 702 0 N4END[15]
rlabel metal3 15072 534 15072 534 0 N4END[1]
rlabel metal2 14976 8148 14976 8148 0 N4END[2]
rlabel metal3 15456 828 15456 828 0 N4END[3]
rlabel metal2 15360 7812 15360 7812 0 N4END[4]
rlabel metal3 15840 996 15840 996 0 N4END[5]
rlabel metal2 15936 7728 15936 7728 0 N4END[6]
rlabel metal3 16224 450 16224 450 0 N4END[7]
rlabel metal3 16416 2634 16416 2634 0 N4END[8]
rlabel metal3 16608 1416 16608 1416 0 N4END[9]
rlabel metal3 17952 1470 17952 1470 0 NN4END[0]
rlabel metal2 20544 6426 20544 6426 0 NN4END[10]
rlabel metal3 20064 534 20064 534 0 NN4END[11]
rlabel metal3 20256 702 20256 702 0 NN4END[12]
rlabel metal3 20448 702 20448 702 0 NN4END[13]
rlabel metal4 19296 4032 19296 4032 0 NN4END[14]
rlabel metal3 20832 912 20832 912 0 NN4END[15]
rlabel metal3 18192 5460 18192 5460 0 NN4END[1]
rlabel metal3 18336 660 18336 660 0 NN4END[2]
rlabel metal3 18528 576 18528 576 0 NN4END[3]
rlabel metal3 18720 1584 18720 1584 0 NN4END[4]
rlabel metal3 18912 660 18912 660 0 NN4END[5]
rlabel metal3 19104 324 19104 324 0 NN4END[6]
rlabel metal3 19296 576 19296 576 0 NN4END[7]
rlabel metal2 17280 3948 17280 3948 0 NN4END[8]
rlabel metal5 19680 4452 19680 4452 0 NN4END[9]
rlabel metal3 21216 828 21216 828 0 S1BEG[0]
rlabel metal3 21408 1206 21408 1206 0 S1BEG[1]
rlabel metal3 21600 702 21600 702 0 S1BEG[2]
rlabel metal3 21792 660 21792 660 0 S1BEG[3]
rlabel metal3 21984 744 21984 744 0 S2BEG[0]
rlabel metal2 21840 3024 21840 3024 0 S2BEG[1]
rlabel metal3 22368 744 22368 744 0 S2BEG[2]
rlabel metal2 22080 3108 22080 3108 0 S2BEG[3]
rlabel metal3 22752 1290 22752 1290 0 S2BEG[4]
rlabel metal3 22944 1248 22944 1248 0 S2BEG[5]
rlabel metal2 22464 2058 22464 2058 0 S2BEG[6]
rlabel metal2 21312 1638 21312 1638 0 S2BEG[7]
rlabel metal2 23544 3948 23544 3948 0 S2BEGb[0]
rlabel metal3 23712 870 23712 870 0 S2BEGb[1]
rlabel metal2 23928 3948 23928 3948 0 S2BEGb[2]
rlabel metal3 24096 1206 24096 1206 0 S2BEGb[3]
rlabel metal2 24312 3192 24312 3192 0 S2BEGb[4]
rlabel metal3 24480 1248 24480 1248 0 S2BEGb[5]
rlabel metal3 24672 828 24672 828 0 S2BEGb[6]
rlabel metal3 24864 786 24864 786 0 S2BEGb[7]
rlabel metal2 25248 3864 25248 3864 0 S4BEG[0]
rlabel metal3 26976 450 26976 450 0 S4BEG[10]
rlabel metal2 28680 3948 28680 3948 0 S4BEG[11]
rlabel metal2 32448 1554 32448 1554 0 S4BEG[12]
rlabel metal3 27552 534 27552 534 0 S4BEG[13]
rlabel metal3 33216 1260 33216 1260 0 S4BEG[14]
rlabel metal2 28560 5292 28560 5292 0 S4BEG[15]
rlabel metal2 25584 3780 25584 3780 0 S4BEG[1]
rlabel metal3 25440 1038 25440 1038 0 S4BEG[2]
rlabel metal3 25632 744 25632 744 0 S4BEG[3]
rlabel metal3 25824 828 25824 828 0 S4BEG[4]
rlabel metal2 26568 4704 26568 4704 0 S4BEG[5]
rlabel metal2 26736 4620 26736 4620 0 S4BEG[6]
rlabel metal2 26736 4368 26736 4368 0 S4BEG[7]
rlabel metal3 26592 366 26592 366 0 S4BEG[8]
rlabel metal4 27600 5460 27600 5460 0 S4BEG[9]
rlabel metal3 33504 1302 33504 1302 0 SS4BEG[0]
rlabel metal3 30048 366 30048 366 0 SS4BEG[10]
rlabel metal3 30240 828 30240 828 0 SS4BEG[11]
rlabel metal3 36192 1302 36192 1302 0 SS4BEG[12]
rlabel metal2 34656 3066 34656 3066 0 SS4BEG[13]
rlabel metal3 30816 3558 30816 3558 0 SS4BEG[14]
rlabel metal3 34416 3192 34416 3192 0 SS4BEG[15]
rlabel metal2 28728 6300 28728 6300 0 SS4BEG[1]
rlabel metal2 29016 6216 29016 6216 0 SS4BEG[2]
rlabel metal2 29472 3780 29472 3780 0 SS4BEG[3]
rlabel metal2 29184 4704 29184 4704 0 SS4BEG[4]
rlabel metal2 29160 7728 29160 7728 0 SS4BEG[5]
rlabel metal3 29280 912 29280 912 0 SS4BEG[6]
rlabel metal2 29544 7728 29544 7728 0 SS4BEG[7]
rlabel metal3 29664 240 29664 240 0 SS4BEG[8]
rlabel metal3 29856 660 29856 660 0 SS4BEG[9]
rlabel metal2 40416 4284 40416 4284 0 UserCLK
rlabel metal2 19704 8904 19704 8904 0 UserCLKo
rlabel metal2 8640 7392 8640 7392 0 _000_
rlabel metal3 7104 10122 7104 10122 0 _001_
rlabel via1 7688 6395 7688 6395 0 _002_
rlabel metal2 8016 6426 8016 6426 0 _003_
rlabel metal2 8156 6426 8156 6426 0 _004_
rlabel metal2 6036 5712 6036 5712 0 _005_
rlabel metal2 6240 4326 6240 4326 0 _006_
rlabel metal2 6432 4200 6432 4200 0 _007_
rlabel metal2 6048 4284 6048 4284 0 _008_
rlabel metal2 5493 4200 5493 4200 0 _009_
rlabel metal2 5664 4242 5664 4242 0 _010_
rlabel metal3 5856 4998 5856 4998 0 _011_
rlabel metal2 6144 5544 6144 5544 0 _012_
rlabel metal3 6912 5082 6912 5082 0 _013_
rlabel metal2 7128 4872 7128 4872 0 _014_
rlabel metal2 6645 5712 6645 5712 0 _015_
rlabel metal2 6240 5754 6240 5754 0 _016_
rlabel via1 10858 7213 10858 7213 0 _017_
rlabel metal2 10656 7434 10656 7434 0 _018_
rlabel metal2 10464 7266 10464 7266 0 _019_
rlabel metal2 11061 7224 11061 7224 0 _020_
rlabel metal2 10176 7728 10176 7728 0 _021_
rlabel metal2 10032 6216 10032 6216 0 _022_
rlabel metal2 10389 6384 10389 6384 0 _023_
rlabel metal2 9270 7266 9270 7266 0 _024_
rlabel metal2 9504 6510 9504 6510 0 _025_
rlabel metal2 10560 6510 10560 6510 0 _026_
rlabel metal2 10896 6468 10896 6468 0 _027_
rlabel metal2 11326 5712 11326 5712 0 _028_
rlabel metal2 11232 5796 11232 5796 0 _029_
rlabel metal2 11259 6384 11259 6384 0 _030_
rlabel metal3 11232 6720 11232 6720 0 _031_
rlabel metal2 7248 7392 7248 7392 0 _032_
rlabel via2 7307 7140 7307 7140 0 _033_
rlabel metal3 7200 8652 7200 8652 0 _034_
rlabel metal2 7632 7308 7632 7308 0 _035_
rlabel via1 7246 7938 7246 7938 0 _036_
rlabel via1 7139 7895 7139 7895 0 _037_
rlabel metal2 6336 7434 6336 7434 0 _038_
rlabel metal2 8184 7896 8184 7896 0 _039_
rlabel metal2 5304 3444 5304 3444 0 _040_
rlabel metal2 6240 3192 6240 3192 0 _041_
rlabel metal2 7083 2688 7083 2688 0 _042_
rlabel metal2 6864 2688 6864 2688 0 _043_
rlabel metal2 6651 2688 6651 2688 0 _044_
rlabel metal2 18624 8736 18624 8736 0 net1
rlabel metal4 22944 2142 22944 2142 0 net10
rlabel metal3 21888 4410 21888 4410 0 net100
rlabel metal2 16584 2100 16584 2100 0 net101
rlabel metal2 23712 9366 23712 9366 0 net102
rlabel metal2 16128 2772 16128 2772 0 net103
rlabel metal2 15552 9408 15552 9408 0 net104
rlabel metal3 34368 5166 34368 5166 0 net105
rlabel metal2 13272 2100 13272 2100 0 net106
rlabel metal2 20256 4074 20256 4074 0 net107
rlabel metal3 18624 6342 18624 6342 0 net108
rlabel metal3 34944 1722 34944 1722 0 net109
rlabel metal4 14400 3486 14400 3486 0 net11
rlabel metal2 21216 9114 21216 9114 0 net110
rlabel metal2 11376 7140 11376 7140 0 net111
rlabel metal2 8400 7812 8400 7812 0 net112
rlabel metal3 8928 9744 8928 9744 0 net113
rlabel metal3 38112 6846 38112 6846 0 net114
rlabel metal3 34752 8274 34752 8274 0 net115
rlabel metal3 14112 8022 14112 8022 0 net116
rlabel metal2 6288 5628 6288 5628 0 net117
rlabel metal3 6816 6216 6816 6216 0 net118
rlabel metal3 14592 10164 14592 10164 0 net119
rlabel metal2 20880 7896 20880 7896 0 net12
rlabel metal3 16992 10710 16992 10710 0 net120
rlabel metal3 15168 8568 15168 8568 0 net121
rlabel metal3 17952 6552 17952 6552 0 net122
rlabel metal3 44160 2184 44160 2184 0 net123
rlabel metal2 42528 9198 42528 9198 0 net124
rlabel metal3 29856 6090 29856 6090 0 net125
rlabel metal3 43584 5838 43584 5838 0 net126
rlabel metal3 43968 5586 43968 5586 0 net127
rlabel metal3 14208 6678 14208 6678 0 net128
rlabel metal3 21600 6720 21600 6720 0 net129
rlabel metal2 13056 6552 13056 6552 0 net13
rlabel metal2 8520 3276 8520 3276 0 net130
rlabel metal3 44736 4914 44736 4914 0 net131
rlabel metal2 17832 6468 17832 6468 0 net132
rlabel metal2 13992 6972 13992 6972 0 net133
rlabel metal2 43776 1764 43776 1764 0 net134
rlabel metal3 2784 5178 2784 5178 0 net135
rlabel metal2 8376 7140 8376 7140 0 net136
rlabel metal2 9672 9240 9672 9240 0 net137
rlabel metal3 9120 9198 9120 9198 0 net138
rlabel metal2 4248 8652 4248 8652 0 net139
rlabel metal3 21984 3150 21984 3150 0 net14
rlabel metal2 2856 4704 2856 4704 0 net140
rlabel metal3 2784 8400 2784 8400 0 net141
rlabel metal3 8640 8148 8640 8148 0 net142
rlabel metal3 42720 7896 42720 7896 0 net143
rlabel metal2 3144 3612 3144 3612 0 net144
rlabel metal2 43632 2604 43632 2604 0 net145
rlabel metal3 11616 7056 11616 7056 0 net146
rlabel metal2 2520 4284 2520 4284 0 net147
rlabel metal2 44544 1974 44544 1974 0 net148
rlabel metal2 44640 1974 44640 1974 0 net149
rlabel metal3 2496 2688 2496 2688 0 net15
rlabel metal2 44016 2520 44016 2520 0 net150
rlabel metal2 44928 2646 44928 2646 0 net151
rlabel metal3 41088 4914 41088 4914 0 net152
rlabel metal2 40704 4074 40704 4074 0 net153
rlabel metal2 41352 2856 41352 2856 0 net154
rlabel metal2 28200 6636 28200 6636 0 net155
rlabel metal2 42264 9660 42264 9660 0 net156
rlabel metal3 41472 9240 41472 9240 0 net157
rlabel metal3 42816 9492 42816 9492 0 net158
rlabel metal2 42408 9576 42408 9576 0 net159
rlabel metal3 8064 7308 8064 7308 0 net16
rlabel metal3 42144 9450 42144 9450 0 net160
rlabel metal3 43008 9702 43008 9702 0 net161
rlabel metal3 41856 9030 41856 9030 0 net162
rlabel metal2 42432 10122 42432 10122 0 net163
rlabel metal2 42816 10248 42816 10248 0 net164
rlabel metal2 43248 10164 43248 10164 0 net165
rlabel metal2 2376 2856 2376 2856 0 net166
rlabel metal2 36408 4704 36408 4704 0 net167
rlabel metal2 37176 6972 37176 6972 0 net168
rlabel metal2 42360 8484 42360 8484 0 net169
rlabel metal3 21888 10038 21888 10038 0 net17
rlabel metal2 37632 10710 37632 10710 0 net170
rlabel metal3 37536 11088 37536 11088 0 net171
rlabel metal2 35712 10290 35712 10290 0 net172
rlabel metal2 42600 9492 42600 9492 0 net173
rlabel metal3 32928 10542 32928 10542 0 net174
rlabel metal3 20064 4998 20064 4998 0 net175
rlabel metal3 17568 2688 17568 2688 0 net176
rlabel metal2 40968 3444 40968 3444 0 net177
rlabel metal2 17664 2646 17664 2646 0 net178
rlabel metal3 21216 5964 21216 5964 0 net179
rlabel metal2 20112 8736 20112 8736 0 net18
rlabel metal2 19344 3486 19344 3486 0 net180
rlabel metal2 21600 5586 21600 5586 0 net181
rlabel metal2 20112 3444 20112 3444 0 net182
rlabel metal2 20880 2688 20880 2688 0 net183
rlabel metal2 20736 2562 20736 2562 0 net184
rlabel metal2 20736 2016 20736 2016 0 net185
rlabel metal3 22752 2814 22752 2814 0 net186
rlabel metal2 23136 7098 23136 7098 0 net187
rlabel metal2 21648 1932 21648 1932 0 net188
rlabel metal2 40056 8148 40056 8148 0 net189
rlabel metal2 1488 9030 1488 9030 0 net19
rlabel metal2 26208 2562 26208 2562 0 net190
rlabel metal3 21696 9072 21696 9072 0 net191
rlabel metal2 18744 6552 18744 6552 0 net192
rlabel metal3 14400 9114 14400 9114 0 net193
rlabel metal2 28008 3192 28008 3192 0 net194
rlabel metal2 25968 4116 25968 4116 0 net195
rlabel metal3 33216 4242 33216 4242 0 net196
rlabel metal2 39912 2856 39912 2856 0 net197
rlabel metal2 39312 1680 39312 1680 0 net198
rlabel metal3 29280 5124 29280 5124 0 net199
rlabel metal2 22752 2688 22752 2688 0 net2
rlabel metal2 2400 4956 2400 4956 0 net20
rlabel metal2 26952 9492 26952 9492 0 net200
rlabel metal2 29952 5124 29952 5124 0 net201
rlabel metal2 25272 3612 25272 3612 0 net202
rlabel metal4 29088 2016 29088 2016 0 net203
rlabel metal2 21216 5292 21216 5292 0 net204
rlabel metal3 20928 2730 20928 2730 0 net205
rlabel metal2 20616 3612 20616 3612 0 net206
rlabel metal2 19848 10416 19848 10416 0 net207
rlabel metal3 21216 7056 21216 7056 0 net208
rlabel metal2 33696 2058 33696 2058 0 net209
rlabel metal2 1752 10416 1752 10416 0 net21
rlabel metal2 28896 5670 28896 5670 0 net210
rlabel metal2 33888 1932 33888 1932 0 net211
rlabel metal3 36096 3906 36096 3906 0 net212
rlabel metal2 38088 4284 38088 4284 0 net213
rlabel metal2 37896 10080 37896 10080 0 net214
rlabel metal2 36384 3444 36384 3444 0 net215
rlabel metal2 32064 6720 32064 6720 0 net216
rlabel metal2 13800 8148 13800 8148 0 net217
rlabel metal2 29568 6384 29568 6384 0 net218
rlabel metal2 29712 6468 29712 6468 0 net219
rlabel metal2 1872 9870 1872 9870 0 net22
rlabel metal3 32064 6342 32064 6342 0 net220
rlabel metal3 8928 6384 8928 6384 0 net221
rlabel metal3 29472 8274 29472 8274 0 net222
rlabel metal4 19584 2856 19584 2856 0 net223
rlabel metal2 9768 5544 9768 5544 0 net224
rlabel metal2 38088 4368 38088 4368 0 net225
rlabel metal2 33504 5586 33504 5586 0 net226
rlabel metal3 21408 7602 21408 7602 0 net227
rlabel metal3 40704 6090 40704 6090 0 net228
rlabel metal3 40992 4494 40992 4494 0 net229
rlabel metal3 2304 7896 2304 7896 0 net23
rlabel metal2 2928 3444 2928 3444 0 net24
rlabel metal2 2280 2100 2280 2100 0 net25
rlabel metal2 15168 10290 15168 10290 0 net26
rlabel metal2 2304 4158 2304 4158 0 net27
rlabel metal2 1752 2100 1752 2100 0 net28
rlabel metal2 2256 2604 2256 2604 0 net29
rlabel metal2 13920 2604 13920 2604 0 net3
rlabel metal2 1512 2520 1512 2520 0 net30
rlabel metal2 2424 3192 2424 3192 0 net31
rlabel metal2 17568 5880 17568 5880 0 net32
rlabel metal2 37920 1932 37920 1932 0 net33
rlabel metal3 2400 3906 2400 3906 0 net34
rlabel metal2 37800 2856 37800 2856 0 net35
rlabel metal2 17952 9870 17952 9870 0 net36
rlabel metal2 5352 3948 5352 3948 0 net37
rlabel metal2 3480 2856 3480 2856 0 net38
rlabel metal2 21648 2688 21648 2688 0 net39
rlabel metal2 1488 3780 1488 3780 0 net4
rlabel metal3 8832 2730 8832 2730 0 net40
rlabel metal2 7521 10248 7521 10248 0 net41
rlabel metal3 13632 6930 13632 6930 0 net42
rlabel metal2 9936 7308 9936 7308 0 net43
rlabel metal3 15840 4032 15840 4032 0 net44
rlabel metal2 14016 8148 14016 8148 0 net45
rlabel metal2 9915 6384 9915 6384 0 net46
rlabel metal3 9312 8190 9312 8190 0 net47
rlabel metal4 13248 4830 13248 4830 0 net48
rlabel metal2 3672 2100 3672 2100 0 net49
rlabel metal2 1872 5166 1872 5166 0 net5
rlabel metal2 13344 4872 13344 4872 0 net50
rlabel metal2 3816 1680 3816 1680 0 net51
rlabel metal2 28416 4662 28416 4662 0 net52
rlabel metal2 4488 2100 4488 2100 0 net53
rlabel metal2 8544 4200 8544 4200 0 net54
rlabel metal3 7200 2730 7200 2730 0 net55
rlabel metal2 14232 7980 14232 7980 0 net56
rlabel metal2 28656 2604 28656 2604 0 net57
rlabel metal4 18096 9576 18096 9576 0 net58
rlabel metal3 16992 6384 16992 6384 0 net59
rlabel metal2 1488 4620 1488 4620 0 net6
rlabel metal3 40608 7014 40608 7014 0 net60
rlabel metal4 17664 2814 17664 2814 0 net61
rlabel metal3 13440 2184 13440 2184 0 net62
rlabel metal2 20544 9660 20544 9660 0 net63
rlabel metal2 15792 2688 15792 2688 0 net64
rlabel metal2 21792 8904 21792 8904 0 net65
rlabel metal3 22944 7770 22944 7770 0 net66
rlabel metal2 35040 9408 35040 9408 0 net67
rlabel metal2 19056 2688 19056 2688 0 net68
rlabel metal2 4248 6216 4248 6216 0 net69
rlabel metal3 2400 5250 2400 5250 0 net7
rlabel metal2 10272 6426 10272 6426 0 net70
rlabel metal2 39456 2688 39456 2688 0 net71
rlabel metal2 14832 10248 14832 10248 0 net72
rlabel metal3 29952 5880 29952 5880 0 net73
rlabel metal2 39168 10206 39168 10206 0 net74
rlabel metal3 28320 8190 28320 8190 0 net75
rlabel metal2 14688 6342 14688 6342 0 net76
rlabel metal2 22584 4368 22584 4368 0 net77
rlabel metal2 20784 10248 20784 10248 0 net78
rlabel metal2 19488 10248 19488 10248 0 net79
rlabel metal2 21216 4872 21216 4872 0 net8
rlabel metal3 16416 10374 16416 10374 0 net80
rlabel metal2 22056 6300 22056 6300 0 net81
rlabel metal2 2112 2520 2112 2520 0 net82
rlabel metal2 41376 7854 41376 7854 0 net83
rlabel metal2 41664 9450 41664 9450 0 net84
rlabel metal2 37056 1848 37056 1848 0 net85
rlabel metal2 30816 4158 30816 4158 0 net86
rlabel metal2 4416 3360 4416 3360 0 net87
rlabel metal2 8640 2646 8640 2646 0 net88
rlabel metal3 2688 3528 2688 3528 0 net89
rlabel metal2 20352 7938 20352 7938 0 net9
rlabel metal2 34608 10248 34608 10248 0 net90
rlabel metal3 30048 6930 30048 6930 0 net91
rlabel metal2 21600 6258 21600 6258 0 net92
rlabel metal2 28512 2688 28512 2688 0 net93
rlabel metal2 8520 1680 8520 1680 0 net94
rlabel metal2 22080 7770 22080 7770 0 net95
rlabel metal2 19296 4956 19296 4956 0 net96
rlabel metal2 20640 9492 20640 9492 0 net97
rlabel metal2 34944 1848 34944 1848 0 net98
rlabel metal2 16008 2100 16008 2100 0 net99
<< properties >>
string FIXED_BBOX 0 0 46368 12180
<< end >>
