module S_EF_DAC8 (Co,
    UserCLK,
    UserCLKo,
    VALUE_top0,
    VALUE_top1,
    VALUE_top2,
    VALUE_top3,
    VALUE_top4,
    VALUE_top5,
    VALUE_top6,
    VALUE_top7,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    NN4BEG,
    S1END,
    S2END,
    S2MID,
    S4END,
    SS4END);
 output Co;
 input UserCLK;
 output UserCLKo;
 output VALUE_top0;
 output VALUE_top1;
 output VALUE_top2;
 output VALUE_top3;
 output VALUE_top4;
 output VALUE_top5;
 output VALUE_top6;
 output VALUE_top7;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 output [15:0] NN4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;
 input [15:0] SS4END;

 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_S_EF_DAC8_switch_matrix.N2BEG0 ;
 wire \Inst_S_EF_DAC8_switch_matrix.N2BEG1 ;
 wire \Inst_S_EF_DAC8_switch_matrix.N2BEG2 ;
 wire \Inst_S_EF_DAC8_switch_matrix.N2BEG3 ;
 wire \Inst_S_EF_DAC8_switch_matrix.N2BEG4 ;
 wire \Inst_S_EF_DAC8_switch_matrix.N2BEG5 ;
 wire \Inst_S_EF_DAC8_switch_matrix.N2BEG6 ;
 wire \Inst_S_EF_DAC8_switch_matrix.N2BEG7 ;
 wire \Inst_S_EF_DAC8_switch_matrix.N2BEGb0 ;
 wire \Inst_S_EF_DAC8_switch_matrix.N2BEGb1 ;
 wire \Inst_S_EF_DAC8_switch_matrix.N2BEGb2 ;
 wire \Inst_S_EF_DAC8_switch_matrix.N2BEGb3 ;
 wire \Inst_S_EF_DAC8_switch_matrix.N2BEGb4 ;
 wire \Inst_S_EF_DAC8_switch_matrix.N2BEGb5 ;
 wire \Inst_S_EF_DAC8_switch_matrix.N2BEGb6 ;
 wire \Inst_S_EF_DAC8_switch_matrix.N2BEGb7 ;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net196;

 sky130_fd_sc_hd__mux4_1 _000_ (.A0(net42),
    .A1(net46),
    .A2(net66),
    .A3(net80),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit30.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit31.Q ),
    .X(net195));
 sky130_fd_sc_hd__mux4_2 _001_ (.A0(net41),
    .A1(net45),
    .A2(net65),
    .A3(net79),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit28.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit29.Q ),
    .X(net194));
 sky130_fd_sc_hd__mux4_1 _002_ (.A0(net40),
    .A1(net44),
    .A2(net64),
    .A3(net78),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit26.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit27.Q ),
    .X(net193));
 sky130_fd_sc_hd__mux4_1 _003_ (.A0(net39),
    .A1(net43),
    .A2(net63),
    .A3(net77),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit24.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit25.Q ),
    .X(net192));
 sky130_fd_sc_hd__mux4_1 _004_ (.A0(net54),
    .A1(net50),
    .A2(net62),
    .A3(net76),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit22.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit23.Q ),
    .X(net191));
 sky130_fd_sc_hd__mux4_2 _005_ (.A0(net53),
    .A1(net49),
    .A2(net61),
    .A3(net75),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit20.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit21.Q ),
    .X(net190));
 sky130_fd_sc_hd__mux4_1 _006_ (.A0(net52),
    .A1(net48),
    .A2(net60),
    .A3(net74),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit18.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit19.Q ),
    .X(net189));
 sky130_fd_sc_hd__mux4_2 _007_ (.A0(net51),
    .A1(net47),
    .A2(net59),
    .A3(net67),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit16.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit17.Q ),
    .X(net188));
 sky130_fd_sc_hd__mux4_1 _008_ (.A0(net43),
    .A1(net59),
    .A2(net67),
    .A3(net81),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit14.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit15.Q ),
    .X(\Inst_S_EF_DAC8_switch_matrix.N2BEGb7 ));
 sky130_fd_sc_hd__mux4_1 _009_ (.A0(net44),
    .A1(net60),
    .A2(net74),
    .A3(net82),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit12.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit13.Q ),
    .X(\Inst_S_EF_DAC8_switch_matrix.N2BEGb6 ));
 sky130_fd_sc_hd__mux4_1 _010_ (.A0(net45),
    .A1(net61),
    .A2(net75),
    .A3(net68),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit10.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit11.Q ),
    .X(\Inst_S_EF_DAC8_switch_matrix.N2BEGb5 ));
 sky130_fd_sc_hd__mux4_1 _011_ (.A0(net46),
    .A1(net62),
    .A2(net76),
    .A3(net69),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit8.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit9.Q ),
    .X(\Inst_S_EF_DAC8_switch_matrix.N2BEGb4 ));
 sky130_fd_sc_hd__mux4_1 _012_ (.A0(net47),
    .A1(net77),
    .A2(net63),
    .A3(net70),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit7.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit6.Q ),
    .X(\Inst_S_EF_DAC8_switch_matrix.N2BEGb3 ));
 sky130_fd_sc_hd__mux4_1 _013_ (.A0(net48),
    .A1(net78),
    .A2(net64),
    .A3(net71),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit5.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit4.Q ),
    .X(\Inst_S_EF_DAC8_switch_matrix.N2BEGb2 ));
 sky130_fd_sc_hd__mux4_1 _014_ (.A0(net49),
    .A1(net79),
    .A2(net65),
    .A3(net72),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit3.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit2.Q ),
    .X(\Inst_S_EF_DAC8_switch_matrix.N2BEGb1 ));
 sky130_fd_sc_hd__mux4_1 _015_ (.A0(net50),
    .A1(net80),
    .A2(net66),
    .A3(net73),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit1.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit0.Q ),
    .X(\Inst_S_EF_DAC8_switch_matrix.N2BEGb0 ));
 sky130_fd_sc_hd__mux4_1 _016_ (.A0(net51),
    .A1(net59),
    .A2(net67),
    .A3(net81),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit30.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit31.Q ),
    .X(\Inst_S_EF_DAC8_switch_matrix.N2BEG7 ));
 sky130_fd_sc_hd__mux4_1 _017_ (.A0(net52),
    .A1(net60),
    .A2(net74),
    .A3(net82),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit29.Q ),
    .X(\Inst_S_EF_DAC8_switch_matrix.N2BEG6 ));
 sky130_fd_sc_hd__mux4_1 _018_ (.A0(net53),
    .A1(net61),
    .A2(net75),
    .A3(net68),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit26.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Inst_S_EF_DAC8_switch_matrix.N2BEG5 ));
 sky130_fd_sc_hd__mux4_1 _019_ (.A0(net54),
    .A1(net62),
    .A2(net76),
    .A3(net69),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit25.Q ),
    .X(\Inst_S_EF_DAC8_switch_matrix.N2BEG4 ));
 sky130_fd_sc_hd__mux4_1 _020_ (.A0(net55),
    .A1(net77),
    .A2(net63),
    .A3(net70),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit23.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit22.Q ),
    .X(\Inst_S_EF_DAC8_switch_matrix.N2BEG3 ));
 sky130_fd_sc_hd__mux4_1 _021_ (.A0(net56),
    .A1(net78),
    .A2(net64),
    .A3(net71),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit21.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit20.Q ),
    .X(\Inst_S_EF_DAC8_switch_matrix.N2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _022_ (.A0(net57),
    .A1(net79),
    .A2(net65),
    .A3(net72),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit19.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit18.Q ),
    .X(\Inst_S_EF_DAC8_switch_matrix.N2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _023_ (.A0(net58),
    .A1(net80),
    .A2(net66),
    .A3(net73),
    .S0(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit17.Q ),
    .S1(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit16.Q ),
    .X(\Inst_S_EF_DAC8_switch_matrix.N2BEG0 ));
 sky130_fd_sc_hd__dlxtp_1 _024_ (.D(net8),
    .GATE(net13),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _025_ (.D(net9),
    .GATE(net14),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _026_ (.D(net10),
    .GATE(net14),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _027_ (.D(net11),
    .GATE(net14),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _028_ (.D(net19),
    .GATE(net13),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _029_ (.D(net20),
    .GATE(net13),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _030_ (.D(net21),
    .GATE(net13),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _031_ (.D(net22),
    .GATE(net13),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _032_ (.D(net23),
    .GATE(net13),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _033_ (.D(net24),
    .GATE(net13),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _034_ (.D(net25),
    .GATE(net14),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _035_ (.D(net26),
    .GATE(net14),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _036_ (.D(net27),
    .GATE(net13),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _037_ (.D(net28),
    .GATE(net13),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _038_ (.D(net30),
    .GATE(net14),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _039_ (.D(net31),
    .GATE(net14),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _040_ (.D(net1),
    .GATE(net15),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _041_ (.D(net12),
    .GATE(net15),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _042_ (.D(net29),
    .GATE(net17),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _043_ (.D(net32),
    .GATE(net17),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _044_ (.D(net33),
    .GATE(net16),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _045_ (.D(net34),
    .GATE(net16),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _046_ (.D(net35),
    .GATE(net15),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _047_ (.D(net36),
    .GATE(net15),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _048_ (.D(net37),
    .GATE(net16),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _049_ (.D(net38),
    .GATE(net16),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _050_ (.D(net2),
    .GATE(net17),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _051_ (.D(net3),
    .GATE(net17),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _052_ (.D(net4),
    .GATE(net16),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _053_ (.D(net5),
    .GATE(net16),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _054_ (.D(net6),
    .GATE(net15),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _055_ (.D(net7),
    .GATE(net15),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _056_ (.D(net8),
    .GATE(net18),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _057_ (.D(net9),
    .GATE(net15),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _058_ (.D(net10),
    .GATE(net16),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _059_ (.D(net11),
    .GATE(net16),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _060_ (.D(net19),
    .GATE(net17),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _061_ (.D(net20),
    .GATE(net18),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _062_ (.D(net21),
    .GATE(net15),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _063_ (.D(net22),
    .GATE(net15),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _064_ (.D(net23),
    .GATE(net15),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _065_ (.D(net24),
    .GATE(net18),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _066_ (.D(net25),
    .GATE(net16),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _067_ (.D(net26),
    .GATE(net16),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _068_ (.D(net27),
    .GATE(net17),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _069_ (.D(net28),
    .GATE(net17),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _070_ (.D(net30),
    .GATE(net17),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _071_ (.D(net31),
    .GATE(net17),
    .Q(\Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit31.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net110));
 sky130_fd_sc_hd__clkbuf_2 _073_ (.A(net1),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 _074_ (.A(net12),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 _075_ (.A(net29),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 _076_ (.A(net32),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 _077_ (.A(net33),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 _078_ (.A(net34),
    .X(net110));
 sky130_fd_sc_hd__buf_1 _079_ (.A(net35),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 _080_ (.A(net36),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 _081_ (.A(net37),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 _082_ (.A(net38),
    .X(net114));
 sky130_fd_sc_hd__buf_1 _083_ (.A(net2),
    .X(net84));
 sky130_fd_sc_hd__buf_1 _084_ (.A(net3),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 _085_ (.A(net4),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 _086_ (.A(net5),
    .X(net87));
 sky130_fd_sc_hd__buf_1 _087_ (.A(net6),
    .X(net88));
 sky130_fd_sc_hd__buf_1 _088_ (.A(net7),
    .X(net89));
 sky130_fd_sc_hd__buf_1 _089_ (.A(net8),
    .X(net90));
 sky130_fd_sc_hd__buf_1 _090_ (.A(net9),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 _091_ (.A(net10),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 _092_ (.A(net11),
    .X(net93));
 sky130_fd_sc_hd__buf_1 _093_ (.A(net19),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 _094_ (.A(net20),
    .X(net96));
 sky130_fd_sc_hd__buf_1 _095_ (.A(net21),
    .X(net97));
 sky130_fd_sc_hd__buf_1 _096_ (.A(net22),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 _097_ (.A(net23),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 _098_ (.A(net24),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 _099_ (.A(net25),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 _100_ (.A(net26),
    .X(net102));
 sky130_fd_sc_hd__buf_1 _101_ (.A(net27),
    .X(net103));
 sky130_fd_sc_hd__buf_1 _102_ (.A(net28),
    .X(net104));
 sky130_fd_sc_hd__buf_1 _103_ (.A(net30),
    .X(net106));
 sky130_fd_sc_hd__buf_1 _104_ (.A(net31),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 _105_ (.A(net17),
    .X(net115));
 sky130_fd_sc_hd__buf_1 _106_ (.A(net13),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 _107_ (.A(FrameStrobe[2]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 _108_ (.A(FrameStrobe[3]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 _109_ (.A(FrameStrobe[4]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 _110_ (.A(FrameStrobe[5]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 _111_ (.A(FrameStrobe[6]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 _112_ (.A(FrameStrobe[7]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 _113_ (.A(FrameStrobe[8]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 _114_ (.A(FrameStrobe[9]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 _115_ (.A(FrameStrobe[10]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 _116_ (.A(FrameStrobe[11]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 _117_ (.A(FrameStrobe[12]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 _118_ (.A(FrameStrobe[13]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 _119_ (.A(FrameStrobe[14]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 _120_ (.A(FrameStrobe[15]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 _121_ (.A(FrameStrobe[16]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 _122_ (.A(FrameStrobe[17]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 _123_ (.A(FrameStrobe[18]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 _124_ (.A(FrameStrobe[19]),
    .X(net125));
 sky130_fd_sc_hd__buf_1 _125_ (.A(net42),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 _126_ (.A(net41),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 _127_ (.A(net40),
    .X(net137));
 sky130_fd_sc_hd__buf_1 _128_ (.A(net39),
    .X(net138));
 sky130_fd_sc_hd__buf_1 _129_ (.A(\Inst_S_EF_DAC8_switch_matrix.N2BEG0 ),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 _130_ (.A(\Inst_S_EF_DAC8_switch_matrix.N2BEG1 ),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 _131_ (.A(\Inst_S_EF_DAC8_switch_matrix.N2BEG2 ),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 _132_ (.A(\Inst_S_EF_DAC8_switch_matrix.N2BEG3 ),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 _133_ (.A(\Inst_S_EF_DAC8_switch_matrix.N2BEG4 ),
    .X(net143));
 sky130_fd_sc_hd__buf_1 _134_ (.A(\Inst_S_EF_DAC8_switch_matrix.N2BEG5 ),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 _135_ (.A(\Inst_S_EF_DAC8_switch_matrix.N2BEG6 ),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 _136_ (.A(\Inst_S_EF_DAC8_switch_matrix.N2BEG7 ),
    .X(net146));
 sky130_fd_sc_hd__buf_1 _137_ (.A(\Inst_S_EF_DAC8_switch_matrix.N2BEGb0 ),
    .X(net147));
 sky130_fd_sc_hd__buf_1 _138_ (.A(\Inst_S_EF_DAC8_switch_matrix.N2BEGb1 ),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 _139_ (.A(\Inst_S_EF_DAC8_switch_matrix.N2BEGb2 ),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 _140_ (.A(\Inst_S_EF_DAC8_switch_matrix.N2BEGb3 ),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 _141_ (.A(\Inst_S_EF_DAC8_switch_matrix.N2BEGb4 ),
    .X(net151));
 sky130_fd_sc_hd__buf_1 _142_ (.A(\Inst_S_EF_DAC8_switch_matrix.N2BEGb5 ),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 _143_ (.A(\Inst_S_EF_DAC8_switch_matrix.N2BEGb6 ),
    .X(net153));
 sky130_fd_sc_hd__buf_1 _144_ (.A(\Inst_S_EF_DAC8_switch_matrix.N2BEGb7 ),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_2 _145_ (.A(S4END[15]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 _146_ (.A(S4END[14]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 _147_ (.A(S4END[13]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_2 _148_ (.A(S4END[12]),
    .X(net164));
 sky130_fd_sc_hd__buf_1 _149_ (.A(S4END[11]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_2 _150_ (.A(S4END[10]),
    .X(net166));
 sky130_fd_sc_hd__buf_1 _151_ (.A(S4END[9]),
    .X(net167));
 sky130_fd_sc_hd__buf_1 _152_ (.A(S4END[8]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 _153_ (.A(net66),
    .X(net169));
 sky130_fd_sc_hd__buf_1 _154_ (.A(net65),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 _155_ (.A(net64),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 _156_ (.A(net63),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 _157_ (.A(net62),
    .X(net158));
 sky130_fd_sc_hd__buf_1 _158_ (.A(net61),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 _159_ (.A(net60),
    .X(net160));
 sky130_fd_sc_hd__buf_1 _160_ (.A(net59),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 _161_ (.A(net73),
    .X(net171));
 sky130_fd_sc_hd__buf_1 _162_ (.A(net72),
    .X(net178));
 sky130_fd_sc_hd__buf_1 _163_ (.A(net71),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 _164_ (.A(net70),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 _165_ (.A(net69),
    .X(net181));
 sky130_fd_sc_hd__buf_1 _166_ (.A(net68),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 _167_ (.A(net82),
    .X(net183));
 sky130_fd_sc_hd__buf_1 _168_ (.A(net81),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 _169_ (.A(net80),
    .X(net185));
 sky130_fd_sc_hd__buf_1 _170_ (.A(net79),
    .X(net186));
 sky130_fd_sc_hd__buf_1 _171_ (.A(net78),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 _172_ (.A(net77),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 _173_ (.A(net76),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 _174_ (.A(net75),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 _175_ (.A(net74),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 _176_ (.A(net67),
    .X(net177));
 sky130_fd_sc_hd__buf_2 _177_ (.A(UserCLK),
    .X(net187));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_121 ();
 sky130_fd_sc_hd__clkbuf_2 fanout13 (.A(FrameStrobe[1]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout14 (.A(FrameStrobe[1]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 fanout15 (.A(net18),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 fanout16 (.A(net18),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 fanout17 (.A(net18),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 fanout18 (.A(FrameStrobe[0]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input1 (.A(FrameData[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(FrameData[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(FrameData[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(FrameData[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(FrameData[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(FrameData[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(FrameData[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(FrameData[16]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(FrameData[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(FrameData[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(FrameData[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(FrameData[1]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(FrameData[20]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input14 (.A(FrameData[21]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input15 (.A(FrameData[22]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input16 (.A(FrameData[23]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input17 (.A(FrameData[24]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input18 (.A(FrameData[25]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input19 (.A(FrameData[26]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input20 (.A(FrameData[27]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(FrameData[28]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(FrameData[29]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(FrameData[2]),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(FrameData[30]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(FrameData[31]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(FrameData[3]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(FrameData[4]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(FrameData[5]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input29 (.A(FrameData[6]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input30 (.A(FrameData[7]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input31 (.A(FrameData[8]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input32 (.A(FrameData[9]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(S1END[0]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input34 (.A(S1END[1]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input35 (.A(S1END[2]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(S1END[3]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input37 (.A(S2END[0]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input38 (.A(S2END[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input39 (.A(S2END[2]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input40 (.A(S2END[3]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input41 (.A(S2END[4]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input42 (.A(S2END[5]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input43 (.A(S2END[6]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input44 (.A(S2END[7]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input45 (.A(S2MID[0]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input46 (.A(S2MID[1]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input47 (.A(S2MID[2]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input48 (.A(S2MID[3]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(S2MID[4]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input50 (.A(S2MID[5]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(S2MID[6]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(S2MID[7]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input53 (.A(S4END[0]),
    .X(net59));
 sky130_fd_sc_hd__dlymetal6s2s_1 input54 (.A(S4END[1]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input55 (.A(S4END[2]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input56 (.A(S4END[3]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input57 (.A(S4END[4]),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 input58 (.A(S4END[5]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input59 (.A(S4END[6]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input60 (.A(S4END[7]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input61 (.A(SS4END[0]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input62 (.A(SS4END[10]),
    .X(net68));
 sky130_fd_sc_hd__dlymetal6s2s_1 input63 (.A(SS4END[11]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input64 (.A(SS4END[12]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(SS4END[13]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 input66 (.A(SS4END[14]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input67 (.A(SS4END[15]),
    .X(net73));
 sky130_fd_sc_hd__dlymetal6s2s_1 input68 (.A(SS4END[1]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 input69 (.A(SS4END[2]),
    .X(net75));
 sky130_fd_sc_hd__dlymetal6s2s_1 input70 (.A(SS4END[3]),
    .X(net76));
 sky130_fd_sc_hd__buf_1 input71 (.A(SS4END[4]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input72 (.A(SS4END[5]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 input73 (.A(SS4END[6]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input74 (.A(SS4END[7]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input75 (.A(SS4END[8]),
    .X(net81));
 sky130_fd_sc_hd__dlymetal6s2s_1 input76 (.A(SS4END[9]),
    .X(net82));
 sky130_fd_sc_hd__buf_2 output77 (.A(net83),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net84),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net85),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net86),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net87),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net88),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net89),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net90),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net91),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net92),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net93),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net94),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net95),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net96),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net97),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net98),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net99),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net100),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net101),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net102),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net103),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net104),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net105),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net106),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net107),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net108),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net109),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net110),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net111),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net112),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net113),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net114),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net115),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net116),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net117),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net118),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net119),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net120),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net121),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net122),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net123),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net124),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net125),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net126),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net127),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net128),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net129),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net130),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net131),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net132),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net133),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net134),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net135),
    .X(N1BEG[0]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net136),
    .X(N1BEG[1]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net137),
    .X(N1BEG[2]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net138),
    .X(N1BEG[3]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net139),
    .X(N2BEG[0]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net140),
    .X(N2BEG[1]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net141),
    .X(N2BEG[2]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net142),
    .X(N2BEG[3]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net143),
    .X(N2BEG[4]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net144),
    .X(N2BEG[5]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net145),
    .X(N2BEG[6]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net146),
    .X(N2BEG[7]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net147),
    .X(N2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net148),
    .X(N2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net149),
    .X(N2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net150),
    .X(N2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net151),
    .X(N2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net152),
    .X(N2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net153),
    .X(N2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net154),
    .X(N2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net155),
    .X(N4BEG[0]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net156),
    .X(N4BEG[10]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net157),
    .X(N4BEG[11]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net158),
    .X(N4BEG[12]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net159),
    .X(N4BEG[13]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net160),
    .X(N4BEG[14]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net161),
    .X(N4BEG[15]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net162),
    .X(N4BEG[1]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net163),
    .X(N4BEG[2]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net164),
    .X(N4BEG[3]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net165),
    .X(N4BEG[4]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net166),
    .X(N4BEG[5]));
 sky130_fd_sc_hd__buf_2 output161 (.A(net167),
    .X(N4BEG[6]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net168),
    .X(N4BEG[7]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net169),
    .X(N4BEG[8]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net170),
    .X(N4BEG[9]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net171),
    .X(NN4BEG[0]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net172),
    .X(NN4BEG[10]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net173),
    .X(NN4BEG[11]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net174),
    .X(NN4BEG[12]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net175),
    .X(NN4BEG[13]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net176),
    .X(NN4BEG[14]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net177),
    .X(NN4BEG[15]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net178),
    .X(NN4BEG[1]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net179),
    .X(NN4BEG[2]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net180),
    .X(NN4BEG[3]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net181),
    .X(NN4BEG[4]));
 sky130_fd_sc_hd__buf_2 output176 (.A(net182),
    .X(NN4BEG[5]));
 sky130_fd_sc_hd__buf_2 output177 (.A(net183),
    .X(NN4BEG[6]));
 sky130_fd_sc_hd__buf_2 output178 (.A(net184),
    .X(NN4BEG[7]));
 sky130_fd_sc_hd__buf_2 output179 (.A(net185),
    .X(NN4BEG[8]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net186),
    .X(NN4BEG[9]));
 sky130_fd_sc_hd__buf_1 output181 (.A(net187),
    .X(UserCLKo));
 sky130_fd_sc_hd__buf_2 output182 (.A(net188),
    .X(VALUE_top0));
 sky130_fd_sc_hd__buf_2 output183 (.A(net189),
    .X(VALUE_top1));
 sky130_fd_sc_hd__buf_2 output184 (.A(net190),
    .X(VALUE_top2));
 sky130_fd_sc_hd__buf_2 output185 (.A(net191),
    .X(VALUE_top3));
 sky130_fd_sc_hd__buf_2 output186 (.A(net192),
    .X(VALUE_top4));
 sky130_fd_sc_hd__buf_2 output187 (.A(net193),
    .X(VALUE_top5));
 sky130_fd_sc_hd__buf_2 output188 (.A(net194),
    .X(VALUE_top6));
 sky130_fd_sc_hd__buf_2 output189 (.A(net195),
    .X(VALUE_top7));
 sky130_fd_sc_hd__conb_1 S_EF_DAC8_190 (.LO(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(FrameStrobe[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(FrameStrobe[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(FrameStrobe[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(FrameStrobe[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(FrameStrobe[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(S4END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(S4END[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net71));
 sky130_fd_sc_hd__decap_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_409 ();
 assign Co = net196;
endmodule
