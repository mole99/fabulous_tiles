VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DSP
  CLASS BLOCK ;
  FOREIGN DSP ;
  ORIGIN 0.000 0.000 ;
  SIZE 196.320 BY 483.840 ;
  PIN Tile_X0Y0_E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 336.220 196.320 336.620 ;
    END
  END Tile_X0Y0_E1BEG[0]
  PIN Tile_X0Y0_E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 337.900 196.320 338.300 ;
    END
  END Tile_X0Y0_E1BEG[1]
  PIN Tile_X0Y0_E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 339.580 196.320 339.980 ;
    END
  END Tile_X0Y0_E1BEG[2]
  PIN Tile_X0Y0_E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 341.260 196.320 341.660 ;
    END
  END Tile_X0Y0_E1BEG[3]
  PIN Tile_X0Y0_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 336.220 0.450 336.620 ;
    END
  END Tile_X0Y0_E1END[0]
  PIN Tile_X0Y0_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 337.900 0.450 338.300 ;
    END
  END Tile_X0Y0_E1END[1]
  PIN Tile_X0Y0_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 339.580 0.450 339.980 ;
    END
  END Tile_X0Y0_E1END[2]
  PIN Tile_X0Y0_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 341.260 0.450 341.660 ;
    END
  END Tile_X0Y0_E1END[3]
  PIN Tile_X0Y0_E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 342.940 196.320 343.340 ;
    END
  END Tile_X0Y0_E2BEG[0]
  PIN Tile_X0Y0_E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 344.620 196.320 345.020 ;
    END
  END Tile_X0Y0_E2BEG[1]
  PIN Tile_X0Y0_E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 346.300 196.320 346.700 ;
    END
  END Tile_X0Y0_E2BEG[2]
  PIN Tile_X0Y0_E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 347.980 196.320 348.380 ;
    END
  END Tile_X0Y0_E2BEG[3]
  PIN Tile_X0Y0_E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 349.660 196.320 350.060 ;
    END
  END Tile_X0Y0_E2BEG[4]
  PIN Tile_X0Y0_E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 351.340 196.320 351.740 ;
    END
  END Tile_X0Y0_E2BEG[5]
  PIN Tile_X0Y0_E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 353.020 196.320 353.420 ;
    END
  END Tile_X0Y0_E2BEG[6]
  PIN Tile_X0Y0_E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 354.700 196.320 355.100 ;
    END
  END Tile_X0Y0_E2BEG[7]
  PIN Tile_X0Y0_E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 356.380 196.320 356.780 ;
    END
  END Tile_X0Y0_E2BEGb[0]
  PIN Tile_X0Y0_E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 358.060 196.320 358.460 ;
    END
  END Tile_X0Y0_E2BEGb[1]
  PIN Tile_X0Y0_E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 359.740 196.320 360.140 ;
    END
  END Tile_X0Y0_E2BEGb[2]
  PIN Tile_X0Y0_E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 361.420 196.320 361.820 ;
    END
  END Tile_X0Y0_E2BEGb[3]
  PIN Tile_X0Y0_E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 363.100 196.320 363.500 ;
    END
  END Tile_X0Y0_E2BEGb[4]
  PIN Tile_X0Y0_E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 364.780 196.320 365.180 ;
    END
  END Tile_X0Y0_E2BEGb[5]
  PIN Tile_X0Y0_E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 366.460 196.320 366.860 ;
    END
  END Tile_X0Y0_E2BEGb[6]
  PIN Tile_X0Y0_E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 368.140 196.320 368.540 ;
    END
  END Tile_X0Y0_E2BEGb[7]
  PIN Tile_X0Y0_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 356.380 0.450 356.780 ;
    END
  END Tile_X0Y0_E2END[0]
  PIN Tile_X0Y0_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 358.060 0.450 358.460 ;
    END
  END Tile_X0Y0_E2END[1]
  PIN Tile_X0Y0_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 359.740 0.450 360.140 ;
    END
  END Tile_X0Y0_E2END[2]
  PIN Tile_X0Y0_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 361.420 0.450 361.820 ;
    END
  END Tile_X0Y0_E2END[3]
  PIN Tile_X0Y0_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 363.100 0.450 363.500 ;
    END
  END Tile_X0Y0_E2END[4]
  PIN Tile_X0Y0_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 364.780 0.450 365.180 ;
    END
  END Tile_X0Y0_E2END[5]
  PIN Tile_X0Y0_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 366.460 0.450 366.860 ;
    END
  END Tile_X0Y0_E2END[6]
  PIN Tile_X0Y0_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 368.140 0.450 368.540 ;
    END
  END Tile_X0Y0_E2END[7]
  PIN Tile_X0Y0_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 342.940 0.450 343.340 ;
    END
  END Tile_X0Y0_E2MID[0]
  PIN Tile_X0Y0_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 344.620 0.450 345.020 ;
    END
  END Tile_X0Y0_E2MID[1]
  PIN Tile_X0Y0_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 346.300 0.450 346.700 ;
    END
  END Tile_X0Y0_E2MID[2]
  PIN Tile_X0Y0_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 347.980 0.450 348.380 ;
    END
  END Tile_X0Y0_E2MID[3]
  PIN Tile_X0Y0_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 349.660 0.450 350.060 ;
    END
  END Tile_X0Y0_E2MID[4]
  PIN Tile_X0Y0_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 351.340 0.450 351.740 ;
    END
  END Tile_X0Y0_E2MID[5]
  PIN Tile_X0Y0_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 353.020 0.450 353.420 ;
    END
  END Tile_X0Y0_E2MID[6]
  PIN Tile_X0Y0_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 354.700 0.450 355.100 ;
    END
  END Tile_X0Y0_E2MID[7]
  PIN Tile_X0Y0_E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 396.700 196.320 397.100 ;
    END
  END Tile_X0Y0_E6BEG[0]
  PIN Tile_X0Y0_E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 413.500 196.320 413.900 ;
    END
  END Tile_X0Y0_E6BEG[10]
  PIN Tile_X0Y0_E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 415.180 196.320 415.580 ;
    END
  END Tile_X0Y0_E6BEG[11]
  PIN Tile_X0Y0_E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 398.380 196.320 398.780 ;
    END
  END Tile_X0Y0_E6BEG[1]
  PIN Tile_X0Y0_E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 400.060 196.320 400.460 ;
    END
  END Tile_X0Y0_E6BEG[2]
  PIN Tile_X0Y0_E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 401.740 196.320 402.140 ;
    END
  END Tile_X0Y0_E6BEG[3]
  PIN Tile_X0Y0_E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 403.420 196.320 403.820 ;
    END
  END Tile_X0Y0_E6BEG[4]
  PIN Tile_X0Y0_E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 405.100 196.320 405.500 ;
    END
  END Tile_X0Y0_E6BEG[5]
  PIN Tile_X0Y0_E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 406.780 196.320 407.180 ;
    END
  END Tile_X0Y0_E6BEG[6]
  PIN Tile_X0Y0_E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 408.460 196.320 408.860 ;
    END
  END Tile_X0Y0_E6BEG[7]
  PIN Tile_X0Y0_E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 410.140 196.320 410.540 ;
    END
  END Tile_X0Y0_E6BEG[8]
  PIN Tile_X0Y0_E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 411.820 196.320 412.220 ;
    END
  END Tile_X0Y0_E6BEG[9]
  PIN Tile_X0Y0_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 396.700 0.450 397.100 ;
    END
  END Tile_X0Y0_E6END[0]
  PIN Tile_X0Y0_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 413.500 0.450 413.900 ;
    END
  END Tile_X0Y0_E6END[10]
  PIN Tile_X0Y0_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 415.180 0.450 415.580 ;
    END
  END Tile_X0Y0_E6END[11]
  PIN Tile_X0Y0_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 398.380 0.450 398.780 ;
    END
  END Tile_X0Y0_E6END[1]
  PIN Tile_X0Y0_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 400.060 0.450 400.460 ;
    END
  END Tile_X0Y0_E6END[2]
  PIN Tile_X0Y0_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 401.740 0.450 402.140 ;
    END
  END Tile_X0Y0_E6END[3]
  PIN Tile_X0Y0_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 403.420 0.450 403.820 ;
    END
  END Tile_X0Y0_E6END[4]
  PIN Tile_X0Y0_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 405.100 0.450 405.500 ;
    END
  END Tile_X0Y0_E6END[5]
  PIN Tile_X0Y0_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 406.780 0.450 407.180 ;
    END
  END Tile_X0Y0_E6END[6]
  PIN Tile_X0Y0_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 408.460 0.450 408.860 ;
    END
  END Tile_X0Y0_E6END[7]
  PIN Tile_X0Y0_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 410.140 0.450 410.540 ;
    END
  END Tile_X0Y0_E6END[8]
  PIN Tile_X0Y0_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 411.820 0.450 412.220 ;
    END
  END Tile_X0Y0_E6END[9]
  PIN Tile_X0Y0_EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 369.820 196.320 370.220 ;
    END
  END Tile_X0Y0_EE4BEG[0]
  PIN Tile_X0Y0_EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 386.620 196.320 387.020 ;
    END
  END Tile_X0Y0_EE4BEG[10]
  PIN Tile_X0Y0_EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 388.300 196.320 388.700 ;
    END
  END Tile_X0Y0_EE4BEG[11]
  PIN Tile_X0Y0_EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 389.980 196.320 390.380 ;
    END
  END Tile_X0Y0_EE4BEG[12]
  PIN Tile_X0Y0_EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 391.660 196.320 392.060 ;
    END
  END Tile_X0Y0_EE4BEG[13]
  PIN Tile_X0Y0_EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 393.340 196.320 393.740 ;
    END
  END Tile_X0Y0_EE4BEG[14]
  PIN Tile_X0Y0_EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 395.020 196.320 395.420 ;
    END
  END Tile_X0Y0_EE4BEG[15]
  PIN Tile_X0Y0_EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 371.500 196.320 371.900 ;
    END
  END Tile_X0Y0_EE4BEG[1]
  PIN Tile_X0Y0_EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 373.180 196.320 373.580 ;
    END
  END Tile_X0Y0_EE4BEG[2]
  PIN Tile_X0Y0_EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 374.860 196.320 375.260 ;
    END
  END Tile_X0Y0_EE4BEG[3]
  PIN Tile_X0Y0_EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 376.540 196.320 376.940 ;
    END
  END Tile_X0Y0_EE4BEG[4]
  PIN Tile_X0Y0_EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 378.220 196.320 378.620 ;
    END
  END Tile_X0Y0_EE4BEG[5]
  PIN Tile_X0Y0_EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 379.900 196.320 380.300 ;
    END
  END Tile_X0Y0_EE4BEG[6]
  PIN Tile_X0Y0_EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 381.580 196.320 381.980 ;
    END
  END Tile_X0Y0_EE4BEG[7]
  PIN Tile_X0Y0_EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 383.260 196.320 383.660 ;
    END
  END Tile_X0Y0_EE4BEG[8]
  PIN Tile_X0Y0_EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 384.940 196.320 385.340 ;
    END
  END Tile_X0Y0_EE4BEG[9]
  PIN Tile_X0Y0_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 369.820 0.450 370.220 ;
    END
  END Tile_X0Y0_EE4END[0]
  PIN Tile_X0Y0_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 386.620 0.450 387.020 ;
    END
  END Tile_X0Y0_EE4END[10]
  PIN Tile_X0Y0_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 388.300 0.450 388.700 ;
    END
  END Tile_X0Y0_EE4END[11]
  PIN Tile_X0Y0_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 389.980 0.450 390.380 ;
    END
  END Tile_X0Y0_EE4END[12]
  PIN Tile_X0Y0_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 391.660 0.450 392.060 ;
    END
  END Tile_X0Y0_EE4END[13]
  PIN Tile_X0Y0_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 393.340 0.450 393.740 ;
    END
  END Tile_X0Y0_EE4END[14]
  PIN Tile_X0Y0_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 395.020 0.450 395.420 ;
    END
  END Tile_X0Y0_EE4END[15]
  PIN Tile_X0Y0_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 371.500 0.450 371.900 ;
    END
  END Tile_X0Y0_EE4END[1]
  PIN Tile_X0Y0_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 373.180 0.450 373.580 ;
    END
  END Tile_X0Y0_EE4END[2]
  PIN Tile_X0Y0_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 374.860 0.450 375.260 ;
    END
  END Tile_X0Y0_EE4END[3]
  PIN Tile_X0Y0_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 376.540 0.450 376.940 ;
    END
  END Tile_X0Y0_EE4END[4]
  PIN Tile_X0Y0_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 378.220 0.450 378.620 ;
    END
  END Tile_X0Y0_EE4END[5]
  PIN Tile_X0Y0_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 379.900 0.450 380.300 ;
    END
  END Tile_X0Y0_EE4END[6]
  PIN Tile_X0Y0_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 381.580 0.450 381.980 ;
    END
  END Tile_X0Y0_EE4END[7]
  PIN Tile_X0Y0_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 383.260 0.450 383.660 ;
    END
  END Tile_X0Y0_EE4END[8]
  PIN Tile_X0Y0_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 384.940 0.450 385.340 ;
    END
  END Tile_X0Y0_EE4END[9]
  PIN Tile_X0Y0_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 416.860 0.450 417.260 ;
    END
  END Tile_X0Y0_FrameData[0]
  PIN Tile_X0Y0_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 433.660 0.450 434.060 ;
    END
  END Tile_X0Y0_FrameData[10]
  PIN Tile_X0Y0_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 435.340 0.450 435.740 ;
    END
  END Tile_X0Y0_FrameData[11]
  PIN Tile_X0Y0_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 437.020 0.450 437.420 ;
    END
  END Tile_X0Y0_FrameData[12]
  PIN Tile_X0Y0_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 438.700 0.450 439.100 ;
    END
  END Tile_X0Y0_FrameData[13]
  PIN Tile_X0Y0_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 440.380 0.450 440.780 ;
    END
  END Tile_X0Y0_FrameData[14]
  PIN Tile_X0Y0_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 442.060 0.450 442.460 ;
    END
  END Tile_X0Y0_FrameData[15]
  PIN Tile_X0Y0_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 443.740 0.450 444.140 ;
    END
  END Tile_X0Y0_FrameData[16]
  PIN Tile_X0Y0_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 445.420 0.450 445.820 ;
    END
  END Tile_X0Y0_FrameData[17]
  PIN Tile_X0Y0_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 447.100 0.450 447.500 ;
    END
  END Tile_X0Y0_FrameData[18]
  PIN Tile_X0Y0_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 448.780 0.450 449.180 ;
    END
  END Tile_X0Y0_FrameData[19]
  PIN Tile_X0Y0_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 418.540 0.450 418.940 ;
    END
  END Tile_X0Y0_FrameData[1]
  PIN Tile_X0Y0_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 450.460 0.450 450.860 ;
    END
  END Tile_X0Y0_FrameData[20]
  PIN Tile_X0Y0_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 452.140 0.450 452.540 ;
    END
  END Tile_X0Y0_FrameData[21]
  PIN Tile_X0Y0_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 453.820 0.450 454.220 ;
    END
  END Tile_X0Y0_FrameData[22]
  PIN Tile_X0Y0_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 455.500 0.450 455.900 ;
    END
  END Tile_X0Y0_FrameData[23]
  PIN Tile_X0Y0_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 457.180 0.450 457.580 ;
    END
  END Tile_X0Y0_FrameData[24]
  PIN Tile_X0Y0_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 458.860 0.450 459.260 ;
    END
  END Tile_X0Y0_FrameData[25]
  PIN Tile_X0Y0_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 460.540 0.450 460.940 ;
    END
  END Tile_X0Y0_FrameData[26]
  PIN Tile_X0Y0_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 462.220 0.450 462.620 ;
    END
  END Tile_X0Y0_FrameData[27]
  PIN Tile_X0Y0_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 463.900 0.450 464.300 ;
    END
  END Tile_X0Y0_FrameData[28]
  PIN Tile_X0Y0_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 465.580 0.450 465.980 ;
    END
  END Tile_X0Y0_FrameData[29]
  PIN Tile_X0Y0_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 420.220 0.450 420.620 ;
    END
  END Tile_X0Y0_FrameData[2]
  PIN Tile_X0Y0_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 467.260 0.450 467.660 ;
    END
  END Tile_X0Y0_FrameData[30]
  PIN Tile_X0Y0_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 468.940 0.450 469.340 ;
    END
  END Tile_X0Y0_FrameData[31]
  PIN Tile_X0Y0_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 421.900 0.450 422.300 ;
    END
  END Tile_X0Y0_FrameData[3]
  PIN Tile_X0Y0_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 423.580 0.450 423.980 ;
    END
  END Tile_X0Y0_FrameData[4]
  PIN Tile_X0Y0_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 425.260 0.450 425.660 ;
    END
  END Tile_X0Y0_FrameData[5]
  PIN Tile_X0Y0_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 426.940 0.450 427.340 ;
    END
  END Tile_X0Y0_FrameData[6]
  PIN Tile_X0Y0_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 428.620 0.450 429.020 ;
    END
  END Tile_X0Y0_FrameData[7]
  PIN Tile_X0Y0_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 430.300 0.450 430.700 ;
    END
  END Tile_X0Y0_FrameData[8]
  PIN Tile_X0Y0_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 431.980 0.450 432.380 ;
    END
  END Tile_X0Y0_FrameData[9]
  PIN Tile_X0Y0_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 416.860 196.320 417.260 ;
    END
  END Tile_X0Y0_FrameData_O[0]
  PIN Tile_X0Y0_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 433.660 196.320 434.060 ;
    END
  END Tile_X0Y0_FrameData_O[10]
  PIN Tile_X0Y0_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 435.340 196.320 435.740 ;
    END
  END Tile_X0Y0_FrameData_O[11]
  PIN Tile_X0Y0_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 437.020 196.320 437.420 ;
    END
  END Tile_X0Y0_FrameData_O[12]
  PIN Tile_X0Y0_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 438.700 196.320 439.100 ;
    END
  END Tile_X0Y0_FrameData_O[13]
  PIN Tile_X0Y0_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 440.380 196.320 440.780 ;
    END
  END Tile_X0Y0_FrameData_O[14]
  PIN Tile_X0Y0_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 442.060 196.320 442.460 ;
    END
  END Tile_X0Y0_FrameData_O[15]
  PIN Tile_X0Y0_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 443.740 196.320 444.140 ;
    END
  END Tile_X0Y0_FrameData_O[16]
  PIN Tile_X0Y0_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 445.420 196.320 445.820 ;
    END
  END Tile_X0Y0_FrameData_O[17]
  PIN Tile_X0Y0_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 447.100 196.320 447.500 ;
    END
  END Tile_X0Y0_FrameData_O[18]
  PIN Tile_X0Y0_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 448.780 196.320 449.180 ;
    END
  END Tile_X0Y0_FrameData_O[19]
  PIN Tile_X0Y0_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 418.540 196.320 418.940 ;
    END
  END Tile_X0Y0_FrameData_O[1]
  PIN Tile_X0Y0_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 450.460 196.320 450.860 ;
    END
  END Tile_X0Y0_FrameData_O[20]
  PIN Tile_X0Y0_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 452.140 196.320 452.540 ;
    END
  END Tile_X0Y0_FrameData_O[21]
  PIN Tile_X0Y0_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 453.820 196.320 454.220 ;
    END
  END Tile_X0Y0_FrameData_O[22]
  PIN Tile_X0Y0_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 455.500 196.320 455.900 ;
    END
  END Tile_X0Y0_FrameData_O[23]
  PIN Tile_X0Y0_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 457.180 196.320 457.580 ;
    END
  END Tile_X0Y0_FrameData_O[24]
  PIN Tile_X0Y0_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 458.860 196.320 459.260 ;
    END
  END Tile_X0Y0_FrameData_O[25]
  PIN Tile_X0Y0_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 460.540 196.320 460.940 ;
    END
  END Tile_X0Y0_FrameData_O[26]
  PIN Tile_X0Y0_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 462.220 196.320 462.620 ;
    END
  END Tile_X0Y0_FrameData_O[27]
  PIN Tile_X0Y0_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 463.900 196.320 464.300 ;
    END
  END Tile_X0Y0_FrameData_O[28]
  PIN Tile_X0Y0_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 465.580 196.320 465.980 ;
    END
  END Tile_X0Y0_FrameData_O[29]
  PIN Tile_X0Y0_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 420.220 196.320 420.620 ;
    END
  END Tile_X0Y0_FrameData_O[2]
  PIN Tile_X0Y0_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 467.260 196.320 467.660 ;
    END
  END Tile_X0Y0_FrameData_O[30]
  PIN Tile_X0Y0_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 468.940 196.320 469.340 ;
    END
  END Tile_X0Y0_FrameData_O[31]
  PIN Tile_X0Y0_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 421.900 196.320 422.300 ;
    END
  END Tile_X0Y0_FrameData_O[3]
  PIN Tile_X0Y0_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 423.580 196.320 423.980 ;
    END
  END Tile_X0Y0_FrameData_O[4]
  PIN Tile_X0Y0_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 425.260 196.320 425.660 ;
    END
  END Tile_X0Y0_FrameData_O[5]
  PIN Tile_X0Y0_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 426.940 196.320 427.340 ;
    END
  END Tile_X0Y0_FrameData_O[6]
  PIN Tile_X0Y0_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 428.620 196.320 429.020 ;
    END
  END Tile_X0Y0_FrameData_O[7]
  PIN Tile_X0Y0_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 430.300 196.320 430.700 ;
    END
  END Tile_X0Y0_FrameData_O[8]
  PIN Tile_X0Y0_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 431.980 196.320 432.380 ;
    END
  END Tile_X0Y0_FrameData_O[9]
  PIN Tile_X0Y0_FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 138.520 483.440 138.920 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[0]
  PIN Tile_X0Y0_FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 148.120 483.440 148.520 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[10]
  PIN Tile_X0Y0_FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 149.080 483.440 149.480 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[11]
  PIN Tile_X0Y0_FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 150.040 483.440 150.440 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[12]
  PIN Tile_X0Y0_FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 151.000 483.440 151.400 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[13]
  PIN Tile_X0Y0_FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 151.960 483.440 152.360 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[14]
  PIN Tile_X0Y0_FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 152.920 483.440 153.320 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[15]
  PIN Tile_X0Y0_FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 153.880 483.440 154.280 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[16]
  PIN Tile_X0Y0_FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 154.840 483.440 155.240 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[17]
  PIN Tile_X0Y0_FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 155.800 483.440 156.200 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[18]
  PIN Tile_X0Y0_FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 156.760 483.440 157.160 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[19]
  PIN Tile_X0Y0_FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 139.480 483.440 139.880 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[1]
  PIN Tile_X0Y0_FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 140.440 483.440 140.840 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[2]
  PIN Tile_X0Y0_FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 141.400 483.440 141.800 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[3]
  PIN Tile_X0Y0_FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 142.360 483.440 142.760 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[4]
  PIN Tile_X0Y0_FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 143.320 483.440 143.720 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[5]
  PIN Tile_X0Y0_FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 144.280 483.440 144.680 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[6]
  PIN Tile_X0Y0_FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 145.240 483.440 145.640 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[7]
  PIN Tile_X0Y0_FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 146.200 483.440 146.600 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[8]
  PIN Tile_X0Y0_FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 147.160 483.440 147.560 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[9]
  PIN Tile_X0Y0_N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 37.720 483.440 38.120 483.840 ;
    END
  END Tile_X0Y0_N1BEG[0]
  PIN Tile_X0Y0_N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 38.680 483.440 39.080 483.840 ;
    END
  END Tile_X0Y0_N1BEG[1]
  PIN Tile_X0Y0_N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 39.640 483.440 40.040 483.840 ;
    END
  END Tile_X0Y0_N1BEG[2]
  PIN Tile_X0Y0_N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.827200 ;
    PORT
      LAYER Metal3 ;
        RECT 40.600 483.440 41.000 483.840 ;
    END
  END Tile_X0Y0_N1BEG[3]
  PIN Tile_X0Y0_N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 41.560 483.440 41.960 483.840 ;
    END
  END Tile_X0Y0_N2BEG[0]
  PIN Tile_X0Y0_N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 42.520 483.440 42.920 483.840 ;
    END
  END Tile_X0Y0_N2BEG[1]
  PIN Tile_X0Y0_N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 43.480 483.440 43.880 483.840 ;
    END
  END Tile_X0Y0_N2BEG[2]
  PIN Tile_X0Y0_N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 44.440 483.440 44.840 483.840 ;
    END
  END Tile_X0Y0_N2BEG[3]
  PIN Tile_X0Y0_N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 45.400 483.440 45.800 483.840 ;
    END
  END Tile_X0Y0_N2BEG[4]
  PIN Tile_X0Y0_N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 46.360 483.440 46.760 483.840 ;
    END
  END Tile_X0Y0_N2BEG[5]
  PIN Tile_X0Y0_N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 47.320 483.440 47.720 483.840 ;
    END
  END Tile_X0Y0_N2BEG[6]
  PIN Tile_X0Y0_N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 48.280 483.440 48.680 483.840 ;
    END
  END Tile_X0Y0_N2BEG[7]
  PIN Tile_X0Y0_N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 49.240 483.440 49.640 483.840 ;
    END
  END Tile_X0Y0_N2BEGb[0]
  PIN Tile_X0Y0_N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 50.200 483.440 50.600 483.840 ;
    END
  END Tile_X0Y0_N2BEGb[1]
  PIN Tile_X0Y0_N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 51.160 483.440 51.560 483.840 ;
    END
  END Tile_X0Y0_N2BEGb[2]
  PIN Tile_X0Y0_N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 52.120 483.440 52.520 483.840 ;
    END
  END Tile_X0Y0_N2BEGb[3]
  PIN Tile_X0Y0_N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.827200 ;
    PORT
      LAYER Metal3 ;
        RECT 53.080 483.440 53.480 483.840 ;
    END
  END Tile_X0Y0_N2BEGb[4]
  PIN Tile_X0Y0_N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 54.040 483.440 54.440 483.840 ;
    END
  END Tile_X0Y0_N2BEGb[5]
  PIN Tile_X0Y0_N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 55.000 483.440 55.400 483.840 ;
    END
  END Tile_X0Y0_N2BEGb[6]
  PIN Tile_X0Y0_N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 55.960 483.440 56.360 483.840 ;
    END
  END Tile_X0Y0_N2BEGb[7]
  PIN Tile_X0Y0_N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 56.920 483.440 57.320 483.840 ;
    END
  END Tile_X0Y0_N4BEG[0]
  PIN Tile_X0Y0_N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 66.520 483.440 66.920 483.840 ;
    END
  END Tile_X0Y0_N4BEG[10]
  PIN Tile_X0Y0_N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 67.480 483.440 67.880 483.840 ;
    END
  END Tile_X0Y0_N4BEG[11]
  PIN Tile_X0Y0_N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 68.440 483.440 68.840 483.840 ;
    END
  END Tile_X0Y0_N4BEG[12]
  PIN Tile_X0Y0_N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 69.400 483.440 69.800 483.840 ;
    END
  END Tile_X0Y0_N4BEG[13]
  PIN Tile_X0Y0_N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 70.360 483.440 70.760 483.840 ;
    END
  END Tile_X0Y0_N4BEG[14]
  PIN Tile_X0Y0_N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 71.320 483.440 71.720 483.840 ;
    END
  END Tile_X0Y0_N4BEG[15]
  PIN Tile_X0Y0_N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 57.880 483.440 58.280 483.840 ;
    END
  END Tile_X0Y0_N4BEG[1]
  PIN Tile_X0Y0_N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 58.840 483.440 59.240 483.840 ;
    END
  END Tile_X0Y0_N4BEG[2]
  PIN Tile_X0Y0_N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 59.800 483.440 60.200 483.840 ;
    END
  END Tile_X0Y0_N4BEG[3]
  PIN Tile_X0Y0_N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 60.760 483.440 61.160 483.840 ;
    END
  END Tile_X0Y0_N4BEG[4]
  PIN Tile_X0Y0_N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 61.720 483.440 62.120 483.840 ;
    END
  END Tile_X0Y0_N4BEG[5]
  PIN Tile_X0Y0_N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 62.680 483.440 63.080 483.840 ;
    END
  END Tile_X0Y0_N4BEG[6]
  PIN Tile_X0Y0_N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 63.640 483.440 64.040 483.840 ;
    END
  END Tile_X0Y0_N4BEG[7]
  PIN Tile_X0Y0_N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 64.600 483.440 65.000 483.840 ;
    END
  END Tile_X0Y0_N4BEG[8]
  PIN Tile_X0Y0_N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 65.560 483.440 65.960 483.840 ;
    END
  END Tile_X0Y0_N4BEG[9]
  PIN Tile_X0Y0_NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 72.280 483.440 72.680 483.840 ;
    END
  END Tile_X0Y0_NN4BEG[0]
  PIN Tile_X0Y0_NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 81.880 483.440 82.280 483.840 ;
    END
  END Tile_X0Y0_NN4BEG[10]
  PIN Tile_X0Y0_NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 82.840 483.440 83.240 483.840 ;
    END
  END Tile_X0Y0_NN4BEG[11]
  PIN Tile_X0Y0_NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 83.800 483.440 84.200 483.840 ;
    END
  END Tile_X0Y0_NN4BEG[12]
  PIN Tile_X0Y0_NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 84.760 483.440 85.160 483.840 ;
    END
  END Tile_X0Y0_NN4BEG[13]
  PIN Tile_X0Y0_NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 85.720 483.440 86.120 483.840 ;
    END
  END Tile_X0Y0_NN4BEG[14]
  PIN Tile_X0Y0_NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 86.680 483.440 87.080 483.840 ;
    END
  END Tile_X0Y0_NN4BEG[15]
  PIN Tile_X0Y0_NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 73.240 483.440 73.640 483.840 ;
    END
  END Tile_X0Y0_NN4BEG[1]
  PIN Tile_X0Y0_NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 74.200 483.440 74.600 483.840 ;
    END
  END Tile_X0Y0_NN4BEG[2]
  PIN Tile_X0Y0_NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 75.160 483.440 75.560 483.840 ;
    END
  END Tile_X0Y0_NN4BEG[3]
  PIN Tile_X0Y0_NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 76.120 483.440 76.520 483.840 ;
    END
  END Tile_X0Y0_NN4BEG[4]
  PIN Tile_X0Y0_NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 77.080 483.440 77.480 483.840 ;
    END
  END Tile_X0Y0_NN4BEG[5]
  PIN Tile_X0Y0_NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 78.040 483.440 78.440 483.840 ;
    END
  END Tile_X0Y0_NN4BEG[6]
  PIN Tile_X0Y0_NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 79.000 483.440 79.400 483.840 ;
    END
  END Tile_X0Y0_NN4BEG[7]
  PIN Tile_X0Y0_NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 79.960 483.440 80.360 483.840 ;
    END
  END Tile_X0Y0_NN4BEG[8]
  PIN Tile_X0Y0_NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 80.920 483.440 81.320 483.840 ;
    END
  END Tile_X0Y0_NN4BEG[9]
  PIN Tile_X0Y0_S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 87.640 483.440 88.040 483.840 ;
    END
  END Tile_X0Y0_S1END[0]
  PIN Tile_X0Y0_S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 88.600 483.440 89.000 483.840 ;
    END
  END Tile_X0Y0_S1END[1]
  PIN Tile_X0Y0_S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 89.560 483.440 89.960 483.840 ;
    END
  END Tile_X0Y0_S1END[2]
  PIN Tile_X0Y0_S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 90.520 483.440 90.920 483.840 ;
    END
  END Tile_X0Y0_S1END[3]
  PIN Tile_X0Y0_S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 99.160 483.440 99.560 483.840 ;
    END
  END Tile_X0Y0_S2END[0]
  PIN Tile_X0Y0_S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 100.120 483.440 100.520 483.840 ;
    END
  END Tile_X0Y0_S2END[1]
  PIN Tile_X0Y0_S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.450800 ;
    PORT
      LAYER Metal3 ;
        RECT 101.080 483.440 101.480 483.840 ;
    END
  END Tile_X0Y0_S2END[2]
  PIN Tile_X0Y0_S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 102.040 483.440 102.440 483.840 ;
    END
  END Tile_X0Y0_S2END[3]
  PIN Tile_X0Y0_S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 103.000 483.440 103.400 483.840 ;
    END
  END Tile_X0Y0_S2END[4]
  PIN Tile_X0Y0_S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 103.960 483.440 104.360 483.840 ;
    END
  END Tile_X0Y0_S2END[5]
  PIN Tile_X0Y0_S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 104.920 483.440 105.320 483.840 ;
    END
  END Tile_X0Y0_S2END[6]
  PIN Tile_X0Y0_S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 105.880 483.440 106.280 483.840 ;
    END
  END Tile_X0Y0_S2END[7]
  PIN Tile_X0Y0_S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 91.480 483.440 91.880 483.840 ;
    END
  END Tile_X0Y0_S2MID[0]
  PIN Tile_X0Y0_S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 92.440 483.440 92.840 483.840 ;
    END
  END Tile_X0Y0_S2MID[1]
  PIN Tile_X0Y0_S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 93.400 483.440 93.800 483.840 ;
    END
  END Tile_X0Y0_S2MID[2]
  PIN Tile_X0Y0_S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 94.360 483.440 94.760 483.840 ;
    END
  END Tile_X0Y0_S2MID[3]
  PIN Tile_X0Y0_S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 95.320 483.440 95.720 483.840 ;
    END
  END Tile_X0Y0_S2MID[4]
  PIN Tile_X0Y0_S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 96.280 483.440 96.680 483.840 ;
    END
  END Tile_X0Y0_S2MID[5]
  PIN Tile_X0Y0_S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 97.240 483.440 97.640 483.840 ;
    END
  END Tile_X0Y0_S2MID[6]
  PIN Tile_X0Y0_S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 98.200 483.440 98.600 483.840 ;
    END
  END Tile_X0Y0_S2MID[7]
  PIN Tile_X0Y0_S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 106.840 483.440 107.240 483.840 ;
    END
  END Tile_X0Y0_S4END[0]
  PIN Tile_X0Y0_S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 116.440 483.440 116.840 483.840 ;
    END
  END Tile_X0Y0_S4END[10]
  PIN Tile_X0Y0_S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 117.400 483.440 117.800 483.840 ;
    END
  END Tile_X0Y0_S4END[11]
  PIN Tile_X0Y0_S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 118.360 483.440 118.760 483.840 ;
    END
  END Tile_X0Y0_S4END[12]
  PIN Tile_X0Y0_S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 119.320 483.440 119.720 483.840 ;
    END
  END Tile_X0Y0_S4END[13]
  PIN Tile_X0Y0_S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 120.280 483.440 120.680 483.840 ;
    END
  END Tile_X0Y0_S4END[14]
  PIN Tile_X0Y0_S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 121.240 483.440 121.640 483.840 ;
    END
  END Tile_X0Y0_S4END[15]
  PIN Tile_X0Y0_S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 107.800 483.440 108.200 483.840 ;
    END
  END Tile_X0Y0_S4END[1]
  PIN Tile_X0Y0_S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 108.760 483.440 109.160 483.840 ;
    END
  END Tile_X0Y0_S4END[2]
  PIN Tile_X0Y0_S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 109.720 483.440 110.120 483.840 ;
    END
  END Tile_X0Y0_S4END[3]
  PIN Tile_X0Y0_S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 110.680 483.440 111.080 483.840 ;
    END
  END Tile_X0Y0_S4END[4]
  PIN Tile_X0Y0_S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 111.640 483.440 112.040 483.840 ;
    END
  END Tile_X0Y0_S4END[5]
  PIN Tile_X0Y0_S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 112.600 483.440 113.000 483.840 ;
    END
  END Tile_X0Y0_S4END[6]
  PIN Tile_X0Y0_S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 113.560 483.440 113.960 483.840 ;
    END
  END Tile_X0Y0_S4END[7]
  PIN Tile_X0Y0_S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 114.520 483.440 114.920 483.840 ;
    END
  END Tile_X0Y0_S4END[8]
  PIN Tile_X0Y0_S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 115.480 483.440 115.880 483.840 ;
    END
  END Tile_X0Y0_S4END[9]
  PIN Tile_X0Y0_SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 122.200 483.440 122.600 483.840 ;
    END
  END Tile_X0Y0_SS4END[0]
  PIN Tile_X0Y0_SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 131.800 483.440 132.200 483.840 ;
    END
  END Tile_X0Y0_SS4END[10]
  PIN Tile_X0Y0_SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 132.760 483.440 133.160 483.840 ;
    END
  END Tile_X0Y0_SS4END[11]
  PIN Tile_X0Y0_SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 133.720 483.440 134.120 483.840 ;
    END
  END Tile_X0Y0_SS4END[12]
  PIN Tile_X0Y0_SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 134.680 483.440 135.080 483.840 ;
    END
  END Tile_X0Y0_SS4END[13]
  PIN Tile_X0Y0_SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 135.640 483.440 136.040 483.840 ;
    END
  END Tile_X0Y0_SS4END[14]
  PIN Tile_X0Y0_SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 136.600 483.440 137.000 483.840 ;
    END
  END Tile_X0Y0_SS4END[15]
  PIN Tile_X0Y0_SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 123.160 483.440 123.560 483.840 ;
    END
  END Tile_X0Y0_SS4END[1]
  PIN Tile_X0Y0_SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 124.120 483.440 124.520 483.840 ;
    END
  END Tile_X0Y0_SS4END[2]
  PIN Tile_X0Y0_SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 125.080 483.440 125.480 483.840 ;
    END
  END Tile_X0Y0_SS4END[3]
  PIN Tile_X0Y0_SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 126.040 483.440 126.440 483.840 ;
    END
  END Tile_X0Y0_SS4END[4]
  PIN Tile_X0Y0_SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 127.000 483.440 127.400 483.840 ;
    END
  END Tile_X0Y0_SS4END[5]
  PIN Tile_X0Y0_SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 127.960 483.440 128.360 483.840 ;
    END
  END Tile_X0Y0_SS4END[6]
  PIN Tile_X0Y0_SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 128.920 483.440 129.320 483.840 ;
    END
  END Tile_X0Y0_SS4END[7]
  PIN Tile_X0Y0_SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 129.880 483.440 130.280 483.840 ;
    END
  END Tile_X0Y0_SS4END[8]
  PIN Tile_X0Y0_SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 130.840 483.440 131.240 483.840 ;
    END
  END Tile_X0Y0_SS4END[9]
  PIN Tile_X0Y0_UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 137.560 483.440 137.960 483.840 ;
    END
  END Tile_X0Y0_UserCLKo
  PIN Tile_X0Y0_W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 255.580 0.450 255.980 ;
    END
  END Tile_X0Y0_W1BEG[0]
  PIN Tile_X0Y0_W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 257.260 0.450 257.660 ;
    END
  END Tile_X0Y0_W1BEG[1]
  PIN Tile_X0Y0_W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 258.940 0.450 259.340 ;
    END
  END Tile_X0Y0_W1BEG[2]
  PIN Tile_X0Y0_W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 260.620 0.450 261.020 ;
    END
  END Tile_X0Y0_W1BEG[3]
  PIN Tile_X0Y0_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 255.580 196.320 255.980 ;
    END
  END Tile_X0Y0_W1END[0]
  PIN Tile_X0Y0_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 257.260 196.320 257.660 ;
    END
  END Tile_X0Y0_W1END[1]
  PIN Tile_X0Y0_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 258.940 196.320 259.340 ;
    END
  END Tile_X0Y0_W1END[2]
  PIN Tile_X0Y0_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 260.620 196.320 261.020 ;
    END
  END Tile_X0Y0_W1END[3]
  PIN Tile_X0Y0_W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 262.300 0.450 262.700 ;
    END
  END Tile_X0Y0_W2BEG[0]
  PIN Tile_X0Y0_W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 263.980 0.450 264.380 ;
    END
  END Tile_X0Y0_W2BEG[1]
  PIN Tile_X0Y0_W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 265.660 0.450 266.060 ;
    END
  END Tile_X0Y0_W2BEG[2]
  PIN Tile_X0Y0_W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 267.340 0.450 267.740 ;
    END
  END Tile_X0Y0_W2BEG[3]
  PIN Tile_X0Y0_W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 269.020 0.450 269.420 ;
    END
  END Tile_X0Y0_W2BEG[4]
  PIN Tile_X0Y0_W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 270.700 0.450 271.100 ;
    END
  END Tile_X0Y0_W2BEG[5]
  PIN Tile_X0Y0_W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 272.380 0.450 272.780 ;
    END
  END Tile_X0Y0_W2BEG[6]
  PIN Tile_X0Y0_W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 274.060 0.450 274.460 ;
    END
  END Tile_X0Y0_W2BEG[7]
  PIN Tile_X0Y0_W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 275.740 0.450 276.140 ;
    END
  END Tile_X0Y0_W2BEGb[0]
  PIN Tile_X0Y0_W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 277.420 0.450 277.820 ;
    END
  END Tile_X0Y0_W2BEGb[1]
  PIN Tile_X0Y0_W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 279.100 0.450 279.500 ;
    END
  END Tile_X0Y0_W2BEGb[2]
  PIN Tile_X0Y0_W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 280.780 0.450 281.180 ;
    END
  END Tile_X0Y0_W2BEGb[3]
  PIN Tile_X0Y0_W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 282.460 0.450 282.860 ;
    END
  END Tile_X0Y0_W2BEGb[4]
  PIN Tile_X0Y0_W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 284.140 0.450 284.540 ;
    END
  END Tile_X0Y0_W2BEGb[5]
  PIN Tile_X0Y0_W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 285.820 0.450 286.220 ;
    END
  END Tile_X0Y0_W2BEGb[6]
  PIN Tile_X0Y0_W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 287.500 0.450 287.900 ;
    END
  END Tile_X0Y0_W2BEGb[7]
  PIN Tile_X0Y0_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 275.740 196.320 276.140 ;
    END
  END Tile_X0Y0_W2END[0]
  PIN Tile_X0Y0_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 277.420 196.320 277.820 ;
    END
  END Tile_X0Y0_W2END[1]
  PIN Tile_X0Y0_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 279.100 196.320 279.500 ;
    END
  END Tile_X0Y0_W2END[2]
  PIN Tile_X0Y0_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 280.780 196.320 281.180 ;
    END
  END Tile_X0Y0_W2END[3]
  PIN Tile_X0Y0_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 282.460 196.320 282.860 ;
    END
  END Tile_X0Y0_W2END[4]
  PIN Tile_X0Y0_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 284.140 196.320 284.540 ;
    END
  END Tile_X0Y0_W2END[5]
  PIN Tile_X0Y0_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 285.820 196.320 286.220 ;
    END
  END Tile_X0Y0_W2END[6]
  PIN Tile_X0Y0_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 287.500 196.320 287.900 ;
    END
  END Tile_X0Y0_W2END[7]
  PIN Tile_X0Y0_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 262.300 196.320 262.700 ;
    END
  END Tile_X0Y0_W2MID[0]
  PIN Tile_X0Y0_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 263.980 196.320 264.380 ;
    END
  END Tile_X0Y0_W2MID[1]
  PIN Tile_X0Y0_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 265.660 196.320 266.060 ;
    END
  END Tile_X0Y0_W2MID[2]
  PIN Tile_X0Y0_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 267.340 196.320 267.740 ;
    END
  END Tile_X0Y0_W2MID[3]
  PIN Tile_X0Y0_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 269.020 196.320 269.420 ;
    END
  END Tile_X0Y0_W2MID[4]
  PIN Tile_X0Y0_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 270.700 196.320 271.100 ;
    END
  END Tile_X0Y0_W2MID[5]
  PIN Tile_X0Y0_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 272.380 196.320 272.780 ;
    END
  END Tile_X0Y0_W2MID[6]
  PIN Tile_X0Y0_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 274.060 196.320 274.460 ;
    END
  END Tile_X0Y0_W2MID[7]
  PIN Tile_X0Y0_W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 316.060 0.450 316.460 ;
    END
  END Tile_X0Y0_W6BEG[0]
  PIN Tile_X0Y0_W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 332.860 0.450 333.260 ;
    END
  END Tile_X0Y0_W6BEG[10]
  PIN Tile_X0Y0_W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 334.540 0.450 334.940 ;
    END
  END Tile_X0Y0_W6BEG[11]
  PIN Tile_X0Y0_W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 317.740 0.450 318.140 ;
    END
  END Tile_X0Y0_W6BEG[1]
  PIN Tile_X0Y0_W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 319.420 0.450 319.820 ;
    END
  END Tile_X0Y0_W6BEG[2]
  PIN Tile_X0Y0_W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 321.100 0.450 321.500 ;
    END
  END Tile_X0Y0_W6BEG[3]
  PIN Tile_X0Y0_W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 322.780 0.450 323.180 ;
    END
  END Tile_X0Y0_W6BEG[4]
  PIN Tile_X0Y0_W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 324.460 0.450 324.860 ;
    END
  END Tile_X0Y0_W6BEG[5]
  PIN Tile_X0Y0_W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 326.140 0.450 326.540 ;
    END
  END Tile_X0Y0_W6BEG[6]
  PIN Tile_X0Y0_W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 327.820 0.450 328.220 ;
    END
  END Tile_X0Y0_W6BEG[7]
  PIN Tile_X0Y0_W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 329.500 0.450 329.900 ;
    END
  END Tile_X0Y0_W6BEG[8]
  PIN Tile_X0Y0_W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 331.180 0.450 331.580 ;
    END
  END Tile_X0Y0_W6BEG[9]
  PIN Tile_X0Y0_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 316.060 196.320 316.460 ;
    END
  END Tile_X0Y0_W6END[0]
  PIN Tile_X0Y0_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 332.860 196.320 333.260 ;
    END
  END Tile_X0Y0_W6END[10]
  PIN Tile_X0Y0_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 334.540 196.320 334.940 ;
    END
  END Tile_X0Y0_W6END[11]
  PIN Tile_X0Y0_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 317.740 196.320 318.140 ;
    END
  END Tile_X0Y0_W6END[1]
  PIN Tile_X0Y0_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 319.420 196.320 319.820 ;
    END
  END Tile_X0Y0_W6END[2]
  PIN Tile_X0Y0_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 321.100 196.320 321.500 ;
    END
  END Tile_X0Y0_W6END[3]
  PIN Tile_X0Y0_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 322.780 196.320 323.180 ;
    END
  END Tile_X0Y0_W6END[4]
  PIN Tile_X0Y0_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 324.460 196.320 324.860 ;
    END
  END Tile_X0Y0_W6END[5]
  PIN Tile_X0Y0_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 326.140 196.320 326.540 ;
    END
  END Tile_X0Y0_W6END[6]
  PIN Tile_X0Y0_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 327.820 196.320 328.220 ;
    END
  END Tile_X0Y0_W6END[7]
  PIN Tile_X0Y0_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 329.500 196.320 329.900 ;
    END
  END Tile_X0Y0_W6END[8]
  PIN Tile_X0Y0_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 331.180 196.320 331.580 ;
    END
  END Tile_X0Y0_W6END[9]
  PIN Tile_X0Y0_WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 289.180 0.450 289.580 ;
    END
  END Tile_X0Y0_WW4BEG[0]
  PIN Tile_X0Y0_WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 305.980 0.450 306.380 ;
    END
  END Tile_X0Y0_WW4BEG[10]
  PIN Tile_X0Y0_WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 307.660 0.450 308.060 ;
    END
  END Tile_X0Y0_WW4BEG[11]
  PIN Tile_X0Y0_WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 309.340 0.450 309.740 ;
    END
  END Tile_X0Y0_WW4BEG[12]
  PIN Tile_X0Y0_WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 311.020 0.450 311.420 ;
    END
  END Tile_X0Y0_WW4BEG[13]
  PIN Tile_X0Y0_WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 312.700 0.450 313.100 ;
    END
  END Tile_X0Y0_WW4BEG[14]
  PIN Tile_X0Y0_WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.827200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 314.380 0.450 314.780 ;
    END
  END Tile_X0Y0_WW4BEG[15]
  PIN Tile_X0Y0_WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 290.860 0.450 291.260 ;
    END
  END Tile_X0Y0_WW4BEG[1]
  PIN Tile_X0Y0_WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 292.540 0.450 292.940 ;
    END
  END Tile_X0Y0_WW4BEG[2]
  PIN Tile_X0Y0_WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 294.220 0.450 294.620 ;
    END
  END Tile_X0Y0_WW4BEG[3]
  PIN Tile_X0Y0_WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 295.900 0.450 296.300 ;
    END
  END Tile_X0Y0_WW4BEG[4]
  PIN Tile_X0Y0_WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 297.580 0.450 297.980 ;
    END
  END Tile_X0Y0_WW4BEG[5]
  PIN Tile_X0Y0_WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 299.260 0.450 299.660 ;
    END
  END Tile_X0Y0_WW4BEG[6]
  PIN Tile_X0Y0_WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 300.940 0.450 301.340 ;
    END
  END Tile_X0Y0_WW4BEG[7]
  PIN Tile_X0Y0_WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 302.620 0.450 303.020 ;
    END
  END Tile_X0Y0_WW4BEG[8]
  PIN Tile_X0Y0_WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 304.300 0.450 304.700 ;
    END
  END Tile_X0Y0_WW4BEG[9]
  PIN Tile_X0Y0_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 289.180 196.320 289.580 ;
    END
  END Tile_X0Y0_WW4END[0]
  PIN Tile_X0Y0_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 305.980 196.320 306.380 ;
    END
  END Tile_X0Y0_WW4END[10]
  PIN Tile_X0Y0_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 307.660 196.320 308.060 ;
    END
  END Tile_X0Y0_WW4END[11]
  PIN Tile_X0Y0_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 309.340 196.320 309.740 ;
    END
  END Tile_X0Y0_WW4END[12]
  PIN Tile_X0Y0_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 311.020 196.320 311.420 ;
    END
  END Tile_X0Y0_WW4END[13]
  PIN Tile_X0Y0_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 312.700 196.320 313.100 ;
    END
  END Tile_X0Y0_WW4END[14]
  PIN Tile_X0Y0_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 314.380 196.320 314.780 ;
    END
  END Tile_X0Y0_WW4END[15]
  PIN Tile_X0Y0_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 290.860 196.320 291.260 ;
    END
  END Tile_X0Y0_WW4END[1]
  PIN Tile_X0Y0_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 292.540 196.320 292.940 ;
    END
  END Tile_X0Y0_WW4END[2]
  PIN Tile_X0Y0_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 294.220 196.320 294.620 ;
    END
  END Tile_X0Y0_WW4END[3]
  PIN Tile_X0Y0_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 295.900 196.320 296.300 ;
    END
  END Tile_X0Y0_WW4END[4]
  PIN Tile_X0Y0_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 297.580 196.320 297.980 ;
    END
  END Tile_X0Y0_WW4END[5]
  PIN Tile_X0Y0_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 299.260 196.320 299.660 ;
    END
  END Tile_X0Y0_WW4END[6]
  PIN Tile_X0Y0_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 300.940 196.320 301.340 ;
    END
  END Tile_X0Y0_WW4END[7]
  PIN Tile_X0Y0_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 302.620 196.320 303.020 ;
    END
  END Tile_X0Y0_WW4END[8]
  PIN Tile_X0Y0_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 304.300 196.320 304.700 ;
    END
  END Tile_X0Y0_WW4END[9]
  PIN Tile_X0Y1_E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 94.300 196.320 94.700 ;
    END
  END Tile_X0Y1_E1BEG[0]
  PIN Tile_X0Y1_E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 95.980 196.320 96.380 ;
    END
  END Tile_X0Y1_E1BEG[1]
  PIN Tile_X0Y1_E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 97.660 196.320 98.060 ;
    END
  END Tile_X0Y1_E1BEG[2]
  PIN Tile_X0Y1_E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 99.340 196.320 99.740 ;
    END
  END Tile_X0Y1_E1BEG[3]
  PIN Tile_X0Y1_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 94.300 0.450 94.700 ;
    END
  END Tile_X0Y1_E1END[0]
  PIN Tile_X0Y1_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 95.980 0.450 96.380 ;
    END
  END Tile_X0Y1_E1END[1]
  PIN Tile_X0Y1_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 97.660 0.450 98.060 ;
    END
  END Tile_X0Y1_E1END[2]
  PIN Tile_X0Y1_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 99.340 0.450 99.740 ;
    END
  END Tile_X0Y1_E1END[3]
  PIN Tile_X0Y1_E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 101.020 196.320 101.420 ;
    END
  END Tile_X0Y1_E2BEG[0]
  PIN Tile_X0Y1_E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 102.700 196.320 103.100 ;
    END
  END Tile_X0Y1_E2BEG[1]
  PIN Tile_X0Y1_E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 104.380 196.320 104.780 ;
    END
  END Tile_X0Y1_E2BEG[2]
  PIN Tile_X0Y1_E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 106.060 196.320 106.460 ;
    END
  END Tile_X0Y1_E2BEG[3]
  PIN Tile_X0Y1_E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 107.740 196.320 108.140 ;
    END
  END Tile_X0Y1_E2BEG[4]
  PIN Tile_X0Y1_E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 109.420 196.320 109.820 ;
    END
  END Tile_X0Y1_E2BEG[5]
  PIN Tile_X0Y1_E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 111.100 196.320 111.500 ;
    END
  END Tile_X0Y1_E2BEG[6]
  PIN Tile_X0Y1_E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.827200 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 112.780 196.320 113.180 ;
    END
  END Tile_X0Y1_E2BEG[7]
  PIN Tile_X0Y1_E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 114.460 196.320 114.860 ;
    END
  END Tile_X0Y1_E2BEGb[0]
  PIN Tile_X0Y1_E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 116.140 196.320 116.540 ;
    END
  END Tile_X0Y1_E2BEGb[1]
  PIN Tile_X0Y1_E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 117.820 196.320 118.220 ;
    END
  END Tile_X0Y1_E2BEGb[2]
  PIN Tile_X0Y1_E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 119.500 196.320 119.900 ;
    END
  END Tile_X0Y1_E2BEGb[3]
  PIN Tile_X0Y1_E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 121.180 196.320 121.580 ;
    END
  END Tile_X0Y1_E2BEGb[4]
  PIN Tile_X0Y1_E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 122.860 196.320 123.260 ;
    END
  END Tile_X0Y1_E2BEGb[5]
  PIN Tile_X0Y1_E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 124.540 196.320 124.940 ;
    END
  END Tile_X0Y1_E2BEGb[6]
  PIN Tile_X0Y1_E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 126.220 196.320 126.620 ;
    END
  END Tile_X0Y1_E2BEGb[7]
  PIN Tile_X0Y1_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 114.460 0.450 114.860 ;
    END
  END Tile_X0Y1_E2END[0]
  PIN Tile_X0Y1_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 116.140 0.450 116.540 ;
    END
  END Tile_X0Y1_E2END[1]
  PIN Tile_X0Y1_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 117.820 0.450 118.220 ;
    END
  END Tile_X0Y1_E2END[2]
  PIN Tile_X0Y1_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 119.500 0.450 119.900 ;
    END
  END Tile_X0Y1_E2END[3]
  PIN Tile_X0Y1_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 121.180 0.450 121.580 ;
    END
  END Tile_X0Y1_E2END[4]
  PIN Tile_X0Y1_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 122.860 0.450 123.260 ;
    END
  END Tile_X0Y1_E2END[5]
  PIN Tile_X0Y1_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 124.540 0.450 124.940 ;
    END
  END Tile_X0Y1_E2END[6]
  PIN Tile_X0Y1_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 126.220 0.450 126.620 ;
    END
  END Tile_X0Y1_E2END[7]
  PIN Tile_X0Y1_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 101.020 0.450 101.420 ;
    END
  END Tile_X0Y1_E2MID[0]
  PIN Tile_X0Y1_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 102.700 0.450 103.100 ;
    END
  END Tile_X0Y1_E2MID[1]
  PIN Tile_X0Y1_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 104.380 0.450 104.780 ;
    END
  END Tile_X0Y1_E2MID[2]
  PIN Tile_X0Y1_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 106.060 0.450 106.460 ;
    END
  END Tile_X0Y1_E2MID[3]
  PIN Tile_X0Y1_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 107.740 0.450 108.140 ;
    END
  END Tile_X0Y1_E2MID[4]
  PIN Tile_X0Y1_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 109.420 0.450 109.820 ;
    END
  END Tile_X0Y1_E2MID[5]
  PIN Tile_X0Y1_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 111.100 0.450 111.500 ;
    END
  END Tile_X0Y1_E2MID[6]
  PIN Tile_X0Y1_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 112.780 0.450 113.180 ;
    END
  END Tile_X0Y1_E2MID[7]
  PIN Tile_X0Y1_E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 154.780 196.320 155.180 ;
    END
  END Tile_X0Y1_E6BEG[0]
  PIN Tile_X0Y1_E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.827200 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 171.580 196.320 171.980 ;
    END
  END Tile_X0Y1_E6BEG[10]
  PIN Tile_X0Y1_E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 173.260 196.320 173.660 ;
    END
  END Tile_X0Y1_E6BEG[11]
  PIN Tile_X0Y1_E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 156.460 196.320 156.860 ;
    END
  END Tile_X0Y1_E6BEG[1]
  PIN Tile_X0Y1_E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 158.140 196.320 158.540 ;
    END
  END Tile_X0Y1_E6BEG[2]
  PIN Tile_X0Y1_E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 159.820 196.320 160.220 ;
    END
  END Tile_X0Y1_E6BEG[3]
  PIN Tile_X0Y1_E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 161.500 196.320 161.900 ;
    END
  END Tile_X0Y1_E6BEG[4]
  PIN Tile_X0Y1_E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 163.180 196.320 163.580 ;
    END
  END Tile_X0Y1_E6BEG[5]
  PIN Tile_X0Y1_E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 164.860 196.320 165.260 ;
    END
  END Tile_X0Y1_E6BEG[6]
  PIN Tile_X0Y1_E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 166.540 196.320 166.940 ;
    END
  END Tile_X0Y1_E6BEG[7]
  PIN Tile_X0Y1_E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 168.220 196.320 168.620 ;
    END
  END Tile_X0Y1_E6BEG[8]
  PIN Tile_X0Y1_E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 169.900 196.320 170.300 ;
    END
  END Tile_X0Y1_E6BEG[9]
  PIN Tile_X0Y1_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 154.780 0.450 155.180 ;
    END
  END Tile_X0Y1_E6END[0]
  PIN Tile_X0Y1_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 171.580 0.450 171.980 ;
    END
  END Tile_X0Y1_E6END[10]
  PIN Tile_X0Y1_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 173.260 0.450 173.660 ;
    END
  END Tile_X0Y1_E6END[11]
  PIN Tile_X0Y1_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 156.460 0.450 156.860 ;
    END
  END Tile_X0Y1_E6END[1]
  PIN Tile_X0Y1_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 158.140 0.450 158.540 ;
    END
  END Tile_X0Y1_E6END[2]
  PIN Tile_X0Y1_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 159.820 0.450 160.220 ;
    END
  END Tile_X0Y1_E6END[3]
  PIN Tile_X0Y1_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 161.500 0.450 161.900 ;
    END
  END Tile_X0Y1_E6END[4]
  PIN Tile_X0Y1_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 163.180 0.450 163.580 ;
    END
  END Tile_X0Y1_E6END[5]
  PIN Tile_X0Y1_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 164.860 0.450 165.260 ;
    END
  END Tile_X0Y1_E6END[6]
  PIN Tile_X0Y1_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 166.540 0.450 166.940 ;
    END
  END Tile_X0Y1_E6END[7]
  PIN Tile_X0Y1_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 168.220 0.450 168.620 ;
    END
  END Tile_X0Y1_E6END[8]
  PIN Tile_X0Y1_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 169.900 0.450 170.300 ;
    END
  END Tile_X0Y1_E6END[9]
  PIN Tile_X0Y1_EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 127.900 196.320 128.300 ;
    END
  END Tile_X0Y1_EE4BEG[0]
  PIN Tile_X0Y1_EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 144.700 196.320 145.100 ;
    END
  END Tile_X0Y1_EE4BEG[10]
  PIN Tile_X0Y1_EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 146.380 196.320 146.780 ;
    END
  END Tile_X0Y1_EE4BEG[11]
  PIN Tile_X0Y1_EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 148.060 196.320 148.460 ;
    END
  END Tile_X0Y1_EE4BEG[12]
  PIN Tile_X0Y1_EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 149.740 196.320 150.140 ;
    END
  END Tile_X0Y1_EE4BEG[13]
  PIN Tile_X0Y1_EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 151.420 196.320 151.820 ;
    END
  END Tile_X0Y1_EE4BEG[14]
  PIN Tile_X0Y1_EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 153.100 196.320 153.500 ;
    END
  END Tile_X0Y1_EE4BEG[15]
  PIN Tile_X0Y1_EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 129.580 196.320 129.980 ;
    END
  END Tile_X0Y1_EE4BEG[1]
  PIN Tile_X0Y1_EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 131.260 196.320 131.660 ;
    END
  END Tile_X0Y1_EE4BEG[2]
  PIN Tile_X0Y1_EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 132.940 196.320 133.340 ;
    END
  END Tile_X0Y1_EE4BEG[3]
  PIN Tile_X0Y1_EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 134.620 196.320 135.020 ;
    END
  END Tile_X0Y1_EE4BEG[4]
  PIN Tile_X0Y1_EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 136.300 196.320 136.700 ;
    END
  END Tile_X0Y1_EE4BEG[5]
  PIN Tile_X0Y1_EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 137.980 196.320 138.380 ;
    END
  END Tile_X0Y1_EE4BEG[6]
  PIN Tile_X0Y1_EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 139.660 196.320 140.060 ;
    END
  END Tile_X0Y1_EE4BEG[7]
  PIN Tile_X0Y1_EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 141.340 196.320 141.740 ;
    END
  END Tile_X0Y1_EE4BEG[8]
  PIN Tile_X0Y1_EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 143.020 196.320 143.420 ;
    END
  END Tile_X0Y1_EE4BEG[9]
  PIN Tile_X0Y1_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 127.900 0.450 128.300 ;
    END
  END Tile_X0Y1_EE4END[0]
  PIN Tile_X0Y1_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 144.700 0.450 145.100 ;
    END
  END Tile_X0Y1_EE4END[10]
  PIN Tile_X0Y1_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 146.380 0.450 146.780 ;
    END
  END Tile_X0Y1_EE4END[11]
  PIN Tile_X0Y1_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 148.060 0.450 148.460 ;
    END
  END Tile_X0Y1_EE4END[12]
  PIN Tile_X0Y1_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 149.740 0.450 150.140 ;
    END
  END Tile_X0Y1_EE4END[13]
  PIN Tile_X0Y1_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 151.420 0.450 151.820 ;
    END
  END Tile_X0Y1_EE4END[14]
  PIN Tile_X0Y1_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 153.100 0.450 153.500 ;
    END
  END Tile_X0Y1_EE4END[15]
  PIN Tile_X0Y1_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 129.580 0.450 129.980 ;
    END
  END Tile_X0Y1_EE4END[1]
  PIN Tile_X0Y1_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 131.260 0.450 131.660 ;
    END
  END Tile_X0Y1_EE4END[2]
  PIN Tile_X0Y1_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 132.940 0.450 133.340 ;
    END
  END Tile_X0Y1_EE4END[3]
  PIN Tile_X0Y1_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 134.620 0.450 135.020 ;
    END
  END Tile_X0Y1_EE4END[4]
  PIN Tile_X0Y1_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 136.300 0.450 136.700 ;
    END
  END Tile_X0Y1_EE4END[5]
  PIN Tile_X0Y1_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 137.980 0.450 138.380 ;
    END
  END Tile_X0Y1_EE4END[6]
  PIN Tile_X0Y1_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 139.660 0.450 140.060 ;
    END
  END Tile_X0Y1_EE4END[7]
  PIN Tile_X0Y1_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 141.340 0.450 141.740 ;
    END
  END Tile_X0Y1_EE4END[8]
  PIN Tile_X0Y1_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 143.020 0.450 143.420 ;
    END
  END Tile_X0Y1_EE4END[9]
  PIN Tile_X0Y1_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 174.940 0.450 175.340 ;
    END
  END Tile_X0Y1_FrameData[0]
  PIN Tile_X0Y1_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 191.740 0.450 192.140 ;
    END
  END Tile_X0Y1_FrameData[10]
  PIN Tile_X0Y1_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 193.420 0.450 193.820 ;
    END
  END Tile_X0Y1_FrameData[11]
  PIN Tile_X0Y1_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 195.100 0.450 195.500 ;
    END
  END Tile_X0Y1_FrameData[12]
  PIN Tile_X0Y1_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 196.780 0.450 197.180 ;
    END
  END Tile_X0Y1_FrameData[13]
  PIN Tile_X0Y1_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 198.460 0.450 198.860 ;
    END
  END Tile_X0Y1_FrameData[14]
  PIN Tile_X0Y1_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 200.140 0.450 200.540 ;
    END
  END Tile_X0Y1_FrameData[15]
  PIN Tile_X0Y1_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 201.820 0.450 202.220 ;
    END
  END Tile_X0Y1_FrameData[16]
  PIN Tile_X0Y1_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 203.500 0.450 203.900 ;
    END
  END Tile_X0Y1_FrameData[17]
  PIN Tile_X0Y1_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 205.180 0.450 205.580 ;
    END
  END Tile_X0Y1_FrameData[18]
  PIN Tile_X0Y1_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 206.860 0.450 207.260 ;
    END
  END Tile_X0Y1_FrameData[19]
  PIN Tile_X0Y1_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 176.620 0.450 177.020 ;
    END
  END Tile_X0Y1_FrameData[1]
  PIN Tile_X0Y1_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 208.540 0.450 208.940 ;
    END
  END Tile_X0Y1_FrameData[20]
  PIN Tile_X0Y1_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 210.220 0.450 210.620 ;
    END
  END Tile_X0Y1_FrameData[21]
  PIN Tile_X0Y1_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 211.900 0.450 212.300 ;
    END
  END Tile_X0Y1_FrameData[22]
  PIN Tile_X0Y1_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 213.580 0.450 213.980 ;
    END
  END Tile_X0Y1_FrameData[23]
  PIN Tile_X0Y1_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 215.260 0.450 215.660 ;
    END
  END Tile_X0Y1_FrameData[24]
  PIN Tile_X0Y1_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 216.940 0.450 217.340 ;
    END
  END Tile_X0Y1_FrameData[25]
  PIN Tile_X0Y1_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 218.620 0.450 219.020 ;
    END
  END Tile_X0Y1_FrameData[26]
  PIN Tile_X0Y1_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 220.300 0.450 220.700 ;
    END
  END Tile_X0Y1_FrameData[27]
  PIN Tile_X0Y1_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 221.980 0.450 222.380 ;
    END
  END Tile_X0Y1_FrameData[28]
  PIN Tile_X0Y1_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 223.660 0.450 224.060 ;
    END
  END Tile_X0Y1_FrameData[29]
  PIN Tile_X0Y1_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 178.300 0.450 178.700 ;
    END
  END Tile_X0Y1_FrameData[2]
  PIN Tile_X0Y1_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 225.340 0.450 225.740 ;
    END
  END Tile_X0Y1_FrameData[30]
  PIN Tile_X0Y1_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 227.020 0.450 227.420 ;
    END
  END Tile_X0Y1_FrameData[31]
  PIN Tile_X0Y1_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 179.980 0.450 180.380 ;
    END
  END Tile_X0Y1_FrameData[3]
  PIN Tile_X0Y1_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 181.660 0.450 182.060 ;
    END
  END Tile_X0Y1_FrameData[4]
  PIN Tile_X0Y1_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 183.340 0.450 183.740 ;
    END
  END Tile_X0Y1_FrameData[5]
  PIN Tile_X0Y1_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 185.020 0.450 185.420 ;
    END
  END Tile_X0Y1_FrameData[6]
  PIN Tile_X0Y1_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 186.700 0.450 187.100 ;
    END
  END Tile_X0Y1_FrameData[7]
  PIN Tile_X0Y1_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 188.380 0.450 188.780 ;
    END
  END Tile_X0Y1_FrameData[8]
  PIN Tile_X0Y1_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 190.060 0.450 190.460 ;
    END
  END Tile_X0Y1_FrameData[9]
  PIN Tile_X0Y1_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 174.940 196.320 175.340 ;
    END
  END Tile_X0Y1_FrameData_O[0]
  PIN Tile_X0Y1_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 191.740 196.320 192.140 ;
    END
  END Tile_X0Y1_FrameData_O[10]
  PIN Tile_X0Y1_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 193.420 196.320 193.820 ;
    END
  END Tile_X0Y1_FrameData_O[11]
  PIN Tile_X0Y1_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 195.100 196.320 195.500 ;
    END
  END Tile_X0Y1_FrameData_O[12]
  PIN Tile_X0Y1_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 196.780 196.320 197.180 ;
    END
  END Tile_X0Y1_FrameData_O[13]
  PIN Tile_X0Y1_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 198.460 196.320 198.860 ;
    END
  END Tile_X0Y1_FrameData_O[14]
  PIN Tile_X0Y1_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 200.140 196.320 200.540 ;
    END
  END Tile_X0Y1_FrameData_O[15]
  PIN Tile_X0Y1_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 201.820 196.320 202.220 ;
    END
  END Tile_X0Y1_FrameData_O[16]
  PIN Tile_X0Y1_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 203.500 196.320 203.900 ;
    END
  END Tile_X0Y1_FrameData_O[17]
  PIN Tile_X0Y1_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 205.180 196.320 205.580 ;
    END
  END Tile_X0Y1_FrameData_O[18]
  PIN Tile_X0Y1_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 206.860 196.320 207.260 ;
    END
  END Tile_X0Y1_FrameData_O[19]
  PIN Tile_X0Y1_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 176.620 196.320 177.020 ;
    END
  END Tile_X0Y1_FrameData_O[1]
  PIN Tile_X0Y1_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 208.540 196.320 208.940 ;
    END
  END Tile_X0Y1_FrameData_O[20]
  PIN Tile_X0Y1_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 210.220 196.320 210.620 ;
    END
  END Tile_X0Y1_FrameData_O[21]
  PIN Tile_X0Y1_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 211.900 196.320 212.300 ;
    END
  END Tile_X0Y1_FrameData_O[22]
  PIN Tile_X0Y1_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 213.580 196.320 213.980 ;
    END
  END Tile_X0Y1_FrameData_O[23]
  PIN Tile_X0Y1_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 215.260 196.320 215.660 ;
    END
  END Tile_X0Y1_FrameData_O[24]
  PIN Tile_X0Y1_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 216.940 196.320 217.340 ;
    END
  END Tile_X0Y1_FrameData_O[25]
  PIN Tile_X0Y1_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 218.620 196.320 219.020 ;
    END
  END Tile_X0Y1_FrameData_O[26]
  PIN Tile_X0Y1_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 220.300 196.320 220.700 ;
    END
  END Tile_X0Y1_FrameData_O[27]
  PIN Tile_X0Y1_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 221.980 196.320 222.380 ;
    END
  END Tile_X0Y1_FrameData_O[28]
  PIN Tile_X0Y1_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 223.660 196.320 224.060 ;
    END
  END Tile_X0Y1_FrameData_O[29]
  PIN Tile_X0Y1_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 178.300 196.320 178.700 ;
    END
  END Tile_X0Y1_FrameData_O[2]
  PIN Tile_X0Y1_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 225.340 196.320 225.740 ;
    END
  END Tile_X0Y1_FrameData_O[30]
  PIN Tile_X0Y1_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 227.020 196.320 227.420 ;
    END
  END Tile_X0Y1_FrameData_O[31]
  PIN Tile_X0Y1_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 179.980 196.320 180.380 ;
    END
  END Tile_X0Y1_FrameData_O[3]
  PIN Tile_X0Y1_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 181.660 196.320 182.060 ;
    END
  END Tile_X0Y1_FrameData_O[4]
  PIN Tile_X0Y1_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 183.340 196.320 183.740 ;
    END
  END Tile_X0Y1_FrameData_O[5]
  PIN Tile_X0Y1_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 185.020 196.320 185.420 ;
    END
  END Tile_X0Y1_FrameData_O[6]
  PIN Tile_X0Y1_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 186.700 196.320 187.100 ;
    END
  END Tile_X0Y1_FrameData_O[7]
  PIN Tile_X0Y1_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 188.380 196.320 188.780 ;
    END
  END Tile_X0Y1_FrameData_O[8]
  PIN Tile_X0Y1_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 190.060 196.320 190.460 ;
    END
  END Tile_X0Y1_FrameData_O[9]
  PIN Tile_X0Y1_FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal3 ;
        RECT 138.520 0.000 138.920 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[0]
  PIN Tile_X0Y1_FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.542100 ;
    PORT
      LAYER Metal3 ;
        RECT 148.120 0.000 148.520 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[10]
  PIN Tile_X0Y1_FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 149.080 0.000 149.480 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[11]
  PIN Tile_X0Y1_FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 150.040 0.000 150.440 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[12]
  PIN Tile_X0Y1_FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 151.000 0.000 151.400 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[13]
  PIN Tile_X0Y1_FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 151.960 0.000 152.360 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[14]
  PIN Tile_X0Y1_FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 152.920 0.000 153.320 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[15]
  PIN Tile_X0Y1_FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 153.880 0.000 154.280 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[16]
  PIN Tile_X0Y1_FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 154.840 0.000 155.240 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[17]
  PIN Tile_X0Y1_FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 155.800 0.000 156.200 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[18]
  PIN Tile_X0Y1_FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 156.760 0.000 157.160 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[19]
  PIN Tile_X0Y1_FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 139.480 0.000 139.880 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[1]
  PIN Tile_X0Y1_FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 140.440 0.000 140.840 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[2]
  PIN Tile_X0Y1_FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.542100 ;
    PORT
      LAYER Metal3 ;
        RECT 141.400 0.000 141.800 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[3]
  PIN Tile_X0Y1_FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.542100 ;
    PORT
      LAYER Metal3 ;
        RECT 142.360 0.000 142.760 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[4]
  PIN Tile_X0Y1_FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal3 ;
        RECT 143.320 0.000 143.720 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[5]
  PIN Tile_X0Y1_FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 144.280 0.000 144.680 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[6]
  PIN Tile_X0Y1_FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.542100 ;
    PORT
      LAYER Metal3 ;
        RECT 145.240 0.000 145.640 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[7]
  PIN Tile_X0Y1_FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 146.200 0.000 146.600 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[8]
  PIN Tile_X0Y1_FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.542100 ;
    PORT
      LAYER Metal3 ;
        RECT 147.160 0.000 147.560 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[9]
  PIN Tile_X0Y1_N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 37.720 0.000 38.120 0.400 ;
    END
  END Tile_X0Y1_N1END[0]
  PIN Tile_X0Y1_N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 38.680 0.000 39.080 0.400 ;
    END
  END Tile_X0Y1_N1END[1]
  PIN Tile_X0Y1_N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 39.640 0.000 40.040 0.400 ;
    END
  END Tile_X0Y1_N1END[2]
  PIN Tile_X0Y1_N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 40.600 0.000 41.000 0.400 ;
    END
  END Tile_X0Y1_N1END[3]
  PIN Tile_X0Y1_N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 49.240 0.000 49.640 0.400 ;
    END
  END Tile_X0Y1_N2END[0]
  PIN Tile_X0Y1_N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 50.200 0.000 50.600 0.400 ;
    END
  END Tile_X0Y1_N2END[1]
  PIN Tile_X0Y1_N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 51.160 0.000 51.560 0.400 ;
    END
  END Tile_X0Y1_N2END[2]
  PIN Tile_X0Y1_N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 52.120 0.000 52.520 0.400 ;
    END
  END Tile_X0Y1_N2END[3]
  PIN Tile_X0Y1_N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 53.080 0.000 53.480 0.400 ;
    END
  END Tile_X0Y1_N2END[4]
  PIN Tile_X0Y1_N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 54.040 0.000 54.440 0.400 ;
    END
  END Tile_X0Y1_N2END[5]
  PIN Tile_X0Y1_N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 55.000 0.000 55.400 0.400 ;
    END
  END Tile_X0Y1_N2END[6]
  PIN Tile_X0Y1_N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 55.960 0.000 56.360 0.400 ;
    END
  END Tile_X0Y1_N2END[7]
  PIN Tile_X0Y1_N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 41.560 0.000 41.960 0.400 ;
    END
  END Tile_X0Y1_N2MID[0]
  PIN Tile_X0Y1_N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 42.520 0.000 42.920 0.400 ;
    END
  END Tile_X0Y1_N2MID[1]
  PIN Tile_X0Y1_N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal3 ;
        RECT 43.480 0.000 43.880 0.400 ;
    END
  END Tile_X0Y1_N2MID[2]
  PIN Tile_X0Y1_N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 44.440 0.000 44.840 0.400 ;
    END
  END Tile_X0Y1_N2MID[3]
  PIN Tile_X0Y1_N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 45.400 0.000 45.800 0.400 ;
    END
  END Tile_X0Y1_N2MID[4]
  PIN Tile_X0Y1_N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 46.360 0.000 46.760 0.400 ;
    END
  END Tile_X0Y1_N2MID[5]
  PIN Tile_X0Y1_N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 47.320 0.000 47.720 0.400 ;
    END
  END Tile_X0Y1_N2MID[6]
  PIN Tile_X0Y1_N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 48.280 0.000 48.680 0.400 ;
    END
  END Tile_X0Y1_N2MID[7]
  PIN Tile_X0Y1_N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 56.920 0.000 57.320 0.400 ;
    END
  END Tile_X0Y1_N4END[0]
  PIN Tile_X0Y1_N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 66.520 0.000 66.920 0.400 ;
    END
  END Tile_X0Y1_N4END[10]
  PIN Tile_X0Y1_N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 67.480 0.000 67.880 0.400 ;
    END
  END Tile_X0Y1_N4END[11]
  PIN Tile_X0Y1_N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 68.440 0.000 68.840 0.400 ;
    END
  END Tile_X0Y1_N4END[12]
  PIN Tile_X0Y1_N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 69.400 0.000 69.800 0.400 ;
    END
  END Tile_X0Y1_N4END[13]
  PIN Tile_X0Y1_N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 70.360 0.000 70.760 0.400 ;
    END
  END Tile_X0Y1_N4END[14]
  PIN Tile_X0Y1_N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 71.320 0.000 71.720 0.400 ;
    END
  END Tile_X0Y1_N4END[15]
  PIN Tile_X0Y1_N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 57.880 0.000 58.280 0.400 ;
    END
  END Tile_X0Y1_N4END[1]
  PIN Tile_X0Y1_N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 58.840 0.000 59.240 0.400 ;
    END
  END Tile_X0Y1_N4END[2]
  PIN Tile_X0Y1_N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 59.800 0.000 60.200 0.400 ;
    END
  END Tile_X0Y1_N4END[3]
  PIN Tile_X0Y1_N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 60.760 0.000 61.160 0.400 ;
    END
  END Tile_X0Y1_N4END[4]
  PIN Tile_X0Y1_N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 61.720 0.000 62.120 0.400 ;
    END
  END Tile_X0Y1_N4END[5]
  PIN Tile_X0Y1_N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.450800 ;
    PORT
      LAYER Metal3 ;
        RECT 62.680 0.000 63.080 0.400 ;
    END
  END Tile_X0Y1_N4END[6]
  PIN Tile_X0Y1_N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 63.640 0.000 64.040 0.400 ;
    END
  END Tile_X0Y1_N4END[7]
  PIN Tile_X0Y1_N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 64.600 0.000 65.000 0.400 ;
    END
  END Tile_X0Y1_N4END[8]
  PIN Tile_X0Y1_N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 65.560 0.000 65.960 0.400 ;
    END
  END Tile_X0Y1_N4END[9]
  PIN Tile_X0Y1_NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 72.280 0.000 72.680 0.400 ;
    END
  END Tile_X0Y1_NN4END[0]
  PIN Tile_X0Y1_NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 81.880 0.000 82.280 0.400 ;
    END
  END Tile_X0Y1_NN4END[10]
  PIN Tile_X0Y1_NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 82.840 0.000 83.240 0.400 ;
    END
  END Tile_X0Y1_NN4END[11]
  PIN Tile_X0Y1_NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 83.800 0.000 84.200 0.400 ;
    END
  END Tile_X0Y1_NN4END[12]
  PIN Tile_X0Y1_NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 84.760 0.000 85.160 0.400 ;
    END
  END Tile_X0Y1_NN4END[13]
  PIN Tile_X0Y1_NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 85.720 0.000 86.120 0.400 ;
    END
  END Tile_X0Y1_NN4END[14]
  PIN Tile_X0Y1_NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 86.680 0.000 87.080 0.400 ;
    END
  END Tile_X0Y1_NN4END[15]
  PIN Tile_X0Y1_NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 73.240 0.000 73.640 0.400 ;
    END
  END Tile_X0Y1_NN4END[1]
  PIN Tile_X0Y1_NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 74.200 0.000 74.600 0.400 ;
    END
  END Tile_X0Y1_NN4END[2]
  PIN Tile_X0Y1_NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 75.160 0.000 75.560 0.400 ;
    END
  END Tile_X0Y1_NN4END[3]
  PIN Tile_X0Y1_NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 76.120 0.000 76.520 0.400 ;
    END
  END Tile_X0Y1_NN4END[4]
  PIN Tile_X0Y1_NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 77.080 0.000 77.480 0.400 ;
    END
  END Tile_X0Y1_NN4END[5]
  PIN Tile_X0Y1_NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 78.040 0.000 78.440 0.400 ;
    END
  END Tile_X0Y1_NN4END[6]
  PIN Tile_X0Y1_NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 79.000 0.000 79.400 0.400 ;
    END
  END Tile_X0Y1_NN4END[7]
  PIN Tile_X0Y1_NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 79.960 0.000 80.360 0.400 ;
    END
  END Tile_X0Y1_NN4END[8]
  PIN Tile_X0Y1_NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 80.920 0.000 81.320 0.400 ;
    END
  END Tile_X0Y1_NN4END[9]
  PIN Tile_X0Y1_S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.827200 ;
    PORT
      LAYER Metal3 ;
        RECT 87.640 0.000 88.040 0.400 ;
    END
  END Tile_X0Y1_S1BEG[0]
  PIN Tile_X0Y1_S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.827200 ;
    PORT
      LAYER Metal3 ;
        RECT 88.600 0.000 89.000 0.400 ;
    END
  END Tile_X0Y1_S1BEG[1]
  PIN Tile_X0Y1_S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 89.560 0.000 89.960 0.400 ;
    END
  END Tile_X0Y1_S1BEG[2]
  PIN Tile_X0Y1_S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 90.520 0.000 90.920 0.400 ;
    END
  END Tile_X0Y1_S1BEG[3]
  PIN Tile_X0Y1_S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 91.480 0.000 91.880 0.400 ;
    END
  END Tile_X0Y1_S2BEG[0]
  PIN Tile_X0Y1_S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 92.440 0.000 92.840 0.400 ;
    END
  END Tile_X0Y1_S2BEG[1]
  PIN Tile_X0Y1_S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 93.400 0.000 93.800 0.400 ;
    END
  END Tile_X0Y1_S2BEG[2]
  PIN Tile_X0Y1_S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 94.360 0.000 94.760 0.400 ;
    END
  END Tile_X0Y1_S2BEG[3]
  PIN Tile_X0Y1_S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 95.320 0.000 95.720 0.400 ;
    END
  END Tile_X0Y1_S2BEG[4]
  PIN Tile_X0Y1_S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 96.280 0.000 96.680 0.400 ;
    END
  END Tile_X0Y1_S2BEG[5]
  PIN Tile_X0Y1_S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 97.240 0.000 97.640 0.400 ;
    END
  END Tile_X0Y1_S2BEG[6]
  PIN Tile_X0Y1_S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 98.200 0.000 98.600 0.400 ;
    END
  END Tile_X0Y1_S2BEG[7]
  PIN Tile_X0Y1_S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 99.160 0.000 99.560 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[0]
  PIN Tile_X0Y1_S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 100.120 0.000 100.520 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[1]
  PIN Tile_X0Y1_S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 101.080 0.000 101.480 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[2]
  PIN Tile_X0Y1_S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 102.040 0.000 102.440 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[3]
  PIN Tile_X0Y1_S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 103.000 0.000 103.400 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[4]
  PIN Tile_X0Y1_S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 103.960 0.000 104.360 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[5]
  PIN Tile_X0Y1_S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 104.920 0.000 105.320 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[6]
  PIN Tile_X0Y1_S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 105.880 0.000 106.280 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[7]
  PIN Tile_X0Y1_S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 106.840 0.000 107.240 0.400 ;
    END
  END Tile_X0Y1_S4BEG[0]
  PIN Tile_X0Y1_S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 116.440 0.000 116.840 0.400 ;
    END
  END Tile_X0Y1_S4BEG[10]
  PIN Tile_X0Y1_S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 117.400 0.000 117.800 0.400 ;
    END
  END Tile_X0Y1_S4BEG[11]
  PIN Tile_X0Y1_S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 118.360 0.000 118.760 0.400 ;
    END
  END Tile_X0Y1_S4BEG[12]
  PIN Tile_X0Y1_S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 119.320 0.000 119.720 0.400 ;
    END
  END Tile_X0Y1_S4BEG[13]
  PIN Tile_X0Y1_S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 120.280 0.000 120.680 0.400 ;
    END
  END Tile_X0Y1_S4BEG[14]
  PIN Tile_X0Y1_S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 121.240 0.000 121.640 0.400 ;
    END
  END Tile_X0Y1_S4BEG[15]
  PIN Tile_X0Y1_S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 107.800 0.000 108.200 0.400 ;
    END
  END Tile_X0Y1_S4BEG[1]
  PIN Tile_X0Y1_S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 108.760 0.000 109.160 0.400 ;
    END
  END Tile_X0Y1_S4BEG[2]
  PIN Tile_X0Y1_S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 109.720 0.000 110.120 0.400 ;
    END
  END Tile_X0Y1_S4BEG[3]
  PIN Tile_X0Y1_S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 110.680 0.000 111.080 0.400 ;
    END
  END Tile_X0Y1_S4BEG[4]
  PIN Tile_X0Y1_S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 111.640 0.000 112.040 0.400 ;
    END
  END Tile_X0Y1_S4BEG[5]
  PIN Tile_X0Y1_S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 112.600 0.000 113.000 0.400 ;
    END
  END Tile_X0Y1_S4BEG[6]
  PIN Tile_X0Y1_S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 113.560 0.000 113.960 0.400 ;
    END
  END Tile_X0Y1_S4BEG[7]
  PIN Tile_X0Y1_S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 114.520 0.000 114.920 0.400 ;
    END
  END Tile_X0Y1_S4BEG[8]
  PIN Tile_X0Y1_S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 115.480 0.000 115.880 0.400 ;
    END
  END Tile_X0Y1_S4BEG[9]
  PIN Tile_X0Y1_SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 122.200 0.000 122.600 0.400 ;
    END
  END Tile_X0Y1_SS4BEG[0]
  PIN Tile_X0Y1_SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.827200 ;
    PORT
      LAYER Metal3 ;
        RECT 131.800 0.000 132.200 0.400 ;
    END
  END Tile_X0Y1_SS4BEG[10]
  PIN Tile_X0Y1_SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.827200 ;
    PORT
      LAYER Metal3 ;
        RECT 132.760 0.000 133.160 0.400 ;
    END
  END Tile_X0Y1_SS4BEG[11]
  PIN Tile_X0Y1_SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 133.720 0.000 134.120 0.400 ;
    END
  END Tile_X0Y1_SS4BEG[12]
  PIN Tile_X0Y1_SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.827200 ;
    PORT
      LAYER Metal3 ;
        RECT 134.680 0.000 135.080 0.400 ;
    END
  END Tile_X0Y1_SS4BEG[13]
  PIN Tile_X0Y1_SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 135.640 0.000 136.040 0.400 ;
    END
  END Tile_X0Y1_SS4BEG[14]
  PIN Tile_X0Y1_SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 136.600 0.000 137.000 0.400 ;
    END
  END Tile_X0Y1_SS4BEG[15]
  PIN Tile_X0Y1_SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 123.160 0.000 123.560 0.400 ;
    END
  END Tile_X0Y1_SS4BEG[1]
  PIN Tile_X0Y1_SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 124.120 0.000 124.520 0.400 ;
    END
  END Tile_X0Y1_SS4BEG[2]
  PIN Tile_X0Y1_SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 125.080 0.000 125.480 0.400 ;
    END
  END Tile_X0Y1_SS4BEG[3]
  PIN Tile_X0Y1_SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 126.040 0.000 126.440 0.400 ;
    END
  END Tile_X0Y1_SS4BEG[4]
  PIN Tile_X0Y1_SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 127.000 0.000 127.400 0.400 ;
    END
  END Tile_X0Y1_SS4BEG[5]
  PIN Tile_X0Y1_SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 127.960 0.000 128.360 0.400 ;
    END
  END Tile_X0Y1_SS4BEG[6]
  PIN Tile_X0Y1_SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 128.920 0.000 129.320 0.400 ;
    END
  END Tile_X0Y1_SS4BEG[7]
  PIN Tile_X0Y1_SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 129.880 0.000 130.280 0.400 ;
    END
  END Tile_X0Y1_SS4BEG[8]
  PIN Tile_X0Y1_SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.827200 ;
    PORT
      LAYER Metal3 ;
        RECT 130.840 0.000 131.240 0.400 ;
    END
  END Tile_X0Y1_SS4BEG[9]
  PIN Tile_X0Y1_UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 12.847899 ;
    PORT
      LAYER Metal3 ;
        RECT 137.560 0.000 137.960 0.400 ;
    END
  END Tile_X0Y1_UserCLK
  PIN Tile_X0Y1_W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 13.660 0.450 14.060 ;
    END
  END Tile_X0Y1_W1BEG[0]
  PIN Tile_X0Y1_W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 15.340 0.450 15.740 ;
    END
  END Tile_X0Y1_W1BEG[1]
  PIN Tile_X0Y1_W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 17.020 0.450 17.420 ;
    END
  END Tile_X0Y1_W1BEG[2]
  PIN Tile_X0Y1_W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 18.700 0.450 19.100 ;
    END
  END Tile_X0Y1_W1BEG[3]
  PIN Tile_X0Y1_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 13.660 196.320 14.060 ;
    END
  END Tile_X0Y1_W1END[0]
  PIN Tile_X0Y1_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 15.340 196.320 15.740 ;
    END
  END Tile_X0Y1_W1END[1]
  PIN Tile_X0Y1_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 17.020 196.320 17.420 ;
    END
  END Tile_X0Y1_W1END[2]
  PIN Tile_X0Y1_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 18.700 196.320 19.100 ;
    END
  END Tile_X0Y1_W1END[3]
  PIN Tile_X0Y1_W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 20.380 0.450 20.780 ;
    END
  END Tile_X0Y1_W2BEG[0]
  PIN Tile_X0Y1_W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 22.060 0.450 22.460 ;
    END
  END Tile_X0Y1_W2BEG[1]
  PIN Tile_X0Y1_W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 23.740 0.450 24.140 ;
    END
  END Tile_X0Y1_W2BEG[2]
  PIN Tile_X0Y1_W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 25.420 0.450 25.820 ;
    END
  END Tile_X0Y1_W2BEG[3]
  PIN Tile_X0Y1_W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 27.100 0.450 27.500 ;
    END
  END Tile_X0Y1_W2BEG[4]
  PIN Tile_X0Y1_W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 28.780 0.450 29.180 ;
    END
  END Tile_X0Y1_W2BEG[5]
  PIN Tile_X0Y1_W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 30.460 0.450 30.860 ;
    END
  END Tile_X0Y1_W2BEG[6]
  PIN Tile_X0Y1_W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 32.140 0.450 32.540 ;
    END
  END Tile_X0Y1_W2BEG[7]
  PIN Tile_X0Y1_W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 33.820 0.450 34.220 ;
    END
  END Tile_X0Y1_W2BEGb[0]
  PIN Tile_X0Y1_W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 35.500 0.450 35.900 ;
    END
  END Tile_X0Y1_W2BEGb[1]
  PIN Tile_X0Y1_W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 37.180 0.450 37.580 ;
    END
  END Tile_X0Y1_W2BEGb[2]
  PIN Tile_X0Y1_W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 38.860 0.450 39.260 ;
    END
  END Tile_X0Y1_W2BEGb[3]
  PIN Tile_X0Y1_W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 40.540 0.450 40.940 ;
    END
  END Tile_X0Y1_W2BEGb[4]
  PIN Tile_X0Y1_W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 42.220 0.450 42.620 ;
    END
  END Tile_X0Y1_W2BEGb[5]
  PIN Tile_X0Y1_W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 43.900 0.450 44.300 ;
    END
  END Tile_X0Y1_W2BEGb[6]
  PIN Tile_X0Y1_W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 45.580 0.450 45.980 ;
    END
  END Tile_X0Y1_W2BEGb[7]
  PIN Tile_X0Y1_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 33.820 196.320 34.220 ;
    END
  END Tile_X0Y1_W2END[0]
  PIN Tile_X0Y1_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 35.500 196.320 35.900 ;
    END
  END Tile_X0Y1_W2END[1]
  PIN Tile_X0Y1_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 37.180 196.320 37.580 ;
    END
  END Tile_X0Y1_W2END[2]
  PIN Tile_X0Y1_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 38.860 196.320 39.260 ;
    END
  END Tile_X0Y1_W2END[3]
  PIN Tile_X0Y1_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 40.540 196.320 40.940 ;
    END
  END Tile_X0Y1_W2END[4]
  PIN Tile_X0Y1_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 42.220 196.320 42.620 ;
    END
  END Tile_X0Y1_W2END[5]
  PIN Tile_X0Y1_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 43.900 196.320 44.300 ;
    END
  END Tile_X0Y1_W2END[6]
  PIN Tile_X0Y1_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 45.580 196.320 45.980 ;
    END
  END Tile_X0Y1_W2END[7]
  PIN Tile_X0Y1_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 20.380 196.320 20.780 ;
    END
  END Tile_X0Y1_W2MID[0]
  PIN Tile_X0Y1_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 22.060 196.320 22.460 ;
    END
  END Tile_X0Y1_W2MID[1]
  PIN Tile_X0Y1_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 23.740 196.320 24.140 ;
    END
  END Tile_X0Y1_W2MID[2]
  PIN Tile_X0Y1_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 25.420 196.320 25.820 ;
    END
  END Tile_X0Y1_W2MID[3]
  PIN Tile_X0Y1_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 27.100 196.320 27.500 ;
    END
  END Tile_X0Y1_W2MID[4]
  PIN Tile_X0Y1_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 28.780 196.320 29.180 ;
    END
  END Tile_X0Y1_W2MID[5]
  PIN Tile_X0Y1_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 30.460 196.320 30.860 ;
    END
  END Tile_X0Y1_W2MID[6]
  PIN Tile_X0Y1_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 32.140 196.320 32.540 ;
    END
  END Tile_X0Y1_W2MID[7]
  PIN Tile_X0Y1_W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 74.140 0.450 74.540 ;
    END
  END Tile_X0Y1_W6BEG[0]
  PIN Tile_X0Y1_W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 90.940 0.450 91.340 ;
    END
  END Tile_X0Y1_W6BEG[10]
  PIN Tile_X0Y1_W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 92.620 0.450 93.020 ;
    END
  END Tile_X0Y1_W6BEG[11]
  PIN Tile_X0Y1_W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 75.820 0.450 76.220 ;
    END
  END Tile_X0Y1_W6BEG[1]
  PIN Tile_X0Y1_W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 77.500 0.450 77.900 ;
    END
  END Tile_X0Y1_W6BEG[2]
  PIN Tile_X0Y1_W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 79.180 0.450 79.580 ;
    END
  END Tile_X0Y1_W6BEG[3]
  PIN Tile_X0Y1_W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 80.860 0.450 81.260 ;
    END
  END Tile_X0Y1_W6BEG[4]
  PIN Tile_X0Y1_W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 82.540 0.450 82.940 ;
    END
  END Tile_X0Y1_W6BEG[5]
  PIN Tile_X0Y1_W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 84.220 0.450 84.620 ;
    END
  END Tile_X0Y1_W6BEG[6]
  PIN Tile_X0Y1_W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 85.900 0.450 86.300 ;
    END
  END Tile_X0Y1_W6BEG[7]
  PIN Tile_X0Y1_W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 87.580 0.450 87.980 ;
    END
  END Tile_X0Y1_W6BEG[8]
  PIN Tile_X0Y1_W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 89.260 0.450 89.660 ;
    END
  END Tile_X0Y1_W6BEG[9]
  PIN Tile_X0Y1_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 74.140 196.320 74.540 ;
    END
  END Tile_X0Y1_W6END[0]
  PIN Tile_X0Y1_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 90.940 196.320 91.340 ;
    END
  END Tile_X0Y1_W6END[10]
  PIN Tile_X0Y1_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 92.620 196.320 93.020 ;
    END
  END Tile_X0Y1_W6END[11]
  PIN Tile_X0Y1_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 75.820 196.320 76.220 ;
    END
  END Tile_X0Y1_W6END[1]
  PIN Tile_X0Y1_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 77.500 196.320 77.900 ;
    END
  END Tile_X0Y1_W6END[2]
  PIN Tile_X0Y1_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 79.180 196.320 79.580 ;
    END
  END Tile_X0Y1_W6END[3]
  PIN Tile_X0Y1_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 80.860 196.320 81.260 ;
    END
  END Tile_X0Y1_W6END[4]
  PIN Tile_X0Y1_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 82.540 196.320 82.940 ;
    END
  END Tile_X0Y1_W6END[5]
  PIN Tile_X0Y1_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 84.220 196.320 84.620 ;
    END
  END Tile_X0Y1_W6END[6]
  PIN Tile_X0Y1_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 85.900 196.320 86.300 ;
    END
  END Tile_X0Y1_W6END[7]
  PIN Tile_X0Y1_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 87.580 196.320 87.980 ;
    END
  END Tile_X0Y1_W6END[8]
  PIN Tile_X0Y1_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 89.260 196.320 89.660 ;
    END
  END Tile_X0Y1_W6END[9]
  PIN Tile_X0Y1_WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 47.260 0.450 47.660 ;
    END
  END Tile_X0Y1_WW4BEG[0]
  PIN Tile_X0Y1_WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 64.060 0.450 64.460 ;
    END
  END Tile_X0Y1_WW4BEG[10]
  PIN Tile_X0Y1_WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 65.740 0.450 66.140 ;
    END
  END Tile_X0Y1_WW4BEG[11]
  PIN Tile_X0Y1_WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 67.420 0.450 67.820 ;
    END
  END Tile_X0Y1_WW4BEG[12]
  PIN Tile_X0Y1_WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 69.100 0.450 69.500 ;
    END
  END Tile_X0Y1_WW4BEG[13]
  PIN Tile_X0Y1_WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 70.780 0.450 71.180 ;
    END
  END Tile_X0Y1_WW4BEG[14]
  PIN Tile_X0Y1_WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 72.460 0.450 72.860 ;
    END
  END Tile_X0Y1_WW4BEG[15]
  PIN Tile_X0Y1_WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 48.940 0.450 49.340 ;
    END
  END Tile_X0Y1_WW4BEG[1]
  PIN Tile_X0Y1_WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 50.620 0.450 51.020 ;
    END
  END Tile_X0Y1_WW4BEG[2]
  PIN Tile_X0Y1_WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 52.300 0.450 52.700 ;
    END
  END Tile_X0Y1_WW4BEG[3]
  PIN Tile_X0Y1_WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 53.980 0.450 54.380 ;
    END
  END Tile_X0Y1_WW4BEG[4]
  PIN Tile_X0Y1_WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 55.660 0.450 56.060 ;
    END
  END Tile_X0Y1_WW4BEG[5]
  PIN Tile_X0Y1_WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 57.340 0.450 57.740 ;
    END
  END Tile_X0Y1_WW4BEG[6]
  PIN Tile_X0Y1_WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 59.020 0.450 59.420 ;
    END
  END Tile_X0Y1_WW4BEG[7]
  PIN Tile_X0Y1_WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 60.700 0.450 61.100 ;
    END
  END Tile_X0Y1_WW4BEG[8]
  PIN Tile_X0Y1_WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 62.380 0.450 62.780 ;
    END
  END Tile_X0Y1_WW4BEG[9]
  PIN Tile_X0Y1_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 47.260 196.320 47.660 ;
    END
  END Tile_X0Y1_WW4END[0]
  PIN Tile_X0Y1_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 64.060 196.320 64.460 ;
    END
  END Tile_X0Y1_WW4END[10]
  PIN Tile_X0Y1_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 65.740 196.320 66.140 ;
    END
  END Tile_X0Y1_WW4END[11]
  PIN Tile_X0Y1_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 67.420 196.320 67.820 ;
    END
  END Tile_X0Y1_WW4END[12]
  PIN Tile_X0Y1_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 69.100 196.320 69.500 ;
    END
  END Tile_X0Y1_WW4END[13]
  PIN Tile_X0Y1_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 70.780 196.320 71.180 ;
    END
  END Tile_X0Y1_WW4END[14]
  PIN Tile_X0Y1_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 72.460 196.320 72.860 ;
    END
  END Tile_X0Y1_WW4END[15]
  PIN Tile_X0Y1_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 48.940 196.320 49.340 ;
    END
  END Tile_X0Y1_WW4END[1]
  PIN Tile_X0Y1_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 50.620 196.320 51.020 ;
    END
  END Tile_X0Y1_WW4END[2]
  PIN Tile_X0Y1_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 52.300 196.320 52.700 ;
    END
  END Tile_X0Y1_WW4END[3]
  PIN Tile_X0Y1_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 53.980 196.320 54.380 ;
    END
  END Tile_X0Y1_WW4END[4]
  PIN Tile_X0Y1_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 55.660 196.320 56.060 ;
    END
  END Tile_X0Y1_WW4END[5]
  PIN Tile_X0Y1_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 57.340 196.320 57.740 ;
    END
  END Tile_X0Y1_WW4END[6]
  PIN Tile_X0Y1_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 59.020 196.320 59.420 ;
    END
  END Tile_X0Y1_WW4END[7]
  PIN Tile_X0Y1_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 60.700 196.320 61.100 ;
    END
  END Tile_X0Y1_WW4END[8]
  PIN Tile_X0Y1_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 195.870 62.380 196.320 62.780 ;
    END
  END Tile_X0Y1_WW4END[9]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 24.460 0.000 26.660 483.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 100.060 0.000 102.260 483.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 175.660 0.000 177.860 483.840 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 18.260 0.000 20.460 483.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 93.860 0.000 96.060 483.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 169.460 0.000 171.660 483.840 ;
    END
  END VPWR
  OBS
      LAYER GatPoly ;
        RECT 5.760 7.410 190.560 476.430 ;
      LAYER Metal1 ;
        RECT 5.760 7.340 190.560 476.500 ;
      LAYER Metal2 ;
        RECT 0.335 469.550 196.195 483.520 ;
        RECT 0.660 468.730 195.660 469.550 ;
        RECT 0.335 467.870 196.195 468.730 ;
        RECT 0.660 467.050 195.660 467.870 ;
        RECT 0.335 466.190 196.195 467.050 ;
        RECT 0.660 465.370 195.660 466.190 ;
        RECT 0.335 464.510 196.195 465.370 ;
        RECT 0.660 463.690 195.660 464.510 ;
        RECT 0.335 462.830 196.195 463.690 ;
        RECT 0.660 462.010 195.660 462.830 ;
        RECT 0.335 461.150 196.195 462.010 ;
        RECT 0.660 460.330 195.660 461.150 ;
        RECT 0.335 459.470 196.195 460.330 ;
        RECT 0.660 458.650 195.660 459.470 ;
        RECT 0.335 457.790 196.195 458.650 ;
        RECT 0.660 456.970 195.660 457.790 ;
        RECT 0.335 456.110 196.195 456.970 ;
        RECT 0.660 455.290 195.660 456.110 ;
        RECT 0.335 454.430 196.195 455.290 ;
        RECT 0.660 453.610 195.660 454.430 ;
        RECT 0.335 452.750 196.195 453.610 ;
        RECT 0.660 451.930 195.660 452.750 ;
        RECT 0.335 451.070 196.195 451.930 ;
        RECT 0.660 450.250 195.660 451.070 ;
        RECT 0.335 449.390 196.195 450.250 ;
        RECT 0.660 448.570 195.660 449.390 ;
        RECT 0.335 447.710 196.195 448.570 ;
        RECT 0.660 446.890 195.660 447.710 ;
        RECT 0.335 446.030 196.195 446.890 ;
        RECT 0.660 445.210 195.660 446.030 ;
        RECT 0.335 444.350 196.195 445.210 ;
        RECT 0.660 443.530 195.660 444.350 ;
        RECT 0.335 442.670 196.195 443.530 ;
        RECT 0.660 441.850 195.660 442.670 ;
        RECT 0.335 440.990 196.195 441.850 ;
        RECT 0.660 440.170 195.660 440.990 ;
        RECT 0.335 439.310 196.195 440.170 ;
        RECT 0.660 438.490 195.660 439.310 ;
        RECT 0.335 437.630 196.195 438.490 ;
        RECT 0.660 436.810 195.660 437.630 ;
        RECT 0.335 435.950 196.195 436.810 ;
        RECT 0.660 435.130 195.660 435.950 ;
        RECT 0.335 434.270 196.195 435.130 ;
        RECT 0.660 433.450 195.660 434.270 ;
        RECT 0.335 432.590 196.195 433.450 ;
        RECT 0.660 431.770 195.660 432.590 ;
        RECT 0.335 430.910 196.195 431.770 ;
        RECT 0.660 430.090 195.660 430.910 ;
        RECT 0.335 429.230 196.195 430.090 ;
        RECT 0.660 428.410 195.660 429.230 ;
        RECT 0.335 427.550 196.195 428.410 ;
        RECT 0.660 426.730 195.660 427.550 ;
        RECT 0.335 425.870 196.195 426.730 ;
        RECT 0.660 425.050 195.660 425.870 ;
        RECT 0.335 424.190 196.195 425.050 ;
        RECT 0.660 423.370 195.660 424.190 ;
        RECT 0.335 422.510 196.195 423.370 ;
        RECT 0.660 421.690 195.660 422.510 ;
        RECT 0.335 420.830 196.195 421.690 ;
        RECT 0.660 420.010 195.660 420.830 ;
        RECT 0.335 419.150 196.195 420.010 ;
        RECT 0.660 418.330 195.660 419.150 ;
        RECT 0.335 417.470 196.195 418.330 ;
        RECT 0.660 416.650 195.660 417.470 ;
        RECT 0.335 415.790 196.195 416.650 ;
        RECT 0.660 414.970 195.660 415.790 ;
        RECT 0.335 414.110 196.195 414.970 ;
        RECT 0.660 413.290 195.660 414.110 ;
        RECT 0.335 412.430 196.195 413.290 ;
        RECT 0.660 411.610 195.660 412.430 ;
        RECT 0.335 410.750 196.195 411.610 ;
        RECT 0.660 409.930 195.660 410.750 ;
        RECT 0.335 409.070 196.195 409.930 ;
        RECT 0.660 408.250 195.660 409.070 ;
        RECT 0.335 407.390 196.195 408.250 ;
        RECT 0.660 406.570 195.660 407.390 ;
        RECT 0.335 405.710 196.195 406.570 ;
        RECT 0.660 404.890 195.660 405.710 ;
        RECT 0.335 404.030 196.195 404.890 ;
        RECT 0.660 403.210 195.660 404.030 ;
        RECT 0.335 402.350 196.195 403.210 ;
        RECT 0.660 401.530 195.660 402.350 ;
        RECT 0.335 400.670 196.195 401.530 ;
        RECT 0.660 399.850 195.660 400.670 ;
        RECT 0.335 398.990 196.195 399.850 ;
        RECT 0.660 398.170 195.660 398.990 ;
        RECT 0.335 397.310 196.195 398.170 ;
        RECT 0.660 396.490 195.660 397.310 ;
        RECT 0.335 395.630 196.195 396.490 ;
        RECT 0.660 394.810 195.660 395.630 ;
        RECT 0.335 393.950 196.195 394.810 ;
        RECT 0.660 393.130 195.660 393.950 ;
        RECT 0.335 392.270 196.195 393.130 ;
        RECT 0.660 391.450 195.660 392.270 ;
        RECT 0.335 390.590 196.195 391.450 ;
        RECT 0.660 389.770 195.660 390.590 ;
        RECT 0.335 388.910 196.195 389.770 ;
        RECT 0.660 388.090 195.660 388.910 ;
        RECT 0.335 387.230 196.195 388.090 ;
        RECT 0.660 386.410 195.660 387.230 ;
        RECT 0.335 385.550 196.195 386.410 ;
        RECT 0.660 384.730 195.660 385.550 ;
        RECT 0.335 383.870 196.195 384.730 ;
        RECT 0.660 383.050 195.660 383.870 ;
        RECT 0.335 382.190 196.195 383.050 ;
        RECT 0.660 381.370 195.660 382.190 ;
        RECT 0.335 380.510 196.195 381.370 ;
        RECT 0.660 379.690 195.660 380.510 ;
        RECT 0.335 378.830 196.195 379.690 ;
        RECT 0.660 378.010 195.660 378.830 ;
        RECT 0.335 377.150 196.195 378.010 ;
        RECT 0.660 376.330 195.660 377.150 ;
        RECT 0.335 375.470 196.195 376.330 ;
        RECT 0.660 374.650 195.660 375.470 ;
        RECT 0.335 373.790 196.195 374.650 ;
        RECT 0.660 372.970 195.660 373.790 ;
        RECT 0.335 372.110 196.195 372.970 ;
        RECT 0.660 371.290 195.660 372.110 ;
        RECT 0.335 370.430 196.195 371.290 ;
        RECT 0.660 369.610 195.660 370.430 ;
        RECT 0.335 368.750 196.195 369.610 ;
        RECT 0.660 367.930 195.660 368.750 ;
        RECT 0.335 367.070 196.195 367.930 ;
        RECT 0.660 366.250 195.660 367.070 ;
        RECT 0.335 365.390 196.195 366.250 ;
        RECT 0.660 364.570 195.660 365.390 ;
        RECT 0.335 363.710 196.195 364.570 ;
        RECT 0.660 362.890 195.660 363.710 ;
        RECT 0.335 362.030 196.195 362.890 ;
        RECT 0.660 361.210 195.660 362.030 ;
        RECT 0.335 360.350 196.195 361.210 ;
        RECT 0.660 359.530 195.660 360.350 ;
        RECT 0.335 358.670 196.195 359.530 ;
        RECT 0.660 357.850 195.660 358.670 ;
        RECT 0.335 356.990 196.195 357.850 ;
        RECT 0.660 356.170 195.660 356.990 ;
        RECT 0.335 355.310 196.195 356.170 ;
        RECT 0.660 354.490 195.660 355.310 ;
        RECT 0.335 353.630 196.195 354.490 ;
        RECT 0.660 352.810 195.660 353.630 ;
        RECT 0.335 351.950 196.195 352.810 ;
        RECT 0.660 351.130 195.660 351.950 ;
        RECT 0.335 350.270 196.195 351.130 ;
        RECT 0.660 349.450 195.660 350.270 ;
        RECT 0.335 348.590 196.195 349.450 ;
        RECT 0.660 347.770 195.660 348.590 ;
        RECT 0.335 346.910 196.195 347.770 ;
        RECT 0.660 346.090 195.660 346.910 ;
        RECT 0.335 345.230 196.195 346.090 ;
        RECT 0.660 344.410 195.660 345.230 ;
        RECT 0.335 343.550 196.195 344.410 ;
        RECT 0.660 342.730 195.660 343.550 ;
        RECT 0.335 341.870 196.195 342.730 ;
        RECT 0.660 341.050 195.660 341.870 ;
        RECT 0.335 340.190 196.195 341.050 ;
        RECT 0.660 339.370 195.660 340.190 ;
        RECT 0.335 338.510 196.195 339.370 ;
        RECT 0.660 337.690 195.660 338.510 ;
        RECT 0.335 336.830 196.195 337.690 ;
        RECT 0.660 336.010 195.660 336.830 ;
        RECT 0.335 335.150 196.195 336.010 ;
        RECT 0.660 334.330 195.660 335.150 ;
        RECT 0.335 333.470 196.195 334.330 ;
        RECT 0.660 332.650 195.660 333.470 ;
        RECT 0.335 331.790 196.195 332.650 ;
        RECT 0.660 330.970 195.660 331.790 ;
        RECT 0.335 330.110 196.195 330.970 ;
        RECT 0.660 329.290 195.660 330.110 ;
        RECT 0.335 328.430 196.195 329.290 ;
        RECT 0.660 327.610 195.660 328.430 ;
        RECT 0.335 326.750 196.195 327.610 ;
        RECT 0.660 325.930 195.660 326.750 ;
        RECT 0.335 325.070 196.195 325.930 ;
        RECT 0.660 324.250 195.660 325.070 ;
        RECT 0.335 323.390 196.195 324.250 ;
        RECT 0.660 322.570 195.660 323.390 ;
        RECT 0.335 321.710 196.195 322.570 ;
        RECT 0.660 320.890 195.660 321.710 ;
        RECT 0.335 320.030 196.195 320.890 ;
        RECT 0.660 319.210 195.660 320.030 ;
        RECT 0.335 318.350 196.195 319.210 ;
        RECT 0.660 317.530 195.660 318.350 ;
        RECT 0.335 316.670 196.195 317.530 ;
        RECT 0.660 315.850 195.660 316.670 ;
        RECT 0.335 314.990 196.195 315.850 ;
        RECT 0.660 314.170 195.660 314.990 ;
        RECT 0.335 313.310 196.195 314.170 ;
        RECT 0.660 312.490 195.660 313.310 ;
        RECT 0.335 311.630 196.195 312.490 ;
        RECT 0.660 310.810 195.660 311.630 ;
        RECT 0.335 309.950 196.195 310.810 ;
        RECT 0.660 309.130 195.660 309.950 ;
        RECT 0.335 308.270 196.195 309.130 ;
        RECT 0.660 307.450 195.660 308.270 ;
        RECT 0.335 306.590 196.195 307.450 ;
        RECT 0.660 305.770 195.660 306.590 ;
        RECT 0.335 304.910 196.195 305.770 ;
        RECT 0.660 304.090 195.660 304.910 ;
        RECT 0.335 303.230 196.195 304.090 ;
        RECT 0.660 302.410 195.660 303.230 ;
        RECT 0.335 301.550 196.195 302.410 ;
        RECT 0.660 300.730 195.660 301.550 ;
        RECT 0.335 299.870 196.195 300.730 ;
        RECT 0.660 299.050 195.660 299.870 ;
        RECT 0.335 298.190 196.195 299.050 ;
        RECT 0.660 297.370 195.660 298.190 ;
        RECT 0.335 296.510 196.195 297.370 ;
        RECT 0.660 295.690 195.660 296.510 ;
        RECT 0.335 294.830 196.195 295.690 ;
        RECT 0.660 294.010 195.660 294.830 ;
        RECT 0.335 293.150 196.195 294.010 ;
        RECT 0.660 292.330 195.660 293.150 ;
        RECT 0.335 291.470 196.195 292.330 ;
        RECT 0.660 290.650 195.660 291.470 ;
        RECT 0.335 289.790 196.195 290.650 ;
        RECT 0.660 288.970 195.660 289.790 ;
        RECT 0.335 288.110 196.195 288.970 ;
        RECT 0.660 287.290 195.660 288.110 ;
        RECT 0.335 286.430 196.195 287.290 ;
        RECT 0.660 285.610 195.660 286.430 ;
        RECT 0.335 284.750 196.195 285.610 ;
        RECT 0.660 283.930 195.660 284.750 ;
        RECT 0.335 283.070 196.195 283.930 ;
        RECT 0.660 282.250 195.660 283.070 ;
        RECT 0.335 281.390 196.195 282.250 ;
        RECT 0.660 280.570 195.660 281.390 ;
        RECT 0.335 279.710 196.195 280.570 ;
        RECT 0.660 278.890 195.660 279.710 ;
        RECT 0.335 278.030 196.195 278.890 ;
        RECT 0.660 277.210 195.660 278.030 ;
        RECT 0.335 276.350 196.195 277.210 ;
        RECT 0.660 275.530 195.660 276.350 ;
        RECT 0.335 274.670 196.195 275.530 ;
        RECT 0.660 273.850 195.660 274.670 ;
        RECT 0.335 272.990 196.195 273.850 ;
        RECT 0.660 272.170 195.660 272.990 ;
        RECT 0.335 271.310 196.195 272.170 ;
        RECT 0.660 270.490 195.660 271.310 ;
        RECT 0.335 269.630 196.195 270.490 ;
        RECT 0.660 268.810 195.660 269.630 ;
        RECT 0.335 267.950 196.195 268.810 ;
        RECT 0.660 267.130 195.660 267.950 ;
        RECT 0.335 266.270 196.195 267.130 ;
        RECT 0.660 265.450 195.660 266.270 ;
        RECT 0.335 264.590 196.195 265.450 ;
        RECT 0.660 263.770 195.660 264.590 ;
        RECT 0.335 262.910 196.195 263.770 ;
        RECT 0.660 262.090 195.660 262.910 ;
        RECT 0.335 261.230 196.195 262.090 ;
        RECT 0.660 260.410 195.660 261.230 ;
        RECT 0.335 259.550 196.195 260.410 ;
        RECT 0.660 258.730 195.660 259.550 ;
        RECT 0.335 257.870 196.195 258.730 ;
        RECT 0.660 257.050 195.660 257.870 ;
        RECT 0.335 256.190 196.195 257.050 ;
        RECT 0.660 255.370 195.660 256.190 ;
        RECT 0.335 227.630 196.195 255.370 ;
        RECT 0.660 226.810 195.660 227.630 ;
        RECT 0.335 225.950 196.195 226.810 ;
        RECT 0.660 225.130 195.660 225.950 ;
        RECT 0.335 224.270 196.195 225.130 ;
        RECT 0.660 223.450 195.660 224.270 ;
        RECT 0.335 222.590 196.195 223.450 ;
        RECT 0.660 221.770 195.660 222.590 ;
        RECT 0.335 220.910 196.195 221.770 ;
        RECT 0.660 220.090 195.660 220.910 ;
        RECT 0.335 219.230 196.195 220.090 ;
        RECT 0.660 218.410 195.660 219.230 ;
        RECT 0.335 217.550 196.195 218.410 ;
        RECT 0.660 216.730 195.660 217.550 ;
        RECT 0.335 215.870 196.195 216.730 ;
        RECT 0.660 215.050 195.660 215.870 ;
        RECT 0.335 214.190 196.195 215.050 ;
        RECT 0.660 213.370 195.660 214.190 ;
        RECT 0.335 212.510 196.195 213.370 ;
        RECT 0.660 211.690 195.660 212.510 ;
        RECT 0.335 210.830 196.195 211.690 ;
        RECT 0.660 210.010 195.660 210.830 ;
        RECT 0.335 209.150 196.195 210.010 ;
        RECT 0.660 208.330 195.660 209.150 ;
        RECT 0.335 207.470 196.195 208.330 ;
        RECT 0.660 206.650 195.660 207.470 ;
        RECT 0.335 205.790 196.195 206.650 ;
        RECT 0.660 204.970 195.660 205.790 ;
        RECT 0.335 204.110 196.195 204.970 ;
        RECT 0.660 203.290 195.660 204.110 ;
        RECT 0.335 202.430 196.195 203.290 ;
        RECT 0.660 201.610 195.660 202.430 ;
        RECT 0.335 200.750 196.195 201.610 ;
        RECT 0.660 199.930 195.660 200.750 ;
        RECT 0.335 199.070 196.195 199.930 ;
        RECT 0.660 198.250 195.660 199.070 ;
        RECT 0.335 197.390 196.195 198.250 ;
        RECT 0.660 196.570 195.660 197.390 ;
        RECT 0.335 195.710 196.195 196.570 ;
        RECT 0.660 194.890 195.660 195.710 ;
        RECT 0.335 194.030 196.195 194.890 ;
        RECT 0.660 193.210 195.660 194.030 ;
        RECT 0.335 192.350 196.195 193.210 ;
        RECT 0.660 191.530 195.660 192.350 ;
        RECT 0.335 190.670 196.195 191.530 ;
        RECT 0.660 189.850 195.660 190.670 ;
        RECT 0.335 188.990 196.195 189.850 ;
        RECT 0.660 188.170 195.660 188.990 ;
        RECT 0.335 187.310 196.195 188.170 ;
        RECT 0.660 186.490 195.660 187.310 ;
        RECT 0.335 185.630 196.195 186.490 ;
        RECT 0.660 184.810 195.660 185.630 ;
        RECT 0.335 183.950 196.195 184.810 ;
        RECT 0.660 183.130 195.660 183.950 ;
        RECT 0.335 182.270 196.195 183.130 ;
        RECT 0.660 181.450 195.660 182.270 ;
        RECT 0.335 180.590 196.195 181.450 ;
        RECT 0.660 179.770 195.660 180.590 ;
        RECT 0.335 178.910 196.195 179.770 ;
        RECT 0.660 178.090 195.660 178.910 ;
        RECT 0.335 177.230 196.195 178.090 ;
        RECT 0.660 176.410 195.660 177.230 ;
        RECT 0.335 175.550 196.195 176.410 ;
        RECT 0.660 174.730 195.660 175.550 ;
        RECT 0.335 173.870 196.195 174.730 ;
        RECT 0.660 173.050 195.660 173.870 ;
        RECT 0.335 172.190 196.195 173.050 ;
        RECT 0.660 171.370 195.660 172.190 ;
        RECT 0.335 170.510 196.195 171.370 ;
        RECT 0.660 169.690 195.660 170.510 ;
        RECT 0.335 168.830 196.195 169.690 ;
        RECT 0.660 168.010 195.660 168.830 ;
        RECT 0.335 167.150 196.195 168.010 ;
        RECT 0.660 166.330 195.660 167.150 ;
        RECT 0.335 165.470 196.195 166.330 ;
        RECT 0.660 164.650 195.660 165.470 ;
        RECT 0.335 163.790 196.195 164.650 ;
        RECT 0.660 162.970 195.660 163.790 ;
        RECT 0.335 162.110 196.195 162.970 ;
        RECT 0.660 161.290 195.660 162.110 ;
        RECT 0.335 160.430 196.195 161.290 ;
        RECT 0.660 159.610 195.660 160.430 ;
        RECT 0.335 158.750 196.195 159.610 ;
        RECT 0.660 157.930 195.660 158.750 ;
        RECT 0.335 157.070 196.195 157.930 ;
        RECT 0.660 156.250 195.660 157.070 ;
        RECT 0.335 155.390 196.195 156.250 ;
        RECT 0.660 154.570 195.660 155.390 ;
        RECT 0.335 153.710 196.195 154.570 ;
        RECT 0.660 152.890 195.660 153.710 ;
        RECT 0.335 152.030 196.195 152.890 ;
        RECT 0.660 151.210 195.660 152.030 ;
        RECT 0.335 150.350 196.195 151.210 ;
        RECT 0.660 149.530 195.660 150.350 ;
        RECT 0.335 148.670 196.195 149.530 ;
        RECT 0.660 147.850 195.660 148.670 ;
        RECT 0.335 146.990 196.195 147.850 ;
        RECT 0.660 146.170 195.660 146.990 ;
        RECT 0.335 145.310 196.195 146.170 ;
        RECT 0.660 144.490 195.660 145.310 ;
        RECT 0.335 143.630 196.195 144.490 ;
        RECT 0.660 142.810 195.660 143.630 ;
        RECT 0.335 141.950 196.195 142.810 ;
        RECT 0.660 141.130 195.660 141.950 ;
        RECT 0.335 140.270 196.195 141.130 ;
        RECT 0.660 139.450 195.660 140.270 ;
        RECT 0.335 138.590 196.195 139.450 ;
        RECT 0.660 137.770 195.660 138.590 ;
        RECT 0.335 136.910 196.195 137.770 ;
        RECT 0.660 136.090 195.660 136.910 ;
        RECT 0.335 135.230 196.195 136.090 ;
        RECT 0.660 134.410 195.660 135.230 ;
        RECT 0.335 133.550 196.195 134.410 ;
        RECT 0.660 132.730 195.660 133.550 ;
        RECT 0.335 131.870 196.195 132.730 ;
        RECT 0.660 131.050 195.660 131.870 ;
        RECT 0.335 130.190 196.195 131.050 ;
        RECT 0.660 129.370 195.660 130.190 ;
        RECT 0.335 128.510 196.195 129.370 ;
        RECT 0.660 127.690 195.660 128.510 ;
        RECT 0.335 126.830 196.195 127.690 ;
        RECT 0.660 126.010 195.660 126.830 ;
        RECT 0.335 125.150 196.195 126.010 ;
        RECT 0.660 124.330 195.660 125.150 ;
        RECT 0.335 123.470 196.195 124.330 ;
        RECT 0.660 122.650 195.660 123.470 ;
        RECT 0.335 121.790 196.195 122.650 ;
        RECT 0.660 120.970 195.660 121.790 ;
        RECT 0.335 120.110 196.195 120.970 ;
        RECT 0.660 119.290 195.660 120.110 ;
        RECT 0.335 118.430 196.195 119.290 ;
        RECT 0.660 117.610 195.660 118.430 ;
        RECT 0.335 116.750 196.195 117.610 ;
        RECT 0.660 115.930 195.660 116.750 ;
        RECT 0.335 115.070 196.195 115.930 ;
        RECT 0.660 114.250 195.660 115.070 ;
        RECT 0.335 113.390 196.195 114.250 ;
        RECT 0.660 112.570 195.660 113.390 ;
        RECT 0.335 111.710 196.195 112.570 ;
        RECT 0.660 110.890 195.660 111.710 ;
        RECT 0.335 110.030 196.195 110.890 ;
        RECT 0.660 109.210 195.660 110.030 ;
        RECT 0.335 108.350 196.195 109.210 ;
        RECT 0.660 107.530 195.660 108.350 ;
        RECT 0.335 106.670 196.195 107.530 ;
        RECT 0.660 105.850 195.660 106.670 ;
        RECT 0.335 104.990 196.195 105.850 ;
        RECT 0.660 104.170 195.660 104.990 ;
        RECT 0.335 103.310 196.195 104.170 ;
        RECT 0.660 102.490 195.660 103.310 ;
        RECT 0.335 101.630 196.195 102.490 ;
        RECT 0.660 100.810 195.660 101.630 ;
        RECT 0.335 99.950 196.195 100.810 ;
        RECT 0.660 99.130 195.660 99.950 ;
        RECT 0.335 98.270 196.195 99.130 ;
        RECT 0.660 97.450 195.660 98.270 ;
        RECT 0.335 96.590 196.195 97.450 ;
        RECT 0.660 95.770 195.660 96.590 ;
        RECT 0.335 94.910 196.195 95.770 ;
        RECT 0.660 94.090 195.660 94.910 ;
        RECT 0.335 93.230 196.195 94.090 ;
        RECT 0.660 92.410 195.660 93.230 ;
        RECT 0.335 91.550 196.195 92.410 ;
        RECT 0.660 90.730 195.660 91.550 ;
        RECT 0.335 89.870 196.195 90.730 ;
        RECT 0.660 89.050 195.660 89.870 ;
        RECT 0.335 88.190 196.195 89.050 ;
        RECT 0.660 87.370 195.660 88.190 ;
        RECT 0.335 86.510 196.195 87.370 ;
        RECT 0.660 85.690 195.660 86.510 ;
        RECT 0.335 84.830 196.195 85.690 ;
        RECT 0.660 84.010 195.660 84.830 ;
        RECT 0.335 83.150 196.195 84.010 ;
        RECT 0.660 82.330 195.660 83.150 ;
        RECT 0.335 81.470 196.195 82.330 ;
        RECT 0.660 80.650 195.660 81.470 ;
        RECT 0.335 79.790 196.195 80.650 ;
        RECT 0.660 78.970 195.660 79.790 ;
        RECT 0.335 78.110 196.195 78.970 ;
        RECT 0.660 77.290 195.660 78.110 ;
        RECT 0.335 76.430 196.195 77.290 ;
        RECT 0.660 75.610 195.660 76.430 ;
        RECT 0.335 74.750 196.195 75.610 ;
        RECT 0.660 73.930 195.660 74.750 ;
        RECT 0.335 73.070 196.195 73.930 ;
        RECT 0.660 72.250 195.660 73.070 ;
        RECT 0.335 71.390 196.195 72.250 ;
        RECT 0.660 70.570 195.660 71.390 ;
        RECT 0.335 69.710 196.195 70.570 ;
        RECT 0.660 68.890 195.660 69.710 ;
        RECT 0.335 68.030 196.195 68.890 ;
        RECT 0.660 67.210 195.660 68.030 ;
        RECT 0.335 66.350 196.195 67.210 ;
        RECT 0.660 65.530 195.660 66.350 ;
        RECT 0.335 64.670 196.195 65.530 ;
        RECT 0.660 63.850 195.660 64.670 ;
        RECT 0.335 62.990 196.195 63.850 ;
        RECT 0.660 62.170 195.660 62.990 ;
        RECT 0.335 61.310 196.195 62.170 ;
        RECT 0.660 60.490 195.660 61.310 ;
        RECT 0.335 59.630 196.195 60.490 ;
        RECT 0.660 58.810 195.660 59.630 ;
        RECT 0.335 57.950 196.195 58.810 ;
        RECT 0.660 57.130 195.660 57.950 ;
        RECT 0.335 56.270 196.195 57.130 ;
        RECT 0.660 55.450 195.660 56.270 ;
        RECT 0.335 54.590 196.195 55.450 ;
        RECT 0.660 53.770 195.660 54.590 ;
        RECT 0.335 52.910 196.195 53.770 ;
        RECT 0.660 52.090 195.660 52.910 ;
        RECT 0.335 51.230 196.195 52.090 ;
        RECT 0.660 50.410 195.660 51.230 ;
        RECT 0.335 49.550 196.195 50.410 ;
        RECT 0.660 48.730 195.660 49.550 ;
        RECT 0.335 47.870 196.195 48.730 ;
        RECT 0.660 47.050 195.660 47.870 ;
        RECT 0.335 46.190 196.195 47.050 ;
        RECT 0.660 45.370 195.660 46.190 ;
        RECT 0.335 44.510 196.195 45.370 ;
        RECT 0.660 43.690 195.660 44.510 ;
        RECT 0.335 42.830 196.195 43.690 ;
        RECT 0.660 42.010 195.660 42.830 ;
        RECT 0.335 41.150 196.195 42.010 ;
        RECT 0.660 40.330 195.660 41.150 ;
        RECT 0.335 39.470 196.195 40.330 ;
        RECT 0.660 38.650 195.660 39.470 ;
        RECT 0.335 37.790 196.195 38.650 ;
        RECT 0.660 36.970 195.660 37.790 ;
        RECT 0.335 36.110 196.195 36.970 ;
        RECT 0.660 35.290 195.660 36.110 ;
        RECT 0.335 34.430 196.195 35.290 ;
        RECT 0.660 33.610 195.660 34.430 ;
        RECT 0.335 32.750 196.195 33.610 ;
        RECT 0.660 31.930 195.660 32.750 ;
        RECT 0.335 31.070 196.195 31.930 ;
        RECT 0.660 30.250 195.660 31.070 ;
        RECT 0.335 29.390 196.195 30.250 ;
        RECT 0.660 28.570 195.660 29.390 ;
        RECT 0.335 27.710 196.195 28.570 ;
        RECT 0.660 26.890 195.660 27.710 ;
        RECT 0.335 26.030 196.195 26.890 ;
        RECT 0.660 25.210 195.660 26.030 ;
        RECT 0.335 24.350 196.195 25.210 ;
        RECT 0.660 23.530 195.660 24.350 ;
        RECT 0.335 22.670 196.195 23.530 ;
        RECT 0.660 21.850 195.660 22.670 ;
        RECT 0.335 20.990 196.195 21.850 ;
        RECT 0.660 20.170 195.660 20.990 ;
        RECT 0.335 19.310 196.195 20.170 ;
        RECT 0.660 18.490 195.660 19.310 ;
        RECT 0.335 17.630 196.195 18.490 ;
        RECT 0.660 16.810 195.660 17.630 ;
        RECT 0.335 15.950 196.195 16.810 ;
        RECT 0.660 15.130 195.660 15.950 ;
        RECT 0.335 14.270 196.195 15.130 ;
        RECT 0.660 13.450 195.660 14.270 ;
        RECT 0.335 0.320 196.195 13.450 ;
      LAYER Metal3 ;
        RECT 0.380 483.230 37.510 483.565 ;
        RECT 38.330 483.230 38.470 483.565 ;
        RECT 39.290 483.230 39.430 483.565 ;
        RECT 40.250 483.230 40.390 483.565 ;
        RECT 41.210 483.230 41.350 483.565 ;
        RECT 42.170 483.230 42.310 483.565 ;
        RECT 43.130 483.230 43.270 483.565 ;
        RECT 44.090 483.230 44.230 483.565 ;
        RECT 45.050 483.230 45.190 483.565 ;
        RECT 46.010 483.230 46.150 483.565 ;
        RECT 46.970 483.230 47.110 483.565 ;
        RECT 47.930 483.230 48.070 483.565 ;
        RECT 48.890 483.230 49.030 483.565 ;
        RECT 49.850 483.230 49.990 483.565 ;
        RECT 50.810 483.230 50.950 483.565 ;
        RECT 51.770 483.230 51.910 483.565 ;
        RECT 52.730 483.230 52.870 483.565 ;
        RECT 53.690 483.230 53.830 483.565 ;
        RECT 54.650 483.230 54.790 483.565 ;
        RECT 55.610 483.230 55.750 483.565 ;
        RECT 56.570 483.230 56.710 483.565 ;
        RECT 57.530 483.230 57.670 483.565 ;
        RECT 58.490 483.230 58.630 483.565 ;
        RECT 59.450 483.230 59.590 483.565 ;
        RECT 60.410 483.230 60.550 483.565 ;
        RECT 61.370 483.230 61.510 483.565 ;
        RECT 62.330 483.230 62.470 483.565 ;
        RECT 63.290 483.230 63.430 483.565 ;
        RECT 64.250 483.230 64.390 483.565 ;
        RECT 65.210 483.230 65.350 483.565 ;
        RECT 66.170 483.230 66.310 483.565 ;
        RECT 67.130 483.230 67.270 483.565 ;
        RECT 68.090 483.230 68.230 483.565 ;
        RECT 69.050 483.230 69.190 483.565 ;
        RECT 70.010 483.230 70.150 483.565 ;
        RECT 70.970 483.230 71.110 483.565 ;
        RECT 71.930 483.230 72.070 483.565 ;
        RECT 72.890 483.230 73.030 483.565 ;
        RECT 73.850 483.230 73.990 483.565 ;
        RECT 74.810 483.230 74.950 483.565 ;
        RECT 75.770 483.230 75.910 483.565 ;
        RECT 76.730 483.230 76.870 483.565 ;
        RECT 77.690 483.230 77.830 483.565 ;
        RECT 78.650 483.230 78.790 483.565 ;
        RECT 79.610 483.230 79.750 483.565 ;
        RECT 80.570 483.230 80.710 483.565 ;
        RECT 81.530 483.230 81.670 483.565 ;
        RECT 82.490 483.230 82.630 483.565 ;
        RECT 83.450 483.230 83.590 483.565 ;
        RECT 84.410 483.230 84.550 483.565 ;
        RECT 85.370 483.230 85.510 483.565 ;
        RECT 86.330 483.230 86.470 483.565 ;
        RECT 87.290 483.230 87.430 483.565 ;
        RECT 88.250 483.230 88.390 483.565 ;
        RECT 89.210 483.230 89.350 483.565 ;
        RECT 90.170 483.230 90.310 483.565 ;
        RECT 91.130 483.230 91.270 483.565 ;
        RECT 92.090 483.230 92.230 483.565 ;
        RECT 93.050 483.230 93.190 483.565 ;
        RECT 94.010 483.230 94.150 483.565 ;
        RECT 94.970 483.230 95.110 483.565 ;
        RECT 95.930 483.230 96.070 483.565 ;
        RECT 96.890 483.230 97.030 483.565 ;
        RECT 97.850 483.230 97.990 483.565 ;
        RECT 98.810 483.230 98.950 483.565 ;
        RECT 99.770 483.230 99.910 483.565 ;
        RECT 100.730 483.230 100.870 483.565 ;
        RECT 101.690 483.230 101.830 483.565 ;
        RECT 102.650 483.230 102.790 483.565 ;
        RECT 103.610 483.230 103.750 483.565 ;
        RECT 104.570 483.230 104.710 483.565 ;
        RECT 105.530 483.230 105.670 483.565 ;
        RECT 106.490 483.230 106.630 483.565 ;
        RECT 107.450 483.230 107.590 483.565 ;
        RECT 108.410 483.230 108.550 483.565 ;
        RECT 109.370 483.230 109.510 483.565 ;
        RECT 110.330 483.230 110.470 483.565 ;
        RECT 111.290 483.230 111.430 483.565 ;
        RECT 112.250 483.230 112.390 483.565 ;
        RECT 113.210 483.230 113.350 483.565 ;
        RECT 114.170 483.230 114.310 483.565 ;
        RECT 115.130 483.230 115.270 483.565 ;
        RECT 116.090 483.230 116.230 483.565 ;
        RECT 117.050 483.230 117.190 483.565 ;
        RECT 118.010 483.230 118.150 483.565 ;
        RECT 118.970 483.230 119.110 483.565 ;
        RECT 119.930 483.230 120.070 483.565 ;
        RECT 120.890 483.230 121.030 483.565 ;
        RECT 121.850 483.230 121.990 483.565 ;
        RECT 122.810 483.230 122.950 483.565 ;
        RECT 123.770 483.230 123.910 483.565 ;
        RECT 124.730 483.230 124.870 483.565 ;
        RECT 125.690 483.230 125.830 483.565 ;
        RECT 126.650 483.230 126.790 483.565 ;
        RECT 127.610 483.230 127.750 483.565 ;
        RECT 128.570 483.230 128.710 483.565 ;
        RECT 129.530 483.230 129.670 483.565 ;
        RECT 130.490 483.230 130.630 483.565 ;
        RECT 131.450 483.230 131.590 483.565 ;
        RECT 132.410 483.230 132.550 483.565 ;
        RECT 133.370 483.230 133.510 483.565 ;
        RECT 134.330 483.230 134.470 483.565 ;
        RECT 135.290 483.230 135.430 483.565 ;
        RECT 136.250 483.230 136.390 483.565 ;
        RECT 137.210 483.230 137.350 483.565 ;
        RECT 138.170 483.230 138.310 483.565 ;
        RECT 139.130 483.230 139.270 483.565 ;
        RECT 140.090 483.230 140.230 483.565 ;
        RECT 141.050 483.230 141.190 483.565 ;
        RECT 142.010 483.230 142.150 483.565 ;
        RECT 142.970 483.230 143.110 483.565 ;
        RECT 143.930 483.230 144.070 483.565 ;
        RECT 144.890 483.230 145.030 483.565 ;
        RECT 145.850 483.230 145.990 483.565 ;
        RECT 146.810 483.230 146.950 483.565 ;
        RECT 147.770 483.230 147.910 483.565 ;
        RECT 148.730 483.230 148.870 483.565 ;
        RECT 149.690 483.230 149.830 483.565 ;
        RECT 150.650 483.230 150.790 483.565 ;
        RECT 151.610 483.230 151.750 483.565 ;
        RECT 152.570 483.230 152.710 483.565 ;
        RECT 153.530 483.230 153.670 483.565 ;
        RECT 154.490 483.230 154.630 483.565 ;
        RECT 155.450 483.230 155.590 483.565 ;
        RECT 156.410 483.230 156.550 483.565 ;
        RECT 157.370 483.230 195.940 483.565 ;
        RECT 0.380 0.610 195.940 483.230 ;
        RECT 0.380 0.275 37.510 0.610 ;
        RECT 38.330 0.275 38.470 0.610 ;
        RECT 39.290 0.275 39.430 0.610 ;
        RECT 40.250 0.275 40.390 0.610 ;
        RECT 41.210 0.275 41.350 0.610 ;
        RECT 42.170 0.275 42.310 0.610 ;
        RECT 43.130 0.275 43.270 0.610 ;
        RECT 44.090 0.275 44.230 0.610 ;
        RECT 45.050 0.275 45.190 0.610 ;
        RECT 46.010 0.275 46.150 0.610 ;
        RECT 46.970 0.275 47.110 0.610 ;
        RECT 47.930 0.275 48.070 0.610 ;
        RECT 48.890 0.275 49.030 0.610 ;
        RECT 49.850 0.275 49.990 0.610 ;
        RECT 50.810 0.275 50.950 0.610 ;
        RECT 51.770 0.275 51.910 0.610 ;
        RECT 52.730 0.275 52.870 0.610 ;
        RECT 53.690 0.275 53.830 0.610 ;
        RECT 54.650 0.275 54.790 0.610 ;
        RECT 55.610 0.275 55.750 0.610 ;
        RECT 56.570 0.275 56.710 0.610 ;
        RECT 57.530 0.275 57.670 0.610 ;
        RECT 58.490 0.275 58.630 0.610 ;
        RECT 59.450 0.275 59.590 0.610 ;
        RECT 60.410 0.275 60.550 0.610 ;
        RECT 61.370 0.275 61.510 0.610 ;
        RECT 62.330 0.275 62.470 0.610 ;
        RECT 63.290 0.275 63.430 0.610 ;
        RECT 64.250 0.275 64.390 0.610 ;
        RECT 65.210 0.275 65.350 0.610 ;
        RECT 66.170 0.275 66.310 0.610 ;
        RECT 67.130 0.275 67.270 0.610 ;
        RECT 68.090 0.275 68.230 0.610 ;
        RECT 69.050 0.275 69.190 0.610 ;
        RECT 70.010 0.275 70.150 0.610 ;
        RECT 70.970 0.275 71.110 0.610 ;
        RECT 71.930 0.275 72.070 0.610 ;
        RECT 72.890 0.275 73.030 0.610 ;
        RECT 73.850 0.275 73.990 0.610 ;
        RECT 74.810 0.275 74.950 0.610 ;
        RECT 75.770 0.275 75.910 0.610 ;
        RECT 76.730 0.275 76.870 0.610 ;
        RECT 77.690 0.275 77.830 0.610 ;
        RECT 78.650 0.275 78.790 0.610 ;
        RECT 79.610 0.275 79.750 0.610 ;
        RECT 80.570 0.275 80.710 0.610 ;
        RECT 81.530 0.275 81.670 0.610 ;
        RECT 82.490 0.275 82.630 0.610 ;
        RECT 83.450 0.275 83.590 0.610 ;
        RECT 84.410 0.275 84.550 0.610 ;
        RECT 85.370 0.275 85.510 0.610 ;
        RECT 86.330 0.275 86.470 0.610 ;
        RECT 87.290 0.275 87.430 0.610 ;
        RECT 88.250 0.275 88.390 0.610 ;
        RECT 89.210 0.275 89.350 0.610 ;
        RECT 90.170 0.275 90.310 0.610 ;
        RECT 91.130 0.275 91.270 0.610 ;
        RECT 92.090 0.275 92.230 0.610 ;
        RECT 93.050 0.275 93.190 0.610 ;
        RECT 94.010 0.275 94.150 0.610 ;
        RECT 94.970 0.275 95.110 0.610 ;
        RECT 95.930 0.275 96.070 0.610 ;
        RECT 96.890 0.275 97.030 0.610 ;
        RECT 97.850 0.275 97.990 0.610 ;
        RECT 98.810 0.275 98.950 0.610 ;
        RECT 99.770 0.275 99.910 0.610 ;
        RECT 100.730 0.275 100.870 0.610 ;
        RECT 101.690 0.275 101.830 0.610 ;
        RECT 102.650 0.275 102.790 0.610 ;
        RECT 103.610 0.275 103.750 0.610 ;
        RECT 104.570 0.275 104.710 0.610 ;
        RECT 105.530 0.275 105.670 0.610 ;
        RECT 106.490 0.275 106.630 0.610 ;
        RECT 107.450 0.275 107.590 0.610 ;
        RECT 108.410 0.275 108.550 0.610 ;
        RECT 109.370 0.275 109.510 0.610 ;
        RECT 110.330 0.275 110.470 0.610 ;
        RECT 111.290 0.275 111.430 0.610 ;
        RECT 112.250 0.275 112.390 0.610 ;
        RECT 113.210 0.275 113.350 0.610 ;
        RECT 114.170 0.275 114.310 0.610 ;
        RECT 115.130 0.275 115.270 0.610 ;
        RECT 116.090 0.275 116.230 0.610 ;
        RECT 117.050 0.275 117.190 0.610 ;
        RECT 118.010 0.275 118.150 0.610 ;
        RECT 118.970 0.275 119.110 0.610 ;
        RECT 119.930 0.275 120.070 0.610 ;
        RECT 120.890 0.275 121.030 0.610 ;
        RECT 121.850 0.275 121.990 0.610 ;
        RECT 122.810 0.275 122.950 0.610 ;
        RECT 123.770 0.275 123.910 0.610 ;
        RECT 124.730 0.275 124.870 0.610 ;
        RECT 125.690 0.275 125.830 0.610 ;
        RECT 126.650 0.275 126.790 0.610 ;
        RECT 127.610 0.275 127.750 0.610 ;
        RECT 128.570 0.275 128.710 0.610 ;
        RECT 129.530 0.275 129.670 0.610 ;
        RECT 130.490 0.275 130.630 0.610 ;
        RECT 131.450 0.275 131.590 0.610 ;
        RECT 132.410 0.275 132.550 0.610 ;
        RECT 133.370 0.275 133.510 0.610 ;
        RECT 134.330 0.275 134.470 0.610 ;
        RECT 135.290 0.275 135.430 0.610 ;
        RECT 136.250 0.275 136.390 0.610 ;
        RECT 137.210 0.275 137.350 0.610 ;
        RECT 138.170 0.275 138.310 0.610 ;
        RECT 139.130 0.275 139.270 0.610 ;
        RECT 140.090 0.275 140.230 0.610 ;
        RECT 141.050 0.275 141.190 0.610 ;
        RECT 142.010 0.275 142.150 0.610 ;
        RECT 142.970 0.275 143.110 0.610 ;
        RECT 143.930 0.275 144.070 0.610 ;
        RECT 144.890 0.275 145.030 0.610 ;
        RECT 145.850 0.275 145.990 0.610 ;
        RECT 146.810 0.275 146.950 0.610 ;
        RECT 147.770 0.275 147.910 0.610 ;
        RECT 148.730 0.275 148.870 0.610 ;
        RECT 149.690 0.275 149.830 0.610 ;
        RECT 150.650 0.275 150.790 0.610 ;
        RECT 151.610 0.275 151.750 0.610 ;
        RECT 152.570 0.275 152.710 0.610 ;
        RECT 153.530 0.275 153.670 0.610 ;
        RECT 154.490 0.275 154.630 0.610 ;
        RECT 155.450 0.275 155.590 0.610 ;
        RECT 156.410 0.275 156.550 0.610 ;
        RECT 157.370 0.275 195.940 0.610 ;
      LAYER Metal4 ;
        RECT 0.335 0.320 195.985 482.680 ;
      LAYER Metal5 ;
        RECT 0.380 0.275 18.050 482.725 ;
        RECT 20.670 0.275 24.250 482.725 ;
        RECT 26.870 0.275 93.650 482.725 ;
        RECT 96.270 0.275 99.850 482.725 ;
        RECT 102.470 0.275 169.250 482.725 ;
        RECT 171.870 0.275 175.450 482.725 ;
        RECT 178.070 0.275 195.940 482.725 ;
  END
END DSP
END LIBRARY

