* NGSPICE file created from N_term_IHP_SRAM.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

.subckt N_term_IHP_SRAM FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1] N1END[2] N1END[3]
+ N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6] N2END[7] N2MID[0]
+ N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3]
+ S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0]
+ S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S4BEG[0] S4BEG[10]
+ S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4]
+ S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] UserCLK UserCLKo VGND VPWR
XFILLER_7_7 VPWR VGND sg13g2_fill_2
XFILLER_9_159 VPWR VGND sg13g2_decap_8
XFILLER_9_104 VPWR VGND sg13g2_decap_8
X_83_ N4END[4] net75 VPWR VGND sg13g2_buf_1
XFILLER_3_56 VPWR VGND sg13g2_decap_8
XFILLER_8_192 VPWR VGND sg13g2_fill_1
XFILLER_10_169 VPWR VGND sg13g2_fill_1
X_66_ N2END[5] net67 VPWR VGND sg13g2_buf_1
XFILLER_5_162 VPWR VGND sg13g2_fill_2
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_2_110 VPWR VGND sg13g2_decap_8
XFILLER_9_11 VPWR VGND sg13g2_decap_8
X_49_ FrameStrobe[17] net41 VPWR VGND sg13g2_buf_1
XFILLER_6_56 VPWR VGND sg13g2_decap_8
XFILLER_6_89 VPWR VGND sg13g2_decap_8
Xoutput42 net42 FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
Xoutput20 net20 FrameData_O[27] VPWR VGND sg13g2_buf_1
Xoutput75 net75 S4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput86 net86 S4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput64 net64 S2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput53 net53 S1BEG[0] VPWR VGND sg13g2_buf_1
Xoutput31 net31 FrameData_O[8] VPWR VGND sg13g2_buf_1
Xoutput7 net7 FrameData_O[15] VPWR VGND sg13g2_buf_1
XFILLER_3_24 VPWR VGND sg13g2_fill_1
X_82_ N4END[5] net74 VPWR VGND sg13g2_buf_1
X_65_ N2END[6] net66 VPWR VGND sg13g2_buf_1
XFILLER_5_141 VPWR VGND sg13g2_decap_8
XFILLER_9_78 VPWR VGND sg13g2_fill_1
XFILLER_9_67 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
X_48_ FrameStrobe[16] net40 VPWR VGND sg13g2_buf_1
XFILLER_6_13 VPWR VGND sg13g2_decap_8
XFILLER_6_35 VPWR VGND sg13g2_decap_8
XFILLER_6_46 VPWR VGND sg13g2_decap_4
XFILLER_6_79 VPWR VGND sg13g2_fill_1
Xoutput21 net21 FrameData_O[28] VPWR VGND sg13g2_buf_1
Xoutput43 net43 FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
Xoutput76 net76 S4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput87 net87 S4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput65 net65 S2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput54 net54 S1BEG[1] VPWR VGND sg13g2_buf_1
Xoutput32 net32 FrameData_O[9] VPWR VGND sg13g2_buf_1
Xoutput8 net8 FrameData_O[16] VPWR VGND sg13g2_buf_1
Xoutput10 net10 FrameData_O[18] VPWR VGND sg13g2_buf_1
X_81_ N4END[6] net88 VPWR VGND sg13g2_buf_1
XFILLER_3_36 VPWR VGND sg13g2_decap_8
XFILLER_10_116 VPWR VGND sg13g2_decap_8
X_64_ N2END[7] net65 VPWR VGND sg13g2_buf_1
XFILLER_5_120 VPWR VGND sg13g2_decap_8
XFILLER_5_175 VPWR VGND sg13g2_decap_4
XFILLER_2_145 VPWR VGND sg13g2_decap_4
XFILLER_2_167 VPWR VGND sg13g2_decap_8
XFILLER_9_46 VPWR VGND sg13g2_decap_8
X_47_ FrameStrobe[15] net39 VPWR VGND sg13g2_buf_1
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_1_80 VPWR VGND sg13g2_fill_1
Xoutput22 net22 FrameData_O[29] VPWR VGND sg13g2_buf_1
Xoutput44 net44 FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
Xoutput33 net33 FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
Xoutput77 net77 S4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput88 net88 S4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput66 net66 S2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput55 net55 S1BEG[2] VPWR VGND sg13g2_buf_1
Xoutput9 net9 FrameData_O[17] VPWR VGND sg13g2_buf_1
Xoutput11 net11 FrameData_O[19] VPWR VGND sg13g2_buf_1
XFILLER_9_118 VPWR VGND sg13g2_decap_4
X_80_ N4END[7] net87 VPWR VGND sg13g2_buf_1
XFILLER_3_15 VPWR VGND sg13g2_decap_8
XFILLER_8_162 VPWR VGND sg13g2_fill_2
XFILLER_8_173 VPWR VGND sg13g2_fill_1
XFILLER_10_139 VPWR VGND sg13g2_fill_2
XFILLER_5_7 VPWR VGND sg13g2_fill_1
X_63_ N2MID[0] net64 VPWR VGND sg13g2_buf_1
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_2_124 VPWR VGND sg13g2_decap_8
X_46_ FrameStrobe[14] net38 VPWR VGND sg13g2_buf_1
XFILLER_9_25 VPWR VGND sg13g2_decap_8
X_29_ FrameData[29] net22 VPWR VGND sg13g2_buf_1
Xoutput34 net34 FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
Xoutput45 net45 FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
Xoutput89 net89 UserCLKo VPWR VGND sg13g2_buf_1
Xoutput23 net23 FrameData_O[2] VPWR VGND sg13g2_buf_1
Xoutput12 net12 FrameData_O[1] VPWR VGND sg13g2_buf_1
Xoutput78 net78 S4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput67 net67 S2BEGb[2] VPWR VGND sg13g2_buf_1
Xoutput56 net56 S1BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_8_130 VPWR VGND sg13g2_decap_8
XFILLER_8_185 VPWR VGND sg13g2_decap_8
XFILLER_5_155 VPWR VGND sg13g2_decap_8
X_62_ N2MID[1] net63 VPWR VGND sg13g2_buf_1
XFILLER_5_188 VPWR VGND sg13g2_fill_1
XFILLER_2_103 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
X_45_ FrameStrobe[13] net37 VPWR VGND sg13g2_buf_1
X_28_ FrameData[28] net21 VPWR VGND sg13g2_buf_1
Xoutput35 net35 FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
Xoutput46 net46 FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
Xoutput24 net24 FrameData_O[30] VPWR VGND sg13g2_buf_1
Xoutput57 net57 S2BEG[0] VPWR VGND sg13g2_buf_1
Xoutput13 net13 FrameData_O[20] VPWR VGND sg13g2_buf_1
Xoutput79 net79 S4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput68 net68 S2BEGb[3] VPWR VGND sg13g2_buf_1
XFILLER_11_4 VPWR VGND sg13g2_decap_4
XFILLER_8_164 VPWR VGND sg13g2_fill_1
XFILLER_5_134 VPWR VGND sg13g2_decap_8
X_61_ N2MID[2] net62 VPWR VGND sg13g2_buf_1
XFILLER_4_71 VPWR VGND sg13g2_decap_8
XFILLER_4_93 VPWR VGND sg13g2_decap_8
X_44_ FrameStrobe[12] net36 VPWR VGND sg13g2_buf_1
X_27_ FrameData[27] net20 VPWR VGND sg13g2_buf_1
XFILLER_6_28 VPWR VGND sg13g2_decap_8
Xoutput36 net36 FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
Xoutput47 net47 FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
Xoutput25 net25 FrameData_O[31] VPWR VGND sg13g2_buf_1
Xoutput69 net69 S2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput58 net58 S2BEG[1] VPWR VGND sg13g2_buf_1
Xoutput14 net14 FrameData_O[21] VPWR VGND sg13g2_buf_1
XFILLER_7_93 VPWR VGND sg13g2_decap_8
XFILLER_3_29 VPWR VGND sg13g2_decap_8
XFILLER_10_109 VPWR VGND sg13g2_decap_8
XFILLER_5_113 VPWR VGND sg13g2_decap_8
XFILLER_5_168 VPWR VGND sg13g2_decap_8
XFILLER_5_179 VPWR VGND sg13g2_fill_1
X_60_ N2MID[3] net61 VPWR VGND sg13g2_buf_1
XFILLER_4_50 VPWR VGND sg13g2_decap_8
XFILLER_9_39 VPWR VGND sg13g2_decap_8
XFILLER_2_138 VPWR VGND sg13g2_decap_8
XFILLER_3_7 VPWR VGND sg13g2_decap_4
X_43_ FrameStrobe[11] net35 VPWR VGND sg13g2_buf_1
X_26_ FrameData[26] net19 VPWR VGND sg13g2_buf_1
XFILLER_1_73 VPWR VGND sg13g2_decap_8
XFILLER_10_93 VPWR VGND sg13g2_decap_8
X_09_ FrameData[9] net32 VPWR VGND sg13g2_buf_1
Xoutput37 net37 FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
Xoutput48 net48 FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
Xoutput15 net15 FrameData_O[22] VPWR VGND sg13g2_buf_1
Xoutput26 net26 FrameData_O[3] VPWR VGND sg13g2_buf_1
Xoutput59 net59 S2BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_7_72 VPWR VGND sg13g2_decap_8
XFILLER_8_144 VPWR VGND sg13g2_fill_2
XFILLER_8_155 VPWR VGND sg13g2_decap_8
XFILLER_4_180 VPWR VGND sg13g2_fill_2
XFILLER_9_18 VPWR VGND sg13g2_decap_8
XFILLER_2_117 VPWR VGND sg13g2_decap_8
X_42_ FrameStrobe[10] net34 VPWR VGND sg13g2_buf_1
XFILLER_1_183 VPWR VGND sg13g2_fill_1
XFILLER_1_172 VPWR VGND sg13g2_decap_8
XFILLER_1_52 VPWR VGND sg13g2_decap_8
X_25_ FrameData[25] net18 VPWR VGND sg13g2_buf_1
XFILLER_10_72 VPWR VGND sg13g2_decap_8
X_08_ FrameData[8] net31 VPWR VGND sg13g2_buf_1
Xoutput38 net38 FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
Xoutput49 net49 FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
Xoutput16 net16 FrameData_O[23] VPWR VGND sg13g2_buf_1
Xoutput27 net27 FrameData_O[4] VPWR VGND sg13g2_buf_1
XFILLER_8_123 VPWR VGND sg13g2_decap_8
XFILLER_8_178 VPWR VGND sg13g2_decap_8
XFILLER_5_148 VPWR VGND sg13g2_fill_2
X_41_ FrameStrobe[9] net52 VPWR VGND sg13g2_buf_1
XFILLER_1_31 VPWR VGND sg13g2_decap_8
X_24_ FrameData[24] net17 VPWR VGND sg13g2_buf_1
XFILLER_10_51 VPWR VGND sg13g2_decap_8
Xoutput39 net39 FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
Xoutput17 net17 FrameData_O[24] VPWR VGND sg13g2_buf_1
Xoutput28 net28 FrameData_O[5] VPWR VGND sg13g2_buf_1
X_07_ FrameData[7] net30 VPWR VGND sg13g2_buf_1
XFILLER_11_8 VPWR VGND sg13g2_fill_1
XFILLER_7_63 VPWR VGND sg13g2_fill_1
XFILLER_8_102 VPWR VGND sg13g2_decap_8
XFILLER_8_146 VPWR VGND sg13g2_fill_1
XFILLER_5_127 VPWR VGND sg13g2_decap_8
XFILLER_4_64 VPWR VGND sg13g2_decap_8
XFILLER_4_86 VPWR VGND sg13g2_decap_8
X_40_ FrameStrobe[8] net51 VPWR VGND sg13g2_buf_1
XFILLER_1_196 VPWR VGND sg13g2_fill_1
XFILLER_8_0 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_fill_2
X_23_ FrameData[23] net16 VPWR VGND sg13g2_buf_1
XFILLER_10_30 VPWR VGND sg13g2_decap_8
Xoutput18 net18 FrameData_O[25] VPWR VGND sg13g2_buf_1
Xoutput29 net29 FrameData_O[6] VPWR VGND sg13g2_buf_1
X_06_ FrameData[6] net29 VPWR VGND sg13g2_buf_1
XFILLER_7_20 VPWR VGND sg13g2_decap_8
XFILLER_7_42 VPWR VGND sg13g2_decap_8
XFILLER_7_86 VPWR VGND sg13g2_decap_8
XFILLER_8_169 VPWR VGND sg13g2_decap_4
XFILLER_5_106 VPWR VGND sg13g2_decap_8
XFILLER_4_21 VPWR VGND sg13g2_decap_8
XFILLER_4_43 VPWR VGND sg13g2_decap_8
XFILLER_4_194 VPWR VGND sg13g2_fill_2
XFILLER_1_66 VPWR VGND sg13g2_decap_8
X_22_ FrameData[22] net15 VPWR VGND sg13g2_buf_1
XFILLER_10_86 VPWR VGND sg13g2_decap_8
X_05_ FrameData[5] net28 VPWR VGND sg13g2_buf_1
Xoutput19 net19 FrameData_O[26] VPWR VGND sg13g2_buf_1
XFILLER_8_137 VPWR VGND sg13g2_decap_8
X_21_ FrameData[21] net14 VPWR VGND sg13g2_buf_1
XFILLER_1_45 VPWR VGND sg13g2_decap_8
XFILLER_10_65 VPWR VGND sg13g2_decap_8
X_04_ FrameData[4] net27 VPWR VGND sg13g2_buf_1
XFILLER_8_116 VPWR VGND sg13g2_decap_8
XFILLER_7_171 VPWR VGND sg13g2_decap_8
XFILLER_4_163 VPWR VGND sg13g2_fill_2
XFILLER_4_196 VPWR VGND sg13g2_fill_1
XFILLER_6_0 VPWR VGND sg13g2_decap_8
XFILLER_1_24 VPWR VGND sg13g2_decap_8
X_20_ FrameData[20] net13 VPWR VGND sg13g2_buf_1
XFILLER_10_44 VPWR VGND sg13g2_decap_8
XFILLER_10_11 VPWR VGND sg13g2_fill_1
X_03_ FrameData[3] net26 VPWR VGND sg13g2_buf_1
XFILLER_7_34 VPWR VGND sg13g2_decap_4
XFILLER_7_56 VPWR VGND sg13g2_decap_8
XFILLER_7_150 VPWR VGND sg13g2_decap_8
XFILLER_4_35 VPWR VGND sg13g2_decap_4
XFILLER_4_57 VPWR VGND sg13g2_decap_8
XFILLER_4_142 VPWR VGND sg13g2_decap_8
XFILLER_1_156 VPWR VGND sg13g2_decap_4
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_10_23 VPWR VGND sg13g2_decap_8
X_79_ N4END[8] net86 VPWR VGND sg13g2_buf_1
X_02_ FrameData[2] net23 VPWR VGND sg13g2_buf_1
XFILLER_7_13 VPWR VGND sg13g2_decap_8
XFILLER_7_79 VPWR VGND sg13g2_decap_8
XFILLER_4_14 VPWR VGND sg13g2_decap_8
XFILLER_4_121 VPWR VGND sg13g2_decap_8
XFILLER_4_176 VPWR VGND sg13g2_decap_4
XFILLER_1_179 VPWR VGND sg13g2_decap_4
XFILLER_1_59 VPWR VGND sg13g2_decap_8
X_78_ N4END[9] net85 VPWR VGND sg13g2_buf_1
XFILLER_10_79 VPWR VGND sg13g2_decap_8
X_01_ FrameData[1] net12 VPWR VGND sg13g2_buf_1
XFILLER_7_185 VPWR VGND sg13g2_fill_1
XFILLER_4_100 VPWR VGND sg13g2_decap_8
XFILLER_1_147 VPWR VGND sg13g2_fill_1
XFILLER_1_38 VPWR VGND sg13g2_decap_8
X_77_ N4END[10] net84 VPWR VGND sg13g2_buf_1
XFILLER_10_58 VPWR VGND sg13g2_decap_8
X_00_ FrameData[0] net1 VPWR VGND sg13g2_buf_1
XFILLER_4_0 VPWR VGND sg13g2_decap_8
XFILLER_8_109 VPWR VGND sg13g2_decap_8
XFILLER_7_142 VPWR VGND sg13g2_decap_4
XFILLER_7_164 VPWR VGND sg13g2_decap_8
XFILLER_4_156 VPWR VGND sg13g2_decap_8
XFILLER_8_7 VPWR VGND sg13g2_fill_1
XFILLER_5_92 VPWR VGND sg13g2_decap_8
XFILLER_1_17 VPWR VGND sg13g2_decap_8
X_76_ N4END[11] net83 VPWR VGND sg13g2_buf_1
XFILLER_10_37 VPWR VGND sg13g2_decap_8
XFILLER_2_82 VPWR VGND sg13g2_decap_8
X_59_ N2MID[4] net60 VPWR VGND sg13g2_buf_1
XFILLER_7_27 VPWR VGND sg13g2_decap_8
XFILLER_7_49 VPWR VGND sg13g2_decap_8
XFILLER_11_183 VPWR VGND sg13g2_fill_2
XFILLER_7_121 VPWR VGND sg13g2_decap_8
XFILLER_7_198 VPWR VGND sg13g2_fill_2
XFILLER_4_28 VPWR VGND sg13g2_decap_8
XFILLER_4_135 VPWR VGND sg13g2_decap_8
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_10_16 VPWR VGND sg13g2_decap_8
X_75_ N4END[12] net82 VPWR VGND sg13g2_buf_1
XFILLER_2_61 VPWR VGND sg13g2_decap_8
X_58_ N2MID[5] net59 VPWR VGND sg13g2_buf_1
XFILLER_11_173 VPWR VGND sg13g2_fill_2
XFILLER_7_100 VPWR VGND sg13g2_decap_8
XFILLER_8_71 VPWR VGND sg13g2_decap_4
XFILLER_4_114 VPWR VGND sg13g2_decap_8
XFILLER_4_169 VPWR VGND sg13g2_decap_8
XFILLER_0_172 VPWR VGND sg13g2_decap_4
XFILLER_5_61 VPWR VGND sg13g2_decap_8
X_74_ N4END[13] net81 VPWR VGND sg13g2_buf_1
X_57_ N2MID[6] net58 VPWR VGND sg13g2_buf_1
XFILLER_11_93 VPWR VGND sg13g2_decap_4
XFILLER_2_0 VPWR VGND sg13g2_decap_8
XFILLER_11_163 VPWR VGND sg13g2_decap_4
XFILLER_7_178 VPWR VGND sg13g2_decap_8
XFILLER_5_40 VPWR VGND sg13g2_decap_8
XFILLER_6_7 VPWR VGND sg13g2_fill_2
X_73_ N4END[14] net80 VPWR VGND sg13g2_buf_1
XFILLER_2_96 VPWR VGND sg13g2_decap_8
X_56_ N2MID[7] net57 VPWR VGND sg13g2_buf_1
XFILLER_11_83 VPWR VGND sg13g2_decap_4
X_39_ FrameStrobe[7] net50 VPWR VGND sg13g2_buf_1
XFILLER_11_153 VPWR VGND sg13g2_decap_4
XFILLER_7_135 VPWR VGND sg13g2_decap_8
XFILLER_7_157 VPWR VGND sg13g2_decap_8
XFILLER_8_62 VPWR VGND sg13g2_decap_4
XFILLER_8_95 VPWR VGND sg13g2_decap_8
XFILLER_4_149 VPWR VGND sg13g2_decap_8
XFILLER_3_160 VPWR VGND sg13g2_decap_8
XFILLER_3_171 VPWR VGND sg13g2_fill_1
XFILLER_5_85 VPWR VGND sg13g2_decap_8
XFILLER_10_0 VPWR VGND sg13g2_decap_8
X_72_ N4END[15] net73 VPWR VGND sg13g2_buf_1
XFILLER_2_31 VPWR VGND sg13g2_decap_8
X_55_ N1END[0] net56 VPWR VGND sg13g2_buf_1
XFILLER_2_75 VPWR VGND sg13g2_decap_8
XFILLER_11_73 VPWR VGND sg13g2_decap_4
X_38_ FrameStrobe[6] net49 VPWR VGND sg13g2_buf_1
XFILLER_11_143 VPWR VGND sg13g2_decap_4
XFILLER_7_114 VPWR VGND sg13g2_decap_8
XFILLER_8_52 VPWR VGND sg13g2_decap_4
XFILLER_8_85 VPWR VGND sg13g2_decap_4
XFILLER_4_128 VPWR VGND sg13g2_decap_8
XFILLER_3_183 VPWR VGND sg13g2_fill_2
XFILLER_3_194 VPWR VGND sg13g2_fill_2
XFILLER_5_31 VPWR VGND sg13g2_decap_4
XFILLER_5_75 VPWR VGND sg13g2_decap_4
X_71_ N2END[0] net72 VPWR VGND sg13g2_buf_1
X_54_ N1END[1] net55 VPWR VGND sg13g2_buf_1
XFILLER_2_54 VPWR VGND sg13g2_decap_8
XFILLER_11_63 VPWR VGND sg13g2_decap_4
X_37_ FrameStrobe[5] net48 VPWR VGND sg13g2_buf_1
XFILLER_11_133 VPWR VGND sg13g2_decap_4
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_6_192 VPWR VGND sg13g2_fill_1
XFILLER_4_107 VPWR VGND sg13g2_decap_8
XFILLER_0_176 VPWR VGND sg13g2_fill_1
XFILLER_0_165 VPWR VGND sg13g2_decap_8
XFILLER_5_54 VPWR VGND sg13g2_decap_8
X_70_ N2END[1] net71 VPWR VGND sg13g2_buf_1
XFILLER_4_7 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_fill_2
X_53_ N1END[2] net54 VPWR VGND sg13g2_buf_1
XFILLER_11_97 VPWR VGND sg13g2_fill_2
XFILLER_11_53 VPWR VGND sg13g2_decap_4
X_36_ FrameStrobe[4] net47 VPWR VGND sg13g2_buf_1
XFILLER_11_167 VPWR VGND sg13g2_fill_2
XFILLER_11_123 VPWR VGND sg13g2_decap_4
XFILLER_6_160 VPWR VGND sg13g2_fill_1
X_19_ FrameData[19] net11 VPWR VGND sg13g2_buf_1
XFILLER_3_185 VPWR VGND sg13g2_fill_1
XFILLER_3_196 VPWR VGND sg13g2_fill_1
XFILLER_5_99 VPWR VGND sg13g2_decap_8
XFILLER_2_45 VPWR VGND sg13g2_decap_4
XFILLER_2_89 VPWR VGND sg13g2_decap_8
X_52_ N1END[3] net53 VPWR VGND sg13g2_buf_1
XFILLER_11_87 VPWR VGND sg13g2_fill_2
XFILLER_11_43 VPWR VGND sg13g2_decap_4
X_35_ FrameStrobe[3] net46 VPWR VGND sg13g2_buf_1
XFILLER_11_157 VPWR VGND sg13g2_fill_2
XFILLER_11_113 VPWR VGND sg13g2_decap_4
XFILLER_7_128 VPWR VGND sg13g2_decap_8
XFILLER_6_183 VPWR VGND sg13g2_decap_4
XFILLER_8_33 VPWR VGND sg13g2_fill_1
XFILLER_8_66 VPWR VGND sg13g2_fill_1
X_18_ FrameData[18] net10 VPWR VGND sg13g2_buf_1
XFILLER_3_131 VPWR VGND sg13g2_fill_2
XFILLER_3_142 VPWR VGND sg13g2_decap_8
XFILLER_5_12 VPWR VGND sg13g2_fill_1
X_51_ FrameStrobe[19] net43 VPWR VGND sg13g2_buf_1
XFILLER_2_24 VPWR VGND sg13g2_decap_8
XFILLER_2_68 VPWR VGND sg13g2_decap_8
XFILLER_11_77 VPWR VGND sg13g2_fill_2
XFILLER_11_33 VPWR VGND sg13g2_decap_4
X_34_ FrameStrobe[2] net45 VPWR VGND sg13g2_buf_1
XFILLER_11_103 VPWR VGND sg13g2_decap_4
XFILLER_11_147 VPWR VGND sg13g2_fill_2
XFILLER_7_107 VPWR VGND sg13g2_decap_8
XFILLER_8_12 VPWR VGND sg13g2_decap_8
XFILLER_8_45 VPWR VGND sg13g2_decap_8
XFILLER_8_56 VPWR VGND sg13g2_fill_2
XFILLER_8_89 VPWR VGND sg13g2_fill_2
X_17_ FrameData[17] net9 VPWR VGND sg13g2_buf_1
XFILLER_3_176 VPWR VGND sg13g2_decap_8
XFILLER_5_24 VPWR VGND sg13g2_decap_8
XFILLER_5_35 VPWR VGND sg13g2_fill_1
XFILLER_5_68 VPWR VGND sg13g2_decap_8
XFILLER_5_79 VPWR VGND sg13g2_fill_2
X_50_ FrameStrobe[18] net42 VPWR VGND sg13g2_buf_1
XFILLER_9_0 VPWR VGND sg13g2_decap_8
XFILLER_11_67 VPWR VGND sg13g2_fill_2
XFILLER_11_23 VPWR VGND sg13g2_decap_4
XFILLER_2_7 VPWR VGND sg13g2_decap_4
X_33_ FrameStrobe[1] net44 VPWR VGND sg13g2_buf_1
XFILLER_9_171 VPWR VGND sg13g2_decap_8
XFILLER_11_137 VPWR VGND sg13g2_fill_2
X_16_ FrameData[16] net8 VPWR VGND sg13g2_buf_1
XFILLER_8_79 VPWR VGND sg13g2_fill_2
XFILLER_3_133 VPWR VGND sg13g2_fill_1
XFILLER_5_47 VPWR VGND sg13g2_decap_8
XFILLER_11_57 VPWR VGND sg13g2_fill_2
XFILLER_11_13 VPWR VGND sg13g2_decap_4
X_32_ FrameStrobe[0] net33 VPWR VGND sg13g2_buf_1
XFILLER_11_127 VPWR VGND sg13g2_fill_2
XFILLER_3_91 VPWR VGND sg13g2_fill_2
XFILLER_6_142 VPWR VGND sg13g2_decap_8
X_15_ FrameData[15] net7 VPWR VGND sg13g2_buf_1
XFILLER_3_123 VPWR VGND sg13g2_decap_4
XFILLER_3_167 VPWR VGND sg13g2_decap_4
XFILLER_9_90 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_fill_2
XFILLER_10_7 VPWR VGND sg13g2_decap_4
XFILLER_2_38 VPWR VGND sg13g2_decap_8
XFILLER_2_49 VPWR VGND sg13g2_fill_1
XFILLER_11_47 VPWR VGND sg13g2_fill_2
X_31_ FrameData[31] net25 VPWR VGND sg13g2_buf_1
XFILLER_11_117 VPWR VGND sg13g2_fill_2
XFILLER_3_70 VPWR VGND sg13g2_decap_8
XFILLER_6_110 VPWR VGND sg13g2_decap_8
XFILLER_6_132 VPWR VGND sg13g2_decap_4
XFILLER_6_176 VPWR VGND sg13g2_decap_8
XFILLER_6_187 VPWR VGND sg13g2_fill_1
XFILLER_8_26 VPWR VGND sg13g2_decap_8
X_14_ FrameData[14] net6 VPWR VGND sg13g2_buf_1
XFILLER_3_102 VPWR VGND sg13g2_decap_4
XFILLER_6_70 VPWR VGND sg13g2_decap_8
XFILLER_2_17 VPWR VGND sg13g2_decap_8
XFILLER_11_37 VPWR VGND sg13g2_fill_2
XFILLER_9_152 VPWR VGND sg13g2_decap_8
X_30_ FrameData[30] net24 VPWR VGND sg13g2_buf_1
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_11_107 VPWR VGND sg13g2_fill_2
XFILLER_3_93 VPWR VGND sg13g2_fill_1
XFILLER_10_162 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_8_38 VPWR VGND sg13g2_decap_8
X_13_ FrameData[13] net5 VPWR VGND sg13g2_buf_1
XFILLER_0_72 VPWR VGND sg13g2_fill_1
XFILLER_5_17 VPWR VGND sg13g2_decap_8
XFILLER_11_27 VPWR VGND sg13g2_fill_2
XFILLER_9_142 VPWR VGND sg13g2_decap_4
XFILLER_3_50 VPWR VGND sg13g2_fill_2
XFILLER_10_141 VPWR VGND sg13g2_fill_1
XFILLER_10_130 VPWR VGND sg13g2_fill_1
XFILLER_10_196 VPWR VGND sg13g2_fill_1
XFILLER_10_174 VPWR VGND sg13g2_fill_2
XFILLER_6_156 VPWR VGND sg13g2_decap_4
X_12_ FrameData[12] net4 VPWR VGND sg13g2_buf_1
XFILLER_2_181 VPWR VGND sg13g2_decap_4
XFILLER_9_60 VPWR VGND sg13g2_decap_8
XFILLER_6_50 VPWR VGND sg13g2_fill_2
Xoutput1 net1 FrameData_O[0] VPWR VGND sg13g2_buf_1
XFILLER_11_17 VPWR VGND sg13g2_fill_2
Xoutput80 net80 S4BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_3_84 VPWR VGND sg13g2_decap_8
X_88_ UserCLK net89 VPWR VGND sg13g2_buf_1
XFILLER_10_153 VPWR VGND sg13g2_decap_4
X_11_ FrameData[11] net3 VPWR VGND sg13g2_buf_1
XFILLER_3_116 VPWR VGND sg13g2_decap_8
XFILLER_3_149 VPWR VGND sg13g2_decap_8
XFILLER_9_83 VPWR VGND sg13g2_decap_8
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_2_160 VPWR VGND sg13g2_fill_2
XFILLER_6_84 VPWR VGND sg13g2_fill_1
Xoutput81 net81 S4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput70 net70 S2BEGb[5] VPWR VGND sg13g2_buf_1
Xoutput2 net2 FrameData_O[10] VPWR VGND sg13g2_buf_1
XFILLER_9_166 VPWR VGND sg13g2_fill_1
XFILLER_9_122 VPWR VGND sg13g2_fill_1
XFILLER_9_111 VPWR VGND sg13g2_decap_8
XFILLER_3_63 VPWR VGND sg13g2_decap_8
X_87_ N4END[0] net79 VPWR VGND sg13g2_buf_1
X_10_ FrameData[10] net2 VPWR VGND sg13g2_buf_1
XFILLER_5_0 VPWR VGND sg13g2_decap_8
XFILLER_6_103 VPWR VGND sg13g2_decap_8
XFILLER_6_125 VPWR VGND sg13g2_decap_8
XFILLER_6_136 VPWR VGND sg13g2_fill_2
XFILLER_6_169 VPWR VGND sg13g2_decap_8
XFILLER_8_19 VPWR VGND sg13g2_decap_8
XFILLER_3_106 VPWR VGND sg13g2_fill_2
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_6_63 VPWR VGND sg13g2_decap_8
XFILLER_6_96 VPWR VGND sg13g2_decap_8
Xoutput82 net82 S4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput71 net71 S2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput60 net60 S2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput3 net3 FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_9_178 VPWR VGND sg13g2_decap_8
X_86_ N4END[1] net78 VPWR VGND sg13g2_buf_1
XFILLER_10_100 VPWR VGND sg13g2_fill_1
X_69_ N2END[2] net70 VPWR VGND sg13g2_buf_1
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_2_162 VPWR VGND sg13g2_fill_1
XFILLER_9_74 VPWR VGND sg13g2_decap_4
XFILLER_6_20 VPWR VGND sg13g2_decap_4
Xoutput50 net50 FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
Xoutput83 net83 S4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput72 net72 S2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput61 net61 S2BEG[4] VPWR VGND sg13g2_buf_1
Xoutput4 net4 FrameData_O[12] VPWR VGND sg13g2_buf_1
XFILLER_9_146 VPWR VGND sg13g2_fill_2
XFILLER_9_135 VPWR VGND sg13g2_decap_8
XFILLER_3_43 VPWR VGND sg13g2_decap_8
X_85_ N4END[2] net77 VPWR VGND sg13g2_buf_1
XFILLER_10_123 VPWR VGND sg13g2_decap_8
XFILLER_6_149 VPWR VGND sg13g2_decap_8
X_68_ N2END[3] net69 VPWR VGND sg13g2_buf_1
XFILLER_2_174 VPWR VGND sg13g2_decap_8
XFILLER_9_97 VPWR VGND sg13g2_decap_8
XFILLER_9_53 VPWR VGND sg13g2_decap_8
XFILLER_7_200 VPWR VGND sg13g2_fill_1
Xoutput40 net40 FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
Xoutput51 net51 FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
Xoutput84 net84 S4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput73 net73 S4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput62 net62 S2BEG[5] VPWR VGND sg13g2_buf_1
Xoutput5 net5 FrameData_O[13] VPWR VGND sg13g2_buf_1
X_84_ N4END[3] net76 VPWR VGND sg13g2_buf_1
XFILLER_3_22 VPWR VGND sg13g2_fill_2
XFILLER_3_77 VPWR VGND sg13g2_decap_8
XFILLER_10_157 VPWR VGND sg13g2_fill_1
XFILLER_10_146 VPWR VGND sg13g2_decap_8
XFILLER_6_117 VPWR VGND sg13g2_decap_4
XFILLER_5_150 VPWR VGND sg13g2_fill_1
X_67_ N2END[4] net68 VPWR VGND sg13g2_buf_1
XFILLER_2_131 VPWR VGND sg13g2_decap_8
XFILLER_2_153 VPWR VGND sg13g2_decap_8
XFILLER_3_0 VPWR VGND sg13g2_decap_8
XFILLER_9_32 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_6_77 VPWR VGND sg13g2_fill_2
Xoutput41 net41 FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
Xoutput52 net52 FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
Xoutput30 net30 FrameData_O[7] VPWR VGND sg13g2_buf_1
Xoutput6 net6 FrameData_O[14] VPWR VGND sg13g2_buf_1
Xoutput74 net74 S4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput85 net85 S4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput63 net63 S2BEG[6] VPWR VGND sg13g2_buf_1
.ends

