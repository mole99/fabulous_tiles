module N_term_single2 (UserCLK,
    UserCLKo,
    VPWR,
    VGND,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1END,
    N2END,
    N2MID,
    N4END,
    NN4END,
    S1BEG,
    S2BEG,
    S2BEGb,
    S4BEG,
    SS4BEG);
 input UserCLK;
 output UserCLKo;
 inout VPWR;
 inout VGND;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] N1END;
 input [7:0] N2END;
 input [7:0] N2MID;
 input [15:0] N4END;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 output [15:0] S4BEG;
 output [15:0] SS4BEG;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;

 sg13g2_buf_1 _000_ (.A(FrameData[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _001_ (.A(FrameData[1]),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _002_ (.A(FrameData[2]),
    .X(net23),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _003_ (.A(FrameData[3]),
    .X(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _004_ (.A(FrameData[4]),
    .X(net27),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _005_ (.A(FrameData[5]),
    .X(net28),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _006_ (.A(FrameData[6]),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _007_ (.A(FrameData[7]),
    .X(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _008_ (.A(FrameData[8]),
    .X(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _009_ (.A(FrameData[9]),
    .X(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _010_ (.A(FrameData[10]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _011_ (.A(FrameData[11]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _012_ (.A(FrameData[12]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _013_ (.A(FrameData[13]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _014_ (.A(FrameData[14]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _015_ (.A(FrameData[15]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _016_ (.A(FrameData[16]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _017_ (.A(FrameData[17]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _018_ (.A(FrameData[18]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _019_ (.A(FrameData[19]),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _020_ (.A(FrameData[20]),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _021_ (.A(FrameData[21]),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _022_ (.A(FrameData[22]),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _023_ (.A(FrameData[23]),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _024_ (.A(FrameData[24]),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _025_ (.A(FrameData[25]),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _026_ (.A(FrameData[26]),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _027_ (.A(FrameData[27]),
    .X(net20),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _028_ (.A(FrameData[28]),
    .X(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _029_ (.A(FrameData[29]),
    .X(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _030_ (.A(FrameData[30]),
    .X(net24),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _031_ (.A(FrameData[31]),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _032_ (.A(FrameStrobe[0]),
    .X(net33),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _033_ (.A(FrameStrobe[1]),
    .X(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _034_ (.A(FrameStrobe[2]),
    .X(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _035_ (.A(FrameStrobe[3]),
    .X(net46),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _036_ (.A(FrameStrobe[4]),
    .X(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _037_ (.A(FrameStrobe[5]),
    .X(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _038_ (.A(FrameStrobe[6]),
    .X(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _039_ (.A(FrameStrobe[7]),
    .X(net50),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _040_ (.A(FrameStrobe[8]),
    .X(net51),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _041_ (.A(FrameStrobe[9]),
    .X(net52),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _042_ (.A(FrameStrobe[10]),
    .X(net34),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _043_ (.A(FrameStrobe[11]),
    .X(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _044_ (.A(FrameStrobe[12]),
    .X(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _045_ (.A(FrameStrobe[13]),
    .X(net37),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _046_ (.A(FrameStrobe[14]),
    .X(net38),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _047_ (.A(FrameStrobe[15]),
    .X(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _048_ (.A(FrameStrobe[16]),
    .X(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _049_ (.A(FrameStrobe[17]),
    .X(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _050_ (.A(FrameStrobe[18]),
    .X(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _051_ (.A(FrameStrobe[19]),
    .X(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _052_ (.A(N1END[3]),
    .X(net53),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _053_ (.A(N1END[2]),
    .X(net54),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _054_ (.A(N1END[1]),
    .X(net55),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _055_ (.A(N1END[0]),
    .X(net56),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _056_ (.A(N2MID[7]),
    .X(net57),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _057_ (.A(N2MID[6]),
    .X(net58),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _058_ (.A(N2MID[5]),
    .X(net59),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _059_ (.A(N2MID[4]),
    .X(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _060_ (.A(N2MID[3]),
    .X(net61),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _061_ (.A(N2MID[2]),
    .X(net62),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _062_ (.A(N2MID[1]),
    .X(net63),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _063_ (.A(N2MID[0]),
    .X(net64),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _064_ (.A(N2END[7]),
    .X(net65),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _065_ (.A(N2END[6]),
    .X(net66),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _066_ (.A(N2END[5]),
    .X(net67),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _067_ (.A(N2END[4]),
    .X(net68),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _068_ (.A(N2END[3]),
    .X(net69),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _069_ (.A(N2END[2]),
    .X(net70),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _070_ (.A(N2END[1]),
    .X(net71),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _071_ (.A(N2END[0]),
    .X(net72),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _072_ (.A(N4END[15]),
    .X(net73),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _073_ (.A(N4END[14]),
    .X(net80),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _074_ (.A(N4END[13]),
    .X(net81),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _075_ (.A(N4END[12]),
    .X(net82),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _076_ (.A(N4END[11]),
    .X(net83),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _077_ (.A(N4END[10]),
    .X(net84),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _078_ (.A(N4END[9]),
    .X(net85),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _079_ (.A(N4END[8]),
    .X(net86),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _080_ (.A(N4END[7]),
    .X(net87),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _081_ (.A(N4END[6]),
    .X(net88),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _082_ (.A(N4END[5]),
    .X(net74),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _083_ (.A(N4END[4]),
    .X(net75),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _084_ (.A(N4END[3]),
    .X(net76),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _085_ (.A(N4END[2]),
    .X(net77),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _086_ (.A(N4END[1]),
    .X(net78),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _087_ (.A(N4END[0]),
    .X(net79),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _088_ (.A(NN4END[15]),
    .X(net89),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _089_ (.A(NN4END[14]),
    .X(net96),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _090_ (.A(NN4END[13]),
    .X(net97),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _091_ (.A(NN4END[12]),
    .X(net98),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _092_ (.A(NN4END[11]),
    .X(net99),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _093_ (.A(NN4END[10]),
    .X(net100),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _094_ (.A(NN4END[9]),
    .X(net101),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _095_ (.A(NN4END[8]),
    .X(net102),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _096_ (.A(NN4END[7]),
    .X(net103),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _097_ (.A(NN4END[6]),
    .X(net104),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _098_ (.A(NN4END[5]),
    .X(net90),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _099_ (.A(NN4END[4]),
    .X(net91),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _100_ (.A(NN4END[3]),
    .X(net92),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _101_ (.A(NN4END[2]),
    .X(net93),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _102_ (.A(NN4END[1]),
    .X(net94),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _103_ (.A(NN4END[0]),
    .X(net95),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _104_ (.A(UserCLK),
    .X(net105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output1 (.A(net1),
    .X(FrameData_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output2 (.A(net2),
    .X(FrameData_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output3 (.A(net3),
    .X(FrameData_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output4 (.A(net4),
    .X(FrameData_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output5 (.A(net5),
    .X(FrameData_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output6 (.A(net6),
    .X(FrameData_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output7 (.A(net7),
    .X(FrameData_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output8 (.A(net8),
    .X(FrameData_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output9 (.A(net9),
    .X(FrameData_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output10 (.A(net10),
    .X(FrameData_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output11 (.A(net11),
    .X(FrameData_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output12 (.A(net12),
    .X(FrameData_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output13 (.A(net13),
    .X(FrameData_O[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output14 (.A(net14),
    .X(FrameData_O[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output15 (.A(net15),
    .X(FrameData_O[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output16 (.A(net16),
    .X(FrameData_O[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net17),
    .X(FrameData_O[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net18),
    .X(FrameData_O[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net19),
    .X(FrameData_O[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net20),
    .X(FrameData_O[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net21),
    .X(FrameData_O[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net22),
    .X(FrameData_O[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output23 (.A(net23),
    .X(FrameData_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output24 (.A(net24),
    .X(FrameData_O[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output25 (.A(net25),
    .X(FrameData_O[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output26 (.A(net26),
    .X(FrameData_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output27 (.A(net27),
    .X(FrameData_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output28 (.A(net28),
    .X(FrameData_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output29 (.A(net29),
    .X(FrameData_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output30 (.A(net30),
    .X(FrameData_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output31 (.A(net31),
    .X(FrameData_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output32 (.A(net32),
    .X(FrameData_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output33 (.A(net33),
    .X(FrameStrobe_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output34 (.A(net34),
    .X(FrameStrobe_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output35 (.A(net35),
    .X(FrameStrobe_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output36 (.A(net36),
    .X(FrameStrobe_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output37 (.A(net37),
    .X(FrameStrobe_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output38 (.A(net38),
    .X(FrameStrobe_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output39 (.A(net39),
    .X(FrameStrobe_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output40 (.A(net40),
    .X(FrameStrobe_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output41 (.A(net41),
    .X(FrameStrobe_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output42 (.A(net42),
    .X(FrameStrobe_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output43 (.A(net43),
    .X(FrameStrobe_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output44 (.A(net44),
    .X(FrameStrobe_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output45 (.A(net45),
    .X(FrameStrobe_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output46 (.A(net46),
    .X(FrameStrobe_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output47 (.A(net47),
    .X(FrameStrobe_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output48 (.A(net48),
    .X(FrameStrobe_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output49 (.A(net49),
    .X(FrameStrobe_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output50 (.A(net50),
    .X(FrameStrobe_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output51 (.A(net51),
    .X(FrameStrobe_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output52 (.A(net52),
    .X(FrameStrobe_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output53 (.A(net53),
    .X(S1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output54 (.A(net54),
    .X(S1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output55 (.A(net55),
    .X(S1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output56 (.A(net56),
    .X(S1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output57 (.A(net57),
    .X(S2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output58 (.A(net58),
    .X(S2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output59 (.A(net59),
    .X(S2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output60 (.A(net60),
    .X(S2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output61 (.A(net61),
    .X(S2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output62 (.A(net62),
    .X(S2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output63 (.A(net63),
    .X(S2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output64 (.A(net64),
    .X(S2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output65 (.A(net65),
    .X(S2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output66 (.A(net66),
    .X(S2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output67 (.A(net67),
    .X(S2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output68 (.A(net68),
    .X(S2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output69 (.A(net69),
    .X(S2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output70 (.A(net70),
    .X(S2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output71 (.A(net71),
    .X(S2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output72 (.A(net72),
    .X(S2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output73 (.A(net73),
    .X(S4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output74 (.A(net74),
    .X(S4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output75 (.A(net75),
    .X(S4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output76 (.A(net76),
    .X(S4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output77 (.A(net77),
    .X(S4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output78 (.A(net78),
    .X(S4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output79 (.A(net79),
    .X(S4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output80 (.A(net80),
    .X(S4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output81 (.A(net81),
    .X(S4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output82 (.A(net82),
    .X(S4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output83 (.A(net83),
    .X(S4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output84 (.A(net84),
    .X(S4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output85 (.A(net85),
    .X(S4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output86 (.A(net86),
    .X(S4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output87 (.A(net87),
    .X(S4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output88 (.A(net88),
    .X(S4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output89 (.A(net89),
    .X(SS4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output90 (.A(net90),
    .X(SS4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output91 (.A(net91),
    .X(SS4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output92 (.A(net92),
    .X(SS4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output93 (.A(net93),
    .X(SS4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output94 (.A(net94),
    .X(SS4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output95 (.A(net95),
    .X(SS4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output96 (.A(net96),
    .X(SS4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output97 (.A(net97),
    .X(SS4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output98 (.A(net98),
    .X(SS4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output99 (.A(net99),
    .X(SS4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output100 (.A(net100),
    .X(SS4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output101 (.A(net101),
    .X(SS4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output102 (.A(net102),
    .X(SS4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output103 (.A(net103),
    .X(SS4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output104 (.A(net104),
    .X(SS4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output105 (.A(net105),
    .X(UserCLKo),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_antennanp ANTENNA_1 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_2 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[5]));
 sg13g2_antennanp ANTENNA_3 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_4 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[7]));
 sg13g2_antennanp ANTENNA_5 (.VDD(VPWR),
    .VSS(VGND),
    .A(net1));
 sg13g2_antennanp ANTENNA_6 (.VDD(VPWR),
    .VSS(VGND),
    .A(net27));
 sg13g2_antennanp ANTENNA_7 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameStrobe[3]));
 sg13g2_antennanp ANTENNA_8 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameStrobe[4]));
 sg13g2_antennanp ANTENNA_9 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_10 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[5]));
 sg13g2_antennanp ANTENNA_11 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_12 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[7]));
 sg13g2_antennanp ANTENNA_13 (.VDD(VPWR),
    .VSS(VGND),
    .A(net1));
 sg13g2_antennanp ANTENNA_14 (.VDD(VPWR),
    .VSS(VGND),
    .A(net22));
 sg13g2_antennanp ANTENNA_15 (.VDD(VPWR),
    .VSS(VGND),
    .A(net27));
 sg13g2_antennanp ANTENNA_16 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[5]));
 sg13g2_antennanp ANTENNA_17 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_18 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[7]));
 sg13g2_antennanp ANTENNA_19 (.VDD(VPWR),
    .VSS(VGND),
    .A(net1));
 sg13g2_antennanp ANTENNA_20 (.VDD(VPWR),
    .VSS(VGND),
    .A(net22));
 sg13g2_antennanp ANTENNA_21 (.VDD(VPWR),
    .VSS(VGND),
    .A(net27));
 sg13g2_antennanp ANTENNA_22 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[5]));
 sg13g2_antennanp ANTENNA_23 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_24 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[7]));
 sg13g2_antennanp ANTENNA_25 (.VDD(VPWR),
    .VSS(VGND),
    .A(net1));
 sg13g2_antennanp ANTENNA_26 (.VDD(VPWR),
    .VSS(VGND),
    .A(net27));
 sg13g2_antennanp ANTENNA_27 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[5]));
 sg13g2_antennanp ANTENNA_28 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_29 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[7]));
 sg13g2_antennanp ANTENNA_30 (.VDD(VPWR),
    .VSS(VGND),
    .A(net1));
 sg13g2_antennanp ANTENNA_31 (.VDD(VPWR),
    .VSS(VGND),
    .A(net27));
 sg13g2_antennanp ANTENNA_32 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[5]));
 sg13g2_antennanp ANTENNA_33 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_34 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[7]));
 sg13g2_antennanp ANTENNA_35 (.VDD(VPWR),
    .VSS(VGND),
    .A(net1));
 sg13g2_antennanp ANTENNA_36 (.VDD(VPWR),
    .VSS(VGND),
    .A(net27));
 sg13g2_antennanp ANTENNA_37 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[5]));
 sg13g2_antennanp ANTENNA_38 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_39 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[7]));
 sg13g2_antennanp ANTENNA_40 (.VDD(VPWR),
    .VSS(VGND),
    .A(net1));
 sg13g2_antennanp ANTENNA_41 (.VDD(VPWR),
    .VSS(VGND),
    .A(net27));
 sg13g2_antennanp ANTENNA_42 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[5]));
 sg13g2_antennanp ANTENNA_43 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_44 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[7]));
 sg13g2_antennanp ANTENNA_45 (.VDD(VPWR),
    .VSS(VGND),
    .A(net1));
 sg13g2_antennanp ANTENNA_46 (.VDD(VPWR),
    .VSS(VGND),
    .A(net27));
 sg13g2_antennanp ANTENNA_47 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[5]));
 sg13g2_antennanp ANTENNA_48 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_49 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[7]));
 sg13g2_antennanp ANTENNA_50 (.VDD(VPWR),
    .VSS(VGND),
    .A(net1));
 sg13g2_antennanp ANTENNA_51 (.VDD(VPWR),
    .VSS(VGND),
    .A(net27));
 sg13g2_antennanp ANTENNA_52 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[5]));
 sg13g2_antennanp ANTENNA_53 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_54 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[7]));
 sg13g2_antennanp ANTENNA_55 (.VDD(VPWR),
    .VSS(VGND),
    .A(net1));
 sg13g2_antennanp ANTENNA_56 (.VDD(VPWR),
    .VSS(VGND),
    .A(net27));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_503 (.VDD(VPWR),
    .VSS(VGND));
endmodule
