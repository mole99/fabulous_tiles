module E_IO (A_I_top,
    A_O_top,
    A_T_top,
    A_config_C_bit0,
    A_config_C_bit1,
    A_config_C_bit2,
    A_config_C_bit3,
    B_I_top,
    B_O_top,
    B_T_top,
    B_config_C_bit0,
    B_config_C_bit1,
    B_config_C_bit2,
    B_config_C_bit3,
    UserCLK,
    UserCLKo,
    E1END,
    E2END,
    E2MID,
    E6END,
    EE4END,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    W1BEG,
    W2BEG,
    W2BEGb,
    W6BEG,
    WW4BEG);
 output A_I_top;
 input A_O_top;
 output A_T_top;
 output A_config_C_bit0;
 output A_config_C_bit1;
 output A_config_C_bit2;
 output A_config_C_bit3;
 output B_I_top;
 input B_O_top;
 output B_T_top;
 output B_config_C_bit0;
 output B_config_C_bit1;
 output B_config_C_bit2;
 output B_config_C_bit3;
 input UserCLK;
 output UserCLKo;
 input [3:0] E1END;
 input [7:0] E2END;
 input [7:0] E2MID;
 input [11:0] E6END;
 input [15:0] EE4END;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] W1BEG;
 output [7:0] W2BEG;
 output [7:0] W2BEGb;
 output [11:0] W6BEG;
 output [15:0] WW4BEG;

 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire \Inst_A_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_B_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_E_IO_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_E_IO_switch_matrix.W1BEG0 ;
 wire \Inst_E_IO_switch_matrix.W1BEG1 ;
 wire \Inst_E_IO_switch_matrix.W1BEG2 ;
 wire \Inst_E_IO_switch_matrix.W1BEG3 ;
 wire \Inst_E_IO_switch_matrix.W2BEG0 ;
 wire \Inst_E_IO_switch_matrix.W2BEG1 ;
 wire \Inst_E_IO_switch_matrix.W2BEG2 ;
 wire \Inst_E_IO_switch_matrix.W2BEG3 ;
 wire \Inst_E_IO_switch_matrix.W2BEG4 ;
 wire \Inst_E_IO_switch_matrix.W2BEG5 ;
 wire \Inst_E_IO_switch_matrix.W2BEG6 ;
 wire \Inst_E_IO_switch_matrix.W2BEG7 ;
 wire \Inst_E_IO_switch_matrix.W2BEGb0 ;
 wire \Inst_E_IO_switch_matrix.W2BEGb1 ;
 wire \Inst_E_IO_switch_matrix.W2BEGb2 ;
 wire \Inst_E_IO_switch_matrix.W2BEGb3 ;
 wire \Inst_E_IO_switch_matrix.W2BEGb4 ;
 wire \Inst_E_IO_switch_matrix.W2BEGb5 ;
 wire \Inst_E_IO_switch_matrix.W2BEGb6 ;
 wire \Inst_E_IO_switch_matrix.W2BEGb7 ;
 wire \Inst_E_IO_switch_matrix.W6BEG0 ;
 wire \Inst_E_IO_switch_matrix.W6BEG1 ;
 wire \Inst_E_IO_switch_matrix.W6BEG10 ;
 wire \Inst_E_IO_switch_matrix.W6BEG11 ;
 wire \Inst_E_IO_switch_matrix.W6BEG2 ;
 wire \Inst_E_IO_switch_matrix.W6BEG3 ;
 wire \Inst_E_IO_switch_matrix.W6BEG4 ;
 wire \Inst_E_IO_switch_matrix.W6BEG5 ;
 wire \Inst_E_IO_switch_matrix.W6BEG6 ;
 wire \Inst_E_IO_switch_matrix.W6BEG7 ;
 wire \Inst_E_IO_switch_matrix.W6BEG8 ;
 wire \Inst_E_IO_switch_matrix.W6BEG9 ;
 wire \Inst_E_IO_switch_matrix.WW4BEG0 ;
 wire \Inst_E_IO_switch_matrix.WW4BEG1 ;
 wire \Inst_E_IO_switch_matrix.WW4BEG10 ;
 wire \Inst_E_IO_switch_matrix.WW4BEG11 ;
 wire \Inst_E_IO_switch_matrix.WW4BEG12 ;
 wire \Inst_E_IO_switch_matrix.WW4BEG13 ;
 wire \Inst_E_IO_switch_matrix.WW4BEG14 ;
 wire \Inst_E_IO_switch_matrix.WW4BEG15 ;
 wire \Inst_E_IO_switch_matrix.WW4BEG2 ;
 wire \Inst_E_IO_switch_matrix.WW4BEG3 ;
 wire \Inst_E_IO_switch_matrix.WW4BEG4 ;
 wire \Inst_E_IO_switch_matrix.WW4BEG5 ;
 wire \Inst_E_IO_switch_matrix.WW4BEG6 ;
 wire \Inst_E_IO_switch_matrix.WW4BEG7 ;
 wire \Inst_E_IO_switch_matrix.WW4BEG8 ;
 wire \Inst_E_IO_switch_matrix.WW4BEG9 ;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire net216;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net215;

 sg13g2_inv_1 _053_ (.Y(_000_),
    .A(\Inst_E_IO_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_inv_1 _054_ (.Y(_001_),
    .A(net7));
 sg13g2_inv_1 _055_ (.Y(_002_),
    .A(\Inst_E_IO_ConfigMem.Inst_frame0_bit20.Q ));
 sg13g2_inv_1 _056_ (.Y(_003_),
    .A(\Inst_E_IO_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_mux4_1 _057_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .A0(net7),
    .A1(net8),
    .A2(net9),
    .A3(net10),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_004_));
 sg13g2_nor2_1 _058_ (.A(\Inst_E_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .B(_004_),
    .Y(_005_));
 sg13g2_nor2_1 _059_ (.A(\Inst_E_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .B(net11),
    .Y(_006_));
 sg13g2_nor2b_1 _060_ (.A(net12),
    .B_N(\Inst_E_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .Y(_007_));
 sg13g2_nor3_1 _061_ (.A(\Inst_E_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .B(_006_),
    .C(_007_),
    .Y(_008_));
 sg13g2_mux2_1 _062_ (.A0(net13),
    .A1(net14),
    .S(\Inst_E_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .X(_009_));
 sg13g2_a21o_1 _063_ (.A2(_009_),
    .A1(\Inst_E_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .B1(_000_),
    .X(_010_));
 sg13g2_o21ai_1 _064_ (.B1(\Inst_E_IO_ConfigMem.Inst_frame0_bit28.Q ),
    .Y(_011_),
    .A1(_008_),
    .A2(_010_));
 sg13g2_mux2_1 _065_ (.A0(net17),
    .A1(net18),
    .S(\Inst_E_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .X(_012_));
 sg13g2_mux2_1 _066_ (.A0(net15),
    .A1(net16),
    .S(\Inst_E_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .X(_013_));
 sg13g2_mux2_1 _067_ (.A0(net21),
    .A1(net22),
    .S(\Inst_E_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .X(_014_));
 sg13g2_mux2_1 _068_ (.A0(net19),
    .A1(net20),
    .S(\Inst_E_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .X(_015_));
 sg13g2_mux4_1 _069_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .A0(_013_),
    .A1(_015_),
    .A2(_012_),
    .A3(_014_),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_016_));
 sg13g2_nand2b_1 _070_ (.Y(_017_),
    .B(_016_),
    .A_N(\Inst_E_IO_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_o21ai_1 _071_ (.B1(_017_),
    .Y(net108),
    .A1(_005_),
    .A2(_011_));
 sg13g2_mux4_1 _072_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .A0(net7),
    .A1(net8),
    .A2(net9),
    .A3(net10),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_018_));
 sg13g2_nor2_1 _073_ (.A(\Inst_E_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .B(_018_),
    .Y(_019_));
 sg13g2_nor2_1 _074_ (.A(net11),
    .B(\Inst_E_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .Y(_020_));
 sg13g2_nor2b_1 _075_ (.A(net12),
    .B_N(\Inst_E_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .Y(_021_));
 sg13g2_nor3_1 _076_ (.A(\Inst_E_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .B(_020_),
    .C(_021_),
    .Y(_022_));
 sg13g2_mux2_1 _077_ (.A0(net13),
    .A1(net14),
    .S(\Inst_E_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_023_));
 sg13g2_a21o_1 _078_ (.A2(_023_),
    .A1(\Inst_E_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .B1(_002_),
    .X(_024_));
 sg13g2_o21ai_1 _079_ (.B1(\Inst_E_IO_ConfigMem.Inst_frame0_bit21.Q ),
    .Y(_025_),
    .A1(_022_),
    .A2(_024_));
 sg13g2_mux2_1 _080_ (.A0(net17),
    .A1(net18),
    .S(\Inst_E_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_026_));
 sg13g2_mux2_1 _081_ (.A0(net15),
    .A1(net16),
    .S(\Inst_E_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_027_));
 sg13g2_mux2_1 _082_ (.A0(net21),
    .A1(net22),
    .S(\Inst_E_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_028_));
 sg13g2_mux2_1 _083_ (.A0(net19),
    .A1(net20),
    .S(\Inst_E_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_029_));
 sg13g2_mux4_1 _084_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .A0(_027_),
    .A1(_029_),
    .A2(_026_),
    .A3(_028_),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_030_));
 sg13g2_nand2b_1 _085_ (.Y(_031_),
    .B(_030_),
    .A_N(\Inst_E_IO_ConfigMem.Inst_frame0_bit21.Q ));
 sg13g2_o21ai_1 _086_ (.B1(_031_),
    .Y(net102),
    .A1(_019_),
    .A2(_025_));
 sg13g2_mux4_1 _087_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame0_bit16.Q ),
    .A0(net3),
    .A1(net35),
    .A2(net23),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame0_bit17.Q ),
    .X(\Inst_E_IO_switch_matrix.W6BEG11 ));
 sg13g2_mux4_1 _088_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame0_bit14.Q ),
    .A0(net4),
    .A1(net42),
    .A2(net26),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame0_bit15.Q ),
    .X(\Inst_E_IO_switch_matrix.W6BEG10 ));
 sg13g2_mux4_1 _089_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame0_bit12.Q ),
    .A0(net45),
    .A1(net38),
    .A2(net29),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame0_bit13.Q ),
    .X(\Inst_E_IO_switch_matrix.W6BEG9 ));
 sg13g2_mux4_1 _090_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame0_bit10.Q ),
    .A0(net46),
    .A1(net39),
    .A2(net30),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame0_bit11.Q ),
    .X(\Inst_E_IO_switch_matrix.W6BEG8 ));
 sg13g2_mux4_1 _091_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame0_bit8.Q ),
    .A0(net3),
    .A1(net49),
    .A2(net33),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame0_bit9.Q ),
    .X(\Inst_E_IO_switch_matrix.W6BEG7 ));
 sg13g2_mux4_1 _092_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame0_bit6.Q ),
    .A0(net4),
    .A1(net50),
    .A2(net34),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame0_bit7.Q ),
    .X(\Inst_E_IO_switch_matrix.W6BEG6 ));
 sg13g2_mux4_1 _093_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(net6),
    .A1(net43),
    .A2(net27),
    .A3(net2),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame0_bit5.Q ),
    .X(\Inst_E_IO_switch_matrix.W6BEG5 ));
 sg13g2_mux4_1 _094_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame0_bit2.Q ),
    .A0(net5),
    .A1(net44),
    .A2(net28),
    .A3(net1),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame0_bit3.Q ),
    .X(\Inst_E_IO_switch_matrix.W6BEG4 ));
 sg13g2_mux4_1 _095_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame0_bit0.Q ),
    .A0(net47),
    .A1(net40),
    .A2(net31),
    .A3(net2),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame0_bit1.Q ),
    .X(\Inst_E_IO_switch_matrix.W6BEG3 ));
 sg13g2_mux4_1 _096_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame1_bit30.Q ),
    .A0(net48),
    .A1(net41),
    .A2(net32),
    .A3(net1),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame1_bit31.Q ),
    .X(\Inst_E_IO_switch_matrix.W6BEG2 ));
 sg13g2_mux4_1 _097_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame1_bit28.Q ),
    .A0(net6),
    .A1(net36),
    .A2(net24),
    .A3(net2),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame1_bit29.Q ),
    .X(\Inst_E_IO_switch_matrix.W6BEG1 ));
 sg13g2_mux4_1 _098_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame1_bit26.Q ),
    .A0(net5),
    .A1(net37),
    .A2(net25),
    .A3(net1),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Inst_E_IO_switch_matrix.W6BEG0 ));
 sg13g2_mux4_1 _099_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame1_bit25.Q ),
    .A0(net16),
    .A1(net20),
    .A2(net18),
    .A3(net22),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame1_bit24.Q ),
    .X(\Inst_E_IO_switch_matrix.WW4BEG15 ));
 sg13g2_mux4_1 _100_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame1_bit23.Q ),
    .A0(net15),
    .A1(net19),
    .A2(net17),
    .A3(net21),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame1_bit22.Q ),
    .X(\Inst_E_IO_switch_matrix.WW4BEG14 ));
 sg13g2_mux4_1 _101_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame1_bit21.Q ),
    .A0(net32),
    .A1(net25),
    .A2(net34),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame1_bit20.Q ),
    .X(\Inst_E_IO_switch_matrix.WW4BEG13 ));
 sg13g2_mux4_1 _102_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame1_bit19.Q ),
    .A0(net26),
    .A1(net30),
    .A2(net28),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame1_bit18.Q ),
    .X(\Inst_E_IO_switch_matrix.WW4BEG12 ));
 sg13g2_mux4_1 _103_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame1_bit17.Q ),
    .A0(net31),
    .A1(net24),
    .A2(net33),
    .A3(net2),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame1_bit16.Q ),
    .X(\Inst_E_IO_switch_matrix.WW4BEG11 ));
 sg13g2_mux4_1 _104_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame1_bit15.Q ),
    .A0(net23),
    .A1(net29),
    .A2(net27),
    .A3(net1),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame1_bit14.Q ),
    .X(\Inst_E_IO_switch_matrix.WW4BEG10 ));
 sg13g2_mux4_1 _105_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame1_bit13.Q ),
    .A0(net26),
    .A1(net30),
    .A2(net28),
    .A3(net32),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame1_bit12.Q ),
    .X(\Inst_E_IO_switch_matrix.WW4BEG9 ));
 sg13g2_mux4_1 _106_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame1_bit11.Q ),
    .A0(net29),
    .A1(net33),
    .A2(net31),
    .A3(net24),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame1_bit10.Q ),
    .X(\Inst_E_IO_switch_matrix.WW4BEG8 ));
 sg13g2_mux4_1 _107_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame1_bit9.Q ),
    .A0(net16),
    .A1(net20),
    .A2(net18),
    .A3(net22),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame1_bit8.Q ),
    .X(\Inst_E_IO_switch_matrix.WW4BEG7 ));
 sg13g2_mux4_1 _108_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame1_bit7.Q ),
    .A0(net15),
    .A1(net19),
    .A2(net17),
    .A3(net21),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame1_bit6.Q ),
    .X(\Inst_E_IO_switch_matrix.WW4BEG6 ));
 sg13g2_mux4_1 _109_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame1_bit4.Q ),
    .A0(net8),
    .A1(net10),
    .A2(net12),
    .A3(net14),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame1_bit5.Q ),
    .X(\Inst_E_IO_switch_matrix.WW4BEG5 ));
 sg13g2_mux4_1 _110_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame1_bit2.Q ),
    .A0(net7),
    .A1(net9),
    .A2(net11),
    .A3(net13),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame1_bit3.Q ),
    .X(\Inst_E_IO_switch_matrix.WW4BEG4 ));
 sg13g2_mux4_1 _111_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame1_bit1.Q ),
    .A0(net32),
    .A1(net25),
    .A2(net34),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame1_bit0.Q ),
    .X(\Inst_E_IO_switch_matrix.WW4BEG3 ));
 sg13g2_mux4_1 _112_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame2_bit31.Q ),
    .A0(net26),
    .A1(net30),
    .A2(net28),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame2_bit30.Q ),
    .X(\Inst_E_IO_switch_matrix.WW4BEG2 ));
 sg13g2_mux4_1 _113_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame2_bit29.Q ),
    .A0(net31),
    .A1(net24),
    .A2(net33),
    .A3(net2),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame2_bit28.Q ),
    .X(\Inst_E_IO_switch_matrix.WW4BEG1 ));
 sg13g2_mux4_1 _114_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame2_bit27.Q ),
    .A0(net23),
    .A1(net29),
    .A2(net27),
    .A3(net1),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame2_bit26.Q ),
    .X(\Inst_E_IO_switch_matrix.WW4BEG0 ));
 sg13g2_mux4_1 _115_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame2_bit24.Q ),
    .A0(net7),
    .A1(net35),
    .A2(net49),
    .A3(net23),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame2_bit25.Q ),
    .X(\Inst_E_IO_switch_matrix.W2BEGb7 ));
 sg13g2_mux4_1 _116_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame2_bit22.Q ),
    .A0(net8),
    .A1(net42),
    .A2(net50),
    .A3(net26),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame2_bit23.Q ),
    .X(\Inst_E_IO_switch_matrix.W2BEGb6 ));
 sg13g2_mux4_1 _117_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame2_bit20.Q ),
    .A0(net9),
    .A1(net43),
    .A2(net36),
    .A3(net27),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame2_bit21.Q ),
    .X(\Inst_E_IO_switch_matrix.W2BEGb5 ));
 sg13g2_mux4_1 _118_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame2_bit18.Q ),
    .A0(net10),
    .A1(net44),
    .A2(net37),
    .A3(net28),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame2_bit19.Q ),
    .X(\Inst_E_IO_switch_matrix.W2BEGb4 ));
 sg13g2_mux4_1 _119_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame2_bit16.Q ),
    .A0(net11),
    .A1(net45),
    .A2(net38),
    .A3(net29),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame2_bit17.Q ),
    .X(\Inst_E_IO_switch_matrix.W2BEGb3 ));
 sg13g2_mux4_1 _120_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame2_bit14.Q ),
    .A0(net12),
    .A1(net46),
    .A2(net39),
    .A3(net30),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame2_bit15.Q ),
    .X(\Inst_E_IO_switch_matrix.W2BEGb2 ));
 sg13g2_mux4_1 _121_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame2_bit12.Q ),
    .A0(net13),
    .A1(net47),
    .A2(net40),
    .A3(net31),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame2_bit13.Q ),
    .X(\Inst_E_IO_switch_matrix.W2BEGb1 ));
 sg13g2_mux4_1 _122_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame2_bit10.Q ),
    .A0(net14),
    .A1(net48),
    .A2(net41),
    .A3(net32),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame2_bit11.Q ),
    .X(\Inst_E_IO_switch_matrix.W2BEGb0 ));
 sg13g2_mux4_1 _123_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame2_bit8.Q ),
    .A0(net15),
    .A1(net35),
    .A2(net49),
    .A3(net23),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame2_bit9.Q ),
    .X(\Inst_E_IO_switch_matrix.W2BEG7 ));
 sg13g2_mux4_1 _124_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame2_bit6.Q ),
    .A0(net16),
    .A1(net42),
    .A2(net50),
    .A3(net26),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame2_bit7.Q ),
    .X(\Inst_E_IO_switch_matrix.W2BEG6 ));
 sg13g2_mux4_1 _125_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame2_bit4.Q ),
    .A0(net17),
    .A1(net43),
    .A2(net36),
    .A3(net27),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame2_bit5.Q ),
    .X(\Inst_E_IO_switch_matrix.W2BEG5 ));
 sg13g2_mux4_1 _126_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame2_bit2.Q ),
    .A0(net18),
    .A1(net44),
    .A2(net37),
    .A3(net28),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame2_bit3.Q ),
    .X(\Inst_E_IO_switch_matrix.W2BEG4 ));
 sg13g2_mux4_1 _127_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame2_bit0.Q ),
    .A0(net19),
    .A1(net45),
    .A2(net38),
    .A3(net29),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame2_bit1.Q ),
    .X(\Inst_E_IO_switch_matrix.W2BEG3 ));
 sg13g2_mux4_1 _128_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame3_bit30.Q ),
    .A0(net20),
    .A1(net46),
    .A2(net39),
    .A3(net30),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame3_bit31.Q ),
    .X(\Inst_E_IO_switch_matrix.W2BEG2 ));
 sg13g2_mux4_1 _129_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame3_bit28.Q ),
    .A0(net21),
    .A1(net47),
    .A2(net40),
    .A3(net31),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame3_bit29.Q ),
    .X(\Inst_E_IO_switch_matrix.W2BEG1 ));
 sg13g2_mux4_1 _130_ (.S0(\Inst_E_IO_ConfigMem.Inst_frame3_bit26.Q ),
    .A0(net22),
    .A1(net48),
    .A2(net41),
    .A3(net32),
    .S1(\Inst_E_IO_ConfigMem.Inst_frame3_bit27.Q ),
    .X(\Inst_E_IO_switch_matrix.W2BEG0 ));
 sg13g2_mux2_1 _131_ (.A0(net3),
    .A1(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S(\Inst_E_IO_ConfigMem.Inst_frame3_bit25.Q ),
    .X(\Inst_E_IO_switch_matrix.W1BEG3 ));
 sg13g2_mux2_1 _132_ (.A0(net4),
    .A1(net2),
    .S(\Inst_E_IO_ConfigMem.Inst_frame3_bit24.Q ),
    .X(\Inst_E_IO_switch_matrix.W1BEG2 ));
 sg13g2_mux2_1 _133_ (.A0(net5),
    .A1(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S(\Inst_E_IO_ConfigMem.Inst_frame3_bit23.Q ),
    .X(\Inst_E_IO_switch_matrix.W1BEG1 ));
 sg13g2_mux2_1 _134_ (.A0(net6),
    .A1(net1),
    .S(\Inst_E_IO_ConfigMem.Inst_frame3_bit22.Q ),
    .X(\Inst_E_IO_switch_matrix.W1BEG0 ));
 sg13g2_nand2b_1 _135_ (.Y(_032_),
    .B(\Inst_E_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .A_N(net8));
 sg13g2_o21ai_1 _136_ (.B1(_032_),
    .Y(_033_),
    .A1(net22),
    .A2(\Inst_E_IO_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_nor2b_1 _137_ (.A(\Inst_E_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .B_N(net10),
    .Y(_034_));
 sg13g2_a21oi_1 _138_ (.A1(\Inst_E_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .A2(_034_),
    .Y(_035_),
    .B1(\Inst_E_IO_ConfigMem.Inst_frame0_bit22.Q ));
 sg13g2_o21ai_1 _139_ (.B1(_035_),
    .Y(_036_),
    .A1(\Inst_E_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .A2(_033_));
 sg13g2_nor3_1 _140_ (.A(_001_),
    .B(\Inst_E_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .C(\Inst_E_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .Y(_037_));
 sg13g2_o21ai_1 _141_ (.B1(\Inst_E_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .Y(_038_),
    .A1(net9),
    .A2(\Inst_E_IO_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_nand2_1 _142_ (.Y(_039_),
    .A(net11),
    .B(\Inst_E_IO_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_nand3_1 _143_ (.B(_038_),
    .C(_039_),
    .A(\Inst_E_IO_ConfigMem.Inst_frame0_bit22.Q ),
    .Y(_040_));
 sg13g2_o21ai_1 _144_ (.B1(_036_),
    .Y(net103),
    .A1(_037_),
    .A2(_040_));
 sg13g2_nor2_1 _145_ (.A(net21),
    .B(\Inst_E_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .Y(_041_));
 sg13g2_a21oi_1 _146_ (.A1(_001_),
    .A2(\Inst_E_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .Y(_042_),
    .B1(_041_));
 sg13g2_nor2_1 _147_ (.A(\Inst_E_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .B(_003_),
    .Y(_043_));
 sg13g2_a221oi_1 _148_ (.B2(net12),
    .C1(\Inst_E_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .B1(_043_),
    .A1(_003_),
    .Y(_044_),
    .A2(_042_));
 sg13g2_nor2b_1 _149_ (.A(\Inst_E_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .B_N(net22),
    .Y(_045_));
 sg13g2_a22oi_1 _150_ (.Y(_046_),
    .B1(_003_),
    .B2(_045_),
    .A2(\Inst_E_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .A1(net11));
 sg13g2_o21ai_1 _151_ (.B1(\Inst_E_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_047_),
    .A1(net13),
    .A2(\Inst_E_IO_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_nand3_1 _152_ (.B(_046_),
    .C(_047_),
    .A(\Inst_E_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_048_));
 sg13g2_nand2b_2 _153_ (.Y(net109),
    .B(_048_),
    .A_N(_044_));
 sg13g2_dlhq_1 _154_ (.D(net56),
    .GATE(net59),
    .Q(net104));
 sg13g2_dlhq_1 _155_ (.D(net57),
    .GATE(net59),
    .Q(net105));
 sg13g2_dlhq_1 _156_ (.D(net58),
    .GATE(net60),
    .Q(net106));
 sg13g2_dlhq_1 _157_ (.D(net78),
    .GATE(net60),
    .Q(net107));
 sg13g2_dlhq_1 _158_ (.D(net79),
    .GATE(net60),
    .Q(net110));
 sg13g2_dlhq_1 _159_ (.D(net80),
    .GATE(net59),
    .Q(net111));
 sg13g2_dlhq_1 _160_ (.D(net82),
    .GATE(net59),
    .Q(net112));
 sg13g2_dlhq_1 _161_ (.D(net83),
    .GATE(net60),
    .Q(net113));
 sg13g2_dlhq_1 _162_ (.D(net84),
    .GATE(net59),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_dlhq_1 _163_ (.D(net85),
    .GATE(net59),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame3_bit23.Q ));
 sg13g2_dlhq_1 _164_ (.D(net86),
    .GATE(net59),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame3_bit24.Q ));
 sg13g2_dlhq_1 _165_ (.D(net87),
    .GATE(net59),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_dlhq_1 _166_ (.D(net88),
    .GATE(net61),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_dlhq_1 _167_ (.D(net89),
    .GATE(net61),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_dlhq_1 _168_ (.D(net90),
    .GATE(net61),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame3_bit28.Q ));
 sg13g2_dlhq_1 _169_ (.D(net91),
    .GATE(net61),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame3_bit29.Q ));
 sg13g2_dlhq_1 _170_ (.D(net93),
    .GATE(net61),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame3_bit30.Q ));
 sg13g2_dlhq_1 _171_ (.D(net94),
    .GATE(net61),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame3_bit31.Q ));
 sg13g2_dlhq_1 _172_ (.D(net51),
    .GATE(net63),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit0.Q ));
 sg13g2_dlhq_1 _173_ (.D(net81),
    .GATE(net63),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit1.Q ));
 sg13g2_dlhq_1 _174_ (.D(net92),
    .GATE(net63),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_dlhq_1 _175_ (.D(net95),
    .GATE(net63),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit3.Q ));
 sg13g2_dlhq_1 _176_ (.D(net96),
    .GATE(net63),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit4.Q ));
 sg13g2_dlhq_1 _177_ (.D(net97),
    .GATE(net63),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_dlhq_1 _178_ (.D(net98),
    .GATE(net62),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_dlhq_1 _179_ (.D(net99),
    .GATE(net62),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_dlhq_1 _180_ (.D(net100),
    .GATE(net62),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit8.Q ));
 sg13g2_dlhq_1 _181_ (.D(net101),
    .GATE(net62),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit9.Q ));
 sg13g2_dlhq_1 _182_ (.D(net52),
    .GATE(net65),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_dlhq_1 _183_ (.D(net53),
    .GATE(net65),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit11.Q ));
 sg13g2_dlhq_1 _184_ (.D(net54),
    .GATE(net65),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_dlhq_1 _185_ (.D(net55),
    .GATE(net65),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_dlhq_1 _186_ (.D(net56),
    .GATE(net65),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_dlhq_1 _187_ (.D(net57),
    .GATE(net65),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_dlhq_1 _188_ (.D(net58),
    .GATE(net63),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_dlhq_1 _189_ (.D(net78),
    .GATE(net63),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit17.Q ));
 sg13g2_dlhq_1 _190_ (.D(net79),
    .GATE(net64),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_dlhq_1 _191_ (.D(net80),
    .GATE(net64),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_dlhq_1 _192_ (.D(net82),
    .GATE(net64),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit20.Q ));
 sg13g2_dlhq_1 _193_ (.D(net83),
    .GATE(net64),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit21.Q ));
 sg13g2_dlhq_1 _194_ (.D(net84),
    .GATE(net62),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_dlhq_1 _195_ (.D(net85),
    .GATE(net62),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit23.Q ));
 sg13g2_dlhq_1 _196_ (.D(net86),
    .GATE(net62),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit24.Q ));
 sg13g2_dlhq_1 _197_ (.D(net87),
    .GATE(net62),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_dlhq_1 _198_ (.D(net88),
    .GATE(net65),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_dlhq_1 _199_ (.D(net89),
    .GATE(net65),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_dlhq_1 _200_ (.D(net90),
    .GATE(net66),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_dlhq_1 _201_ (.D(net91),
    .GATE(net66),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_dlhq_1 _202_ (.D(net93),
    .GATE(net66),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_dlhq_1 _203_ (.D(net94),
    .GATE(net66),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_dlhq_1 _204_ (.D(net51),
    .GATE(net71),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_dlhq_1 _205_ (.D(net81),
    .GATE(net71),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_dlhq_1 _206_ (.D(net92),
    .GATE(net68),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_dlhq_1 _207_ (.D(net95),
    .GATE(net68),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_dlhq_1 _208_ (.D(net96),
    .GATE(net67),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_dlhq_1 _209_ (.D(net97),
    .GATE(net67),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_dlhq_1 _210_ (.D(net98),
    .GATE(net68),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_dlhq_1 _211_ (.D(net99),
    .GATE(net68),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_dlhq_1 _212_ (.D(net100),
    .GATE(net67),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit8.Q ));
 sg13g2_dlhq_1 _213_ (.D(net101),
    .GATE(net67),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit9.Q ));
 sg13g2_dlhq_1 _214_ (.D(net52),
    .GATE(net69),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_dlhq_1 _215_ (.D(net53),
    .GATE(net69),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_dlhq_1 _216_ (.D(net54),
    .GATE(net69),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit12.Q ));
 sg13g2_dlhq_1 _217_ (.D(net55),
    .GATE(net69),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit13.Q ));
 sg13g2_dlhq_1 _218_ (.D(net56),
    .GATE(net67),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit14.Q ));
 sg13g2_dlhq_1 _219_ (.D(net57),
    .GATE(net67),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit15.Q ));
 sg13g2_dlhq_1 _220_ (.D(net58),
    .GATE(net70),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit16.Q ));
 sg13g2_dlhq_1 _221_ (.D(net78),
    .GATE(net70),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit17.Q ));
 sg13g2_dlhq_1 _222_ (.D(net79),
    .GATE(net69),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_dlhq_1 _223_ (.D(net80),
    .GATE(net69),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit19.Q ));
 sg13g2_dlhq_1 _224_ (.D(net82),
    .GATE(net69),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_dlhq_1 _225_ (.D(net83),
    .GATE(net69),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit21.Q ));
 sg13g2_dlhq_1 _226_ (.D(net84),
    .GATE(net68),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_dlhq_1 _227_ (.D(net85),
    .GATE(net68),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit23.Q ));
 sg13g2_dlhq_1 _228_ (.D(net86),
    .GATE(net67),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit24.Q ));
 sg13g2_dlhq_1 _229_ (.D(net87),
    .GATE(net67),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_dlhq_1 _230_ (.D(net88),
    .GATE(net71),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_dlhq_1 _231_ (.D(net89),
    .GATE(net71),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit27.Q ));
 sg13g2_dlhq_1 _232_ (.D(net90),
    .GATE(net70),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit28.Q ));
 sg13g2_dlhq_1 _233_ (.D(net91),
    .GATE(net70),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit29.Q ));
 sg13g2_dlhq_1 _234_ (.D(net93),
    .GATE(net71),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit30.Q ));
 sg13g2_dlhq_1 _235_ (.D(net94),
    .GATE(net71),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame1_bit31.Q ));
 sg13g2_dlhq_1 _236_ (.D(net51),
    .GATE(net76),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit0.Q ));
 sg13g2_dlhq_1 _237_ (.D(net81),
    .GATE(net76),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit1.Q ));
 sg13g2_dlhq_1 _238_ (.D(net92),
    .GATE(net74),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_dlhq_1 _239_ (.D(net95),
    .GATE(net74),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit3.Q ));
 sg13g2_dlhq_1 _240_ (.D(net96),
    .GATE(net73),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_dlhq_1 _241_ (.D(net97),
    .GATE(net73),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit5.Q ));
 sg13g2_dlhq_1 _242_ (.D(net98),
    .GATE(net72),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit6.Q ));
 sg13g2_dlhq_1 _243_ (.D(net99),
    .GATE(net72),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit7.Q ));
 sg13g2_dlhq_1 _244_ (.D(net100),
    .GATE(net72),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_dlhq_1 _245_ (.D(net101),
    .GATE(net72),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit9.Q ));
 sg13g2_dlhq_1 _246_ (.D(net52),
    .GATE(net75),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit10.Q ));
 sg13g2_dlhq_1 _247_ (.D(net53),
    .GATE(net75),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit11.Q ));
 sg13g2_dlhq_1 _248_ (.D(net54),
    .GATE(net75),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit12.Q ));
 sg13g2_dlhq_1 _249_ (.D(net55),
    .GATE(net75),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit13.Q ));
 sg13g2_dlhq_1 _250_ (.D(net56),
    .GATE(net72),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit14.Q ));
 sg13g2_dlhq_1 _251_ (.D(net57),
    .GATE(net72),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit15.Q ));
 sg13g2_dlhq_1 _252_ (.D(net58),
    .GATE(net72),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit16.Q ));
 sg13g2_dlhq_1 _253_ (.D(net78),
    .GATE(net72),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit17.Q ));
 sg13g2_dlhq_1 _254_ (.D(net79),
    .GATE(net73),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_dlhq_1 _255_ (.D(net80),
    .GATE(net73),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_dlhq_1 _256_ (.D(net82),
    .GATE(net73),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit20.Q ));
 sg13g2_dlhq_1 _257_ (.D(net83),
    .GATE(net73),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit21.Q ));
 sg13g2_dlhq_1 _258_ (.D(net84),
    .GATE(net74),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit22.Q ));
 sg13g2_dlhq_1 _259_ (.D(net85),
    .GATE(net73),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_dlhq_1 _260_ (.D(net86),
    .GATE(net73),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_dlhq_1 _261_ (.D(net87),
    .GATE(net76),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_dlhq_1 _262_ (.D(net88),
    .GATE(net75),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_dlhq_1 _263_ (.D(net89),
    .GATE(net75),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_dlhq_1 _264_ (.D(net90),
    .GATE(net77),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_dlhq_1 _265_ (.D(net91),
    .GATE(net77),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_dlhq_1 _266_ (.D(net93),
    .GATE(net75),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_dlhq_1 _267_ (.D(net94),
    .GATE(net75),
    .Q(\Inst_E_IO_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_dfrbp_1 _268_ (.CLK(UserCLK),
    .RESET_B(net215),
    .D(net1),
    .Q_N(_050_),
    .Q(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ));
 sg13g2_dfrbp_1 _269_ (.CLK(UserCLK),
    .RESET_B(net216),
    .D(net2),
    .Q_N(_049_),
    .Q(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ));
 sg13g2_tiehi _269__197 (.L_HI(net216));
 sg13g2_antennanp ANTENNA_1 (.A(net129));
 sg13g2_buf_1 _272_ (.A(net92),
    .X(net136));
 sg13g2_buf_1 _273_ (.A(net95),
    .X(net139));
 sg13g2_buf_1 _274_ (.A(net96),
    .X(net140));
 sg13g2_buf_1 _275_ (.A(net97),
    .X(net141));
 sg13g2_buf_2 _276_ (.A(net98),
    .X(net142));
 sg13g2_buf_2 _277_ (.A(net99),
    .X(net143));
 sg13g2_buf_1 _278_ (.A(net100),
    .X(net144));
 sg13g2_buf_2 _279_ (.A(net101),
    .X(net145));
 sg13g2_buf_1 _280_ (.A(net52),
    .X(net115));
 sg13g2_buf_1 _281_ (.A(net53),
    .X(net116));
 sg13g2_buf_1 _282_ (.A(net54),
    .X(net117));
 sg13g2_buf_1 _283_ (.A(net55),
    .X(net118));
 sg13g2_buf_2 _284_ (.A(net56),
    .X(net119));
 sg13g2_buf_2 _285_ (.A(net57),
    .X(net120));
 sg13g2_buf_1 _286_ (.A(net58),
    .X(net121));
 sg13g2_buf_1 _287_ (.A(net78),
    .X(net122));
 sg13g2_buf_1 _288_ (.A(net79),
    .X(net123));
 sg13g2_buf_2 _289_ (.A(net80),
    .X(net124));
 sg13g2_buf_2 _290_ (.A(net82),
    .X(net126));
 sg13g2_buf_1 _291_ (.A(net83),
    .X(net127));
 sg13g2_buf_2 _292_ (.A(net84),
    .X(net128));
 sg13g2_buf_2 _293_ (.A(net85),
    .X(net129));
 sg13g2_buf_2 _294_ (.A(net86),
    .X(net130));
 sg13g2_buf_2 _295_ (.A(net87),
    .X(net131));
 sg13g2_buf_2 _296_ (.A(net88),
    .X(net132));
 sg13g2_buf_2 _297_ (.A(net89),
    .X(net133));
 sg13g2_buf_1 _298_ (.A(net90),
    .X(net134));
 sg13g2_buf_1 _299_ (.A(net91),
    .X(net135));
 sg13g2_buf_2 _300_ (.A(net93),
    .X(net137));
 sg13g2_buf_2 _301_ (.A(net94),
    .X(net138));
 sg13g2_buf_1 _302_ (.A(net77),
    .X(net146));
 sg13g2_buf_1 _303_ (.A(net70),
    .X(net157));
 sg13g2_buf_1 _304_ (.A(net66),
    .X(net158));
 sg13g2_buf_1 _305_ (.A(net61),
    .X(net159));
 sg13g2_buf_1 _306_ (.A(FrameStrobe[4]),
    .X(net160));
 sg13g2_buf_1 _307_ (.A(FrameStrobe[5]),
    .X(net161));
 sg13g2_buf_1 _308_ (.A(FrameStrobe[6]),
    .X(net162));
 sg13g2_buf_1 _309_ (.A(FrameStrobe[7]),
    .X(net163));
 sg13g2_buf_1 _310_ (.A(FrameStrobe[8]),
    .X(net164));
 sg13g2_buf_1 _311_ (.A(FrameStrobe[9]),
    .X(net165));
 sg13g2_buf_1 _312_ (.A(FrameStrobe[10]),
    .X(net147));
 sg13g2_buf_1 _313_ (.A(FrameStrobe[11]),
    .X(net148));
 sg13g2_buf_1 _314_ (.A(FrameStrobe[12]),
    .X(net149));
 sg13g2_buf_1 _315_ (.A(FrameStrobe[13]),
    .X(net150));
 sg13g2_buf_1 _316_ (.A(FrameStrobe[14]),
    .X(net151));
 sg13g2_buf_1 _317_ (.A(FrameStrobe[15]),
    .X(net152));
 sg13g2_buf_1 _318_ (.A(FrameStrobe[16]),
    .X(net153));
 sg13g2_buf_1 _319_ (.A(FrameStrobe[17]),
    .X(net154));
 sg13g2_buf_1 _320_ (.A(FrameStrobe[18]),
    .X(net155));
 sg13g2_buf_1 _321_ (.A(FrameStrobe[19]),
    .X(net156));
 sg13g2_buf_1 _322_ (.A(UserCLK),
    .X(net166));
 sg13g2_buf_1 _323_ (.A(\Inst_E_IO_switch_matrix.W1BEG0 ),
    .X(net167));
 sg13g2_buf_1 _324_ (.A(\Inst_E_IO_switch_matrix.W1BEG1 ),
    .X(net168));
 sg13g2_buf_1 _325_ (.A(\Inst_E_IO_switch_matrix.W1BEG2 ),
    .X(net169));
 sg13g2_buf_1 _326_ (.A(\Inst_E_IO_switch_matrix.W1BEG3 ),
    .X(net170));
 sg13g2_buf_2 _327_ (.A(\Inst_E_IO_switch_matrix.W2BEG0 ),
    .X(net171));
 sg13g2_buf_2 _328_ (.A(\Inst_E_IO_switch_matrix.W2BEG1 ),
    .X(net172));
 sg13g2_buf_2 _329_ (.A(\Inst_E_IO_switch_matrix.W2BEG2 ),
    .X(net173));
 sg13g2_buf_2 _330_ (.A(\Inst_E_IO_switch_matrix.W2BEG3 ),
    .X(net174));
 sg13g2_buf_1 _331_ (.A(\Inst_E_IO_switch_matrix.W2BEG4 ),
    .X(net175));
 sg13g2_buf_2 _332_ (.A(\Inst_E_IO_switch_matrix.W2BEG5 ),
    .X(net176));
 sg13g2_buf_1 _333_ (.A(\Inst_E_IO_switch_matrix.W2BEG6 ),
    .X(net177));
 sg13g2_buf_1 _334_ (.A(\Inst_E_IO_switch_matrix.W2BEG7 ),
    .X(net178));
 sg13g2_buf_2 _335_ (.A(\Inst_E_IO_switch_matrix.W2BEGb0 ),
    .X(net179));
 sg13g2_buf_2 _336_ (.A(\Inst_E_IO_switch_matrix.W2BEGb1 ),
    .X(net180));
 sg13g2_buf_2 _337_ (.A(\Inst_E_IO_switch_matrix.W2BEGb2 ),
    .X(net181));
 sg13g2_buf_2 _338_ (.A(\Inst_E_IO_switch_matrix.W2BEGb3 ),
    .X(net182));
 sg13g2_buf_2 _339_ (.A(\Inst_E_IO_switch_matrix.W2BEGb4 ),
    .X(net183));
 sg13g2_buf_1 _340_ (.A(\Inst_E_IO_switch_matrix.W2BEGb5 ),
    .X(net184));
 sg13g2_buf_1 _341_ (.A(\Inst_E_IO_switch_matrix.W2BEGb6 ),
    .X(net185));
 sg13g2_buf_1 _342_ (.A(\Inst_E_IO_switch_matrix.W2BEGb7 ),
    .X(net186));
 sg13g2_buf_2 _343_ (.A(\Inst_E_IO_switch_matrix.W6BEG0 ),
    .X(net187));
 sg13g2_buf_2 _344_ (.A(\Inst_E_IO_switch_matrix.W6BEG1 ),
    .X(net190));
 sg13g2_buf_2 _345_ (.A(\Inst_E_IO_switch_matrix.W6BEG2 ),
    .X(net191));
 sg13g2_buf_2 _346_ (.A(\Inst_E_IO_switch_matrix.W6BEG3 ),
    .X(net192));
 sg13g2_buf_1 _347_ (.A(\Inst_E_IO_switch_matrix.W6BEG4 ),
    .X(net193));
 sg13g2_buf_1 _348_ (.A(\Inst_E_IO_switch_matrix.W6BEG5 ),
    .X(net194));
 sg13g2_buf_1 _349_ (.A(\Inst_E_IO_switch_matrix.W6BEG6 ),
    .X(net195));
 sg13g2_buf_1 _350_ (.A(\Inst_E_IO_switch_matrix.W6BEG7 ),
    .X(net196));
 sg13g2_buf_2 _351_ (.A(\Inst_E_IO_switch_matrix.W6BEG8 ),
    .X(net197));
 sg13g2_buf_2 _352_ (.A(\Inst_E_IO_switch_matrix.W6BEG9 ),
    .X(net198));
 sg13g2_buf_1 _353_ (.A(\Inst_E_IO_switch_matrix.W6BEG10 ),
    .X(net188));
 sg13g2_buf_1 _354_ (.A(\Inst_E_IO_switch_matrix.W6BEG11 ),
    .X(net189));
 sg13g2_buf_2 _355_ (.A(\Inst_E_IO_switch_matrix.WW4BEG0 ),
    .X(net199));
 sg13g2_buf_2 _356_ (.A(\Inst_E_IO_switch_matrix.WW4BEG1 ),
    .X(net206));
 sg13g2_buf_2 _357_ (.A(\Inst_E_IO_switch_matrix.WW4BEG2 ),
    .X(net207));
 sg13g2_buf_2 _358_ (.A(\Inst_E_IO_switch_matrix.WW4BEG3 ),
    .X(net208));
 sg13g2_buf_1 _359_ (.A(\Inst_E_IO_switch_matrix.WW4BEG4 ),
    .X(net209));
 sg13g2_buf_1 _360_ (.A(\Inst_E_IO_switch_matrix.WW4BEG5 ),
    .X(net210));
 sg13g2_buf_1 _361_ (.A(\Inst_E_IO_switch_matrix.WW4BEG6 ),
    .X(net211));
 sg13g2_buf_1 _362_ (.A(\Inst_E_IO_switch_matrix.WW4BEG7 ),
    .X(net212));
 sg13g2_buf_2 _363_ (.A(\Inst_E_IO_switch_matrix.WW4BEG8 ),
    .X(net213));
 sg13g2_buf_2 _364_ (.A(\Inst_E_IO_switch_matrix.WW4BEG9 ),
    .X(net214));
 sg13g2_buf_2 _365_ (.A(\Inst_E_IO_switch_matrix.WW4BEG10 ),
    .X(net200));
 sg13g2_buf_2 _366_ (.A(\Inst_E_IO_switch_matrix.WW4BEG11 ),
    .X(net201));
 sg13g2_buf_2 _367_ (.A(\Inst_E_IO_switch_matrix.WW4BEG12 ),
    .X(net202));
 sg13g2_buf_2 _368_ (.A(\Inst_E_IO_switch_matrix.WW4BEG13 ),
    .X(net203));
 sg13g2_buf_1 _369_ (.A(\Inst_E_IO_switch_matrix.WW4BEG14 ),
    .X(net204));
 sg13g2_buf_1 _370_ (.A(\Inst_E_IO_switch_matrix.WW4BEG15 ),
    .X(net205));
 sg13g2_buf_2 _371_ (.A(net51),
    .X(net114));
 sg13g2_buf_2 _372_ (.A(net81),
    .X(net125));
 sg13g2_buf_2 fanout59 (.A(net60),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(net61),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(FrameStrobe[3]),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(net64),
    .X(net62));
 sg13g2_buf_4 fanout63 (.X(net63),
    .A(net64));
 sg13g2_buf_2 fanout64 (.A(FrameStrobe[2]),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(FrameStrobe[2]),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(FrameStrobe[2]),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(FrameStrobe[1]),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(FrameStrobe[1]),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(net71),
    .X(net69));
 sg13g2_buf_1 fanout70 (.A(net71),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(FrameStrobe[1]),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(net74),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(net74),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(FrameStrobe[0]),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(net76),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(net77),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(FrameStrobe[0]),
    .X(net77));
 sg13g2_buf_4 input1 (.X(net1),
    .A(A_O_top));
 sg13g2_buf_4 input2 (.X(net2),
    .A(B_O_top));
 sg13g2_buf_1 input3 (.A(E1END[0]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(E1END[1]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(E1END[2]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(E1END[3]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(E2END[0]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(E2END[1]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(E2END[2]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(E2END[3]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(E2END[4]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(E2END[5]),
    .X(net12));
 sg13g2_buf_2 input13 (.A(E2END[6]),
    .X(net13));
 sg13g2_buf_2 input14 (.A(E2END[7]),
    .X(net14));
 sg13g2_buf_2 input15 (.A(E2MID[0]),
    .X(net15));
 sg13g2_buf_2 input16 (.A(E2MID[1]),
    .X(net16));
 sg13g2_buf_2 input17 (.A(E2MID[2]),
    .X(net17));
 sg13g2_buf_2 input18 (.A(E2MID[3]),
    .X(net18));
 sg13g2_buf_2 input19 (.A(E2MID[4]),
    .X(net19));
 sg13g2_buf_2 input20 (.A(E2MID[5]),
    .X(net20));
 sg13g2_buf_2 input21 (.A(E2MID[6]),
    .X(net21));
 sg13g2_buf_2 input22 (.A(E2MID[7]),
    .X(net22));
 sg13g2_buf_2 input23 (.A(E6END[0]),
    .X(net23));
 sg13g2_buf_1 input24 (.A(E6END[10]),
    .X(net24));
 sg13g2_buf_1 input25 (.A(E6END[11]),
    .X(net25));
 sg13g2_buf_4 input26 (.X(net26),
    .A(E6END[1]));
 sg13g2_buf_2 input27 (.A(E6END[2]),
    .X(net27));
 sg13g2_buf_2 input28 (.A(E6END[3]),
    .X(net28));
 sg13g2_buf_2 input29 (.A(E6END[4]),
    .X(net29));
 sg13g2_buf_2 input30 (.A(E6END[5]),
    .X(net30));
 sg13g2_buf_2 input31 (.A(E6END[6]),
    .X(net31));
 sg13g2_buf_2 input32 (.A(E6END[7]),
    .X(net32));
 sg13g2_buf_4 input33 (.X(net33),
    .A(E6END[8]));
 sg13g2_buf_2 input34 (.A(E6END[9]),
    .X(net34));
 sg13g2_buf_2 input35 (.A(EE4END[0]),
    .X(net35));
 sg13g2_buf_2 input36 (.A(EE4END[10]),
    .X(net36));
 sg13g2_buf_2 input37 (.A(EE4END[11]),
    .X(net37));
 sg13g2_buf_1 input38 (.A(EE4END[12]),
    .X(net38));
 sg13g2_buf_1 input39 (.A(EE4END[13]),
    .X(net39));
 sg13g2_buf_1 input40 (.A(EE4END[14]),
    .X(net40));
 sg13g2_buf_1 input41 (.A(EE4END[15]),
    .X(net41));
 sg13g2_buf_2 input42 (.A(EE4END[1]),
    .X(net42));
 sg13g2_buf_1 input43 (.A(EE4END[2]),
    .X(net43));
 sg13g2_buf_2 input44 (.A(EE4END[3]),
    .X(net44));
 sg13g2_buf_1 input45 (.A(EE4END[4]),
    .X(net45));
 sg13g2_buf_1 input46 (.A(EE4END[5]),
    .X(net46));
 sg13g2_buf_2 input47 (.A(EE4END[6]),
    .X(net47));
 sg13g2_buf_1 input48 (.A(EE4END[7]),
    .X(net48));
 sg13g2_buf_2 input49 (.A(EE4END[8]),
    .X(net49));
 sg13g2_buf_2 input50 (.A(EE4END[9]),
    .X(net50));
 sg13g2_buf_1 input51 (.A(FrameData[0]),
    .X(net51));
 sg13g2_buf_1 input52 (.A(FrameData[10]),
    .X(net52));
 sg13g2_buf_1 input53 (.A(FrameData[11]),
    .X(net53));
 sg13g2_buf_1 input54 (.A(FrameData[12]),
    .X(net54));
 sg13g2_buf_1 input55 (.A(FrameData[13]),
    .X(net55));
 sg13g2_buf_4 input56 (.X(net56),
    .A(FrameData[14]));
 sg13g2_buf_4 input57 (.X(net57),
    .A(FrameData[15]));
 sg13g2_buf_4 input58 (.X(net58),
    .A(FrameData[16]));
 sg13g2_buf_4 input59 (.X(net78),
    .A(FrameData[17]));
 sg13g2_buf_2 input60 (.A(FrameData[18]),
    .X(net79));
 sg13g2_buf_4 input61 (.X(net80),
    .A(FrameData[19]));
 sg13g2_buf_1 input62 (.A(FrameData[1]),
    .X(net81));
 sg13g2_buf_4 input63 (.X(net82),
    .A(FrameData[20]));
 sg13g2_buf_2 input64 (.A(FrameData[21]),
    .X(net83));
 sg13g2_buf_4 input65 (.X(net84),
    .A(FrameData[22]));
 sg13g2_buf_4 input66 (.X(net85),
    .A(FrameData[23]));
 sg13g2_buf_4 input67 (.X(net86),
    .A(FrameData[24]));
 sg13g2_buf_4 input68 (.X(net87),
    .A(FrameData[25]));
 sg13g2_buf_2 input69 (.A(FrameData[26]),
    .X(net88));
 sg13g2_buf_2 input70 (.A(FrameData[27]),
    .X(net89));
 sg13g2_buf_1 input71 (.A(FrameData[28]),
    .X(net90));
 sg13g2_buf_1 input72 (.A(FrameData[29]),
    .X(net91));
 sg13g2_buf_2 input73 (.A(FrameData[2]),
    .X(net92));
 sg13g2_buf_2 input74 (.A(FrameData[30]),
    .X(net93));
 sg13g2_buf_2 input75 (.A(FrameData[31]),
    .X(net94));
 sg13g2_buf_2 input76 (.A(FrameData[3]),
    .X(net95));
 sg13g2_buf_2 input77 (.A(FrameData[4]),
    .X(net96));
 sg13g2_buf_2 input78 (.A(FrameData[5]),
    .X(net97));
 sg13g2_buf_2 input79 (.A(FrameData[6]),
    .X(net98));
 sg13g2_buf_4 input80 (.X(net99),
    .A(FrameData[7]));
 sg13g2_buf_2 input81 (.A(FrameData[8]),
    .X(net100));
 sg13g2_buf_2 input82 (.A(FrameData[9]),
    .X(net101));
 sg13g2_buf_1 output83 (.A(net102),
    .X(A_I_top));
 sg13g2_buf_1 output84 (.A(net103),
    .X(A_T_top));
 sg13g2_buf_1 output85 (.A(net104),
    .X(A_config_C_bit0));
 sg13g2_buf_1 output86 (.A(net105),
    .X(A_config_C_bit1));
 sg13g2_buf_1 output87 (.A(net106),
    .X(A_config_C_bit2));
 sg13g2_buf_1 output88 (.A(net107),
    .X(A_config_C_bit3));
 sg13g2_buf_1 output89 (.A(net108),
    .X(B_I_top));
 sg13g2_buf_1 output90 (.A(net109),
    .X(B_T_top));
 sg13g2_buf_1 output91 (.A(net110),
    .X(B_config_C_bit0));
 sg13g2_buf_1 output92 (.A(net111),
    .X(B_config_C_bit1));
 sg13g2_buf_1 output93 (.A(net112),
    .X(B_config_C_bit2));
 sg13g2_buf_1 output94 (.A(net113),
    .X(B_config_C_bit3));
 sg13g2_buf_1 output95 (.A(net114),
    .X(FrameData_O[0]));
 sg13g2_buf_1 output96 (.A(net115),
    .X(FrameData_O[10]));
 sg13g2_buf_1 output97 (.A(net116),
    .X(FrameData_O[11]));
 sg13g2_buf_1 output98 (.A(net117),
    .X(FrameData_O[12]));
 sg13g2_buf_1 output99 (.A(net118),
    .X(FrameData_O[13]));
 sg13g2_buf_1 output100 (.A(net119),
    .X(FrameData_O[14]));
 sg13g2_buf_1 output101 (.A(net120),
    .X(FrameData_O[15]));
 sg13g2_buf_1 output102 (.A(net121),
    .X(FrameData_O[16]));
 sg13g2_buf_1 output103 (.A(net122),
    .X(FrameData_O[17]));
 sg13g2_buf_1 output104 (.A(net123),
    .X(FrameData_O[18]));
 sg13g2_buf_1 output105 (.A(net124),
    .X(FrameData_O[19]));
 sg13g2_buf_1 output106 (.A(net125),
    .X(FrameData_O[1]));
 sg13g2_buf_1 output107 (.A(net126),
    .X(FrameData_O[20]));
 sg13g2_buf_1 output108 (.A(net127),
    .X(FrameData_O[21]));
 sg13g2_buf_1 output109 (.A(net128),
    .X(FrameData_O[22]));
 sg13g2_buf_1 output110 (.A(net129),
    .X(FrameData_O[23]));
 sg13g2_buf_1 output111 (.A(net130),
    .X(FrameData_O[24]));
 sg13g2_buf_1 output112 (.A(net131),
    .X(FrameData_O[25]));
 sg13g2_buf_1 output113 (.A(net132),
    .X(FrameData_O[26]));
 sg13g2_buf_1 output114 (.A(net133),
    .X(FrameData_O[27]));
 sg13g2_buf_1 output115 (.A(net134),
    .X(FrameData_O[28]));
 sg13g2_buf_1 output116 (.A(net135),
    .X(FrameData_O[29]));
 sg13g2_buf_1 output117 (.A(net136),
    .X(FrameData_O[2]));
 sg13g2_buf_1 output118 (.A(net137),
    .X(FrameData_O[30]));
 sg13g2_buf_1 output119 (.A(net138),
    .X(FrameData_O[31]));
 sg13g2_buf_1 output120 (.A(net139),
    .X(FrameData_O[3]));
 sg13g2_buf_1 output121 (.A(net140),
    .X(FrameData_O[4]));
 sg13g2_buf_1 output122 (.A(net141),
    .X(FrameData_O[5]));
 sg13g2_buf_1 output123 (.A(net142),
    .X(FrameData_O[6]));
 sg13g2_buf_1 output124 (.A(net143),
    .X(FrameData_O[7]));
 sg13g2_buf_1 output125 (.A(net144),
    .X(FrameData_O[8]));
 sg13g2_buf_1 output126 (.A(net145),
    .X(FrameData_O[9]));
 sg13g2_buf_1 output127 (.A(net146),
    .X(FrameStrobe_O[0]));
 sg13g2_buf_1 output128 (.A(net147),
    .X(FrameStrobe_O[10]));
 sg13g2_buf_1 output129 (.A(net148),
    .X(FrameStrobe_O[11]));
 sg13g2_buf_1 output130 (.A(net149),
    .X(FrameStrobe_O[12]));
 sg13g2_buf_1 output131 (.A(net150),
    .X(FrameStrobe_O[13]));
 sg13g2_buf_1 output132 (.A(net151),
    .X(FrameStrobe_O[14]));
 sg13g2_buf_1 output133 (.A(net152),
    .X(FrameStrobe_O[15]));
 sg13g2_buf_1 output134 (.A(net153),
    .X(FrameStrobe_O[16]));
 sg13g2_buf_1 output135 (.A(net154),
    .X(FrameStrobe_O[17]));
 sg13g2_buf_1 output136 (.A(net155),
    .X(FrameStrobe_O[18]));
 sg13g2_buf_1 output137 (.A(net156),
    .X(FrameStrobe_O[19]));
 sg13g2_buf_1 output138 (.A(net157),
    .X(FrameStrobe_O[1]));
 sg13g2_buf_1 output139 (.A(net158),
    .X(FrameStrobe_O[2]));
 sg13g2_buf_1 output140 (.A(net159),
    .X(FrameStrobe_O[3]));
 sg13g2_buf_1 output141 (.A(net160),
    .X(FrameStrobe_O[4]));
 sg13g2_buf_1 output142 (.A(net161),
    .X(FrameStrobe_O[5]));
 sg13g2_buf_1 output143 (.A(net162),
    .X(FrameStrobe_O[6]));
 sg13g2_buf_1 output144 (.A(net163),
    .X(FrameStrobe_O[7]));
 sg13g2_buf_1 output145 (.A(net164),
    .X(FrameStrobe_O[8]));
 sg13g2_buf_1 output146 (.A(net165),
    .X(FrameStrobe_O[9]));
 sg13g2_buf_1 output147 (.A(net166),
    .X(UserCLKo));
 sg13g2_buf_1 output148 (.A(net167),
    .X(W1BEG[0]));
 sg13g2_buf_1 output149 (.A(net168),
    .X(W1BEG[1]));
 sg13g2_buf_1 output150 (.A(net169),
    .X(W1BEG[2]));
 sg13g2_buf_1 output151 (.A(net170),
    .X(W1BEG[3]));
 sg13g2_buf_1 output152 (.A(net171),
    .X(W2BEG[0]));
 sg13g2_buf_1 output153 (.A(net172),
    .X(W2BEG[1]));
 sg13g2_buf_1 output154 (.A(net173),
    .X(W2BEG[2]));
 sg13g2_buf_1 output155 (.A(net174),
    .X(W2BEG[3]));
 sg13g2_buf_1 output156 (.A(net175),
    .X(W2BEG[4]));
 sg13g2_buf_1 output157 (.A(net176),
    .X(W2BEG[5]));
 sg13g2_buf_1 output158 (.A(net177),
    .X(W2BEG[6]));
 sg13g2_buf_1 output159 (.A(net178),
    .X(W2BEG[7]));
 sg13g2_buf_1 output160 (.A(net179),
    .X(W2BEGb[0]));
 sg13g2_buf_1 output161 (.A(net180),
    .X(W2BEGb[1]));
 sg13g2_buf_1 output162 (.A(net181),
    .X(W2BEGb[2]));
 sg13g2_buf_1 output163 (.A(net182),
    .X(W2BEGb[3]));
 sg13g2_buf_1 output164 (.A(net183),
    .X(W2BEGb[4]));
 sg13g2_buf_1 output165 (.A(net184),
    .X(W2BEGb[5]));
 sg13g2_buf_1 output166 (.A(net185),
    .X(W2BEGb[6]));
 sg13g2_buf_1 output167 (.A(net186),
    .X(W2BEGb[7]));
 sg13g2_buf_1 output168 (.A(net187),
    .X(W6BEG[0]));
 sg13g2_buf_1 output169 (.A(net188),
    .X(W6BEG[10]));
 sg13g2_buf_1 output170 (.A(net189),
    .X(W6BEG[11]));
 sg13g2_buf_1 output171 (.A(net190),
    .X(W6BEG[1]));
 sg13g2_buf_1 output172 (.A(net191),
    .X(W6BEG[2]));
 sg13g2_buf_1 output173 (.A(net192),
    .X(W6BEG[3]));
 sg13g2_buf_1 output174 (.A(net193),
    .X(W6BEG[4]));
 sg13g2_buf_1 output175 (.A(net194),
    .X(W6BEG[5]));
 sg13g2_buf_1 output176 (.A(net195),
    .X(W6BEG[6]));
 sg13g2_buf_1 output177 (.A(net196),
    .X(W6BEG[7]));
 sg13g2_buf_1 output178 (.A(net197),
    .X(W6BEG[8]));
 sg13g2_buf_1 output179 (.A(net198),
    .X(W6BEG[9]));
 sg13g2_buf_1 output180 (.A(net199),
    .X(WW4BEG[0]));
 sg13g2_buf_1 output181 (.A(net200),
    .X(WW4BEG[10]));
 sg13g2_buf_1 output182 (.A(net201),
    .X(WW4BEG[11]));
 sg13g2_buf_1 output183 (.A(net202),
    .X(WW4BEG[12]));
 sg13g2_buf_1 output184 (.A(net203),
    .X(WW4BEG[13]));
 sg13g2_buf_1 output185 (.A(net204),
    .X(WW4BEG[14]));
 sg13g2_buf_1 output186 (.A(net205),
    .X(WW4BEG[15]));
 sg13g2_buf_1 output187 (.A(net206),
    .X(WW4BEG[1]));
 sg13g2_buf_1 output188 (.A(net207),
    .X(WW4BEG[2]));
 sg13g2_buf_1 output189 (.A(net208),
    .X(WW4BEG[3]));
 sg13g2_buf_1 output190 (.A(net209),
    .X(WW4BEG[4]));
 sg13g2_buf_1 output191 (.A(net210),
    .X(WW4BEG[5]));
 sg13g2_buf_1 output192 (.A(net211),
    .X(WW4BEG[6]));
 sg13g2_buf_1 output193 (.A(net212),
    .X(WW4BEG[7]));
 sg13g2_buf_1 output194 (.A(net213),
    .X(WW4BEG[8]));
 sg13g2_buf_1 output195 (.A(net214),
    .X(WW4BEG[9]));
 sg13g2_tiehi _268__196 (.L_HI(net215));
 sg13g2_antennanp ANTENNA_2 (.A(FrameStrobe[10]));
 sg13g2_antennanp ANTENNA_3 (.A(FrameStrobe[11]));
 sg13g2_antennanp ANTENNA_4 (.A(FrameStrobe[12]));
 sg13g2_antennanp ANTENNA_5 (.A(FrameStrobe[14]));
 sg13g2_antennanp ANTENNA_6 (.A(FrameStrobe[16]));
 sg13g2_antennanp ANTENNA_7 (.A(FrameStrobe[18]));
 sg13g2_antennanp ANTENNA_8 (.A(FrameStrobe[19]));
 sg13g2_antennanp ANTENNA_9 (.A(FrameStrobe[3]));
 sg13g2_antennanp ANTENNA_10 (.A(FrameStrobe[4]));
 sg13g2_antennanp ANTENNA_11 (.A(FrameStrobe[6]));
 sg13g2_antennanp ANTENNA_12 (.A(FrameStrobe[7]));
 sg13g2_antennanp ANTENNA_13 (.A(FrameStrobe[8]));
 sg13g2_antennanp ANTENNA_14 (.A(FrameStrobe[9]));
 sg13g2_antennanp ANTENNA_15 (.A(net174));
 sg13g2_antennanp ANTENNA_16 (.A(net180));
 sg13g2_antennanp ANTENNA_17 (.A(net182));
 sg13g2_antennanp ANTENNA_18 (.A(net206));
 sg13g2_antennanp ANTENNA_19 (.A(FrameStrobe[10]));
 sg13g2_antennanp ANTENNA_20 (.A(FrameStrobe[11]));
 sg13g2_antennanp ANTENNA_21 (.A(FrameStrobe[12]));
 sg13g2_antennanp ANTENNA_22 (.A(FrameStrobe[14]));
 sg13g2_antennanp ANTENNA_23 (.A(FrameStrobe[16]));
 sg13g2_antennanp ANTENNA_24 (.A(FrameStrobe[18]));
 sg13g2_antennanp ANTENNA_25 (.A(FrameStrobe[19]));
 sg13g2_antennanp ANTENNA_26 (.A(FrameStrobe[3]));
 sg13g2_antennanp ANTENNA_27 (.A(FrameStrobe[4]));
 sg13g2_antennanp ANTENNA_28 (.A(FrameStrobe[6]));
 sg13g2_antennanp ANTENNA_29 (.A(FrameStrobe[7]));
 sg13g2_antennanp ANTENNA_30 (.A(FrameStrobe[8]));
 sg13g2_antennanp ANTENNA_31 (.A(FrameStrobe[9]));
 sg13g2_antennanp ANTENNA_32 (.A(net174));
 sg13g2_antennanp ANTENNA_33 (.A(net180));
 sg13g2_antennanp ANTENNA_34 (.A(net182));
 sg13g2_antennanp ANTENNA_35 (.A(net206));
 sg13g2_antennanp ANTENNA_36 (.A(FrameStrobe[10]));
 sg13g2_antennanp ANTENNA_37 (.A(FrameStrobe[11]));
 sg13g2_antennanp ANTENNA_38 (.A(FrameStrobe[12]));
 sg13g2_antennanp ANTENNA_39 (.A(FrameStrobe[14]));
 sg13g2_antennanp ANTENNA_40 (.A(FrameStrobe[16]));
 sg13g2_antennanp ANTENNA_41 (.A(FrameStrobe[18]));
 sg13g2_antennanp ANTENNA_42 (.A(FrameStrobe[19]));
 sg13g2_antennanp ANTENNA_43 (.A(FrameStrobe[3]));
 sg13g2_antennanp ANTENNA_44 (.A(FrameStrobe[4]));
 sg13g2_antennanp ANTENNA_45 (.A(FrameStrobe[6]));
 sg13g2_antennanp ANTENNA_46 (.A(FrameStrobe[7]));
 sg13g2_antennanp ANTENNA_47 (.A(FrameStrobe[8]));
 sg13g2_antennanp ANTENNA_48 (.A(FrameStrobe[9]));
 sg13g2_antennanp ANTENNA_49 (.A(net174));
 sg13g2_antennanp ANTENNA_50 (.A(net180));
 sg13g2_antennanp ANTENNA_51 (.A(net182));
 sg13g2_antennanp ANTENNA_52 (.A(net206));
 sg13g2_antennanp ANTENNA_53 (.A(FrameStrobe[10]));
 sg13g2_antennanp ANTENNA_54 (.A(FrameStrobe[11]));
 sg13g2_antennanp ANTENNA_55 (.A(FrameStrobe[12]));
 sg13g2_antennanp ANTENNA_56 (.A(FrameStrobe[14]));
 sg13g2_antennanp ANTENNA_57 (.A(FrameStrobe[16]));
 sg13g2_antennanp ANTENNA_58 (.A(FrameStrobe[18]));
 sg13g2_antennanp ANTENNA_59 (.A(FrameStrobe[19]));
 sg13g2_antennanp ANTENNA_60 (.A(FrameStrobe[3]));
 sg13g2_antennanp ANTENNA_61 (.A(FrameStrobe[4]));
 sg13g2_antennanp ANTENNA_62 (.A(FrameStrobe[6]));
 sg13g2_antennanp ANTENNA_63 (.A(FrameStrobe[7]));
 sg13g2_antennanp ANTENNA_64 (.A(FrameStrobe[8]));
 sg13g2_antennanp ANTENNA_65 (.A(FrameStrobe[9]));
 sg13g2_antennanp ANTENNA_66 (.A(net174));
 sg13g2_antennanp ANTENNA_67 (.A(net180));
 sg13g2_antennanp ANTENNA_68 (.A(net182));
 sg13g2_antennanp ANTENNA_69 (.A(net206));
 sg13g2_antennanp ANTENNA_70 (.A(FrameStrobe[10]));
 sg13g2_antennanp ANTENNA_71 (.A(FrameStrobe[11]));
 sg13g2_antennanp ANTENNA_72 (.A(FrameStrobe[12]));
 sg13g2_antennanp ANTENNA_73 (.A(FrameStrobe[14]));
 sg13g2_antennanp ANTENNA_74 (.A(FrameStrobe[16]));
 sg13g2_antennanp ANTENNA_75 (.A(FrameStrobe[18]));
 sg13g2_antennanp ANTENNA_76 (.A(FrameStrobe[19]));
 sg13g2_antennanp ANTENNA_77 (.A(FrameStrobe[3]));
 sg13g2_antennanp ANTENNA_78 (.A(FrameStrobe[4]));
 sg13g2_antennanp ANTENNA_79 (.A(FrameStrobe[6]));
 sg13g2_antennanp ANTENNA_80 (.A(FrameStrobe[7]));
 sg13g2_antennanp ANTENNA_81 (.A(FrameStrobe[8]));
 sg13g2_antennanp ANTENNA_82 (.A(FrameStrobe[9]));
 sg13g2_antennanp ANTENNA_83 (.A(net174));
 sg13g2_antennanp ANTENNA_84 (.A(net180));
 sg13g2_antennanp ANTENNA_85 (.A(net182));
 sg13g2_antennanp ANTENNA_86 (.A(net206));
 sg13g2_antennanp ANTENNA_87 (.A(FrameStrobe[10]));
 sg13g2_antennanp ANTENNA_88 (.A(FrameStrobe[11]));
 sg13g2_antennanp ANTENNA_89 (.A(FrameStrobe[12]));
 sg13g2_antennanp ANTENNA_90 (.A(FrameStrobe[14]));
 sg13g2_antennanp ANTENNA_91 (.A(FrameStrobe[16]));
 sg13g2_antennanp ANTENNA_92 (.A(FrameStrobe[18]));
 sg13g2_antennanp ANTENNA_93 (.A(FrameStrobe[19]));
 sg13g2_antennanp ANTENNA_94 (.A(FrameStrobe[3]));
 sg13g2_antennanp ANTENNA_95 (.A(FrameStrobe[4]));
 sg13g2_antennanp ANTENNA_96 (.A(FrameStrobe[6]));
 sg13g2_antennanp ANTENNA_97 (.A(FrameStrobe[7]));
 sg13g2_antennanp ANTENNA_98 (.A(FrameStrobe[8]));
 sg13g2_antennanp ANTENNA_99 (.A(FrameStrobe[9]));
 sg13g2_antennanp ANTENNA_100 (.A(net174));
 sg13g2_antennanp ANTENNA_101 (.A(net180));
 sg13g2_antennanp ANTENNA_102 (.A(net182));
 sg13g2_antennanp ANTENNA_103 (.A(net206));
 sg13g2_antennanp ANTENNA_104 (.A(FrameStrobe[10]));
 sg13g2_antennanp ANTENNA_105 (.A(FrameStrobe[11]));
 sg13g2_antennanp ANTENNA_106 (.A(FrameStrobe[12]));
 sg13g2_antennanp ANTENNA_107 (.A(FrameStrobe[16]));
 sg13g2_antennanp ANTENNA_108 (.A(FrameStrobe[18]));
 sg13g2_antennanp ANTENNA_109 (.A(FrameStrobe[19]));
 sg13g2_antennanp ANTENNA_110 (.A(FrameStrobe[3]));
 sg13g2_antennanp ANTENNA_111 (.A(FrameStrobe[4]));
 sg13g2_antennanp ANTENNA_112 (.A(FrameStrobe[6]));
 sg13g2_antennanp ANTENNA_113 (.A(FrameStrobe[7]));
 sg13g2_antennanp ANTENNA_114 (.A(FrameStrobe[9]));
 sg13g2_antennanp ANTENNA_115 (.A(net174));
 sg13g2_antennanp ANTENNA_116 (.A(net180));
 sg13g2_antennanp ANTENNA_117 (.A(net182));
 sg13g2_antennanp ANTENNA_118 (.A(net206));
 sg13g2_antennanp ANTENNA_119 (.A(FrameStrobe[10]));
 sg13g2_antennanp ANTENNA_120 (.A(FrameStrobe[11]));
 sg13g2_antennanp ANTENNA_121 (.A(FrameStrobe[12]));
 sg13g2_antennanp ANTENNA_122 (.A(FrameStrobe[16]));
 sg13g2_antennanp ANTENNA_123 (.A(FrameStrobe[17]));
 sg13g2_antennanp ANTENNA_124 (.A(FrameStrobe[18]));
 sg13g2_antennanp ANTENNA_125 (.A(FrameStrobe[19]));
 sg13g2_antennanp ANTENNA_126 (.A(FrameStrobe[3]));
 sg13g2_antennanp ANTENNA_127 (.A(FrameStrobe[4]));
 sg13g2_antennanp ANTENNA_128 (.A(FrameStrobe[6]));
 sg13g2_antennanp ANTENNA_129 (.A(net174));
 sg13g2_antennanp ANTENNA_130 (.A(net180));
 sg13g2_antennanp ANTENNA_131 (.A(net182));
 sg13g2_antennanp ANTENNA_132 (.A(net206));
 sg13g2_antennanp ANTENNA_133 (.A(FrameStrobe[10]));
 sg13g2_antennanp ANTENNA_134 (.A(FrameStrobe[16]));
 sg13g2_antennanp ANTENNA_135 (.A(FrameStrobe[17]));
 sg13g2_antennanp ANTENNA_136 (.A(FrameStrobe[18]));
 sg13g2_antennanp ANTENNA_137 (.A(FrameStrobe[19]));
 sg13g2_antennanp ANTENNA_138 (.A(FrameStrobe[3]));
 sg13g2_antennanp ANTENNA_139 (.A(FrameStrobe[4]));
 sg13g2_antennanp ANTENNA_140 (.A(FrameStrobe[9]));
 sg13g2_antennanp ANTENNA_141 (.A(net174));
 sg13g2_antennanp ANTENNA_142 (.A(net180));
 sg13g2_antennanp ANTENNA_143 (.A(net182));
 sg13g2_antennanp ANTENNA_144 (.A(net206));
 sg13g2_antennanp ANTENNA_145 (.A(FrameStrobe[10]));
 sg13g2_antennanp ANTENNA_146 (.A(FrameStrobe[17]));
 sg13g2_antennanp ANTENNA_147 (.A(FrameStrobe[18]));
 sg13g2_antennanp ANTENNA_148 (.A(FrameStrobe[19]));
 sg13g2_antennanp ANTENNA_149 (.A(FrameStrobe[4]));
 sg13g2_antennanp ANTENNA_150 (.A(FrameStrobe[6]));
 sg13g2_antennanp ANTENNA_151 (.A(FrameStrobe[9]));
 sg13g2_antennanp ANTENNA_152 (.A(net174));
 sg13g2_antennanp ANTENNA_153 (.A(net180));
 sg13g2_antennanp ANTENNA_154 (.A(net182));
 sg13g2_antennanp ANTENNA_155 (.A(net206));
 sg13g2_decap_8 FILLER_0_52 ();
 sg13g2_decap_8 FILLER_0_59 ();
 sg13g2_decap_8 FILLER_0_66 ();
 sg13g2_decap_8 FILLER_0_73 ();
 sg13g2_decap_8 FILLER_0_80 ();
 sg13g2_decap_4 FILLER_0_87 ();
 sg13g2_fill_1 FILLER_1_7 ();
 sg13g2_fill_1 FILLER_1_24 ();
 sg13g2_fill_2 FILLER_1_31 ();
 sg13g2_decap_8 FILLER_1_57 ();
 sg13g2_decap_8 FILLER_1_64 ();
 sg13g2_decap_8 FILLER_1_71 ();
 sg13g2_decap_8 FILLER_1_78 ();
 sg13g2_decap_8 FILLER_1_85 ();
 sg13g2_fill_2 FILLER_1_92 ();
 sg13g2_fill_1 FILLER_1_94 ();
 sg13g2_fill_1 FILLER_2_3 ();
 sg13g2_decap_8 FILLER_2_64 ();
 sg13g2_decap_8 FILLER_2_71 ();
 sg13g2_decap_8 FILLER_2_78 ();
 sg13g2_decap_8 FILLER_2_85 ();
 sg13g2_fill_2 FILLER_2_92 ();
 sg13g2_fill_1 FILLER_2_94 ();
 sg13g2_fill_2 FILLER_3_3 ();
 sg13g2_fill_2 FILLER_3_27 ();
 sg13g2_fill_1 FILLER_3_46 ();
 sg13g2_decap_8 FILLER_3_67 ();
 sg13g2_decap_8 FILLER_3_74 ();
 sg13g2_decap_8 FILLER_3_81 ();
 sg13g2_fill_2 FILLER_3_88 ();
 sg13g2_fill_1 FILLER_3_90 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_12 ();
 sg13g2_fill_1 FILLER_4_31 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_fill_1 FILLER_4_98 ();
 sg13g2_fill_2 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_55 ();
 sg13g2_decap_8 FILLER_5_86 ();
 sg13g2_fill_2 FILLER_5_93 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_fill_2 FILLER_7_30 ();
 sg13g2_fill_2 FILLER_7_49 ();
 sg13g2_decap_4 FILLER_7_68 ();
 sg13g2_fill_2 FILLER_7_93 ();
 sg13g2_fill_1 FILLER_8_37 ();
 sg13g2_decap_8 FILLER_8_60 ();
 sg13g2_decap_4 FILLER_8_77 ();
 sg13g2_fill_1 FILLER_8_98 ();
 sg13g2_fill_1 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_28 ();
 sg13g2_fill_2 FILLER_9_46 ();
 sg13g2_fill_2 FILLER_9_58 ();
 sg13g2_fill_1 FILLER_9_77 ();
 sg13g2_fill_2 FILLER_10_46 ();
 sg13g2_fill_1 FILLER_10_48 ();
 sg13g2_fill_2 FILLER_10_96 ();
 sg13g2_fill_1 FILLER_10_98 ();
 sg13g2_fill_2 FILLER_11_8 ();
 sg13g2_fill_1 FILLER_11_10 ();
 sg13g2_fill_2 FILLER_11_28 ();
 sg13g2_fill_1 FILLER_11_30 ();
 sg13g2_decap_8 FILLER_11_60 ();
 sg13g2_decap_4 FILLER_11_67 ();
 sg13g2_fill_1 FILLER_11_79 ();
 sg13g2_fill_2 FILLER_11_88 ();
 sg13g2_fill_1 FILLER_11_90 ();
 sg13g2_fill_2 FILLER_12_8 ();
 sg13g2_fill_2 FILLER_12_31 ();
 sg13g2_fill_1 FILLER_12_50 ();
 sg13g2_fill_1 FILLER_12_72 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_2 ();
 sg13g2_fill_1 FILLER_13_29 ();
 sg13g2_fill_1 FILLER_13_51 ();
 sg13g2_decap_4 FILLER_14_46 ();
 sg13g2_fill_1 FILLER_14_50 ();
 sg13g2_decap_4 FILLER_14_55 ();
 sg13g2_decap_8 FILLER_14_64 ();
 sg13g2_fill_1 FILLER_14_71 ();
 sg13g2_fill_1 FILLER_14_77 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_53 ();
 sg13g2_fill_2 FILLER_15_57 ();
 sg13g2_fill_2 FILLER_15_73 ();
 sg13g2_fill_2 FILLER_15_96 ();
 sg13g2_fill_1 FILLER_15_98 ();
 sg13g2_fill_1 FILLER_16_12 ();
 sg13g2_fill_2 FILLER_16_42 ();
 sg13g2_fill_1 FILLER_16_44 ();
 sg13g2_fill_1 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_54 ();
 sg13g2_fill_2 FILLER_16_61 ();
 sg13g2_fill_1 FILLER_16_90 ();
 sg13g2_fill_1 FILLER_17_33 ();
 sg13g2_fill_2 FILLER_17_93 ();
 sg13g2_decap_8 FILLER_18_44 ();
 sg13g2_decap_4 FILLER_18_68 ();
 sg13g2_fill_2 FILLER_18_72 ();
 sg13g2_fill_1 FILLER_19_5 ();
 sg13g2_fill_1 FILLER_19_27 ();
 sg13g2_fill_2 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_61 ();
 sg13g2_fill_2 FILLER_19_97 ();
 sg13g2_fill_1 FILLER_20_52 ();
 sg13g2_fill_2 FILLER_20_57 ();
 sg13g2_fill_1 FILLER_21_5 ();
 sg13g2_fill_1 FILLER_21_27 ();
 sg13g2_decap_8 FILLER_21_57 ();
 sg13g2_fill_2 FILLER_21_64 ();
 sg13g2_fill_1 FILLER_21_66 ();
 sg13g2_fill_2 FILLER_21_92 ();
 sg13g2_fill_1 FILLER_21_94 ();
 sg13g2_fill_2 FILLER_22_5 ();
 sg13g2_fill_2 FILLER_22_68 ();
 sg13g2_fill_2 FILLER_22_96 ();
 sg13g2_fill_1 FILLER_22_98 ();
 sg13g2_fill_2 FILLER_23_39 ();
 sg13g2_fill_2 FILLER_24_97 ();
 sg13g2_fill_1 FILLER_25_5 ();
 sg13g2_fill_2 FILLER_25_97 ();
 sg13g2_fill_2 FILLER_26_5 ();
 sg13g2_fill_2 FILLER_26_55 ();
 sg13g2_fill_1 FILLER_27_27 ();
 sg13g2_fill_2 FILLER_27_49 ();
 sg13g2_fill_1 FILLER_27_74 ();
 sg13g2_fill_2 FILLER_28_44 ();
 sg13g2_fill_1 FILLER_28_59 ();
 sg13g2_fill_2 FILLER_28_68 ();
 sg13g2_fill_2 FILLER_29_72 ();
 sg13g2_fill_2 FILLER_29_97 ();
 sg13g2_fill_2 FILLER_30_17 ();
 sg13g2_fill_1 FILLER_30_29 ();
 sg13g2_fill_1 FILLER_30_81 ();
 sg13g2_fill_1 FILLER_31_17 ();
 sg13g2_fill_2 FILLER_31_48 ();
 sg13g2_fill_2 FILLER_31_67 ();
 sg13g2_fill_1 FILLER_32_5 ();
 sg13g2_fill_1 FILLER_32_23 ();
 sg13g2_fill_2 FILLER_32_89 ();
 sg13g2_fill_1 FILLER_33_81 ();
 sg13g2_fill_1 FILLER_34_51 ();
 sg13g2_fill_2 FILLER_34_97 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_65 ();
 sg13g2_fill_1 FILLER_36_10 ();
 sg13g2_fill_2 FILLER_36_33 ();
 sg13g2_fill_2 FILLER_36_64 ();
 sg13g2_fill_1 FILLER_36_83 ();
 sg13g2_fill_2 FILLER_36_93 ();
 sg13g2_fill_1 FILLER_37_17 ();
 sg13g2_fill_2 FILLER_37_76 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_19 ();
 sg13g2_fill_2 FILLER_38_86 ();
 sg13g2_fill_2 FILLER_38_97 ();
 sg13g2_fill_2 FILLER_39_58 ();
 sg13g2_fill_2 FILLER_39_97 ();
 sg13g2_fill_2 FILLER_40_79 ();
 sg13g2_fill_2 FILLER_41_51 ();
 sg13g2_fill_1 FILLER_42_68 ();
 sg13g2_fill_1 FILLER_42_98 ();
 sg13g2_fill_2 FILLER_44_71 ();
 sg13g2_fill_1 FILLER_45_61 ();
 sg13g2_fill_1 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_39 ();
 sg13g2_fill_1 FILLER_46_61 ();
 sg13g2_fill_1 FILLER_46_83 ();
 sg13g2_fill_2 FILLER_46_89 ();
 sg13g2_fill_2 FILLER_47_49 ();
 sg13g2_fill_2 FILLER_47_97 ();
 sg13g2_fill_2 FILLER_48_29 ();
 sg13g2_fill_1 FILLER_48_48 ();
 sg13g2_fill_1 FILLER_48_59 ();
 sg13g2_fill_2 FILLER_48_77 ();
 sg13g2_fill_2 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_98 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_19 ();
 sg13g2_fill_2 FILLER_50_67 ();
 sg13g2_fill_1 FILLER_51_8 ();
 sg13g2_fill_2 FILLER_51_89 ();
 sg13g2_fill_2 FILLER_52_44 ();
 sg13g2_fill_2 FILLER_53_52 ();
 sg13g2_fill_1 FILLER_54_20 ();
 sg13g2_fill_2 FILLER_54_73 ();
 sg13g2_fill_1 FILLER_54_84 ();
 sg13g2_fill_1 FILLER_55_16 ();
 sg13g2_fill_1 FILLER_55_29 ();
 sg13g2_fill_1 FILLER_55_37 ();
 sg13g2_fill_2 FILLER_55_45 ();
 sg13g2_fill_2 FILLER_55_59 ();
 sg13g2_fill_2 FILLER_55_79 ();
 sg13g2_fill_1 FILLER_55_84 ();
 sg13g2_fill_2 FILLER_56_23 ();
 sg13g2_fill_1 FILLER_56_37 ();
 sg13g2_fill_2 FILLER_56_50 ();
 sg13g2_fill_1 FILLER_56_60 ();
 sg13g2_fill_2 FILLER_56_79 ();
 sg13g2_fill_2 FILLER_56_89 ();
 sg13g2_fill_2 FILLER_57_8 ();
 sg13g2_fill_1 FILLER_57_28 ();
 sg13g2_fill_2 FILLER_57_93 ();
endmodule
