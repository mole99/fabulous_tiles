magic
tech sky130A
magscale 1 2
timestamp 1740383322
<< viali >>
rect 3433 8585 3467 8619
rect 4169 8585 4203 8619
rect 4537 8585 4571 8619
rect 5273 8585 5307 8619
rect 5641 8585 5675 8619
rect 6469 8585 6503 8619
rect 6837 8585 6871 8619
rect 7205 8585 7239 8619
rect 9321 8585 9355 8619
rect 10057 8585 10091 8619
rect 10885 8585 10919 8619
rect 11161 8585 11195 8619
rect 12173 8585 12207 8619
rect 12817 8585 12851 8619
rect 13185 8585 13219 8619
rect 13829 8585 13863 8619
rect 14933 8585 14967 8619
rect 15301 8585 15335 8619
rect 16405 8585 16439 8619
rect 17049 8585 17083 8619
rect 18843 8585 18877 8619
rect 21281 8585 21315 8619
rect 24409 8585 24443 8619
rect 24869 8585 24903 8619
rect 25789 8585 25823 8619
rect 29193 8585 29227 8619
rect 31585 8585 31619 8619
rect 33241 8585 33275 8619
rect 33885 8585 33919 8619
rect 35541 8585 35575 8619
rect 36645 8585 36679 8619
rect 37749 8585 37783 8619
rect 38485 8585 38519 8619
rect 39037 8585 39071 8619
rect 2329 8449 2363 8483
rect 3617 8449 3651 8483
rect 3801 8449 3835 8483
rect 4353 8449 4387 8483
rect 4721 8449 4755 8483
rect 5089 8449 5123 8483
rect 5457 8449 5491 8483
rect 5825 8449 5859 8483
rect 6193 8449 6227 8483
rect 6653 8449 6687 8483
rect 7021 8449 7055 8483
rect 7389 8449 7423 8483
rect 7757 8449 7791 8483
rect 9505 8449 9539 8483
rect 9873 8449 9907 8483
rect 10241 8449 10275 8483
rect 10333 8449 10367 8483
rect 10701 8449 10735 8483
rect 11345 8449 11379 8483
rect 11897 8449 11931 8483
rect 11989 8449 12023 8483
rect 12357 8449 12391 8483
rect 13001 8449 13035 8483
rect 13369 8449 13403 8483
rect 13461 8449 13495 8483
rect 13645 8449 13679 8483
rect 14289 8449 14323 8483
rect 14657 8449 14691 8483
rect 14749 8449 14783 8483
rect 15117 8449 15151 8483
rect 15761 8449 15795 8483
rect 16129 8449 16163 8483
rect 16221 8449 16255 8483
rect 17233 8449 17267 8483
rect 17877 8449 17911 8483
rect 18153 8449 18187 8483
rect 19073 8449 19107 8483
rect 19533 8449 19567 8483
rect 20729 8449 20763 8483
rect 21465 8449 21499 8483
rect 22017 8449 22051 8483
rect 22109 8449 22143 8483
rect 22385 8449 22419 8483
rect 22845 8449 22879 8483
rect 23397 8449 23431 8483
rect 24041 8449 24075 8483
rect 24593 8449 24627 8483
rect 24685 8449 24719 8483
rect 25145 8449 25179 8483
rect 25421 8449 25455 8483
rect 25697 8449 25731 8483
rect 25973 8449 26007 8483
rect 26249 8449 26283 8483
rect 26341 8449 26375 8483
rect 26801 8449 26835 8483
rect 27169 8449 27203 8483
rect 27445 8449 27479 8483
rect 27537 8449 27571 8483
rect 27997 8449 28031 8483
rect 28273 8449 28307 8483
rect 28365 8449 28399 8483
rect 28825 8449 28859 8483
rect 29101 8449 29135 8483
rect 29377 8449 29411 8483
rect 29837 8449 29871 8483
rect 30665 8449 30699 8483
rect 30941 8449 30975 8483
rect 31217 8449 31251 8483
rect 31493 8449 31527 8483
rect 31769 8449 31803 8483
rect 32413 8449 32447 8483
rect 33057 8449 33091 8483
rect 33701 8449 33735 8483
rect 34069 8449 34103 8483
rect 34437 8449 34471 8483
rect 34989 8449 35023 8483
rect 35357 8449 35391 8483
rect 35725 8449 35759 8483
rect 35817 8449 35851 8483
rect 36461 8449 36495 8483
rect 36829 8449 36863 8483
rect 37289 8449 37323 8483
rect 37933 8449 37967 8483
rect 38025 8449 38059 8483
rect 38669 8449 38703 8483
rect 39129 8449 39163 8483
rect 39221 8449 39255 8483
rect 1409 8381 1443 8415
rect 1685 8381 1719 8415
rect 2605 8381 2639 8415
rect 7481 8381 7515 8415
rect 16865 8381 16899 8415
rect 19257 8381 19291 8415
rect 20821 8381 20855 8415
rect 20913 8381 20947 8415
rect 23489 8381 23523 8415
rect 23581 8381 23615 8415
rect 29561 8381 29595 8415
rect 32137 8381 32171 8415
rect 3985 8313 4019 8347
rect 4905 8313 4939 8347
rect 6009 8313 6043 8347
rect 10517 8313 10551 8347
rect 11713 8313 11747 8347
rect 12541 8313 12575 8347
rect 14105 8313 14139 8347
rect 14473 8313 14507 8347
rect 15577 8313 15611 8347
rect 15945 8313 15979 8347
rect 20269 8313 20303 8347
rect 21833 8313 21867 8347
rect 22293 8313 22327 8347
rect 22569 8313 22603 8347
rect 22661 8313 22695 8347
rect 24961 8313 24995 8347
rect 26065 8313 26099 8347
rect 27721 8313 27755 8347
rect 28089 8313 28123 8347
rect 28549 8313 28583 8347
rect 31033 8313 31067 8347
rect 33517 8313 33551 8347
rect 34253 8313 34287 8347
rect 34805 8313 34839 8347
rect 35173 8313 35207 8347
rect 36277 8313 36311 8347
rect 38209 8313 38243 8347
rect 39405 8313 39439 8347
rect 8493 8245 8527 8279
rect 9689 8245 9723 8279
rect 20361 8245 20395 8279
rect 23029 8245 23063 8279
rect 23857 8245 23891 8279
rect 25237 8245 25271 8279
rect 25513 8245 25547 8279
rect 26525 8245 26559 8279
rect 26617 8245 26651 8279
rect 26985 8245 27019 8279
rect 27261 8245 27295 8279
rect 27813 8245 27847 8279
rect 28641 8245 28675 8279
rect 28917 8245 28951 8279
rect 30481 8245 30515 8279
rect 30757 8245 30791 8279
rect 31309 8245 31343 8279
rect 36001 8245 36035 8279
rect 37473 8245 37507 8279
rect 3433 8041 3467 8075
rect 3893 8041 3927 8075
rect 4261 8041 4295 8075
rect 4813 8041 4847 8075
rect 5365 8041 5399 8075
rect 5825 8041 5859 8075
rect 6193 8041 6227 8075
rect 6837 8041 6871 8075
rect 7481 8041 7515 8075
rect 10149 8041 10183 8075
rect 15577 8041 15611 8075
rect 19717 8041 19751 8075
rect 24961 8041 24995 8075
rect 26249 8041 26283 8075
rect 33241 8041 33275 8075
rect 33793 8041 33827 8075
rect 34805 8041 34839 8075
rect 35725 8041 35759 8075
rect 36277 8041 36311 8075
rect 36921 8041 36955 8075
rect 37289 8041 37323 8075
rect 38209 8041 38243 8075
rect 38669 8041 38703 8075
rect 2605 7973 2639 8007
rect 7113 7973 7147 8007
rect 9965 7973 9999 8007
rect 11805 7973 11839 8007
rect 12725 7973 12759 8007
rect 16865 7973 16899 8007
rect 20637 7973 20671 8007
rect 22109 7973 22143 8007
rect 27445 7973 27479 8007
rect 28365 7973 28399 8007
rect 32413 7973 32447 8007
rect 35081 7973 35115 8007
rect 38025 7973 38059 8007
rect 1409 7905 1443 7939
rect 2973 7905 3007 7939
rect 10425 7905 10459 7939
rect 13277 7905 13311 7939
rect 15117 7905 15151 7939
rect 15853 7905 15887 7939
rect 17693 7905 17727 7939
rect 18245 7905 18279 7939
rect 19993 7905 20027 7939
rect 20177 7905 20211 7939
rect 21030 7905 21064 7939
rect 21189 7905 21223 7939
rect 22385 7905 22419 7939
rect 22569 7905 22603 7939
rect 23029 7905 23063 7939
rect 23305 7905 23339 7939
rect 23443 7905 23477 7939
rect 25237 7905 25271 7939
rect 30757 7905 30791 7939
rect 1685 7837 1719 7871
rect 2789 7837 2823 7871
rect 3065 7837 3099 7871
rect 3617 7837 3651 7871
rect 4077 7837 4111 7871
rect 4445 7837 4479 7871
rect 4997 7837 5031 7871
rect 5549 7837 5583 7871
rect 6009 7837 6043 7871
rect 6377 7837 6411 7871
rect 6561 7837 6595 7871
rect 6653 7837 6687 7871
rect 7297 7837 7331 7871
rect 7665 7837 7699 7871
rect 7757 7837 7791 7871
rect 8033 7837 8067 7871
rect 8953 7837 8987 7871
rect 9229 7837 9263 7871
rect 10333 7837 10367 7871
rect 10701 7837 10735 7871
rect 11989 7837 12023 7871
rect 12081 7837 12115 7871
rect 12265 7837 12299 7871
rect 13001 7837 13035 7871
rect 13118 7837 13152 7871
rect 14841 7837 14875 7871
rect 15393 7837 15427 7871
rect 15761 7837 15795 7871
rect 16129 7837 16163 7871
rect 17509 7837 17543 7871
rect 17969 7837 18003 7871
rect 18521 7837 18555 7871
rect 19441 7813 19475 7847
rect 19901 7833 19935 7867
rect 20913 7837 20947 7871
rect 22293 7837 22327 7871
rect 23581 7837 23615 7871
rect 24225 7837 24259 7871
rect 24593 7837 24627 7871
rect 24685 7837 24719 7871
rect 25145 7837 25179 7871
rect 25513 7837 25547 7871
rect 27077 7837 27111 7871
rect 27353 7837 27387 7871
rect 27629 7837 27663 7871
rect 29101 7837 29135 7871
rect 29377 7837 29411 7871
rect 29653 7837 29687 7871
rect 29929 7837 29963 7871
rect 31033 7837 31067 7871
rect 32045 7837 32079 7871
rect 32321 7837 32355 7871
rect 32597 7837 32631 7871
rect 32873 7837 32907 7871
rect 33149 7837 33183 7871
rect 33425 7837 33459 7871
rect 33977 7837 34011 7871
rect 34161 7837 34195 7871
rect 34989 7837 35023 7871
rect 35265 7837 35299 7871
rect 35357 7837 35391 7871
rect 35909 7837 35943 7871
rect 36461 7837 36495 7871
rect 36737 7837 36771 7871
rect 37105 7837 37139 7871
rect 37565 7837 37599 7871
rect 37841 7837 37875 7871
rect 38393 7837 38427 7871
rect 38485 7837 38519 7871
rect 38853 7837 38887 7871
rect 39221 7837 39255 7871
rect 2421 7769 2455 7803
rect 13921 7769 13955 7803
rect 27997 7769 28031 7803
rect 3249 7701 3283 7735
rect 6561 7701 6595 7735
rect 8769 7701 8803 7735
rect 11437 7701 11471 7735
rect 14105 7701 14139 7735
rect 15209 7701 15243 7735
rect 17141 7701 17175 7735
rect 17601 7701 17635 7735
rect 18153 7701 18187 7735
rect 19625 7701 19659 7735
rect 21833 7701 21867 7735
rect 24409 7701 24443 7735
rect 24869 7701 24903 7735
rect 26341 7701 26375 7735
rect 28089 7701 28123 7735
rect 30665 7701 30699 7735
rect 31769 7701 31803 7735
rect 31861 7701 31895 7735
rect 32137 7701 32171 7735
rect 32689 7701 32723 7735
rect 32965 7701 32999 7735
rect 34345 7701 34379 7735
rect 35541 7701 35575 7735
rect 37381 7701 37415 7735
rect 39037 7701 39071 7735
rect 39405 7701 39439 7735
rect 1593 7497 1627 7531
rect 5365 7497 5399 7531
rect 5825 7497 5859 7531
rect 7297 7497 7331 7531
rect 11897 7497 11931 7531
rect 13369 7497 13403 7531
rect 13645 7497 13679 7531
rect 14013 7497 14047 7531
rect 15025 7497 15059 7531
rect 15301 7497 15335 7531
rect 16221 7497 16255 7531
rect 17049 7497 17083 7531
rect 17325 7497 17359 7531
rect 17693 7497 17727 7531
rect 18337 7497 18371 7531
rect 18613 7497 18647 7531
rect 19073 7497 19107 7531
rect 20453 7497 20487 7531
rect 21005 7497 21039 7531
rect 22109 7497 22143 7531
rect 23213 7497 23247 7531
rect 24133 7497 24167 7531
rect 27169 7497 27203 7531
rect 31217 7497 31251 7531
rect 31493 7497 31527 7531
rect 32137 7497 32171 7531
rect 32505 7497 32539 7531
rect 35541 7497 35575 7531
rect 37473 7497 37507 7531
rect 38301 7497 38335 7531
rect 38669 7497 38703 7531
rect 39037 7497 39071 7531
rect 39405 7497 39439 7531
rect 1869 7429 1903 7463
rect 2605 7429 2639 7463
rect 3157 7429 3191 7463
rect 6745 7429 6779 7463
rect 12817 7429 12851 7463
rect 14473 7429 14507 7463
rect 23765 7429 23799 7463
rect 1501 7361 1535 7395
rect 2237 7361 2271 7395
rect 2973 7361 3007 7395
rect 5181 7361 5215 7395
rect 6837 7361 6871 7395
rect 7481 7361 7515 7395
rect 7757 7361 7791 7395
rect 8677 7361 8711 7395
rect 8953 7361 8987 7395
rect 9873 7361 9907 7395
rect 10241 7361 10275 7395
rect 11345 7361 11379 7395
rect 11989 7361 12023 7395
rect 12725 7361 12759 7395
rect 13185 7361 13219 7395
rect 13829 7361 13863 7395
rect 14381 7361 14415 7395
rect 15209 7361 15243 7395
rect 15485 7361 15519 7395
rect 16037 7361 16071 7395
rect 16957 7361 16991 7395
rect 17233 7361 17267 7395
rect 18153 7361 18187 7395
rect 18797 7361 18831 7395
rect 18889 7361 18923 7395
rect 19165 7361 19199 7395
rect 19720 7361 19754 7395
rect 20729 7361 20763 7395
rect 21189 7361 21223 7395
rect 21925 7361 21959 7395
rect 22477 7361 22511 7395
rect 23673 7361 23707 7395
rect 25145 7361 25179 7395
rect 26985 7361 27019 7395
rect 27537 7361 27571 7395
rect 28457 7361 28491 7395
rect 29101 7361 29135 7395
rect 29837 7361 29871 7395
rect 30573 7361 30607 7395
rect 31033 7361 31067 7395
rect 31309 7361 31343 7395
rect 31769 7361 31803 7395
rect 35357 7361 35391 7395
rect 37657 7361 37691 7395
rect 37749 7361 37783 7395
rect 38117 7361 38151 7395
rect 38485 7361 38519 7395
rect 38853 7361 38887 7395
rect 39221 7361 39255 7395
rect 2421 7293 2455 7327
rect 5917 7293 5951 7327
rect 6101 7293 6135 7327
rect 6929 7293 6963 7327
rect 8815 7293 8849 7327
rect 9689 7293 9723 7327
rect 9965 7293 9999 7327
rect 12081 7293 12115 7327
rect 12909 7293 12943 7327
rect 14565 7293 14599 7327
rect 17785 7293 17819 7327
rect 17877 7293 17911 7327
rect 19441 7293 19475 7327
rect 22201 7293 22235 7327
rect 23581 7293 23615 7327
rect 27261 7293 27295 7327
rect 30665 7293 30699 7327
rect 30757 7293 30791 7327
rect 32597 7293 32631 7327
rect 32689 7293 32723 7327
rect 2053 7225 2087 7259
rect 6377 7225 6411 7259
rect 8033 7225 8067 7259
rect 9229 7225 9263 7259
rect 10977 7225 11011 7259
rect 11161 7225 11195 7259
rect 12357 7225 12391 7259
rect 20913 7225 20947 7259
rect 28273 7225 28307 7259
rect 29285 7225 29319 7259
rect 31585 7225 31619 7259
rect 37933 7225 37967 7259
rect 2697 7157 2731 7191
rect 5457 7157 5491 7191
rect 7849 7157 7883 7191
rect 11529 7157 11563 7191
rect 16773 7157 16807 7191
rect 18337 7157 18371 7191
rect 19349 7157 19383 7191
rect 25329 7157 25363 7191
rect 28641 7157 28675 7191
rect 30021 7157 30055 7191
rect 30205 7157 30239 7191
rect 4905 6953 4939 6987
rect 8769 6953 8803 6987
rect 10057 6953 10091 6987
rect 11253 6953 11287 6987
rect 15209 6953 15243 6987
rect 16129 6953 16163 6987
rect 37841 6953 37875 6987
rect 20545 6885 20579 6919
rect 22293 6885 22327 6919
rect 25145 6885 25179 6919
rect 12265 6817 12299 6851
rect 14565 6817 14599 6851
rect 14749 6817 14783 6851
rect 16865 6817 16899 6851
rect 17049 6817 17083 6851
rect 17417 6817 17451 6851
rect 17877 6817 17911 6851
rect 18270 6817 18304 6851
rect 21189 6817 21223 6851
rect 30113 6817 30147 6851
rect 31677 6817 31711 6851
rect 32321 6817 32355 6851
rect 32597 6817 32631 6851
rect 1409 6749 1443 6783
rect 1685 6749 1719 6783
rect 3893 6749 3927 6783
rect 4169 6749 4203 6783
rect 5549 6749 5583 6783
rect 6469 6749 6503 6783
rect 7757 6749 7791 6783
rect 8033 6749 8067 6783
rect 9222 6749 9256 6783
rect 9413 6749 9447 6783
rect 10241 6749 10275 6783
rect 10609 6749 10643 6783
rect 10701 6749 10735 6783
rect 11437 6749 11471 6783
rect 11529 6749 11563 6783
rect 13185 6749 13219 6783
rect 16313 6749 16347 6783
rect 16773 6749 16807 6783
rect 17233 6749 17267 6783
rect 18153 6749 18187 6783
rect 18429 6749 18463 6783
rect 19533 6749 19567 6783
rect 19809 6749 19843 6783
rect 21097 6749 21131 6783
rect 23029 6749 23063 6783
rect 23305 6749 23339 6783
rect 25329 6749 25363 6783
rect 28825 6749 28859 6783
rect 29929 6749 29963 6783
rect 30573 6749 30607 6783
rect 31401 6749 31435 6783
rect 31861 6749 31895 6783
rect 32735 6749 32769 6783
rect 32873 6749 32907 6783
rect 37657 6749 37691 6783
rect 38117 6749 38151 6783
rect 38393 6749 38427 6783
rect 38485 6749 38519 6783
rect 38853 6749 38887 6783
rect 39221 6749 39255 6783
rect 14841 6681 14875 6715
rect 5733 6613 5767 6647
rect 6653 6613 6687 6647
rect 9045 6613 9079 6647
rect 9597 6613 9631 6647
rect 10425 6613 10459 6647
rect 10885 6613 10919 6647
rect 11713 6613 11747 6647
rect 12449 6613 12483 6647
rect 12541 6613 12575 6647
rect 12909 6613 12943 6647
rect 13001 6613 13035 6647
rect 16405 6613 16439 6647
rect 19073 6613 19107 6647
rect 20637 6613 20671 6647
rect 21005 6613 21039 6647
rect 28641 6613 28675 6647
rect 29561 6613 29595 6647
rect 30021 6613 30055 6647
rect 30389 6613 30423 6647
rect 31217 6613 31251 6647
rect 33517 6613 33551 6647
rect 38025 6613 38059 6647
rect 38209 6613 38243 6647
rect 38669 6613 38703 6647
rect 39037 6613 39071 6647
rect 39405 6613 39439 6647
rect 5733 6409 5767 6443
rect 7757 6409 7791 6443
rect 11989 6409 12023 6443
rect 17693 6409 17727 6443
rect 18153 6409 18187 6443
rect 20269 6409 20303 6443
rect 22385 6409 22419 6443
rect 23489 6409 23523 6443
rect 28733 6409 28767 6443
rect 31125 6409 31159 6443
rect 32137 6409 32171 6443
rect 33241 6409 33275 6443
rect 35725 6409 35759 6443
rect 38577 6409 38611 6443
rect 39405 6409 39439 6443
rect 3709 6341 3743 6375
rect 4445 6341 4479 6375
rect 18521 6341 18555 6375
rect 1501 6273 1535 6307
rect 1777 6273 1811 6307
rect 4629 6273 4663 6307
rect 4721 6273 4755 6307
rect 4997 6273 5031 6307
rect 7021 6273 7055 6307
rect 7849 6273 7883 6307
rect 8401 6273 8435 6307
rect 9413 6273 9447 6307
rect 10517 6273 10551 6307
rect 12725 6273 12759 6307
rect 13001 6273 13035 6307
rect 13185 6273 13219 6307
rect 13461 6273 13495 6307
rect 15485 6273 15519 6307
rect 16129 6273 16163 6307
rect 16957 6273 16991 6307
rect 18061 6273 18095 6307
rect 18613 6273 18647 6307
rect 20177 6273 20211 6307
rect 20913 6273 20947 6307
rect 21189 6273 21223 6307
rect 23121 6273 23155 6307
rect 24225 6273 24259 6307
rect 24501 6273 24535 6307
rect 25053 6273 25087 6307
rect 26249 6273 26283 6307
rect 27261 6273 27295 6307
rect 28917 6273 28951 6307
rect 29653 6273 29687 6307
rect 29929 6273 29963 6307
rect 31493 6273 31527 6307
rect 32321 6273 32355 6307
rect 33977 6273 34011 6307
rect 34529 6273 34563 6307
rect 34805 6273 34839 6307
rect 35817 6273 35851 6307
rect 38761 6273 38795 6307
rect 38853 6273 38887 6307
rect 39221 6273 39255 6307
rect 1685 6205 1719 6239
rect 6745 6205 6779 6239
rect 9137 6205 9171 6239
rect 10241 6205 10275 6239
rect 14289 6205 14323 6239
rect 14473 6205 14507 6239
rect 15209 6205 15243 6239
rect 15347 6205 15381 6239
rect 16681 6205 16715 6239
rect 18705 6205 18739 6239
rect 20085 6205 20119 6239
rect 23397 6205 23431 6239
rect 24777 6205 24811 6239
rect 26341 6205 26375 6239
rect 26433 6205 26467 6239
rect 26985 6205 27019 6239
rect 29791 6205 29825 6239
rect 30665 6205 30699 6239
rect 30849 6205 30883 6239
rect 31585 6205 31619 6239
rect 31769 6205 31803 6239
rect 34253 6205 34287 6239
rect 3893 6137 3927 6171
rect 14197 6137 14231 6171
rect 14933 6137 14967 6171
rect 20637 6137 20671 6171
rect 21005 6137 21039 6171
rect 25789 6137 25823 6171
rect 27997 6137 28031 6171
rect 30205 6137 30239 6171
rect 1961 6069 1995 6103
rect 8033 6069 8067 6103
rect 8493 6069 8527 6103
rect 10149 6069 10183 6103
rect 11253 6069 11287 6103
rect 17877 6069 17911 6103
rect 20729 6069 20763 6103
rect 25881 6069 25915 6103
rect 29009 6069 29043 6103
rect 35541 6069 35575 6103
rect 39037 6069 39071 6103
rect 1593 5865 1627 5899
rect 2145 5865 2179 5899
rect 15117 5865 15151 5899
rect 21833 5865 21867 5899
rect 24409 5865 24443 5899
rect 28641 5865 28675 5899
rect 32229 5865 32263 5899
rect 36001 5865 36035 5899
rect 39405 5865 39439 5899
rect 5089 5797 5123 5831
rect 9321 5797 9355 5831
rect 28549 5797 28583 5831
rect 39037 5797 39071 5831
rect 6285 5729 6319 5763
rect 11989 5729 12023 5763
rect 12725 5729 12759 5763
rect 12909 5729 12943 5763
rect 27537 5729 27571 5763
rect 29193 5729 29227 5763
rect 30481 5729 30515 5763
rect 30941 5729 30975 5763
rect 31493 5729 31527 5763
rect 32781 5729 32815 5763
rect 35449 5729 35483 5763
rect 1409 5661 1443 5695
rect 1685 5661 1719 5695
rect 1961 5661 1995 5695
rect 4537 5661 4571 5695
rect 4813 5661 4847 5695
rect 4905 5661 4939 5695
rect 6561 5661 6595 5695
rect 9137 5661 9171 5695
rect 10517 5661 10551 5695
rect 11161 5661 11195 5695
rect 11897 5661 11931 5695
rect 14105 5661 14139 5695
rect 14381 5661 14415 5695
rect 20821 5661 20855 5695
rect 21097 5661 21131 5695
rect 25145 5661 25179 5695
rect 25421 5661 25455 5695
rect 26433 5661 26467 5695
rect 26709 5661 26743 5695
rect 27813 5661 27847 5695
rect 30297 5661 30331 5695
rect 31217 5661 31251 5695
rect 31334 5661 31368 5695
rect 32137 5661 32171 5695
rect 32689 5661 32723 5695
rect 38209 5661 38243 5695
rect 38853 5661 38887 5695
rect 39221 5661 39255 5695
rect 11805 5593 11839 5627
rect 35633 5593 35667 5627
rect 1869 5525 1903 5559
rect 3801 5525 3835 5559
rect 7297 5525 7331 5559
rect 10609 5525 10643 5559
rect 11345 5525 11379 5559
rect 11437 5525 11471 5559
rect 12265 5525 12299 5559
rect 12633 5525 12667 5559
rect 27445 5525 27479 5559
rect 29009 5525 29043 5559
rect 29101 5525 29135 5559
rect 32597 5525 32631 5559
rect 35541 5525 35575 5559
rect 38025 5525 38059 5559
rect 2329 5321 2363 5355
rect 6469 5321 6503 5355
rect 11621 5321 11655 5355
rect 16865 5321 16899 5355
rect 27997 5321 28031 5355
rect 38577 5321 38611 5355
rect 39405 5321 39439 5355
rect 1869 5253 1903 5287
rect 2053 5253 2087 5287
rect 26157 5253 26191 5287
rect 1501 5185 1535 5219
rect 2237 5185 2271 5219
rect 2789 5185 2823 5219
rect 5457 5185 5491 5219
rect 6653 5185 6687 5219
rect 7573 5185 7607 5219
rect 8401 5185 8435 5219
rect 8664 5185 8698 5219
rect 9965 5185 9999 5219
rect 10609 5185 10643 5219
rect 11805 5185 11839 5219
rect 11989 5185 12023 5219
rect 12173 5185 12207 5219
rect 14657 5185 14691 5219
rect 15761 5185 15795 5219
rect 16681 5185 16715 5219
rect 17233 5185 17267 5219
rect 18245 5185 18279 5219
rect 18981 5185 19015 5219
rect 19257 5185 19291 5219
rect 19901 5185 19935 5219
rect 20177 5185 20211 5219
rect 21097 5185 21131 5219
rect 22109 5185 22143 5219
rect 22661 5185 22695 5219
rect 25145 5185 25179 5219
rect 27261 5185 27295 5219
rect 28181 5185 28215 5219
rect 28825 5185 28859 5219
rect 32137 5185 32171 5219
rect 32321 5185 32355 5219
rect 35725 5185 35759 5219
rect 38761 5185 38795 5219
rect 38853 5185 38887 5219
rect 39221 5185 39255 5219
rect 2513 5117 2547 5151
rect 5181 5117 5215 5151
rect 7297 5117 7331 5151
rect 10333 5117 10367 5151
rect 12909 5117 12943 5151
rect 13047 5117 13081 5151
rect 13185 5117 13219 5151
rect 14381 5117 14415 5151
rect 15485 5117 15519 5151
rect 16957 5117 16991 5151
rect 18061 5117 18095 5151
rect 19119 5117 19153 5151
rect 22385 5117 22419 5151
rect 26985 5117 27019 5151
rect 28549 5117 28583 5151
rect 6193 5049 6227 5083
rect 11345 5049 11379 5083
rect 12633 5049 12667 5083
rect 15393 5049 15427 5083
rect 16497 5049 16531 5083
rect 18705 5049 18739 5083
rect 19993 5049 20027 5083
rect 26341 5049 26375 5083
rect 1593 4981 1627 5015
rect 3525 4981 3559 5015
rect 8309 4981 8343 5015
rect 9413 4981 9447 5015
rect 10149 4981 10183 5015
rect 13829 4981 13863 5015
rect 17969 4981 18003 5015
rect 21281 4981 21315 5015
rect 22293 4981 22327 5015
rect 23397 4981 23431 5015
rect 24961 4981 24995 5015
rect 28365 4981 28399 5015
rect 29561 4981 29595 5015
rect 35541 4981 35575 5015
rect 39037 4981 39071 5015
rect 7021 4777 7055 4811
rect 8125 4777 8159 4811
rect 10793 4777 10827 4811
rect 10977 4777 11011 4811
rect 12173 4777 12207 4811
rect 14749 4777 14783 4811
rect 16865 4777 16899 4811
rect 25605 4777 25639 4811
rect 27261 4777 27295 4811
rect 28917 4777 28951 4811
rect 35909 4777 35943 4811
rect 38301 4777 38335 4811
rect 39405 4777 39439 4811
rect 1685 4709 1719 4743
rect 3065 4709 3099 4743
rect 6929 4709 6963 4743
rect 21281 4709 21315 4743
rect 25513 4709 25547 4743
rect 33885 4709 33919 4743
rect 34805 4709 34839 4743
rect 35081 4709 35115 4743
rect 38577 4709 38611 4743
rect 39037 4709 39071 4743
rect 5917 4641 5951 4675
rect 7573 4641 7607 4675
rect 15853 4641 15887 4675
rect 19533 4641 19567 4675
rect 19993 4641 20027 4675
rect 20386 4641 20420 4675
rect 20545 4641 20579 4675
rect 22293 4641 22327 4675
rect 22385 4641 22419 4675
rect 22569 4641 22603 4675
rect 23029 4641 23063 4675
rect 23305 4641 23339 4675
rect 23443 4641 23477 4675
rect 26065 4641 26099 4675
rect 26157 4641 26191 4675
rect 29929 4641 29963 4675
rect 31769 4641 31803 4675
rect 32413 4641 32447 4675
rect 32689 4641 32723 4675
rect 32806 4641 32840 4675
rect 35633 4641 35667 4675
rect 36461 4641 36495 4675
rect 1777 4573 1811 4607
rect 2053 4573 2087 4607
rect 2329 4573 2363 4607
rect 4537 4573 4571 4607
rect 4813 4573 4847 4607
rect 6193 4573 6227 4607
rect 8309 4573 8343 4607
rect 10703 4573 10737 4607
rect 11161 4573 11195 4607
rect 12909 4573 12943 4607
rect 13185 4573 13219 4607
rect 15485 4573 15519 4607
rect 15761 4573 15795 4607
rect 16129 4573 16163 4607
rect 17417 4573 17451 4607
rect 17693 4573 17727 4607
rect 19349 4573 19383 4607
rect 20269 4573 20303 4607
rect 22017 4573 22051 4607
rect 23581 4573 23615 4607
rect 24501 4573 24535 4607
rect 24777 4573 24811 4607
rect 25973 4573 26007 4607
rect 27077 4573 27111 4607
rect 27353 4573 27387 4607
rect 27905 4573 27939 4607
rect 28181 4573 28215 4607
rect 29009 4573 29043 4607
rect 30205 4573 30239 4607
rect 31953 4573 31987 4607
rect 32965 4573 32999 4607
rect 33701 4573 33735 4607
rect 34989 4573 35023 4607
rect 35449 4573 35483 4607
rect 38485 4573 38519 4607
rect 38761 4573 38795 4607
rect 38853 4573 38887 4607
rect 39221 4573 39255 4607
rect 1501 4505 1535 4539
rect 7389 4505 7423 4539
rect 31033 4505 31067 4539
rect 31217 4505 31251 4539
rect 36277 4505 36311 4539
rect 1961 4437 1995 4471
rect 3801 4437 3835 4471
rect 7481 4437 7515 4471
rect 18429 4437 18463 4471
rect 21189 4437 21223 4471
rect 24225 4437 24259 4471
rect 27537 4437 27571 4471
rect 29193 4437 29227 4471
rect 30941 4437 30975 4471
rect 33609 4437 33643 4471
rect 35541 4437 35575 4471
rect 36369 4437 36403 4471
rect 1961 4233 1995 4267
rect 3065 4233 3099 4267
rect 8493 4233 8527 4267
rect 11161 4233 11195 4267
rect 19165 4233 19199 4267
rect 22937 4233 22971 4267
rect 24961 4233 24995 4267
rect 25421 4233 25455 4267
rect 30849 4233 30883 4267
rect 31953 4233 31987 4267
rect 34805 4233 34839 4267
rect 35909 4233 35943 4267
rect 1501 4165 1535 4199
rect 19073 4165 19107 4199
rect 20177 4165 20211 4199
rect 25329 4165 25363 4199
rect 30389 4165 30423 4199
rect 30481 4165 30515 4199
rect 1777 4097 1811 4131
rect 2145 4097 2179 4131
rect 2421 4097 2455 4131
rect 4169 4097 4203 4131
rect 4328 4097 4362 4131
rect 4445 4097 4479 4131
rect 5181 4097 5215 4131
rect 6377 4097 6411 4131
rect 7573 4097 7607 4131
rect 8861 4097 8895 4131
rect 8953 4097 8987 4131
rect 10379 4097 10413 4131
rect 13185 4097 13219 4131
rect 14197 4097 14231 4131
rect 15669 4097 15703 4131
rect 18613 4097 18647 4131
rect 19165 4097 19199 4131
rect 20085 4097 20119 4131
rect 20821 4097 20855 4131
rect 22569 4097 22603 4131
rect 23673 4097 23707 4131
rect 24869 4097 24903 4131
rect 27721 4097 27755 4131
rect 31217 4097 31251 4131
rect 33517 4097 33551 4131
rect 34069 4097 34103 4131
rect 35173 4097 35207 4131
rect 37565 4097 37599 4131
rect 38853 4097 38887 4131
rect 39221 4097 39255 4131
rect 3157 4029 3191 4063
rect 3341 4029 3375 4063
rect 4721 4029 4755 4063
rect 5365 4029 5399 4063
rect 6561 4029 6595 4063
rect 7021 4029 7055 4063
rect 7297 4029 7331 4063
rect 7435 4029 7469 4063
rect 9045 4029 9079 4063
rect 9321 4029 9355 4063
rect 9505 4029 9539 4063
rect 10241 4029 10275 4063
rect 10517 4029 10551 4063
rect 13921 4029 13955 4063
rect 19257 4029 19291 4063
rect 19993 4029 20027 4063
rect 22845 4029 22879 4063
rect 23949 4029 23983 4063
rect 25605 4029 25639 4063
rect 27997 4029 28031 4063
rect 30297 4029 30331 4063
rect 30941 4029 30975 4063
rect 33793 4029 33827 4063
rect 34897 4029 34931 4063
rect 1685 3961 1719 3995
rect 2329 3961 2363 3995
rect 2605 3961 2639 3995
rect 2697 3961 2731 3995
rect 8217 3961 8251 3995
rect 9965 3961 9999 3995
rect 14933 3961 14967 3995
rect 18705 3961 18739 3995
rect 20545 3961 20579 3995
rect 20637 3961 20671 3995
rect 21833 3961 21867 3995
rect 37749 3961 37783 3995
rect 39405 3961 39439 3995
rect 3525 3893 3559 3927
rect 13369 3893 13403 3927
rect 15853 3893 15887 3927
rect 18429 3893 18463 3927
rect 24685 3893 24719 3927
rect 26985 3893 27019 3927
rect 33701 3893 33735 3927
rect 39037 3893 39071 3927
rect 2881 3689 2915 3723
rect 12541 3689 12575 3723
rect 17233 3689 17267 3723
rect 20177 3689 20211 3723
rect 26985 3689 27019 3723
rect 34713 3689 34747 3723
rect 36001 3689 36035 3723
rect 39405 3689 39439 3723
rect 2789 3621 2823 3655
rect 8217 3621 8251 3655
rect 9597 3621 9631 3655
rect 11713 3621 11747 3655
rect 12173 3621 12207 3655
rect 15209 3621 15243 3655
rect 29193 3621 29227 3655
rect 31493 3621 31527 3655
rect 39037 3621 39071 3655
rect 1685 3553 1719 3587
rect 3341 3553 3375 3587
rect 3433 3553 3467 3587
rect 5917 3553 5951 3587
rect 6745 3553 6779 3587
rect 7205 3553 7239 3587
rect 8953 3553 8987 3587
rect 9137 3553 9171 3587
rect 9873 3553 9907 3587
rect 10149 3553 10183 3587
rect 11069 3553 11103 3587
rect 13553 3553 13587 3587
rect 17141 3553 17175 3587
rect 19441 3553 19475 3587
rect 23765 3553 23799 3587
rect 31079 3553 31113 3587
rect 31953 3553 31987 3587
rect 1409 3485 1443 3519
rect 2329 3485 2363 3519
rect 2605 3485 2639 3519
rect 3249 3485 3283 3519
rect 4997 3485 5031 3519
rect 5733 3485 5767 3519
rect 6561 3485 6595 3519
rect 7481 3485 7515 3519
rect 10011 3485 10045 3519
rect 11161 3485 11195 3519
rect 11253 3485 11287 3519
rect 11897 3485 11931 3519
rect 11989 3485 12023 3519
rect 13277 3485 13311 3519
rect 15393 3485 15427 3519
rect 16865 3485 16899 3519
rect 17417 3485 17451 3519
rect 17785 3485 17819 3519
rect 19717 3485 19751 3519
rect 20361 3485 20395 3519
rect 22109 3485 22143 3519
rect 23489 3485 23523 3519
rect 25973 3485 26007 3519
rect 26249 3485 26283 3519
rect 27261 3485 27295 3519
rect 27537 3485 27571 3519
rect 30941 3485 30975 3519
rect 31217 3485 31251 3519
rect 32137 3485 32171 3519
rect 34897 3485 34931 3519
rect 34989 3485 35023 3519
rect 36185 3485 36219 3519
rect 38853 3485 38887 3519
rect 39221 3485 39255 3519
rect 5825 3417 5859 3451
rect 29009 3417 29043 3451
rect 2513 3349 2547 3383
rect 3341 3349 3375 3383
rect 5181 3349 5215 3383
rect 5365 3349 5399 3383
rect 6193 3349 6227 3383
rect 6653 3349 6687 3383
rect 10793 3349 10827 3383
rect 11161 3349 11195 3383
rect 11621 3349 11655 3383
rect 16129 3349 16163 3383
rect 17601 3349 17635 3383
rect 19625 3349 19659 3383
rect 20085 3349 20119 3383
rect 22293 3349 22327 3383
rect 22753 3349 22787 3383
rect 28273 3349 28307 3383
rect 30297 3349 30331 3383
rect 35173 3349 35207 3383
rect 3709 3145 3743 3179
rect 4353 3145 4387 3179
rect 4813 3145 4847 3179
rect 5917 3145 5951 3179
rect 11529 3145 11563 3179
rect 11897 3145 11931 3179
rect 17785 3145 17819 3179
rect 18153 3145 18187 3179
rect 20729 3145 20763 3179
rect 23121 3145 23155 3179
rect 25789 3145 25823 3179
rect 26341 3145 26375 3179
rect 27629 3145 27663 3179
rect 30389 3145 30423 3179
rect 31309 3145 31343 3179
rect 34069 3145 34103 3179
rect 38209 3145 38243 3179
rect 39405 3145 39439 3179
rect 11989 3077 12023 3111
rect 2421 3009 2455 3043
rect 2973 3009 3007 3043
rect 3249 3009 3283 3043
rect 3525 3009 3559 3043
rect 3801 3009 3835 3043
rect 4537 3009 4571 3043
rect 4629 3009 4663 3043
rect 5181 3009 5215 3043
rect 6929 3009 6963 3043
rect 9229 3009 9263 3043
rect 9505 3009 9539 3043
rect 10563 3009 10597 3043
rect 10701 3009 10735 3043
rect 13185 3009 13219 3043
rect 13645 3009 13679 3043
rect 14841 3009 14875 3043
rect 16037 3009 16071 3043
rect 16129 3009 16163 3043
rect 16957 3009 16991 3043
rect 19441 3009 19475 3043
rect 19993 3009 20027 3043
rect 22569 3009 22603 3043
rect 22845 3009 22879 3043
rect 22937 3009 22971 3043
rect 25053 3009 25087 3043
rect 25881 3009 25915 3043
rect 26157 3009 26191 3043
rect 27445 3009 27479 3043
rect 29653 3009 29687 3043
rect 30849 3009 30883 3043
rect 31493 3009 31527 3043
rect 33701 3009 33735 3043
rect 33977 3009 34011 3043
rect 34253 3009 34287 3043
rect 38393 3009 38427 3043
rect 38485 3009 38519 3043
rect 38853 3009 38887 3043
rect 39221 3009 39255 3043
rect 1409 2941 1443 2975
rect 1685 2941 1719 2975
rect 3157 2941 3191 2975
rect 4905 2941 4939 2975
rect 6653 2941 6687 2975
rect 9689 2941 9723 2975
rect 10425 2941 10459 2975
rect 12173 2941 12207 2975
rect 13461 2941 13495 2975
rect 14565 2941 14599 2975
rect 16221 2941 16255 2975
rect 16681 2941 16715 2975
rect 18245 2941 18279 2975
rect 18337 2941 18371 2975
rect 19717 2941 19751 2975
rect 24777 2941 24811 2975
rect 29377 2941 29411 2975
rect 30941 2941 30975 2975
rect 31033 2941 31067 2975
rect 3433 2873 3467 2907
rect 7665 2873 7699 2907
rect 10149 2873 10183 2907
rect 12449 2873 12483 2907
rect 13829 2873 13863 2907
rect 15577 2873 15611 2907
rect 15669 2873 15703 2907
rect 17693 2873 17727 2907
rect 26065 2873 26099 2907
rect 2513 2805 2547 2839
rect 3985 2805 4019 2839
rect 4353 2805 4387 2839
rect 9413 2805 9447 2839
rect 11345 2805 11379 2839
rect 19625 2805 19659 2839
rect 21833 2805 21867 2839
rect 30481 2805 30515 2839
rect 32965 2805 32999 2839
rect 38669 2805 38703 2839
rect 39037 2805 39071 2839
rect 5917 2601 5951 2635
rect 10333 2601 10367 2635
rect 11345 2601 11379 2635
rect 12633 2601 12667 2635
rect 17049 2601 17083 2635
rect 23673 2601 23707 2635
rect 31677 2601 31711 2635
rect 33333 2601 33367 2635
rect 39405 2601 39439 2635
rect 23029 2533 23063 2567
rect 23305 2533 23339 2567
rect 23949 2533 23983 2567
rect 39037 2533 39071 2567
rect 2329 2465 2363 2499
rect 2605 2465 2639 2499
rect 4813 2465 4847 2499
rect 4905 2465 4939 2499
rect 7389 2465 7423 2499
rect 10793 2465 10827 2499
rect 17509 2465 17543 2499
rect 17693 2465 17727 2499
rect 20361 2465 20395 2499
rect 22017 2465 22051 2499
rect 31125 2465 31159 2499
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 3433 2397 3467 2431
rect 4537 2397 4571 2431
rect 5181 2397 5215 2431
rect 6009 2397 6043 2431
rect 6837 2397 6871 2431
rect 7205 2397 7239 2431
rect 7481 2397 7515 2431
rect 8033 2397 8067 2431
rect 9505 2397 9539 2431
rect 10057 2397 10091 2431
rect 10517 2397 10551 2431
rect 10977 2397 11011 2431
rect 12449 2397 12483 2431
rect 13461 2397 13495 2431
rect 14105 2397 14139 2431
rect 14933 2397 14967 2431
rect 15669 2397 15703 2431
rect 16129 2397 16163 2431
rect 16681 2397 16715 2431
rect 18153 2397 18187 2431
rect 18337 2397 18371 2431
rect 19073 2397 19107 2431
rect 20085 2397 20119 2431
rect 20821 2397 20855 2431
rect 20913 2397 20947 2431
rect 21557 2397 21591 2431
rect 22293 2397 22327 2431
rect 23121 2397 23155 2431
rect 23489 2397 23523 2431
rect 24133 2397 24167 2431
rect 24409 2397 24443 2431
rect 30481 2397 30515 2431
rect 37749 2397 37783 2431
rect 38117 2397 38151 2431
rect 38485 2397 38519 2431
rect 38853 2397 38887 2431
rect 39221 2397 39255 2431
rect 6469 2329 6503 2363
rect 6653 2329 6687 2363
rect 7021 2329 7055 2363
rect 9045 2329 9079 2363
rect 9229 2329 9263 2363
rect 11805 2329 11839 2363
rect 11989 2329 12023 2363
rect 33241 2329 33275 2363
rect 3525 2261 3559 2295
rect 6193 2261 6227 2295
rect 7665 2261 7699 2295
rect 8217 2261 8251 2295
rect 9689 2261 9723 2295
rect 10241 2261 10275 2295
rect 10885 2261 10919 2295
rect 13277 2261 13311 2295
rect 14289 2261 14323 2295
rect 14749 2261 14783 2295
rect 15485 2261 15519 2295
rect 16313 2261 16347 2295
rect 16865 2261 16899 2295
rect 17417 2261 17451 2295
rect 17969 2261 18003 2295
rect 18521 2261 18555 2295
rect 18889 2261 18923 2295
rect 19349 2261 19383 2295
rect 20637 2261 20671 2295
rect 21097 2261 21131 2295
rect 21373 2261 21407 2295
rect 24593 2261 24627 2295
rect 30297 2261 30331 2295
rect 31217 2261 31251 2295
rect 31309 2261 31343 2295
rect 37933 2261 37967 2295
rect 38301 2261 38335 2295
rect 38669 2261 38703 2295
<< metal1 >>
rect 10594 10820 10600 10872
rect 10652 10860 10658 10872
rect 17218 10860 17224 10872
rect 10652 10832 17224 10860
rect 10652 10820 10658 10832
rect 17218 10820 17224 10832
rect 17276 10820 17282 10872
rect 10778 10684 10784 10736
rect 10836 10724 10842 10736
rect 17402 10724 17408 10736
rect 10836 10696 17408 10724
rect 10836 10684 10842 10696
rect 17402 10684 17408 10696
rect 17460 10684 17466 10736
rect 8570 10412 8576 10464
rect 8628 10452 8634 10464
rect 36446 10452 36452 10464
rect 8628 10424 36452 10452
rect 8628 10412 8634 10424
rect 36446 10412 36452 10424
rect 36504 10412 36510 10464
rect 4246 10344 4252 10396
rect 4304 10384 4310 10396
rect 29822 10384 29828 10396
rect 4304 10356 29828 10384
rect 4304 10344 4310 10356
rect 29822 10344 29828 10356
rect 29880 10344 29886 10396
rect 17218 10276 17224 10328
rect 17276 10316 17282 10328
rect 17276 10288 31754 10316
rect 17276 10276 17282 10288
rect 4154 10208 4160 10260
rect 4212 10248 4218 10260
rect 25222 10248 25228 10260
rect 4212 10220 25228 10248
rect 4212 10208 4218 10220
rect 25222 10208 25228 10220
rect 25280 10208 25286 10260
rect 25590 10208 25596 10260
rect 25648 10248 25654 10260
rect 26510 10248 26516 10260
rect 25648 10220 26516 10248
rect 25648 10208 25654 10220
rect 26510 10208 26516 10220
rect 26568 10208 26574 10260
rect 31726 10248 31754 10288
rect 37642 10248 37648 10260
rect 31726 10220 37648 10248
rect 37642 10208 37648 10220
rect 37700 10208 37706 10260
rect 11882 10140 11888 10192
rect 11940 10180 11946 10192
rect 28994 10180 29000 10192
rect 11940 10152 29000 10180
rect 11940 10140 11946 10152
rect 28994 10140 29000 10152
rect 29052 10140 29058 10192
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 17218 10112 17224 10124
rect 6972 10084 17224 10112
rect 6972 10072 6978 10084
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 17402 10072 17408 10124
rect 17460 10112 17466 10124
rect 30374 10112 30380 10124
rect 17460 10084 30380 10112
rect 17460 10072 17466 10084
rect 30374 10072 30380 10084
rect 30432 10072 30438 10124
rect 8662 10004 8668 10056
rect 8720 10044 8726 10056
rect 30742 10044 30748 10056
rect 8720 10016 30748 10044
rect 8720 10004 8726 10016
rect 30742 10004 30748 10016
rect 30800 10004 30806 10056
rect 2590 9936 2596 9988
rect 2648 9976 2654 9988
rect 24578 9976 24584 9988
rect 2648 9948 24584 9976
rect 2648 9936 2654 9948
rect 24578 9936 24584 9948
rect 24636 9936 24642 9988
rect 14734 9868 14740 9920
rect 14792 9908 14798 9920
rect 15102 9908 15108 9920
rect 14792 9880 15108 9908
rect 14792 9868 14798 9880
rect 15102 9868 15108 9880
rect 15160 9868 15166 9920
rect 17218 9868 17224 9920
rect 17276 9908 17282 9920
rect 31478 9908 31484 9920
rect 17276 9880 31484 9908
rect 17276 9868 17282 9880
rect 31478 9868 31484 9880
rect 31536 9868 31542 9920
rect 9950 9800 9956 9852
rect 10008 9840 10014 9852
rect 29546 9840 29552 9852
rect 10008 9812 29552 9840
rect 10008 9800 10014 9812
rect 29546 9800 29552 9812
rect 29604 9800 29610 9852
rect 10870 9732 10876 9784
rect 10928 9772 10934 9784
rect 11790 9772 11796 9784
rect 10928 9744 11796 9772
rect 10928 9732 10934 9744
rect 11790 9732 11796 9744
rect 11848 9732 11854 9784
rect 12158 9732 12164 9784
rect 12216 9772 12222 9784
rect 13078 9772 13084 9784
rect 12216 9744 13084 9772
rect 12216 9732 12222 9744
rect 13078 9732 13084 9744
rect 13136 9732 13142 9784
rect 14458 9732 14464 9784
rect 14516 9772 14522 9784
rect 21542 9772 21548 9784
rect 14516 9744 21548 9772
rect 14516 9732 14522 9744
rect 21542 9732 21548 9744
rect 21600 9732 21606 9784
rect 25866 9732 25872 9784
rect 25924 9772 25930 9784
rect 27430 9772 27436 9784
rect 25924 9744 27436 9772
rect 25924 9732 25930 9744
rect 27430 9732 27436 9744
rect 27488 9732 27494 9784
rect 10042 9664 10048 9716
rect 10100 9704 10106 9716
rect 11238 9704 11244 9716
rect 10100 9676 11244 9704
rect 10100 9664 10106 9676
rect 11238 9664 11244 9676
rect 11296 9664 11302 9716
rect 11698 9664 11704 9716
rect 11756 9704 11762 9716
rect 12894 9704 12900 9716
rect 11756 9676 12900 9704
rect 11756 9664 11762 9676
rect 12894 9664 12900 9676
rect 12952 9664 12958 9716
rect 19426 9704 19432 9716
rect 13004 9676 19432 9704
rect 13004 9648 13032 9676
rect 19426 9664 19432 9676
rect 19484 9664 19490 9716
rect 20346 9664 20352 9716
rect 20404 9704 20410 9716
rect 20806 9704 20812 9716
rect 20404 9676 20812 9704
rect 20404 9664 20410 9676
rect 20806 9664 20812 9676
rect 20864 9664 20870 9716
rect 31754 9664 31760 9716
rect 31812 9664 31818 9716
rect 4522 9596 4528 9648
rect 4580 9636 4586 9648
rect 12434 9636 12440 9648
rect 4580 9608 12440 9636
rect 4580 9596 4586 9608
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 12986 9596 12992 9648
rect 13044 9596 13050 9648
rect 15562 9596 15568 9648
rect 15620 9636 15626 9648
rect 15620 9608 22094 9636
rect 15620 9596 15626 9608
rect 5258 9528 5264 9580
rect 5316 9568 5322 9580
rect 12250 9568 12256 9580
rect 5316 9540 12256 9568
rect 5316 9528 5322 9540
rect 12250 9528 12256 9540
rect 12308 9528 12314 9580
rect 13078 9528 13084 9580
rect 13136 9568 13142 9580
rect 16574 9568 16580 9580
rect 13136 9540 16580 9568
rect 13136 9528 13142 9540
rect 16574 9528 16580 9540
rect 16632 9528 16638 9580
rect 17034 9528 17040 9580
rect 17092 9568 17098 9580
rect 19702 9568 19708 9580
rect 17092 9540 19708 9568
rect 17092 9528 17098 9540
rect 19702 9528 19708 9540
rect 19760 9528 19766 9580
rect 22066 9568 22094 9608
rect 28074 9596 28080 9648
rect 28132 9636 28138 9648
rect 28902 9636 28908 9648
rect 28132 9608 28908 9636
rect 28132 9596 28138 9608
rect 28902 9596 28908 9608
rect 28960 9596 28966 9648
rect 30006 9596 30012 9648
rect 30064 9636 30070 9648
rect 31570 9636 31576 9648
rect 30064 9608 31576 9636
rect 30064 9596 30070 9608
rect 31570 9596 31576 9608
rect 31628 9596 31634 9648
rect 28718 9568 28724 9580
rect 22066 9540 28724 9568
rect 28718 9528 28724 9540
rect 28776 9528 28782 9580
rect 31772 9512 31800 9664
rect 31846 9596 31852 9648
rect 31904 9636 31910 9648
rect 32674 9636 32680 9648
rect 31904 9608 32680 9636
rect 31904 9596 31910 9608
rect 32674 9596 32680 9608
rect 32732 9596 32738 9648
rect 7282 9460 7288 9512
rect 7340 9500 7346 9512
rect 7926 9500 7932 9512
rect 7340 9472 7932 9500
rect 7340 9460 7346 9472
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 28442 9500 28448 9512
rect 15488 9472 28448 9500
rect 6362 9392 6368 9444
rect 6420 9432 6426 9444
rect 14090 9432 14096 9444
rect 6420 9404 14096 9432
rect 6420 9392 6426 9404
rect 14090 9392 14096 9404
rect 14148 9392 14154 9444
rect 5626 9324 5632 9376
rect 5684 9364 5690 9376
rect 11606 9364 11612 9376
rect 5684 9336 11612 9364
rect 5684 9324 5690 9336
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 12710 9324 12716 9376
rect 12768 9364 12774 9376
rect 15488 9364 15516 9472
rect 28442 9460 28448 9472
rect 28500 9460 28506 9512
rect 31754 9460 31760 9512
rect 31812 9460 31818 9512
rect 18046 9392 18052 9444
rect 18104 9432 18110 9444
rect 18104 9404 28994 9432
rect 18104 9392 18110 9404
rect 12768 9336 15516 9364
rect 12768 9324 12774 9336
rect 16942 9324 16948 9376
rect 17000 9364 17006 9376
rect 26694 9364 26700 9376
rect 17000 9336 26700 9364
rect 17000 9324 17006 9336
rect 26694 9324 26700 9336
rect 26752 9324 26758 9376
rect 28966 9364 28994 9404
rect 31938 9364 31944 9376
rect 28966 9336 31944 9364
rect 31938 9324 31944 9336
rect 31996 9324 32002 9376
rect 2682 9256 2688 9308
rect 2740 9296 2746 9308
rect 10318 9296 10324 9308
rect 2740 9268 10324 9296
rect 2740 9256 2746 9268
rect 10318 9256 10324 9268
rect 10376 9256 10382 9308
rect 11330 9256 11336 9308
rect 11388 9296 11394 9308
rect 22186 9296 22192 9308
rect 11388 9268 22192 9296
rect 11388 9256 11394 9268
rect 22186 9256 22192 9268
rect 22244 9256 22250 9308
rect 24854 9256 24860 9308
rect 24912 9296 24918 9308
rect 32858 9296 32864 9308
rect 24912 9268 32864 9296
rect 24912 9256 24918 9268
rect 32858 9256 32864 9268
rect 32916 9256 32922 9308
rect 1670 9188 1676 9240
rect 1728 9228 1734 9240
rect 9674 9228 9680 9240
rect 1728 9200 9680 9228
rect 1728 9188 1734 9200
rect 9674 9188 9680 9200
rect 9732 9188 9738 9240
rect 11422 9188 11428 9240
rect 11480 9228 11486 9240
rect 11480 9200 13032 9228
rect 11480 9188 11486 9200
rect 3602 9120 3608 9172
rect 3660 9160 3666 9172
rect 8478 9160 8484 9172
rect 3660 9132 8484 9160
rect 3660 9120 3666 9132
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 13004 9160 13032 9200
rect 13354 9188 13360 9240
rect 13412 9228 13418 9240
rect 19610 9228 19616 9240
rect 13412 9200 19616 9228
rect 13412 9188 13418 9200
rect 19610 9188 19616 9200
rect 19668 9188 19674 9240
rect 19702 9188 19708 9240
rect 19760 9228 19766 9240
rect 31018 9228 31024 9240
rect 19760 9200 31024 9228
rect 19760 9188 19766 9200
rect 31018 9188 31024 9200
rect 31076 9188 31082 9240
rect 25774 9160 25780 9172
rect 9646 9132 12940 9160
rect 13004 9132 25780 9160
rect 5350 9052 5356 9104
rect 5408 9092 5414 9104
rect 9646 9092 9674 9132
rect 5408 9064 9674 9092
rect 5408 9052 5414 9064
rect 9766 9052 9772 9104
rect 9824 9092 9830 9104
rect 10134 9092 10140 9104
rect 9824 9064 10140 9092
rect 9824 9052 9830 9064
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 11238 9052 11244 9104
rect 11296 9092 11302 9104
rect 12912 9092 12940 9132
rect 25774 9120 25780 9132
rect 25832 9120 25838 9172
rect 25866 9120 25872 9172
rect 25924 9160 25930 9172
rect 28074 9160 28080 9172
rect 25924 9132 28080 9160
rect 25924 9120 25930 9132
rect 28074 9120 28080 9132
rect 28132 9120 28138 9172
rect 32398 9160 32404 9172
rect 31726 9132 32404 9160
rect 14642 9092 14648 9104
rect 11296 9064 12848 9092
rect 12912 9064 14648 9092
rect 11296 9052 11302 9064
rect 10226 8984 10232 9036
rect 10284 9024 10290 9036
rect 12710 9024 12716 9036
rect 10284 8996 12716 9024
rect 10284 8984 10290 8996
rect 12710 8984 12716 8996
rect 12768 8984 12774 9036
rect 12820 9024 12848 9064
rect 14642 9052 14648 9064
rect 14700 9052 14706 9104
rect 17862 9052 17868 9104
rect 17920 9092 17926 9104
rect 18506 9092 18512 9104
rect 17920 9064 18512 9092
rect 17920 9052 17926 9064
rect 18506 9052 18512 9064
rect 18564 9052 18570 9104
rect 18782 9052 18788 9104
rect 18840 9092 18846 9104
rect 22646 9092 22652 9104
rect 18840 9064 22652 9092
rect 18840 9052 18846 9064
rect 22646 9052 22652 9064
rect 22704 9052 22710 9104
rect 30282 9092 30288 9104
rect 22756 9064 30288 9092
rect 16022 9024 16028 9036
rect 12820 8996 16028 9024
rect 16022 8984 16028 8996
rect 16080 8984 16086 9036
rect 16298 8984 16304 9036
rect 16356 9024 16362 9036
rect 21910 9024 21916 9036
rect 16356 8996 21916 9024
rect 16356 8984 16362 8996
rect 21910 8984 21916 8996
rect 21968 8984 21974 9036
rect 22094 8984 22100 9036
rect 22152 9024 22158 9036
rect 22756 9024 22784 9064
rect 30282 9052 30288 9064
rect 30340 9052 30346 9104
rect 22152 8996 22784 9024
rect 22152 8984 22158 8996
rect 23198 8984 23204 9036
rect 23256 9024 23262 9036
rect 30466 9024 30472 9036
rect 23256 8996 30472 9024
rect 23256 8984 23262 8996
rect 30466 8984 30472 8996
rect 30524 8984 30530 9036
rect 7006 8916 7012 8968
rect 7064 8956 7070 8968
rect 15470 8956 15476 8968
rect 7064 8928 15476 8956
rect 7064 8916 7070 8928
rect 15470 8916 15476 8928
rect 15528 8916 15534 8968
rect 19518 8916 19524 8968
rect 19576 8956 19582 8968
rect 23216 8956 23244 8984
rect 31726 8956 31754 9132
rect 32398 9120 32404 9132
rect 32456 9120 32462 9172
rect 19576 8928 23244 8956
rect 26896 8928 31754 8956
rect 19576 8916 19582 8928
rect 5902 8848 5908 8900
rect 5960 8888 5966 8900
rect 10502 8888 10508 8900
rect 5960 8860 10508 8888
rect 5960 8848 5966 8860
rect 10502 8848 10508 8860
rect 10560 8848 10566 8900
rect 11790 8848 11796 8900
rect 11848 8888 11854 8900
rect 13538 8888 13544 8900
rect 11848 8860 13544 8888
rect 11848 8848 11854 8860
rect 13538 8848 13544 8860
rect 13596 8848 13602 8900
rect 13814 8848 13820 8900
rect 13872 8888 13878 8900
rect 26896 8888 26924 8928
rect 35342 8916 35348 8968
rect 35400 8956 35406 8968
rect 36538 8956 36544 8968
rect 35400 8928 36544 8956
rect 35400 8916 35406 8928
rect 36538 8916 36544 8928
rect 36596 8916 36602 8968
rect 13872 8860 26924 8888
rect 13872 8848 13878 8860
rect 30374 8848 30380 8900
rect 30432 8888 30438 8900
rect 38930 8888 38936 8900
rect 30432 8860 38936 8888
rect 30432 8848 30438 8860
rect 38930 8848 38936 8860
rect 38988 8848 38994 8900
rect 5810 8780 5816 8832
rect 5868 8820 5874 8832
rect 12986 8820 12992 8832
rect 5868 8792 12992 8820
rect 5868 8780 5874 8792
rect 12986 8780 12992 8792
rect 13044 8780 13050 8832
rect 13262 8780 13268 8832
rect 13320 8820 13326 8832
rect 19334 8820 19340 8832
rect 13320 8792 19340 8820
rect 13320 8780 13326 8792
rect 19334 8780 19340 8792
rect 19392 8780 19398 8832
rect 21910 8780 21916 8832
rect 21968 8820 21974 8832
rect 26602 8820 26608 8832
rect 21968 8792 26608 8820
rect 21968 8780 21974 8792
rect 26602 8780 26608 8792
rect 26660 8780 26666 8832
rect 26970 8780 26976 8832
rect 27028 8820 27034 8832
rect 28258 8820 28264 8832
rect 27028 8792 28264 8820
rect 27028 8780 27034 8792
rect 28258 8780 28264 8792
rect 28316 8780 28322 8832
rect 28626 8780 28632 8832
rect 28684 8820 28690 8832
rect 30650 8820 30656 8832
rect 28684 8792 30656 8820
rect 28684 8780 28690 8792
rect 30650 8780 30656 8792
rect 30708 8780 30714 8832
rect 33042 8780 33048 8832
rect 33100 8820 33106 8832
rect 33778 8820 33784 8832
rect 33100 8792 33784 8820
rect 33100 8780 33106 8792
rect 33778 8780 33784 8792
rect 33836 8780 33842 8832
rect 33870 8780 33876 8832
rect 33928 8820 33934 8832
rect 34330 8820 34336 8832
rect 33928 8792 34336 8820
rect 33928 8780 33934 8792
rect 34330 8780 34336 8792
rect 34388 8780 34394 8832
rect 34514 8780 34520 8832
rect 34572 8820 34578 8832
rect 36998 8820 37004 8832
rect 34572 8792 37004 8820
rect 34572 8780 34578 8792
rect 36998 8780 37004 8792
rect 37056 8780 37062 8832
rect 1104 8730 39836 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 39010 8730
rect 39062 8678 39074 8730
rect 39126 8678 39138 8730
rect 39190 8678 39202 8730
rect 39254 8678 39266 8730
rect 39318 8678 39836 8730
rect 1104 8656 39836 8678
rect 3421 8619 3479 8625
rect 3421 8585 3433 8619
rect 3467 8616 3479 8619
rect 3786 8616 3792 8628
rect 3467 8588 3792 8616
rect 3467 8585 3479 8588
rect 3421 8579 3479 8585
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 4157 8619 4215 8625
rect 4157 8585 4169 8619
rect 4203 8616 4215 8619
rect 4338 8616 4344 8628
rect 4203 8588 4344 8616
rect 4203 8585 4215 8588
rect 4157 8579 4215 8585
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 4525 8619 4583 8625
rect 4525 8585 4537 8619
rect 4571 8616 4583 8619
rect 4890 8616 4896 8628
rect 4571 8588 4896 8616
rect 4571 8585 4583 8588
rect 4525 8579 4583 8585
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 5261 8619 5319 8625
rect 5261 8585 5273 8619
rect 5307 8585 5319 8619
rect 5261 8579 5319 8585
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8616 5687 8619
rect 6270 8616 6276 8628
rect 5675 8588 6276 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 1302 8508 1308 8560
rect 1360 8548 1366 8560
rect 5276 8548 5304 8579
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 6457 8619 6515 8625
rect 6457 8585 6469 8619
rect 6503 8585 6515 8619
rect 6457 8579 6515 8585
rect 5994 8548 6000 8560
rect 1360 8520 3832 8548
rect 5276 8520 6000 8548
rect 1360 8508 1366 8520
rect 474 8440 480 8492
rect 532 8480 538 8492
rect 2317 8483 2375 8489
rect 2317 8480 2329 8483
rect 532 8452 2329 8480
rect 532 8440 538 8452
rect 2317 8449 2329 8452
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 3602 8440 3608 8492
rect 3660 8440 3666 8492
rect 3804 8489 3832 8520
rect 5994 8508 6000 8520
rect 6052 8508 6058 8560
rect 6472 8548 6500 8579
rect 6638 8576 6644 8628
rect 6696 8616 6702 8628
rect 6825 8619 6883 8625
rect 6825 8616 6837 8619
rect 6696 8588 6837 8616
rect 6696 8576 6702 8588
rect 6825 8585 6837 8588
rect 6871 8585 6883 8619
rect 6825 8579 6883 8585
rect 7193 8619 7251 8625
rect 7193 8585 7205 8619
rect 7239 8616 7251 8619
rect 8846 8616 8852 8628
rect 7239 8588 8852 8616
rect 7239 8585 7251 8588
rect 7193 8579 7251 8585
rect 8846 8576 8852 8588
rect 8904 8576 8910 8628
rect 9309 8619 9367 8625
rect 9309 8585 9321 8619
rect 9355 8616 9367 8619
rect 9674 8616 9680 8628
rect 9355 8588 9680 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 9950 8616 9956 8628
rect 9784 8588 9956 8616
rect 7282 8548 7288 8560
rect 6472 8520 7288 8548
rect 7282 8508 7288 8520
rect 7340 8508 7346 8560
rect 8478 8508 8484 8560
rect 8536 8548 8542 8560
rect 8536 8520 9674 8548
rect 8536 8508 8542 8520
rect 9646 8492 9674 8520
rect 3789 8483 3847 8489
rect 3789 8449 3801 8483
rect 3835 8449 3847 8483
rect 3789 8443 3847 8449
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 4522 8480 4528 8492
rect 4387 8452 4528 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 4706 8440 4712 8492
rect 4764 8440 4770 8492
rect 5074 8440 5080 8492
rect 5132 8440 5138 8492
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8480 5503 8483
rect 5626 8480 5632 8492
rect 5491 8452 5632 8480
rect 5491 8449 5503 8452
rect 5445 8443 5503 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5810 8440 5816 8492
rect 5868 8440 5874 8492
rect 6178 8440 6184 8492
rect 6236 8440 6242 8492
rect 6638 8440 6644 8492
rect 6696 8440 6702 8492
rect 7006 8440 7012 8492
rect 7064 8440 7070 8492
rect 7374 8440 7380 8492
rect 7432 8440 7438 8492
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8480 7803 8483
rect 7834 8480 7840 8492
rect 7791 8452 7840 8480
rect 7791 8449 7803 8452
rect 7745 8443 7803 8449
rect 7834 8440 7840 8452
rect 7892 8480 7898 8492
rect 9214 8480 9220 8492
rect 7892 8452 9220 8480
rect 7892 8440 7898 8452
rect 9214 8440 9220 8452
rect 9272 8440 9278 8492
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 9646 8452 9680 8492
rect 9674 8440 9680 8452
rect 9732 8440 9738 8492
rect 750 8372 756 8424
rect 808 8412 814 8424
rect 1397 8415 1455 8421
rect 1397 8412 1409 8415
rect 808 8384 1409 8412
rect 808 8372 814 8384
rect 1397 8381 1409 8384
rect 1443 8381 1455 8415
rect 1397 8375 1455 8381
rect 1670 8372 1676 8424
rect 1728 8372 1734 8424
rect 2593 8415 2651 8421
rect 2593 8381 2605 8415
rect 2639 8412 2651 8415
rect 4798 8412 4804 8424
rect 2639 8384 4804 8412
rect 2639 8381 2651 8384
rect 2593 8375 2651 8381
rect 4798 8372 4804 8384
rect 4856 8372 4862 8424
rect 6822 8412 6828 8424
rect 6012 8384 6828 8412
rect 3786 8304 3792 8356
rect 3844 8344 3850 8356
rect 3973 8347 4031 8353
rect 3973 8344 3985 8347
rect 3844 8316 3985 8344
rect 3844 8304 3850 8316
rect 3973 8313 3985 8316
rect 4019 8313 4031 8347
rect 3973 8307 4031 8313
rect 4893 8347 4951 8353
rect 4893 8313 4905 8347
rect 4939 8344 4951 8347
rect 5442 8344 5448 8356
rect 4939 8316 5448 8344
rect 4939 8313 4951 8316
rect 4893 8307 4951 8313
rect 5442 8304 5448 8316
rect 5500 8304 5506 8356
rect 6012 8353 6040 8384
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 7190 8372 7196 8424
rect 7248 8412 7254 8424
rect 7469 8415 7527 8421
rect 7469 8412 7481 8415
rect 7248 8384 7481 8412
rect 7248 8372 7254 8384
rect 7469 8381 7481 8384
rect 7515 8381 7527 8415
rect 9784 8412 9812 8588
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 10042 8576 10048 8628
rect 10100 8576 10106 8628
rect 10870 8576 10876 8628
rect 10928 8576 10934 8628
rect 11149 8619 11207 8625
rect 11149 8585 11161 8619
rect 11195 8616 11207 8619
rect 12066 8616 12072 8628
rect 11195 8588 12072 8616
rect 11195 8585 11207 8588
rect 11149 8579 11207 8585
rect 12066 8576 12072 8588
rect 12124 8576 12130 8628
rect 12158 8576 12164 8628
rect 12216 8576 12222 8628
rect 12802 8576 12808 8628
rect 12860 8576 12866 8628
rect 13170 8576 13176 8628
rect 13228 8576 13234 8628
rect 13817 8619 13875 8625
rect 13817 8585 13829 8619
rect 13863 8616 13875 8619
rect 14550 8616 14556 8628
rect 13863 8588 14556 8616
rect 13863 8585 13875 8588
rect 13817 8579 13875 8585
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 14642 8576 14648 8628
rect 14700 8616 14706 8628
rect 14700 8588 14872 8616
rect 14700 8576 14706 8588
rect 11238 8548 11244 8560
rect 10060 8520 11244 8548
rect 9861 8483 9919 8489
rect 9861 8449 9873 8483
rect 9907 8480 9919 8483
rect 10060 8480 10088 8520
rect 11238 8508 11244 8520
rect 11296 8508 11302 8560
rect 13078 8548 13084 8560
rect 11900 8520 13084 8548
rect 9907 8452 10088 8480
rect 9907 8449 9919 8452
rect 9861 8443 9919 8449
rect 10226 8440 10232 8492
rect 10284 8440 10290 8492
rect 10318 8440 10324 8492
rect 10376 8440 10382 8492
rect 10502 8440 10508 8492
rect 10560 8480 10566 8492
rect 10689 8484 10747 8489
rect 10612 8483 10747 8484
rect 10612 8480 10701 8483
rect 10560 8456 10701 8480
rect 10560 8452 10640 8456
rect 10560 8440 10566 8452
rect 10689 8449 10701 8456
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 11330 8440 11336 8492
rect 11388 8440 11394 8492
rect 11900 8489 11928 8520
rect 13078 8508 13084 8520
rect 13136 8508 13142 8560
rect 13538 8508 13544 8560
rect 13596 8548 13602 8560
rect 14844 8548 14872 8588
rect 14918 8576 14924 8628
rect 14976 8576 14982 8628
rect 15289 8619 15347 8625
rect 15289 8585 15301 8619
rect 15335 8616 15347 8619
rect 16206 8616 16212 8628
rect 15335 8588 16212 8616
rect 15335 8585 15347 8588
rect 15289 8579 15347 8585
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 16390 8576 16396 8628
rect 16448 8576 16454 8628
rect 17037 8619 17095 8625
rect 17037 8585 17049 8619
rect 17083 8616 17095 8619
rect 17310 8616 17316 8628
rect 17083 8588 17316 8616
rect 17083 8585 17095 8588
rect 17037 8579 17095 8585
rect 17310 8576 17316 8588
rect 17368 8576 17374 8628
rect 17678 8576 17684 8628
rect 17736 8616 17742 8628
rect 18831 8619 18889 8625
rect 18831 8616 18843 8619
rect 17736 8588 18843 8616
rect 17736 8576 17742 8588
rect 18831 8585 18843 8588
rect 18877 8616 18889 8619
rect 18877 8588 19334 8616
rect 18877 8585 18889 8588
rect 18831 8579 18889 8585
rect 13596 8520 14780 8548
rect 14844 8520 15148 8548
rect 13596 8508 13602 8520
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8449 11943 8483
rect 11885 8443 11943 8449
rect 11977 8483 12035 8489
rect 11977 8449 11989 8483
rect 12023 8449 12035 8483
rect 11977 8443 12035 8449
rect 7469 8375 7527 8381
rect 9600 8384 9812 8412
rect 5997 8347 6055 8353
rect 5997 8313 6009 8347
rect 6043 8313 6055 8347
rect 5997 8307 6055 8313
rect 7466 8236 7472 8288
rect 7524 8276 7530 8288
rect 8202 8276 8208 8288
rect 7524 8248 8208 8276
rect 7524 8236 7530 8248
rect 8202 8236 8208 8248
rect 8260 8236 8266 8288
rect 8478 8236 8484 8288
rect 8536 8236 8542 8288
rect 8938 8236 8944 8288
rect 8996 8276 9002 8288
rect 9600 8276 9628 8384
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 11992 8412 12020 8443
rect 12250 8440 12256 8492
rect 12308 8480 12314 8492
rect 12345 8483 12403 8489
rect 12345 8480 12357 8483
rect 12308 8452 12357 8480
rect 12308 8440 12314 8452
rect 12345 8449 12357 8452
rect 12391 8449 12403 8483
rect 12345 8443 12403 8449
rect 12989 8483 13047 8489
rect 12989 8449 13001 8483
rect 13035 8480 13047 8483
rect 13262 8480 13268 8492
rect 13035 8452 13268 8480
rect 13035 8449 13047 8452
rect 12989 8443 13047 8449
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 13354 8440 13360 8492
rect 13412 8440 13418 8492
rect 13449 8483 13507 8489
rect 13449 8449 13461 8483
rect 13495 8480 13507 8483
rect 13630 8480 13636 8492
rect 13495 8452 13636 8480
rect 13495 8449 13507 8452
rect 13449 8443 13507 8449
rect 13630 8440 13636 8452
rect 13688 8440 13694 8492
rect 14274 8440 14280 8492
rect 14332 8440 14338 8492
rect 14752 8489 14780 8520
rect 15120 8489 15148 8520
rect 15838 8508 15844 8560
rect 15896 8548 15902 8560
rect 15896 8520 16252 8548
rect 15896 8508 15902 8520
rect 14645 8483 14703 8489
rect 14645 8449 14657 8483
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 14737 8483 14795 8489
rect 14737 8449 14749 8483
rect 14783 8449 14795 8483
rect 14737 8443 14795 8449
rect 15105 8483 15163 8489
rect 15105 8449 15117 8483
rect 15151 8449 15163 8483
rect 15105 8443 15163 8449
rect 11296 8384 12020 8412
rect 11296 8372 11302 8384
rect 12434 8372 12440 8424
rect 12492 8412 12498 8424
rect 13170 8412 13176 8424
rect 12492 8384 13176 8412
rect 12492 8372 12498 8384
rect 13170 8372 13176 8384
rect 13228 8372 13234 8424
rect 13538 8372 13544 8424
rect 13596 8412 13602 8424
rect 14366 8412 14372 8424
rect 13596 8384 14372 8412
rect 13596 8372 13602 8384
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 14660 8412 14688 8443
rect 15746 8440 15752 8492
rect 15804 8440 15810 8492
rect 16114 8440 16120 8492
rect 16172 8440 16178 8492
rect 16224 8489 16252 8520
rect 17494 8508 17500 8560
rect 17552 8548 17558 8560
rect 19306 8548 19334 8588
rect 19702 8576 19708 8628
rect 19760 8616 19766 8628
rect 21174 8616 21180 8628
rect 19760 8588 21180 8616
rect 19760 8576 19766 8588
rect 21174 8576 21180 8588
rect 21232 8576 21238 8628
rect 21269 8619 21327 8625
rect 21269 8585 21281 8619
rect 21315 8616 21327 8619
rect 21542 8616 21548 8628
rect 21315 8588 21548 8616
rect 21315 8585 21327 8588
rect 21269 8579 21327 8585
rect 21542 8576 21548 8588
rect 21600 8576 21606 8628
rect 22002 8576 22008 8628
rect 22060 8616 22066 8628
rect 22060 8588 22416 8616
rect 22060 8576 22066 8588
rect 21634 8548 21640 8560
rect 17552 8520 17908 8548
rect 19306 8520 21640 8548
rect 17552 8508 17558 8520
rect 16209 8483 16267 8489
rect 16209 8449 16221 8483
rect 16255 8449 16267 8483
rect 16209 8443 16267 8449
rect 17221 8483 17279 8489
rect 17221 8449 17233 8483
rect 17267 8480 17279 8483
rect 17770 8480 17776 8492
rect 17267 8452 17776 8480
rect 17267 8449 17279 8452
rect 17221 8443 17279 8449
rect 17770 8440 17776 8452
rect 17828 8440 17834 8492
rect 17880 8489 17908 8520
rect 21634 8508 21640 8520
rect 21692 8508 21698 8560
rect 21726 8508 21732 8560
rect 21784 8548 21790 8560
rect 21784 8520 22140 8548
rect 21784 8508 21790 8520
rect 17865 8483 17923 8489
rect 17865 8449 17877 8483
rect 17911 8449 17923 8483
rect 17865 8443 17923 8449
rect 18138 8440 18144 8492
rect 18196 8440 18202 8492
rect 18690 8440 18696 8492
rect 18748 8480 18754 8492
rect 19061 8483 19119 8489
rect 19061 8480 19073 8483
rect 18748 8452 19073 8480
rect 18748 8440 18754 8452
rect 19061 8449 19073 8452
rect 19107 8449 19119 8483
rect 19521 8483 19579 8489
rect 19521 8480 19533 8483
rect 19061 8443 19119 8449
rect 19168 8452 19533 8480
rect 15378 8412 15384 8424
rect 14660 8384 15384 8412
rect 15378 8372 15384 8384
rect 15436 8372 15442 8424
rect 16482 8412 16488 8424
rect 15856 8384 16488 8412
rect 10505 8347 10563 8353
rect 10505 8313 10517 8347
rect 10551 8344 10563 8347
rect 11514 8344 11520 8356
rect 10551 8316 11520 8344
rect 10551 8313 10563 8316
rect 10505 8307 10563 8313
rect 11514 8304 11520 8316
rect 11572 8304 11578 8356
rect 11698 8304 11704 8356
rect 11756 8304 11762 8356
rect 12529 8347 12587 8353
rect 12529 8313 12541 8347
rect 12575 8344 12587 8347
rect 13722 8344 13728 8356
rect 12575 8316 13728 8344
rect 12575 8313 12587 8316
rect 12529 8307 12587 8313
rect 13722 8304 13728 8316
rect 13780 8304 13786 8356
rect 14090 8304 14096 8356
rect 14148 8304 14154 8356
rect 14461 8347 14519 8353
rect 14461 8313 14473 8347
rect 14507 8344 14519 8347
rect 14734 8344 14740 8356
rect 14507 8316 14740 8344
rect 14507 8313 14519 8316
rect 14461 8307 14519 8313
rect 14734 8304 14740 8316
rect 14792 8304 14798 8356
rect 14918 8304 14924 8356
rect 14976 8344 14982 8356
rect 15565 8347 15623 8353
rect 14976 8316 15424 8344
rect 14976 8304 14982 8316
rect 8996 8248 9628 8276
rect 9677 8279 9735 8285
rect 8996 8236 9002 8248
rect 9677 8245 9689 8279
rect 9723 8276 9735 8279
rect 10686 8276 10692 8288
rect 9723 8248 10692 8276
rect 9723 8245 9735 8248
rect 9677 8239 9735 8245
rect 10686 8236 10692 8248
rect 10744 8236 10750 8288
rect 11330 8236 11336 8288
rect 11388 8276 11394 8288
rect 13538 8276 13544 8288
rect 11388 8248 13544 8276
rect 11388 8236 11394 8248
rect 13538 8236 13544 8248
rect 13596 8236 13602 8288
rect 13630 8236 13636 8288
rect 13688 8276 13694 8288
rect 15286 8276 15292 8288
rect 13688 8248 15292 8276
rect 13688 8236 13694 8248
rect 15286 8236 15292 8248
rect 15344 8236 15350 8288
rect 15396 8276 15424 8316
rect 15565 8313 15577 8347
rect 15611 8344 15623 8347
rect 15856 8344 15884 8384
rect 16482 8372 16488 8384
rect 16540 8372 16546 8424
rect 16853 8415 16911 8421
rect 16853 8381 16865 8415
rect 16899 8412 16911 8415
rect 17586 8412 17592 8424
rect 16899 8384 17592 8412
rect 16899 8381 16911 8384
rect 16853 8375 16911 8381
rect 17586 8372 17592 8384
rect 17644 8372 17650 8424
rect 15611 8316 15884 8344
rect 15933 8347 15991 8353
rect 15611 8313 15623 8316
rect 15565 8307 15623 8313
rect 15933 8313 15945 8347
rect 15979 8344 15991 8347
rect 16758 8344 16764 8356
rect 15979 8316 16764 8344
rect 15979 8313 15991 8316
rect 15933 8307 15991 8313
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 19168 8344 19196 8452
rect 19521 8449 19533 8452
rect 19567 8449 19579 8483
rect 19521 8443 19579 8449
rect 20530 8440 20536 8492
rect 20588 8480 20594 8492
rect 20717 8483 20775 8489
rect 20717 8480 20729 8483
rect 20588 8452 20729 8480
rect 20588 8440 20594 8452
rect 20717 8449 20729 8452
rect 20763 8449 20775 8483
rect 20717 8443 20775 8449
rect 21358 8440 21364 8492
rect 21416 8480 21422 8492
rect 21453 8483 21511 8489
rect 21453 8480 21465 8483
rect 21416 8452 21465 8480
rect 21416 8440 21422 8452
rect 21453 8449 21465 8452
rect 21499 8449 21511 8483
rect 21453 8443 21511 8449
rect 21542 8440 21548 8492
rect 21600 8480 21606 8492
rect 22112 8489 22140 8520
rect 22388 8489 22416 8588
rect 22554 8576 22560 8628
rect 22612 8616 22618 8628
rect 22612 8588 24164 8616
rect 22612 8576 22618 8588
rect 22462 8508 22468 8560
rect 22520 8548 22526 8560
rect 22520 8520 24072 8548
rect 22520 8508 22526 8520
rect 22005 8483 22063 8489
rect 22005 8480 22017 8483
rect 21600 8452 22017 8480
rect 21600 8440 21606 8452
rect 22005 8449 22017 8452
rect 22051 8449 22063 8483
rect 22005 8443 22063 8449
rect 22097 8483 22155 8489
rect 22097 8449 22109 8483
rect 22143 8449 22155 8483
rect 22097 8443 22155 8449
rect 22373 8483 22431 8489
rect 22373 8449 22385 8483
rect 22419 8449 22431 8483
rect 22373 8443 22431 8449
rect 22833 8483 22891 8489
rect 22833 8449 22845 8483
rect 22879 8449 22891 8483
rect 22833 8443 22891 8449
rect 19245 8415 19303 8421
rect 19245 8381 19257 8415
rect 19291 8381 19303 8415
rect 19245 8375 19303 8381
rect 16868 8316 19196 8344
rect 16868 8276 16896 8316
rect 15396 8248 16896 8276
rect 18782 8236 18788 8288
rect 18840 8276 18846 8288
rect 19260 8276 19288 8375
rect 20070 8372 20076 8424
rect 20128 8412 20134 8424
rect 20809 8415 20867 8421
rect 20809 8412 20821 8415
rect 20128 8384 20821 8412
rect 20128 8372 20134 8384
rect 20809 8381 20821 8384
rect 20855 8381 20867 8415
rect 20809 8375 20867 8381
rect 20901 8415 20959 8421
rect 20901 8381 20913 8415
rect 20947 8381 20959 8415
rect 20901 8375 20959 8381
rect 20257 8347 20315 8353
rect 20257 8313 20269 8347
rect 20303 8344 20315 8347
rect 20622 8344 20628 8356
rect 20303 8316 20628 8344
rect 20303 8313 20315 8316
rect 20257 8307 20315 8313
rect 20622 8304 20628 8316
rect 20680 8304 20686 8356
rect 18840 8248 19288 8276
rect 18840 8236 18846 8248
rect 20346 8236 20352 8288
rect 20404 8236 20410 8288
rect 20438 8236 20444 8288
rect 20496 8276 20502 8288
rect 20916 8276 20944 8375
rect 20990 8372 20996 8424
rect 21048 8412 21054 8424
rect 22848 8412 22876 8443
rect 23106 8440 23112 8492
rect 23164 8480 23170 8492
rect 24044 8489 24072 8520
rect 23385 8483 23443 8489
rect 23385 8480 23397 8483
rect 23164 8452 23397 8480
rect 23164 8440 23170 8452
rect 23385 8449 23397 8452
rect 23431 8449 23443 8483
rect 23385 8443 23443 8449
rect 24029 8483 24087 8489
rect 24029 8449 24041 8483
rect 24075 8449 24087 8483
rect 24136 8480 24164 8588
rect 24394 8576 24400 8628
rect 24452 8576 24458 8628
rect 24854 8576 24860 8628
rect 24912 8576 24918 8628
rect 25774 8576 25780 8628
rect 25832 8576 25838 8628
rect 26510 8576 26516 8628
rect 26568 8616 26574 8628
rect 27154 8616 27160 8628
rect 26568 8588 27160 8616
rect 26568 8576 26574 8588
rect 27154 8576 27160 8588
rect 27212 8576 27218 8628
rect 27522 8576 27528 8628
rect 27580 8616 27586 8628
rect 27580 8588 28856 8616
rect 27580 8576 27586 8588
rect 24486 8508 24492 8560
rect 24544 8548 24550 8560
rect 24544 8520 26004 8548
rect 24544 8508 24550 8520
rect 24581 8483 24639 8489
rect 24581 8480 24593 8483
rect 24136 8452 24593 8480
rect 24029 8443 24087 8449
rect 24581 8449 24593 8452
rect 24627 8449 24639 8483
rect 24581 8443 24639 8449
rect 24670 8440 24676 8492
rect 24728 8440 24734 8492
rect 25130 8440 25136 8492
rect 25188 8440 25194 8492
rect 25406 8440 25412 8492
rect 25464 8440 25470 8492
rect 25976 8489 26004 8520
rect 26142 8508 26148 8560
rect 26200 8548 26206 8560
rect 26200 8520 27292 8548
rect 26200 8508 26206 8520
rect 25685 8483 25743 8489
rect 25685 8449 25697 8483
rect 25731 8449 25743 8483
rect 25685 8443 25743 8449
rect 25961 8483 26019 8489
rect 25961 8449 25973 8483
rect 26007 8449 26019 8483
rect 25961 8443 26019 8449
rect 21048 8384 22876 8412
rect 21048 8372 21054 8384
rect 23290 8372 23296 8424
rect 23348 8412 23354 8424
rect 23477 8415 23535 8421
rect 23477 8412 23489 8415
rect 23348 8384 23489 8412
rect 23348 8372 23354 8384
rect 23477 8381 23489 8384
rect 23523 8381 23535 8415
rect 23477 8375 23535 8381
rect 23566 8372 23572 8424
rect 23624 8372 23630 8424
rect 23658 8372 23664 8424
rect 23716 8412 23722 8424
rect 25700 8412 25728 8443
rect 26234 8440 26240 8492
rect 26292 8440 26298 8492
rect 26326 8440 26332 8492
rect 26384 8440 26390 8492
rect 26786 8440 26792 8492
rect 26844 8440 26850 8492
rect 27062 8480 27068 8492
rect 26896 8452 27068 8480
rect 23716 8384 25728 8412
rect 23716 8372 23722 8384
rect 25774 8372 25780 8424
rect 25832 8412 25838 8424
rect 26896 8412 26924 8452
rect 27062 8440 27068 8452
rect 27120 8440 27126 8492
rect 27154 8440 27160 8492
rect 27212 8440 27218 8492
rect 25832 8384 26924 8412
rect 27264 8412 27292 8520
rect 27338 8508 27344 8560
rect 27396 8548 27402 8560
rect 27396 8520 28396 8548
rect 27396 8508 27402 8520
rect 27430 8440 27436 8492
rect 27488 8440 27494 8492
rect 27525 8483 27583 8489
rect 27525 8449 27537 8483
rect 27571 8449 27583 8483
rect 27985 8483 28043 8489
rect 27985 8480 27997 8483
rect 27525 8443 27583 8449
rect 27632 8452 27997 8480
rect 27540 8412 27568 8443
rect 27264 8384 27568 8412
rect 25832 8372 25838 8384
rect 21821 8347 21879 8353
rect 21821 8313 21833 8347
rect 21867 8344 21879 8347
rect 21910 8344 21916 8356
rect 21867 8316 21916 8344
rect 21867 8313 21879 8316
rect 21821 8307 21879 8313
rect 21910 8304 21916 8316
rect 21968 8304 21974 8356
rect 22094 8304 22100 8356
rect 22152 8344 22158 8356
rect 22281 8347 22339 8353
rect 22281 8344 22293 8347
rect 22152 8316 22293 8344
rect 22152 8304 22158 8316
rect 22281 8313 22293 8316
rect 22327 8313 22339 8347
rect 22281 8307 22339 8313
rect 22370 8304 22376 8356
rect 22428 8344 22434 8356
rect 22557 8347 22615 8353
rect 22557 8344 22569 8347
rect 22428 8316 22569 8344
rect 22428 8304 22434 8316
rect 22557 8313 22569 8316
rect 22603 8313 22615 8347
rect 22557 8307 22615 8313
rect 22646 8304 22652 8356
rect 22704 8304 22710 8356
rect 22830 8304 22836 8356
rect 22888 8344 22894 8356
rect 24949 8347 25007 8353
rect 24949 8344 24961 8347
rect 22888 8316 24961 8344
rect 22888 8304 22894 8316
rect 24949 8313 24961 8316
rect 24995 8313 25007 8347
rect 26053 8347 26111 8353
rect 26053 8344 26065 8347
rect 24949 8307 25007 8313
rect 25056 8316 26065 8344
rect 20496 8248 20944 8276
rect 20496 8236 20502 8248
rect 22002 8236 22008 8288
rect 22060 8276 22066 8288
rect 23017 8279 23075 8285
rect 23017 8276 23029 8279
rect 22060 8248 23029 8276
rect 22060 8236 22066 8248
rect 23017 8245 23029 8248
rect 23063 8245 23075 8279
rect 23017 8239 23075 8245
rect 23842 8236 23848 8288
rect 23900 8236 23906 8288
rect 24762 8236 24768 8288
rect 24820 8276 24826 8288
rect 25056 8276 25084 8316
rect 26053 8313 26065 8316
rect 26099 8313 26111 8347
rect 26053 8307 26111 8313
rect 26418 8304 26424 8356
rect 26476 8344 26482 8356
rect 27632 8344 27660 8452
rect 27985 8449 27997 8452
rect 28031 8449 28043 8483
rect 27985 8443 28043 8449
rect 28258 8440 28264 8492
rect 28316 8440 28322 8492
rect 28368 8489 28396 8520
rect 28828 8489 28856 8588
rect 28994 8576 29000 8628
rect 29052 8616 29058 8628
rect 29181 8619 29239 8625
rect 29181 8616 29193 8619
rect 29052 8588 29193 8616
rect 29052 8576 29058 8588
rect 29181 8585 29193 8588
rect 29227 8585 29239 8619
rect 29181 8579 29239 8585
rect 29730 8576 29736 8628
rect 29788 8616 29794 8628
rect 31573 8619 31631 8625
rect 29788 8588 31524 8616
rect 29788 8576 29794 8588
rect 28902 8508 28908 8560
rect 28960 8548 28966 8560
rect 28960 8520 29408 8548
rect 28960 8508 28966 8520
rect 29380 8489 29408 8520
rect 29454 8508 29460 8560
rect 29512 8548 29518 8560
rect 29512 8520 31248 8548
rect 29512 8508 29518 8520
rect 28353 8483 28411 8489
rect 28353 8449 28365 8483
rect 28399 8449 28411 8483
rect 28353 8443 28411 8449
rect 28813 8483 28871 8489
rect 28813 8449 28825 8483
rect 28859 8449 28871 8483
rect 28813 8443 28871 8449
rect 29089 8483 29147 8489
rect 29089 8449 29101 8483
rect 29135 8449 29147 8483
rect 29089 8443 29147 8449
rect 29365 8483 29423 8489
rect 29365 8449 29377 8483
rect 29411 8449 29423 8483
rect 29365 8443 29423 8449
rect 27798 8372 27804 8424
rect 27856 8412 27862 8424
rect 29104 8412 29132 8443
rect 29822 8440 29828 8492
rect 29880 8440 29886 8492
rect 30650 8440 30656 8492
rect 30708 8440 30714 8492
rect 30926 8440 30932 8492
rect 30984 8440 30990 8492
rect 31220 8489 31248 8520
rect 31496 8489 31524 8588
rect 31573 8585 31585 8619
rect 31619 8616 31631 8619
rect 31938 8616 31944 8628
rect 31619 8588 31944 8616
rect 31619 8585 31631 8588
rect 31573 8579 31631 8585
rect 31938 8576 31944 8588
rect 31996 8576 32002 8628
rect 32490 8576 32496 8628
rect 32548 8616 32554 8628
rect 33229 8619 33287 8625
rect 33229 8616 33241 8619
rect 32548 8588 33241 8616
rect 32548 8576 32554 8588
rect 33229 8585 33241 8588
rect 33275 8585 33287 8619
rect 33229 8579 33287 8585
rect 33778 8576 33784 8628
rect 33836 8616 33842 8628
rect 33873 8619 33931 8625
rect 33873 8616 33885 8619
rect 33836 8588 33885 8616
rect 33836 8576 33842 8588
rect 33873 8585 33885 8588
rect 33919 8585 33931 8619
rect 33873 8579 33931 8585
rect 34146 8576 34152 8628
rect 34204 8616 34210 8628
rect 34204 8588 34652 8616
rect 34204 8576 34210 8588
rect 31662 8508 31668 8560
rect 31720 8548 31726 8560
rect 34514 8548 34520 8560
rect 31720 8520 32444 8548
rect 31720 8508 31726 8520
rect 31205 8483 31263 8489
rect 31205 8449 31217 8483
rect 31251 8449 31263 8483
rect 31205 8443 31263 8449
rect 31481 8483 31539 8489
rect 31481 8449 31493 8483
rect 31527 8449 31539 8483
rect 31481 8443 31539 8449
rect 31570 8440 31576 8492
rect 31628 8480 31634 8492
rect 32416 8489 32444 8520
rect 34440 8520 34520 8548
rect 31757 8483 31815 8489
rect 31757 8480 31769 8483
rect 31628 8452 31769 8480
rect 31628 8440 31634 8452
rect 31757 8449 31769 8452
rect 31803 8449 31815 8483
rect 31757 8443 31815 8449
rect 32401 8483 32459 8489
rect 32401 8449 32413 8483
rect 32447 8449 32459 8483
rect 32401 8443 32459 8449
rect 33045 8483 33103 8489
rect 33045 8449 33057 8483
rect 33091 8449 33103 8483
rect 33045 8443 33103 8449
rect 33689 8483 33747 8489
rect 33689 8449 33701 8483
rect 33735 8480 33747 8483
rect 33778 8480 33784 8492
rect 33735 8452 33784 8480
rect 33735 8449 33747 8452
rect 33689 8443 33747 8449
rect 27856 8384 29132 8412
rect 27856 8372 27862 8384
rect 29178 8372 29184 8424
rect 29236 8412 29242 8424
rect 29549 8415 29607 8421
rect 29549 8412 29561 8415
rect 29236 8384 29561 8412
rect 29236 8372 29242 8384
rect 29549 8381 29561 8384
rect 29595 8381 29607 8415
rect 31294 8412 31300 8424
rect 29549 8375 29607 8381
rect 29840 8384 31300 8412
rect 26476 8316 27660 8344
rect 26476 8304 26482 8316
rect 27706 8304 27712 8356
rect 27764 8304 27770 8356
rect 28074 8304 28080 8356
rect 28132 8304 28138 8356
rect 28537 8347 28595 8353
rect 28537 8313 28549 8347
rect 28583 8344 28595 8347
rect 29840 8344 29868 8384
rect 31294 8372 31300 8384
rect 31352 8372 31358 8424
rect 31386 8372 31392 8424
rect 31444 8412 31450 8424
rect 32125 8415 32183 8421
rect 32125 8412 32137 8415
rect 31444 8384 32137 8412
rect 31444 8372 31450 8384
rect 32125 8381 32137 8384
rect 32171 8381 32183 8415
rect 33066 8412 33094 8443
rect 33778 8440 33784 8452
rect 33836 8440 33842 8492
rect 34440 8489 34468 8520
rect 34514 8508 34520 8520
rect 34572 8508 34578 8560
rect 34057 8483 34115 8489
rect 34057 8449 34069 8483
rect 34103 8480 34115 8483
rect 34425 8483 34483 8489
rect 34103 8452 34376 8480
rect 34103 8449 34115 8452
rect 34057 8443 34115 8449
rect 32125 8375 32183 8381
rect 32232 8384 33094 8412
rect 28583 8316 29868 8344
rect 28583 8313 28595 8316
rect 28537 8307 28595 8313
rect 29914 8304 29920 8356
rect 29972 8344 29978 8356
rect 31021 8347 31079 8353
rect 31021 8344 31033 8347
rect 29972 8316 31033 8344
rect 29972 8304 29978 8316
rect 31021 8313 31033 8316
rect 31067 8313 31079 8347
rect 31021 8307 31079 8313
rect 31202 8304 31208 8356
rect 31260 8344 31266 8356
rect 32232 8344 32260 8384
rect 33410 8372 33416 8424
rect 33468 8412 33474 8424
rect 34348 8412 34376 8452
rect 34425 8449 34437 8483
rect 34471 8449 34483 8483
rect 34425 8443 34483 8449
rect 34514 8412 34520 8424
rect 33468 8384 34284 8412
rect 34348 8384 34520 8412
rect 33468 8372 33474 8384
rect 31260 8316 32260 8344
rect 31260 8304 31266 8316
rect 32766 8304 32772 8356
rect 32824 8344 32830 8356
rect 34256 8353 34284 8384
rect 34514 8372 34520 8384
rect 34572 8372 34578 8424
rect 34624 8412 34652 8588
rect 34698 8576 34704 8628
rect 34756 8616 34762 8628
rect 35529 8619 35587 8625
rect 35529 8616 35541 8619
rect 34756 8588 35541 8616
rect 34756 8576 34762 8588
rect 35529 8585 35541 8588
rect 35575 8585 35587 8619
rect 35529 8579 35587 8585
rect 35802 8576 35808 8628
rect 35860 8616 35866 8628
rect 36633 8619 36691 8625
rect 36633 8616 36645 8619
rect 35860 8588 36645 8616
rect 35860 8576 35866 8588
rect 36633 8585 36645 8588
rect 36679 8585 36691 8619
rect 36633 8579 36691 8585
rect 36906 8576 36912 8628
rect 36964 8616 36970 8628
rect 37737 8619 37795 8625
rect 37737 8616 37749 8619
rect 36964 8588 37749 8616
rect 36964 8576 36970 8588
rect 37737 8585 37749 8588
rect 37783 8585 37795 8619
rect 37737 8579 37795 8585
rect 38473 8619 38531 8625
rect 38473 8585 38485 8619
rect 38519 8585 38531 8619
rect 38473 8579 38531 8585
rect 37090 8548 37096 8560
rect 34992 8520 37096 8548
rect 34992 8489 35020 8520
rect 37090 8508 37096 8520
rect 37148 8508 37154 8560
rect 37458 8508 37464 8560
rect 37516 8548 37522 8560
rect 38488 8548 38516 8579
rect 38930 8576 38936 8628
rect 38988 8616 38994 8628
rect 39025 8619 39083 8625
rect 39025 8616 39037 8619
rect 38988 8588 39037 8616
rect 38988 8576 38994 8588
rect 39025 8585 39037 8588
rect 39071 8585 39083 8619
rect 39025 8579 39083 8585
rect 37516 8520 38516 8548
rect 37516 8508 37522 8520
rect 34977 8483 35035 8489
rect 34977 8449 34989 8483
rect 35023 8449 35035 8483
rect 34977 8443 35035 8449
rect 35342 8440 35348 8492
rect 35400 8440 35406 8492
rect 35710 8440 35716 8492
rect 35768 8440 35774 8492
rect 35802 8440 35808 8492
rect 35860 8440 35866 8492
rect 36449 8483 36507 8489
rect 36449 8449 36461 8483
rect 36495 8480 36507 8483
rect 36722 8480 36728 8492
rect 36495 8452 36728 8480
rect 36495 8449 36507 8452
rect 36449 8443 36507 8449
rect 36722 8440 36728 8452
rect 36780 8440 36786 8492
rect 36814 8440 36820 8492
rect 36872 8440 36878 8492
rect 37274 8440 37280 8492
rect 37332 8440 37338 8492
rect 37826 8440 37832 8492
rect 37884 8480 37890 8492
rect 37921 8483 37979 8489
rect 37921 8480 37933 8483
rect 37884 8452 37933 8480
rect 37884 8440 37890 8452
rect 37921 8449 37933 8452
rect 37967 8449 37979 8483
rect 37921 8443 37979 8449
rect 38013 8483 38071 8489
rect 38013 8449 38025 8483
rect 38059 8449 38071 8483
rect 38013 8443 38071 8449
rect 34624 8384 35204 8412
rect 33505 8347 33563 8353
rect 33505 8344 33517 8347
rect 32824 8316 33517 8344
rect 32824 8304 32830 8316
rect 33505 8313 33517 8316
rect 33551 8313 33563 8347
rect 33505 8307 33563 8313
rect 34241 8347 34299 8353
rect 34241 8313 34253 8347
rect 34287 8313 34299 8347
rect 34241 8307 34299 8313
rect 34330 8304 34336 8356
rect 34388 8344 34394 8356
rect 34793 8347 34851 8353
rect 34793 8344 34805 8347
rect 34388 8316 34805 8344
rect 34388 8304 34394 8316
rect 34793 8313 34805 8316
rect 34839 8313 34851 8347
rect 34793 8307 34851 8313
rect 34974 8304 34980 8356
rect 35032 8344 35038 8356
rect 35176 8353 35204 8384
rect 35618 8372 35624 8424
rect 35676 8412 35682 8424
rect 38028 8412 38056 8443
rect 38562 8440 38568 8492
rect 38620 8480 38626 8492
rect 38657 8483 38715 8489
rect 38657 8480 38669 8483
rect 38620 8452 38669 8480
rect 38620 8440 38626 8452
rect 38657 8449 38669 8452
rect 38703 8449 38715 8483
rect 38657 8443 38715 8449
rect 39117 8483 39175 8489
rect 39117 8449 39129 8483
rect 39163 8480 39175 8483
rect 39209 8483 39267 8489
rect 39209 8480 39221 8483
rect 39163 8452 39221 8480
rect 39163 8449 39175 8452
rect 39117 8443 39175 8449
rect 39209 8449 39221 8452
rect 39255 8449 39267 8483
rect 39209 8443 39267 8449
rect 35676 8384 38056 8412
rect 35676 8372 35682 8384
rect 35161 8347 35219 8353
rect 35032 8316 35112 8344
rect 35032 8304 35038 8316
rect 24820 8248 25084 8276
rect 24820 8236 24826 8248
rect 25222 8236 25228 8288
rect 25280 8236 25286 8288
rect 25498 8236 25504 8288
rect 25556 8236 25562 8288
rect 26510 8236 26516 8288
rect 26568 8236 26574 8288
rect 26602 8236 26608 8288
rect 26660 8236 26666 8288
rect 26694 8236 26700 8288
rect 26752 8276 26758 8288
rect 26973 8279 27031 8285
rect 26973 8276 26985 8279
rect 26752 8248 26985 8276
rect 26752 8236 26758 8248
rect 26973 8245 26985 8248
rect 27019 8245 27031 8279
rect 26973 8239 27031 8245
rect 27062 8236 27068 8288
rect 27120 8276 27126 8288
rect 27249 8279 27307 8285
rect 27249 8276 27261 8279
rect 27120 8248 27261 8276
rect 27120 8236 27126 8248
rect 27249 8245 27261 8248
rect 27295 8245 27307 8279
rect 27249 8239 27307 8245
rect 27801 8279 27859 8285
rect 27801 8245 27813 8279
rect 27847 8276 27859 8279
rect 27890 8276 27896 8288
rect 27847 8248 27896 8276
rect 27847 8245 27859 8248
rect 27801 8239 27859 8245
rect 27890 8236 27896 8248
rect 27948 8236 27954 8288
rect 28629 8279 28687 8285
rect 28629 8245 28641 8279
rect 28675 8276 28687 8279
rect 28718 8276 28724 8288
rect 28675 8248 28724 8276
rect 28675 8245 28687 8248
rect 28629 8239 28687 8245
rect 28718 8236 28724 8248
rect 28776 8236 28782 8288
rect 28810 8236 28816 8288
rect 28868 8276 28874 8288
rect 28905 8279 28963 8285
rect 28905 8276 28917 8279
rect 28868 8248 28917 8276
rect 28868 8236 28874 8248
rect 28905 8245 28917 8248
rect 28951 8245 28963 8279
rect 28905 8239 28963 8245
rect 30466 8236 30472 8288
rect 30524 8236 30530 8288
rect 30742 8236 30748 8288
rect 30800 8236 30806 8288
rect 30926 8236 30932 8288
rect 30984 8276 30990 8288
rect 31297 8279 31355 8285
rect 31297 8276 31309 8279
rect 30984 8248 31309 8276
rect 30984 8236 30990 8248
rect 31297 8245 31309 8248
rect 31343 8245 31355 8279
rect 31297 8239 31355 8245
rect 31662 8236 31668 8288
rect 31720 8276 31726 8288
rect 34882 8276 34888 8288
rect 31720 8248 34888 8276
rect 31720 8236 31726 8248
rect 34882 8236 34888 8248
rect 34940 8236 34946 8288
rect 35084 8276 35112 8316
rect 35161 8313 35173 8347
rect 35207 8313 35219 8347
rect 35161 8307 35219 8313
rect 35250 8304 35256 8356
rect 35308 8344 35314 8356
rect 36265 8347 36323 8353
rect 36265 8344 36277 8347
rect 35308 8316 36277 8344
rect 35308 8304 35314 8316
rect 36265 8313 36277 8316
rect 36311 8313 36323 8347
rect 36265 8307 36323 8313
rect 36354 8304 36360 8356
rect 36412 8344 36418 8356
rect 36412 8316 37136 8344
rect 36412 8304 36418 8316
rect 35989 8279 36047 8285
rect 35989 8276 36001 8279
rect 35084 8248 36001 8276
rect 35989 8245 36001 8248
rect 36035 8245 36047 8279
rect 37108 8276 37136 8316
rect 37182 8304 37188 8356
rect 37240 8344 37246 8356
rect 38197 8347 38255 8353
rect 38197 8344 38209 8347
rect 37240 8316 38209 8344
rect 37240 8304 37246 8316
rect 38197 8313 38209 8316
rect 38243 8313 38255 8347
rect 38197 8307 38255 8313
rect 39390 8304 39396 8356
rect 39448 8304 39454 8356
rect 37461 8279 37519 8285
rect 37461 8276 37473 8279
rect 37108 8248 37473 8276
rect 35989 8239 36047 8245
rect 37461 8245 37473 8248
rect 37507 8245 37519 8279
rect 37461 8239 37519 8245
rect 1104 8186 39836 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 37950 8186
rect 38002 8134 38014 8186
rect 38066 8134 38078 8186
rect 38130 8134 38142 8186
rect 38194 8134 38206 8186
rect 38258 8134 39836 8186
rect 1104 8112 39836 8134
rect 3418 8032 3424 8084
rect 3476 8032 3482 8084
rect 3510 8032 3516 8084
rect 3568 8072 3574 8084
rect 3881 8075 3939 8081
rect 3881 8072 3893 8075
rect 3568 8044 3893 8072
rect 3568 8032 3574 8044
rect 3881 8041 3893 8044
rect 3927 8041 3939 8075
rect 3881 8035 3939 8041
rect 4062 8032 4068 8084
rect 4120 8072 4126 8084
rect 4249 8075 4307 8081
rect 4249 8072 4261 8075
rect 4120 8044 4261 8072
rect 4120 8032 4126 8044
rect 4249 8041 4261 8044
rect 4295 8041 4307 8075
rect 4249 8035 4307 8041
rect 4614 8032 4620 8084
rect 4672 8072 4678 8084
rect 4801 8075 4859 8081
rect 4801 8072 4813 8075
rect 4672 8044 4813 8072
rect 4672 8032 4678 8044
rect 4801 8041 4813 8044
rect 4847 8041 4859 8075
rect 4801 8035 4859 8041
rect 5166 8032 5172 8084
rect 5224 8072 5230 8084
rect 5353 8075 5411 8081
rect 5353 8072 5365 8075
rect 5224 8044 5365 8072
rect 5224 8032 5230 8044
rect 5353 8041 5365 8044
rect 5399 8041 5411 8075
rect 5353 8035 5411 8041
rect 5718 8032 5724 8084
rect 5776 8072 5782 8084
rect 5813 8075 5871 8081
rect 5813 8072 5825 8075
rect 5776 8044 5825 8072
rect 5776 8032 5782 8044
rect 5813 8041 5825 8044
rect 5859 8041 5871 8075
rect 5813 8035 5871 8041
rect 6181 8075 6239 8081
rect 6181 8041 6193 8075
rect 6227 8072 6239 8075
rect 6546 8072 6552 8084
rect 6227 8044 6552 8072
rect 6227 8041 6239 8044
rect 6181 8035 6239 8041
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 6730 8032 6736 8084
rect 6788 8072 6794 8084
rect 6825 8075 6883 8081
rect 6825 8072 6837 8075
rect 6788 8044 6837 8072
rect 6788 8032 6794 8044
rect 6825 8041 6837 8044
rect 6871 8041 6883 8075
rect 6825 8035 6883 8041
rect 7466 8032 7472 8084
rect 7524 8032 7530 8084
rect 8938 8072 8944 8084
rect 7760 8044 8944 8072
rect 2590 7964 2596 8016
rect 2648 7964 2654 8016
rect 5074 7964 5080 8016
rect 5132 8004 5138 8016
rect 7101 8007 7159 8013
rect 5132 7976 6960 8004
rect 5132 7964 5138 7976
rect 658 7896 664 7948
rect 716 7936 722 7948
rect 1397 7939 1455 7945
rect 1397 7936 1409 7939
rect 716 7908 1409 7936
rect 716 7896 722 7908
rect 1397 7905 1409 7908
rect 1443 7905 1455 7939
rect 1397 7899 1455 7905
rect 2961 7939 3019 7945
rect 2961 7905 2973 7939
rect 3007 7936 3019 7939
rect 6822 7936 6828 7948
rect 3007 7908 6828 7936
rect 3007 7905 3019 7908
rect 2961 7899 3019 7905
rect 6822 7896 6828 7908
rect 6880 7896 6886 7948
rect 6932 7936 6960 7976
rect 7101 7973 7113 8007
rect 7147 8004 7159 8007
rect 7650 8004 7656 8016
rect 7147 7976 7656 8004
rect 7147 7973 7159 7976
rect 7101 7967 7159 7973
rect 7650 7964 7656 7976
rect 7708 7964 7714 8016
rect 7760 7936 7788 8044
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 10137 8075 10195 8081
rect 10137 8041 10149 8075
rect 10183 8072 10195 8075
rect 10410 8072 10416 8084
rect 10183 8044 10416 8072
rect 10183 8041 10195 8044
rect 10137 8035 10195 8041
rect 10410 8032 10416 8044
rect 10468 8032 10474 8084
rect 10520 8044 12756 8072
rect 9953 8007 10011 8013
rect 9953 7973 9965 8007
rect 9999 8004 10011 8007
rect 10520 8004 10548 8044
rect 9999 7976 10548 8004
rect 11793 8007 11851 8013
rect 9999 7973 10011 7976
rect 9953 7967 10011 7973
rect 11793 7973 11805 8007
rect 11839 8004 11851 8007
rect 12342 8004 12348 8016
rect 11839 7976 12348 8004
rect 11839 7973 11851 7976
rect 11793 7967 11851 7973
rect 12342 7964 12348 7976
rect 12400 7964 12406 8016
rect 12728 8013 12756 8044
rect 12802 8032 12808 8084
rect 12860 8072 12866 8084
rect 13262 8072 13268 8084
rect 12860 8044 13268 8072
rect 12860 8032 12866 8044
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 13354 8032 13360 8084
rect 13412 8072 13418 8084
rect 13412 8044 14044 8072
rect 13412 8032 13418 8044
rect 12713 8007 12771 8013
rect 12713 7973 12725 8007
rect 12759 7973 12771 8007
rect 14016 8004 14044 8044
rect 14090 8032 14096 8084
rect 14148 8072 14154 8084
rect 15565 8075 15623 8081
rect 14148 8044 15240 8072
rect 14148 8032 14154 8044
rect 14366 8004 14372 8016
rect 14016 7976 14372 8004
rect 12713 7967 12771 7973
rect 14366 7964 14372 7976
rect 14424 7964 14430 8016
rect 6932 7908 7788 7936
rect 8662 7896 8668 7948
rect 8720 7936 8726 7948
rect 8846 7936 8852 7948
rect 8720 7908 8852 7936
rect 8720 7896 8726 7908
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 10226 7896 10232 7948
rect 10284 7936 10290 7948
rect 10413 7939 10471 7945
rect 10413 7936 10425 7939
rect 10284 7908 10425 7936
rect 10284 7896 10290 7908
rect 10413 7905 10425 7908
rect 10459 7905 10471 7939
rect 10413 7899 10471 7905
rect 11514 7896 11520 7948
rect 11572 7936 11578 7948
rect 13265 7939 13323 7945
rect 13265 7936 13277 7939
rect 11572 7908 13277 7936
rect 11572 7896 11578 7908
rect 13265 7905 13277 7908
rect 13311 7905 13323 7939
rect 13265 7899 13323 7905
rect 15102 7896 15108 7948
rect 15160 7896 15166 7948
rect 15212 7936 15240 8044
rect 15565 8041 15577 8075
rect 15611 8072 15623 8075
rect 15654 8072 15660 8084
rect 15611 8044 15660 8072
rect 15611 8041 15623 8044
rect 15565 8035 15623 8041
rect 15654 8032 15660 8044
rect 15712 8032 15718 8084
rect 19426 8072 19432 8084
rect 17880 8044 19432 8072
rect 16853 8007 16911 8013
rect 16853 7973 16865 8007
rect 16899 8004 16911 8007
rect 16899 7976 17724 8004
rect 16899 7973 16911 7976
rect 16853 7967 16911 7973
rect 15654 7936 15660 7948
rect 15212 7908 15660 7936
rect 15654 7896 15660 7908
rect 15712 7936 15718 7948
rect 17696 7945 17724 7976
rect 15841 7939 15899 7945
rect 15841 7936 15853 7939
rect 15712 7908 15853 7936
rect 15712 7896 15718 7908
rect 15841 7905 15853 7908
rect 15887 7905 15899 7939
rect 15841 7899 15899 7905
rect 17681 7939 17739 7945
rect 17681 7905 17693 7939
rect 17727 7905 17739 7939
rect 17681 7899 17739 7905
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 1719 7840 2728 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 382 7760 388 7812
rect 440 7800 446 7812
rect 2409 7803 2467 7809
rect 2409 7800 2421 7803
rect 440 7772 2421 7800
rect 440 7760 446 7772
rect 2409 7769 2421 7772
rect 2455 7769 2467 7803
rect 2700 7800 2728 7840
rect 2774 7828 2780 7880
rect 2832 7828 2838 7880
rect 2866 7828 2872 7880
rect 2924 7868 2930 7880
rect 3053 7871 3111 7877
rect 3053 7868 3065 7871
rect 2924 7840 3065 7868
rect 2924 7828 2930 7840
rect 3053 7837 3065 7840
rect 3099 7837 3111 7871
rect 3053 7831 3111 7837
rect 3602 7828 3608 7880
rect 3660 7828 3666 7880
rect 3970 7828 3976 7880
rect 4028 7868 4034 7880
rect 4065 7871 4123 7877
rect 4065 7868 4077 7871
rect 4028 7840 4077 7868
rect 4028 7828 4034 7840
rect 4065 7837 4077 7840
rect 4111 7837 4123 7871
rect 4065 7831 4123 7837
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7868 4491 7871
rect 4890 7868 4896 7880
rect 4479 7840 4896 7868
rect 4479 7837 4491 7840
rect 4433 7831 4491 7837
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 4982 7828 4988 7880
rect 5040 7828 5046 7880
rect 5534 7828 5540 7880
rect 5592 7828 5598 7880
rect 5994 7828 6000 7880
rect 6052 7828 6058 7880
rect 6362 7828 6368 7880
rect 6420 7828 6426 7880
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7868 6607 7871
rect 6641 7871 6699 7877
rect 6641 7868 6653 7871
rect 6595 7840 6653 7868
rect 6595 7837 6607 7840
rect 6549 7831 6607 7837
rect 6641 7837 6653 7840
rect 6687 7837 6699 7871
rect 6641 7831 6699 7837
rect 7282 7828 7288 7880
rect 7340 7828 7346 7880
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 7432 7840 7665 7868
rect 7432 7828 7438 7840
rect 7653 7837 7665 7840
rect 7699 7837 7711 7871
rect 7653 7831 7711 7837
rect 7742 7828 7748 7880
rect 7800 7828 7806 7880
rect 8018 7828 8024 7880
rect 8076 7828 8082 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8588 7840 8953 7868
rect 7558 7800 7564 7812
rect 2700 7772 7564 7800
rect 2409 7763 2467 7769
rect 7558 7760 7564 7772
rect 7616 7760 7622 7812
rect 8386 7760 8392 7812
rect 8444 7800 8450 7812
rect 8588 7800 8616 7840
rect 8941 7837 8953 7840
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 9214 7828 9220 7880
rect 9272 7828 9278 7880
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7838 10379 7871
rect 10367 7837 10456 7838
rect 10321 7831 10456 7837
rect 10336 7812 10456 7831
rect 10686 7828 10692 7880
rect 10744 7868 10750 7880
rect 11146 7868 11152 7880
rect 10744 7840 11152 7868
rect 10744 7828 10750 7840
rect 11146 7828 11152 7840
rect 11204 7868 11210 7880
rect 11204 7840 11928 7868
rect 11204 7828 11210 7840
rect 9950 7800 9956 7812
rect 8444 7772 8616 7800
rect 8956 7772 9956 7800
rect 8444 7760 8450 7772
rect 1210 7692 1216 7744
rect 1268 7732 1274 7744
rect 1946 7732 1952 7744
rect 1268 7704 1952 7732
rect 1268 7692 1274 7704
rect 1946 7692 1952 7704
rect 2004 7692 2010 7744
rect 3237 7735 3295 7741
rect 3237 7701 3249 7735
rect 3283 7732 3295 7735
rect 4430 7732 4436 7744
rect 3283 7704 4436 7732
rect 3283 7701 3295 7704
rect 3237 7695 3295 7701
rect 4430 7692 4436 7704
rect 4488 7692 4494 7744
rect 6549 7735 6607 7741
rect 6549 7701 6561 7735
rect 6595 7732 6607 7735
rect 6638 7732 6644 7744
rect 6595 7704 6644 7732
rect 6595 7701 6607 7704
rect 6549 7695 6607 7701
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 6730 7692 6736 7744
rect 6788 7732 6794 7744
rect 8662 7732 8668 7744
rect 6788 7704 8668 7732
rect 6788 7692 6794 7704
rect 8662 7692 8668 7704
rect 8720 7692 8726 7744
rect 8757 7735 8815 7741
rect 8757 7701 8769 7735
rect 8803 7732 8815 7735
rect 8956 7732 8984 7772
rect 9950 7760 9956 7772
rect 10008 7760 10014 7812
rect 10336 7810 10416 7812
rect 10410 7760 10416 7810
rect 10468 7760 10474 7812
rect 8803 7704 8984 7732
rect 8803 7701 8815 7704
rect 8757 7695 8815 7701
rect 9030 7692 9036 7744
rect 9088 7732 9094 7744
rect 11146 7732 11152 7744
rect 9088 7704 11152 7732
rect 9088 7692 9094 7704
rect 11146 7692 11152 7704
rect 11204 7692 11210 7744
rect 11422 7692 11428 7744
rect 11480 7692 11486 7744
rect 11900 7732 11928 7840
rect 11974 7828 11980 7880
rect 12032 7828 12038 7880
rect 12066 7828 12072 7880
rect 12124 7828 12130 7880
rect 12250 7828 12256 7880
rect 12308 7828 12314 7880
rect 12986 7828 12992 7880
rect 13044 7828 13050 7880
rect 13078 7828 13084 7880
rect 13136 7877 13142 7880
rect 13136 7871 13164 7877
rect 13152 7837 13164 7871
rect 14829 7871 14887 7877
rect 14829 7868 14841 7871
rect 13136 7831 13164 7837
rect 13832 7840 14841 7868
rect 13136 7828 13142 7831
rect 13832 7732 13860 7840
rect 14829 7837 14841 7840
rect 14875 7868 14887 7871
rect 14918 7868 14924 7880
rect 14875 7840 14924 7868
rect 14875 7837 14887 7840
rect 14829 7831 14887 7837
rect 14918 7828 14924 7840
rect 14976 7828 14982 7880
rect 15381 7871 15439 7877
rect 15381 7868 15393 7871
rect 15028 7840 15393 7868
rect 13909 7803 13967 7809
rect 13909 7769 13921 7803
rect 13955 7800 13967 7803
rect 15028 7800 15056 7840
rect 15381 7837 15393 7840
rect 15427 7837 15439 7871
rect 15381 7831 15439 7837
rect 15749 7871 15807 7877
rect 15749 7837 15761 7871
rect 15795 7864 15807 7871
rect 16117 7871 16175 7877
rect 15795 7837 15976 7864
rect 15749 7836 15976 7837
rect 15749 7831 15807 7836
rect 15948 7800 15976 7836
rect 16117 7837 16129 7871
rect 16163 7868 16175 7871
rect 16206 7868 16212 7880
rect 16163 7840 16212 7868
rect 16163 7837 16175 7840
rect 16117 7831 16175 7837
rect 16206 7828 16212 7840
rect 16264 7828 16270 7880
rect 17497 7871 17555 7877
rect 17497 7837 17509 7871
rect 17543 7868 17555 7871
rect 17880 7868 17908 8044
rect 19426 8032 19432 8044
rect 19484 8032 19490 8084
rect 19702 8032 19708 8084
rect 19760 8032 19766 8084
rect 19886 8032 19892 8084
rect 19944 8072 19950 8084
rect 20346 8072 20352 8084
rect 19944 8044 20352 8072
rect 19944 8032 19950 8044
rect 20346 8032 20352 8044
rect 20404 8032 20410 8084
rect 23106 8032 23112 8084
rect 23164 8072 23170 8084
rect 24949 8075 25007 8081
rect 24949 8072 24961 8075
rect 23164 8044 24961 8072
rect 23164 8032 23170 8044
rect 18966 8004 18972 8016
rect 17972 7976 18972 8004
rect 17972 7877 18000 7976
rect 18966 7964 18972 7976
rect 19024 7964 19030 8016
rect 20530 8004 20536 8016
rect 19352 7976 20208 8004
rect 18233 7939 18291 7945
rect 18233 7905 18245 7939
rect 18279 7936 18291 7939
rect 18414 7936 18420 7948
rect 18279 7908 18420 7936
rect 18279 7905 18291 7908
rect 18233 7899 18291 7905
rect 18414 7896 18420 7908
rect 18472 7896 18478 7948
rect 17543 7840 17908 7868
rect 17957 7871 18015 7877
rect 17543 7837 17555 7840
rect 17497 7831 17555 7837
rect 17957 7837 17969 7871
rect 18003 7837 18015 7871
rect 17957 7831 18015 7837
rect 18506 7828 18512 7880
rect 18564 7828 18570 7880
rect 18966 7828 18972 7880
rect 19024 7868 19030 7880
rect 19242 7868 19248 7880
rect 19024 7840 19248 7868
rect 19024 7828 19030 7840
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 17402 7800 17408 7812
rect 13955 7772 15056 7800
rect 15120 7772 15700 7800
rect 15948 7772 17408 7800
rect 13955 7769 13967 7772
rect 13909 7763 13967 7769
rect 11900 7704 13860 7732
rect 14093 7735 14151 7741
rect 14093 7701 14105 7735
rect 14139 7732 14151 7735
rect 14182 7732 14188 7744
rect 14139 7704 14188 7732
rect 14139 7701 14151 7704
rect 14093 7695 14151 7701
rect 14182 7692 14188 7704
rect 14240 7692 14246 7744
rect 14366 7692 14372 7744
rect 14424 7732 14430 7744
rect 15120 7732 15148 7772
rect 14424 7704 15148 7732
rect 14424 7692 14430 7704
rect 15194 7692 15200 7744
rect 15252 7692 15258 7744
rect 15672 7732 15700 7772
rect 17402 7760 17408 7772
rect 17460 7760 17466 7812
rect 18322 7760 18328 7812
rect 18380 7800 18386 7812
rect 19352 7800 19380 7976
rect 20180 7945 20208 7976
rect 20272 7976 20536 8004
rect 19981 7939 20039 7945
rect 19981 7905 19993 7939
rect 20027 7936 20039 7939
rect 20165 7939 20223 7945
rect 20027 7908 20116 7936
rect 20027 7905 20039 7908
rect 19981 7899 20039 7905
rect 19794 7868 19800 7880
rect 19429 7847 19487 7853
rect 19429 7813 19441 7847
rect 19475 7844 19487 7847
rect 19628 7844 19800 7868
rect 19475 7840 19800 7844
rect 19475 7816 19656 7840
rect 19794 7828 19800 7840
rect 19852 7828 19858 7880
rect 19886 7828 19892 7880
rect 19944 7864 19950 7880
rect 20088 7868 20116 7908
rect 20165 7905 20177 7939
rect 20211 7905 20223 7939
rect 20165 7899 20223 7905
rect 20272 7868 20300 7976
rect 20530 7964 20536 7976
rect 20588 7964 20594 8016
rect 20622 7964 20628 8016
rect 20680 7964 20686 8016
rect 21634 7964 21640 8016
rect 21692 7964 21698 8016
rect 22097 8007 22155 8013
rect 22097 7973 22109 8007
rect 22143 8004 22155 8007
rect 22186 8004 22192 8016
rect 22143 7976 22192 8004
rect 22143 7973 22155 7976
rect 22097 7967 22155 7973
rect 22186 7964 22192 7976
rect 22244 7964 22250 8016
rect 22296 7976 22600 8004
rect 21018 7939 21076 7945
rect 21018 7936 21030 7939
rect 20364 7908 21030 7936
rect 20364 7880 20392 7908
rect 21018 7905 21030 7908
rect 21064 7905 21076 7939
rect 21018 7899 21076 7905
rect 21177 7939 21235 7945
rect 21177 7905 21189 7939
rect 21223 7936 21235 7939
rect 21542 7936 21548 7948
rect 21223 7908 21548 7936
rect 21223 7905 21235 7908
rect 21177 7899 21235 7905
rect 21542 7896 21548 7908
rect 21600 7896 21606 7948
rect 21652 7936 21680 7964
rect 22296 7936 22324 7976
rect 22572 7948 22600 7976
rect 21652 7908 22324 7936
rect 22373 7939 22431 7945
rect 22373 7905 22385 7939
rect 22419 7936 22431 7939
rect 22419 7908 22508 7936
rect 22419 7905 22431 7908
rect 22373 7899 22431 7905
rect 19944 7836 19985 7864
rect 20088 7840 20300 7868
rect 19944 7828 19950 7836
rect 19889 7827 19947 7828
rect 19475 7813 19487 7816
rect 19429 7807 19487 7813
rect 18380 7772 19380 7800
rect 18380 7760 18386 7772
rect 16206 7732 16212 7744
rect 15672 7704 16212 7732
rect 16206 7692 16212 7704
rect 16264 7732 16270 7744
rect 16390 7732 16396 7744
rect 16264 7704 16396 7732
rect 16264 7692 16270 7704
rect 16390 7692 16396 7704
rect 16448 7692 16454 7744
rect 17129 7735 17187 7741
rect 17129 7701 17141 7735
rect 17175 7732 17187 7735
rect 17218 7732 17224 7744
rect 17175 7704 17224 7732
rect 17175 7701 17187 7704
rect 17129 7695 17187 7701
rect 17218 7692 17224 7704
rect 17276 7692 17282 7744
rect 17586 7692 17592 7744
rect 17644 7692 17650 7744
rect 18141 7735 18199 7741
rect 18141 7701 18153 7735
rect 18187 7732 18199 7735
rect 19334 7732 19340 7744
rect 18187 7704 19340 7732
rect 18187 7701 18199 7704
rect 18141 7695 18199 7701
rect 19334 7692 19340 7704
rect 19392 7692 19398 7744
rect 19613 7735 19671 7741
rect 19613 7701 19625 7735
rect 19659 7732 19671 7735
rect 20088 7732 20116 7840
rect 20346 7828 20352 7880
rect 20404 7828 20410 7880
rect 20898 7828 20904 7880
rect 20956 7828 20962 7880
rect 22002 7828 22008 7880
rect 22060 7868 22066 7880
rect 22281 7871 22339 7877
rect 22281 7868 22293 7871
rect 22060 7840 22293 7868
rect 22060 7828 22066 7840
rect 22281 7837 22293 7840
rect 22327 7837 22339 7871
rect 22281 7831 22339 7837
rect 22094 7760 22100 7812
rect 22152 7800 22158 7812
rect 22370 7800 22376 7812
rect 22152 7772 22376 7800
rect 22152 7760 22158 7772
rect 22370 7760 22376 7772
rect 22428 7800 22434 7812
rect 22480 7800 22508 7908
rect 22554 7896 22560 7948
rect 22612 7896 22618 7948
rect 22922 7896 22928 7948
rect 22980 7936 22986 7948
rect 23017 7939 23075 7945
rect 23017 7936 23029 7939
rect 22980 7908 23029 7936
rect 22980 7896 22986 7908
rect 23017 7905 23029 7908
rect 23063 7905 23075 7939
rect 23017 7899 23075 7905
rect 23106 7896 23112 7948
rect 23164 7936 23170 7948
rect 23293 7939 23351 7945
rect 23293 7936 23305 7939
rect 23164 7908 23305 7936
rect 23164 7896 23170 7908
rect 23293 7905 23305 7908
rect 23339 7905 23351 7939
rect 23293 7899 23351 7905
rect 23431 7939 23489 7945
rect 23431 7905 23443 7939
rect 23477 7936 23489 7939
rect 23952 7936 23980 8044
rect 24949 8041 24961 8044
rect 24995 8041 25007 8075
rect 24949 8035 25007 8041
rect 26237 8075 26295 8081
rect 26237 8041 26249 8075
rect 26283 8072 26295 8075
rect 30374 8072 30380 8084
rect 26283 8044 30380 8072
rect 26283 8041 26295 8044
rect 26237 8035 26295 8041
rect 30374 8032 30380 8044
rect 30432 8032 30438 8084
rect 30466 8032 30472 8084
rect 30524 8072 30530 8084
rect 31662 8072 31668 8084
rect 30524 8044 31668 8072
rect 30524 8032 30530 8044
rect 31662 8032 31668 8044
rect 31720 8032 31726 8084
rect 32306 8032 32312 8084
rect 32364 8072 32370 8084
rect 33229 8075 33287 8081
rect 33229 8072 33241 8075
rect 32364 8044 33241 8072
rect 32364 8032 32370 8044
rect 33229 8041 33241 8044
rect 33275 8041 33287 8075
rect 33229 8035 33287 8041
rect 33594 8032 33600 8084
rect 33652 8072 33658 8084
rect 33781 8075 33839 8081
rect 33781 8072 33793 8075
rect 33652 8044 33793 8072
rect 33652 8032 33658 8044
rect 33781 8041 33793 8044
rect 33827 8041 33839 8075
rect 33781 8035 33839 8041
rect 34422 8032 34428 8084
rect 34480 8072 34486 8084
rect 34793 8075 34851 8081
rect 34793 8072 34805 8075
rect 34480 8044 34805 8072
rect 34480 8032 34486 8044
rect 34793 8041 34805 8044
rect 34839 8041 34851 8075
rect 34793 8035 34851 8041
rect 35526 8032 35532 8084
rect 35584 8072 35590 8084
rect 35713 8075 35771 8081
rect 35713 8072 35725 8075
rect 35584 8044 35725 8072
rect 35584 8032 35590 8044
rect 35713 8041 35725 8044
rect 35759 8041 35771 8075
rect 35713 8035 35771 8041
rect 36078 8032 36084 8084
rect 36136 8072 36142 8084
rect 36265 8075 36323 8081
rect 36265 8072 36277 8075
rect 36136 8044 36277 8072
rect 36136 8032 36142 8044
rect 36265 8041 36277 8044
rect 36311 8041 36323 8075
rect 36265 8035 36323 8041
rect 36630 8032 36636 8084
rect 36688 8072 36694 8084
rect 36909 8075 36967 8081
rect 36909 8072 36921 8075
rect 36688 8044 36921 8072
rect 36688 8032 36694 8044
rect 36909 8041 36921 8044
rect 36955 8041 36967 8075
rect 36909 8035 36967 8041
rect 37274 8032 37280 8084
rect 37332 8032 37338 8084
rect 37826 8032 37832 8084
rect 37884 8072 37890 8084
rect 38197 8075 38255 8081
rect 38197 8072 38209 8075
rect 37884 8044 38209 8072
rect 37884 8032 37890 8044
rect 38197 8041 38209 8044
rect 38243 8041 38255 8075
rect 38197 8035 38255 8041
rect 38654 8032 38660 8084
rect 38712 8032 38718 8084
rect 24026 7964 24032 8016
rect 24084 7964 24090 8016
rect 27430 7964 27436 8016
rect 27488 7964 27494 8016
rect 28353 8007 28411 8013
rect 28353 7973 28365 8007
rect 28399 7973 28411 8007
rect 28353 7967 28411 7973
rect 23477 7908 23980 7936
rect 24044 7936 24072 7964
rect 24044 7908 24716 7936
rect 23477 7905 23489 7908
rect 23431 7899 23489 7905
rect 23566 7828 23572 7880
rect 23624 7828 23630 7880
rect 24213 7871 24271 7877
rect 24213 7837 24225 7871
rect 24259 7868 24271 7871
rect 24394 7868 24400 7880
rect 24259 7840 24400 7868
rect 24259 7837 24271 7840
rect 24213 7831 24271 7837
rect 24394 7828 24400 7840
rect 24452 7828 24458 7880
rect 24578 7828 24584 7880
rect 24636 7828 24642 7880
rect 24688 7877 24716 7908
rect 24854 7896 24860 7948
rect 24912 7936 24918 7948
rect 25225 7939 25283 7945
rect 25225 7936 25237 7939
rect 24912 7908 25237 7936
rect 24912 7896 24918 7908
rect 25225 7905 25237 7908
rect 25271 7905 25283 7939
rect 28368 7936 28396 7967
rect 32398 7964 32404 8016
rect 32456 7964 32462 8016
rect 35069 8007 35127 8013
rect 35069 8004 35081 8007
rect 34992 7976 35081 8004
rect 30745 7939 30803 7945
rect 30745 7936 30757 7939
rect 25225 7899 25283 7905
rect 27448 7908 28396 7936
rect 30300 7908 30757 7936
rect 24673 7871 24731 7877
rect 24673 7837 24685 7871
rect 24719 7837 24731 7871
rect 24673 7831 24731 7837
rect 25133 7871 25191 7877
rect 25133 7837 25145 7871
rect 25179 7837 25191 7871
rect 25133 7831 25191 7837
rect 25148 7800 25176 7831
rect 22428 7772 22508 7800
rect 24228 7772 25176 7800
rect 25240 7800 25268 7899
rect 25501 7871 25559 7877
rect 25501 7837 25513 7871
rect 25547 7868 25559 7871
rect 25590 7868 25596 7880
rect 25547 7840 25596 7868
rect 25547 7837 25559 7840
rect 25501 7831 25559 7837
rect 25590 7828 25596 7840
rect 25648 7828 25654 7880
rect 26786 7828 26792 7880
rect 26844 7868 26850 7880
rect 27065 7871 27123 7877
rect 27065 7868 27077 7871
rect 26844 7840 27077 7868
rect 26844 7828 26850 7840
rect 27065 7837 27077 7840
rect 27111 7837 27123 7871
rect 27065 7831 27123 7837
rect 27154 7828 27160 7880
rect 27212 7868 27218 7880
rect 27338 7868 27344 7880
rect 27212 7840 27344 7868
rect 27212 7828 27218 7840
rect 27338 7828 27344 7840
rect 27396 7828 27402 7880
rect 25240 7772 26464 7800
rect 22428 7760 22434 7772
rect 24228 7744 24256 7772
rect 19659 7704 20116 7732
rect 21821 7735 21879 7741
rect 19659 7701 19671 7704
rect 19613 7695 19671 7701
rect 21821 7701 21833 7735
rect 21867 7732 21879 7735
rect 22002 7732 22008 7744
rect 21867 7704 22008 7732
rect 21867 7701 21879 7704
rect 21821 7695 21879 7701
rect 22002 7692 22008 7704
rect 22060 7692 22066 7744
rect 22186 7692 22192 7744
rect 22244 7732 22250 7744
rect 22830 7732 22836 7744
rect 22244 7704 22836 7732
rect 22244 7692 22250 7704
rect 22830 7692 22836 7704
rect 22888 7692 22894 7744
rect 24210 7692 24216 7744
rect 24268 7692 24274 7744
rect 24302 7692 24308 7744
rect 24360 7732 24366 7744
rect 24397 7735 24455 7741
rect 24397 7732 24409 7735
rect 24360 7704 24409 7732
rect 24360 7692 24366 7704
rect 24397 7701 24409 7704
rect 24443 7701 24455 7735
rect 24397 7695 24455 7701
rect 24857 7735 24915 7741
rect 24857 7701 24869 7735
rect 24903 7732 24915 7735
rect 25406 7732 25412 7744
rect 24903 7704 25412 7732
rect 24903 7701 24915 7704
rect 24857 7695 24915 7701
rect 25406 7692 25412 7704
rect 25464 7692 25470 7744
rect 26326 7692 26332 7744
rect 26384 7692 26390 7744
rect 26436 7732 26464 7772
rect 26602 7760 26608 7812
rect 26660 7800 26666 7812
rect 27448 7800 27476 7908
rect 27614 7828 27620 7880
rect 27672 7828 27678 7880
rect 29086 7828 29092 7880
rect 29144 7828 29150 7880
rect 29362 7828 29368 7880
rect 29420 7828 29426 7880
rect 29454 7828 29460 7880
rect 29512 7868 29518 7880
rect 29641 7871 29699 7877
rect 29641 7868 29653 7871
rect 29512 7840 29653 7868
rect 29512 7828 29518 7840
rect 29641 7837 29653 7840
rect 29687 7837 29699 7871
rect 29641 7831 29699 7837
rect 29822 7828 29828 7880
rect 29880 7868 29886 7880
rect 29917 7871 29975 7877
rect 29917 7868 29929 7871
rect 29880 7840 29929 7868
rect 29880 7828 29886 7840
rect 29917 7837 29929 7840
rect 29963 7837 29975 7871
rect 30300 7868 30328 7908
rect 30745 7905 30757 7908
rect 30791 7905 30803 7939
rect 30745 7899 30803 7905
rect 31846 7896 31852 7948
rect 31904 7936 31910 7948
rect 31904 7908 33180 7936
rect 31904 7896 31910 7908
rect 29917 7831 29975 7837
rect 30024 7864 30144 7868
rect 30208 7864 30328 7868
rect 30024 7840 30328 7864
rect 31021 7871 31079 7877
rect 26660 7772 27476 7800
rect 26660 7760 26666 7772
rect 27798 7760 27804 7812
rect 27856 7800 27862 7812
rect 27985 7803 28043 7809
rect 27985 7800 27997 7803
rect 27856 7772 27997 7800
rect 27856 7760 27862 7772
rect 27985 7769 27997 7772
rect 28031 7769 28043 7803
rect 27985 7763 28043 7769
rect 28534 7760 28540 7812
rect 28592 7800 28598 7812
rect 30024 7800 30052 7840
rect 30116 7836 30236 7840
rect 31021 7837 31033 7871
rect 31067 7868 31079 7871
rect 31386 7868 31392 7880
rect 31067 7840 31392 7868
rect 31067 7837 31079 7840
rect 31021 7831 31079 7837
rect 31386 7828 31392 7840
rect 31444 7828 31450 7880
rect 31754 7828 31760 7880
rect 31812 7868 31818 7880
rect 32033 7871 32091 7877
rect 32033 7868 32045 7871
rect 31812 7840 32045 7868
rect 31812 7828 31818 7840
rect 32033 7837 32045 7840
rect 32079 7837 32091 7871
rect 32033 7831 32091 7837
rect 32309 7871 32367 7877
rect 32309 7837 32321 7871
rect 32355 7837 32367 7871
rect 32309 7831 32367 7837
rect 28592 7772 30052 7800
rect 30576 7772 31064 7800
rect 28592 7760 28598 7772
rect 28077 7735 28135 7741
rect 28077 7732 28089 7735
rect 26436 7704 28089 7732
rect 28077 7701 28089 7704
rect 28123 7732 28135 7735
rect 28994 7732 29000 7744
rect 28123 7704 29000 7732
rect 28123 7701 28135 7704
rect 28077 7695 28135 7701
rect 28994 7692 29000 7704
rect 29052 7732 29058 7744
rect 30576 7732 30604 7772
rect 29052 7704 30604 7732
rect 30653 7735 30711 7741
rect 29052 7692 29058 7704
rect 30653 7701 30665 7735
rect 30699 7732 30711 7735
rect 30742 7732 30748 7744
rect 30699 7704 30748 7732
rect 30699 7701 30711 7704
rect 30653 7695 30711 7701
rect 30742 7692 30748 7704
rect 30800 7692 30806 7744
rect 31036 7732 31064 7772
rect 31110 7760 31116 7812
rect 31168 7800 31174 7812
rect 32324 7800 32352 7831
rect 32398 7828 32404 7880
rect 32456 7868 32462 7880
rect 32585 7871 32643 7877
rect 32585 7868 32597 7871
rect 32456 7840 32597 7868
rect 32456 7828 32462 7840
rect 32585 7837 32597 7840
rect 32631 7837 32643 7871
rect 32585 7831 32643 7837
rect 32674 7828 32680 7880
rect 32732 7868 32738 7880
rect 33152 7877 33180 7908
rect 32861 7871 32919 7877
rect 32861 7868 32873 7871
rect 32732 7840 32873 7868
rect 32732 7828 32738 7840
rect 32861 7837 32873 7840
rect 32907 7837 32919 7871
rect 32861 7831 32919 7837
rect 33137 7871 33195 7877
rect 33137 7837 33149 7871
rect 33183 7837 33195 7871
rect 33137 7831 33195 7837
rect 33413 7871 33471 7877
rect 33413 7837 33425 7871
rect 33459 7868 33471 7871
rect 33870 7868 33876 7880
rect 33459 7840 33876 7868
rect 33459 7837 33471 7840
rect 33413 7831 33471 7837
rect 33870 7828 33876 7840
rect 33928 7828 33934 7880
rect 33965 7871 34023 7877
rect 33965 7837 33977 7871
rect 34011 7837 34023 7871
rect 33965 7831 34023 7837
rect 31168 7772 32352 7800
rect 33980 7800 34008 7831
rect 34146 7828 34152 7880
rect 34204 7828 34210 7880
rect 34992 7877 35020 7976
rect 35069 7973 35081 7976
rect 35115 7973 35127 8007
rect 35069 7967 35127 7973
rect 35342 7964 35348 8016
rect 35400 8004 35406 8016
rect 35400 7976 37228 8004
rect 35400 7964 35406 7976
rect 36078 7936 36084 7948
rect 35084 7908 36084 7936
rect 34977 7871 35035 7877
rect 34977 7837 34989 7871
rect 35023 7837 35035 7871
rect 34977 7831 35035 7837
rect 35084 7800 35112 7908
rect 36078 7896 36084 7908
rect 36136 7896 36142 7948
rect 36170 7896 36176 7948
rect 36228 7936 36234 7948
rect 36228 7908 37136 7936
rect 36228 7896 36234 7908
rect 35158 7828 35164 7880
rect 35216 7868 35222 7880
rect 35253 7871 35311 7877
rect 35253 7868 35265 7871
rect 35216 7840 35265 7868
rect 35216 7828 35222 7840
rect 35253 7837 35265 7840
rect 35299 7837 35311 7871
rect 35253 7831 35311 7837
rect 35345 7871 35403 7877
rect 35345 7837 35357 7871
rect 35391 7868 35403 7871
rect 35526 7868 35532 7880
rect 35391 7840 35532 7868
rect 35391 7837 35403 7840
rect 35345 7831 35403 7837
rect 35526 7828 35532 7840
rect 35584 7828 35590 7880
rect 35894 7828 35900 7880
rect 35952 7828 35958 7880
rect 36354 7828 36360 7880
rect 36412 7868 36418 7880
rect 36449 7871 36507 7877
rect 36449 7868 36461 7871
rect 36412 7840 36461 7868
rect 36412 7828 36418 7840
rect 36449 7837 36461 7840
rect 36495 7837 36507 7871
rect 36449 7831 36507 7837
rect 36630 7828 36636 7880
rect 36688 7868 36694 7880
rect 37108 7877 37136 7908
rect 36725 7871 36783 7877
rect 36725 7868 36737 7871
rect 36688 7840 36737 7868
rect 36688 7828 36694 7840
rect 36725 7837 36737 7840
rect 36771 7837 36783 7871
rect 36725 7831 36783 7837
rect 37093 7871 37151 7877
rect 37093 7837 37105 7871
rect 37139 7837 37151 7871
rect 37200 7868 37228 7976
rect 37734 7964 37740 8016
rect 37792 8004 37798 8016
rect 38013 8007 38071 8013
rect 38013 8004 38025 8007
rect 37792 7976 38025 8004
rect 37792 7964 37798 7976
rect 38013 7973 38025 7976
rect 38059 7973 38071 8007
rect 38013 7967 38071 7973
rect 37366 7896 37372 7948
rect 37424 7936 37430 7948
rect 37424 7908 38424 7936
rect 37424 7896 37430 7908
rect 37553 7871 37611 7877
rect 37553 7868 37565 7871
rect 37200 7840 37565 7868
rect 37093 7831 37151 7837
rect 37553 7837 37565 7840
rect 37599 7837 37611 7871
rect 37553 7831 37611 7837
rect 37826 7828 37832 7880
rect 37884 7828 37890 7880
rect 38396 7877 38424 7908
rect 38381 7871 38439 7877
rect 38381 7837 38393 7871
rect 38427 7837 38439 7871
rect 38381 7831 38439 7837
rect 38470 7828 38476 7880
rect 38528 7828 38534 7880
rect 38838 7828 38844 7880
rect 38896 7828 38902 7880
rect 39209 7871 39267 7877
rect 39209 7837 39221 7871
rect 39255 7837 39267 7871
rect 39209 7831 39267 7837
rect 33980 7772 35112 7800
rect 31168 7760 31174 7772
rect 37458 7760 37464 7812
rect 37516 7800 37522 7812
rect 39224 7800 39252 7831
rect 37516 7772 39252 7800
rect 37516 7760 37522 7772
rect 31662 7732 31668 7744
rect 31036 7704 31668 7732
rect 31662 7692 31668 7704
rect 31720 7692 31726 7744
rect 31754 7692 31760 7744
rect 31812 7692 31818 7744
rect 31846 7692 31852 7744
rect 31904 7692 31910 7744
rect 32122 7692 32128 7744
rect 32180 7692 32186 7744
rect 32674 7692 32680 7744
rect 32732 7692 32738 7744
rect 32950 7692 32956 7744
rect 33008 7692 33014 7744
rect 34330 7692 34336 7744
rect 34388 7692 34394 7744
rect 35529 7735 35587 7741
rect 35529 7701 35541 7735
rect 35575 7732 35587 7735
rect 35618 7732 35624 7744
rect 35575 7704 35624 7732
rect 35575 7701 35587 7704
rect 35529 7695 35587 7701
rect 35618 7692 35624 7704
rect 35676 7692 35682 7744
rect 36354 7692 36360 7744
rect 36412 7732 36418 7744
rect 37369 7735 37427 7741
rect 37369 7732 37381 7735
rect 36412 7704 37381 7732
rect 36412 7692 36418 7704
rect 37369 7701 37381 7704
rect 37415 7701 37427 7735
rect 37369 7695 37427 7701
rect 37550 7692 37556 7744
rect 37608 7732 37614 7744
rect 38194 7732 38200 7744
rect 37608 7704 38200 7732
rect 37608 7692 37614 7704
rect 38194 7692 38200 7704
rect 38252 7692 38258 7744
rect 38930 7692 38936 7744
rect 38988 7732 38994 7744
rect 39025 7735 39083 7741
rect 39025 7732 39037 7735
rect 38988 7704 39037 7732
rect 38988 7692 38994 7704
rect 39025 7701 39037 7704
rect 39071 7701 39083 7735
rect 39025 7695 39083 7701
rect 39390 7692 39396 7744
rect 39448 7692 39454 7744
rect 1104 7642 39836 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 39010 7642
rect 39062 7590 39074 7642
rect 39126 7590 39138 7642
rect 39190 7590 39202 7642
rect 39254 7590 39266 7642
rect 39318 7590 39836 7642
rect 1104 7568 39836 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7528 1639 7531
rect 5258 7528 5264 7540
rect 1627 7500 5264 7528
rect 1627 7497 1639 7500
rect 1581 7491 1639 7497
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 5350 7488 5356 7540
rect 5408 7488 5414 7540
rect 5813 7531 5871 7537
rect 5813 7497 5825 7531
rect 5859 7528 5871 7531
rect 5859 7500 7052 7528
rect 5859 7497 5871 7500
rect 5813 7491 5871 7497
rect 934 7420 940 7472
rect 992 7460 998 7472
rect 1857 7463 1915 7469
rect 1857 7460 1869 7463
rect 992 7432 1869 7460
rect 992 7420 998 7432
rect 1857 7429 1869 7432
rect 1903 7429 1915 7463
rect 1857 7423 1915 7429
rect 1946 7420 1952 7472
rect 2004 7460 2010 7472
rect 2593 7463 2651 7469
rect 2593 7460 2605 7463
rect 2004 7432 2605 7460
rect 2004 7420 2010 7432
rect 2593 7429 2605 7432
rect 2639 7429 2651 7463
rect 2593 7423 2651 7429
rect 3145 7463 3203 7469
rect 3145 7429 3157 7463
rect 3191 7460 3203 7463
rect 4154 7460 4160 7472
rect 3191 7432 4160 7460
rect 3191 7429 3203 7432
rect 3145 7423 3203 7429
rect 4154 7420 4160 7432
rect 4212 7420 4218 7472
rect 4890 7420 4896 7472
rect 4948 7460 4954 7472
rect 6086 7460 6092 7472
rect 4948 7432 6092 7460
rect 4948 7420 4954 7432
rect 6086 7420 6092 7432
rect 6144 7420 6150 7472
rect 6730 7420 6736 7472
rect 6788 7420 6794 7472
rect 7024 7460 7052 7500
rect 7098 7488 7104 7540
rect 7156 7528 7162 7540
rect 7285 7531 7343 7537
rect 7285 7528 7297 7531
rect 7156 7500 7297 7528
rect 7156 7488 7162 7500
rect 7285 7497 7297 7500
rect 7331 7497 7343 7531
rect 7285 7491 7343 7497
rect 7558 7488 7564 7540
rect 7616 7528 7622 7540
rect 7616 7500 9720 7528
rect 7616 7488 7622 7500
rect 9692 7460 9720 7500
rect 9950 7488 9956 7540
rect 10008 7528 10014 7540
rect 11330 7528 11336 7540
rect 10008 7500 11336 7528
rect 10008 7488 10014 7500
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 11422 7488 11428 7540
rect 11480 7528 11486 7540
rect 11885 7531 11943 7537
rect 11480 7500 11836 7528
rect 11480 7488 11486 7500
rect 11606 7460 11612 7472
rect 7024 7432 8156 7460
rect 9692 7432 11612 7460
rect 750 7352 756 7404
rect 808 7392 814 7404
rect 1489 7395 1547 7401
rect 1489 7392 1501 7395
rect 808 7364 1501 7392
rect 808 7352 814 7364
rect 1489 7361 1501 7364
rect 1535 7361 1547 7395
rect 1489 7355 1547 7361
rect 2225 7395 2283 7401
rect 2225 7361 2237 7395
rect 2271 7361 2283 7395
rect 2225 7355 2283 7361
rect 1118 7284 1124 7336
rect 1176 7324 1182 7336
rect 2240 7324 2268 7355
rect 2958 7352 2964 7404
rect 3016 7352 3022 7404
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7361 5227 7395
rect 6825 7395 6883 7401
rect 6825 7392 6837 7395
rect 5169 7355 5227 7361
rect 5920 7364 6837 7392
rect 1176 7296 2268 7324
rect 2409 7327 2467 7333
rect 1176 7284 1182 7296
rect 2409 7293 2421 7327
rect 2455 7324 2467 7327
rect 5074 7324 5080 7336
rect 2455 7296 5080 7324
rect 2455 7293 2467 7296
rect 2409 7287 2467 7293
rect 5074 7284 5080 7296
rect 5132 7284 5138 7336
rect 2041 7259 2099 7265
rect 2041 7225 2053 7259
rect 2087 7256 2099 7259
rect 3602 7256 3608 7268
rect 2087 7228 3608 7256
rect 2087 7225 2099 7228
rect 2041 7219 2099 7225
rect 3602 7216 3608 7228
rect 3660 7216 3666 7268
rect 5184 7256 5212 7355
rect 5810 7284 5816 7336
rect 5868 7324 5874 7336
rect 5920 7333 5948 7364
rect 6825 7361 6837 7364
rect 6871 7361 6883 7395
rect 6825 7355 6883 7361
rect 7098 7352 7104 7404
rect 7156 7392 7162 7404
rect 7469 7395 7527 7401
rect 7469 7392 7481 7395
rect 7156 7364 7481 7392
rect 7156 7352 7162 7364
rect 7469 7361 7481 7364
rect 7515 7361 7527 7395
rect 7469 7355 7527 7361
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7392 7803 7395
rect 8018 7392 8024 7404
rect 7791 7364 8024 7392
rect 7791 7361 7803 7364
rect 7745 7355 7803 7361
rect 5905 7327 5963 7333
rect 5905 7324 5917 7327
rect 5868 7296 5917 7324
rect 5868 7284 5874 7296
rect 5905 7293 5917 7296
rect 5951 7293 5963 7327
rect 5905 7287 5963 7293
rect 6086 7284 6092 7336
rect 6144 7284 6150 7336
rect 6917 7327 6975 7333
rect 6917 7293 6929 7327
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 6365 7259 6423 7265
rect 6365 7256 6377 7259
rect 5184 7228 6377 7256
rect 6365 7225 6377 7228
rect 6411 7225 6423 7259
rect 6365 7219 6423 7225
rect 6454 7216 6460 7268
rect 6512 7256 6518 7268
rect 6932 7256 6960 7287
rect 7006 7284 7012 7336
rect 7064 7324 7070 7336
rect 7760 7324 7788 7355
rect 8018 7352 8024 7364
rect 8076 7352 8082 7404
rect 7064 7296 7788 7324
rect 8128 7324 8156 7432
rect 11606 7420 11612 7432
rect 11664 7420 11670 7472
rect 8662 7352 8668 7404
rect 8720 7352 8726 7404
rect 8938 7352 8944 7404
rect 8996 7352 9002 7404
rect 9766 7392 9772 7404
rect 9508 7364 9772 7392
rect 8803 7327 8861 7333
rect 8803 7324 8815 7327
rect 8128 7296 8815 7324
rect 7064 7284 7070 7296
rect 8803 7293 8815 7296
rect 8849 7324 8861 7327
rect 9508 7324 9536 7364
rect 9766 7352 9772 7364
rect 9824 7352 9830 7404
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7392 9919 7395
rect 10134 7392 10140 7404
rect 9907 7364 10140 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 10134 7352 10140 7364
rect 10192 7352 10198 7404
rect 10229 7395 10287 7401
rect 10229 7361 10241 7395
rect 10275 7392 10287 7395
rect 10275 7364 10640 7392
rect 10275 7361 10287 7364
rect 10229 7355 10287 7361
rect 8849 7296 9536 7324
rect 8849 7293 8861 7296
rect 8803 7287 8861 7293
rect 9674 7284 9680 7336
rect 9732 7284 9738 7336
rect 9950 7284 9956 7336
rect 10008 7284 10014 7336
rect 6512 7228 6960 7256
rect 6512 7216 6518 7228
rect 7742 7216 7748 7268
rect 7800 7256 7806 7268
rect 8021 7259 8079 7265
rect 8021 7256 8033 7259
rect 7800 7228 8033 7256
rect 7800 7216 7806 7228
rect 8021 7225 8033 7228
rect 8067 7225 8079 7259
rect 8021 7219 8079 7225
rect 9217 7259 9275 7265
rect 9217 7225 9229 7259
rect 9263 7225 9275 7259
rect 9217 7219 9275 7225
rect 2685 7191 2743 7197
rect 2685 7157 2697 7191
rect 2731 7188 2743 7191
rect 2866 7188 2872 7200
rect 2731 7160 2872 7188
rect 2731 7157 2743 7160
rect 2685 7151 2743 7157
rect 2866 7148 2872 7160
rect 2924 7148 2930 7200
rect 5445 7191 5503 7197
rect 5445 7157 5457 7191
rect 5491 7188 5503 7191
rect 5534 7188 5540 7200
rect 5491 7160 5540 7188
rect 5491 7157 5503 7160
rect 5445 7151 5503 7157
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 5994 7148 6000 7200
rect 6052 7188 6058 7200
rect 7098 7188 7104 7200
rect 6052 7160 7104 7188
rect 6052 7148 6058 7160
rect 7098 7148 7104 7160
rect 7156 7148 7162 7200
rect 7374 7148 7380 7200
rect 7432 7188 7438 7200
rect 7837 7191 7895 7197
rect 7837 7188 7849 7191
rect 7432 7160 7849 7188
rect 7432 7148 7438 7160
rect 7837 7157 7849 7160
rect 7883 7157 7895 7191
rect 7837 7151 7895 7157
rect 8478 7148 8484 7200
rect 8536 7188 8542 7200
rect 9232 7188 9260 7219
rect 9490 7216 9496 7268
rect 9548 7256 9554 7268
rect 9968 7256 9996 7284
rect 9548 7228 9996 7256
rect 9548 7216 9554 7228
rect 8536 7160 9260 7188
rect 8536 7148 8542 7160
rect 9306 7148 9312 7200
rect 9364 7188 9370 7200
rect 10612 7188 10640 7364
rect 11330 7352 11336 7404
rect 11388 7352 11394 7404
rect 11514 7392 11520 7404
rect 11440 7364 11520 7392
rect 11440 7324 11468 7364
rect 11514 7352 11520 7364
rect 11572 7352 11578 7404
rect 10980 7296 11468 7324
rect 11808 7324 11836 7500
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 12526 7528 12532 7540
rect 11931 7500 12532 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 12618 7488 12624 7540
rect 12676 7528 12682 7540
rect 13357 7531 13415 7537
rect 13357 7528 13369 7531
rect 12676 7500 13369 7528
rect 12676 7488 12682 7500
rect 13357 7497 13369 7500
rect 13403 7497 13415 7531
rect 13357 7491 13415 7497
rect 13446 7488 13452 7540
rect 13504 7528 13510 7540
rect 13633 7531 13691 7537
rect 13633 7528 13645 7531
rect 13504 7500 13645 7528
rect 13504 7488 13510 7500
rect 13633 7497 13645 7500
rect 13679 7497 13691 7531
rect 13633 7491 13691 7497
rect 14001 7531 14059 7537
rect 14001 7497 14013 7531
rect 14047 7528 14059 7531
rect 14274 7528 14280 7540
rect 14047 7500 14280 7528
rect 14047 7497 14059 7500
rect 14001 7491 14059 7497
rect 14274 7488 14280 7500
rect 14332 7488 14338 7540
rect 14826 7488 14832 7540
rect 14884 7528 14890 7540
rect 15013 7531 15071 7537
rect 15013 7528 15025 7531
rect 14884 7500 15025 7528
rect 14884 7488 14890 7500
rect 15013 7497 15025 7500
rect 15059 7497 15071 7531
rect 15013 7491 15071 7497
rect 15289 7531 15347 7537
rect 15289 7497 15301 7531
rect 15335 7528 15347 7531
rect 15470 7528 15476 7540
rect 15335 7500 15476 7528
rect 15335 7497 15347 7500
rect 15289 7491 15347 7497
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 15930 7488 15936 7540
rect 15988 7528 15994 7540
rect 16209 7531 16267 7537
rect 16209 7528 16221 7531
rect 15988 7500 16221 7528
rect 15988 7488 15994 7500
rect 16209 7497 16221 7500
rect 16255 7497 16267 7531
rect 17037 7531 17095 7537
rect 17037 7528 17049 7531
rect 16209 7491 16267 7497
rect 16408 7500 17049 7528
rect 12805 7463 12863 7469
rect 12805 7460 12817 7463
rect 12452 7432 12817 7460
rect 12452 7404 12480 7432
rect 12805 7429 12817 7432
rect 12851 7460 12863 7463
rect 13078 7460 13084 7472
rect 12851 7432 13084 7460
rect 12851 7429 12863 7432
rect 12805 7423 12863 7429
rect 13078 7420 13084 7432
rect 13136 7420 13142 7472
rect 13262 7420 13268 7472
rect 13320 7460 13326 7472
rect 14461 7463 14519 7469
rect 14461 7460 14473 7463
rect 13320 7432 14473 7460
rect 13320 7420 13326 7432
rect 14461 7429 14473 7432
rect 14507 7429 14519 7463
rect 14461 7423 14519 7429
rect 15746 7420 15752 7472
rect 15804 7460 15810 7472
rect 16408 7460 16436 7500
rect 17037 7497 17049 7500
rect 17083 7497 17095 7531
rect 17037 7491 17095 7497
rect 17313 7531 17371 7537
rect 17313 7497 17325 7531
rect 17359 7497 17371 7531
rect 17313 7491 17371 7497
rect 17681 7531 17739 7537
rect 17681 7497 17693 7531
rect 17727 7528 17739 7531
rect 18046 7528 18052 7540
rect 17727 7500 18052 7528
rect 17727 7497 17739 7500
rect 17681 7491 17739 7497
rect 17328 7460 17356 7491
rect 18046 7488 18052 7500
rect 18104 7488 18110 7540
rect 18322 7488 18328 7540
rect 18380 7488 18386 7540
rect 18601 7531 18659 7537
rect 18601 7497 18613 7531
rect 18647 7497 18659 7531
rect 18601 7491 18659 7497
rect 19061 7531 19119 7537
rect 19061 7497 19073 7531
rect 19107 7528 19119 7531
rect 19518 7528 19524 7540
rect 19107 7500 19524 7528
rect 19107 7497 19119 7500
rect 19061 7491 19119 7497
rect 15804 7432 16436 7460
rect 16960 7432 17356 7460
rect 15804 7420 15810 7432
rect 11977 7395 12035 7401
rect 11977 7361 11989 7395
rect 12023 7392 12035 7395
rect 12434 7392 12440 7404
rect 12023 7364 12440 7392
rect 12023 7361 12035 7364
rect 11977 7355 12035 7361
rect 12434 7352 12440 7364
rect 12492 7352 12498 7404
rect 12618 7352 12624 7404
rect 12676 7392 12682 7404
rect 12713 7395 12771 7401
rect 12713 7392 12725 7395
rect 12676 7364 12725 7392
rect 12676 7352 12682 7364
rect 12713 7361 12725 7364
rect 12759 7361 12771 7395
rect 13173 7395 13231 7401
rect 13173 7392 13185 7395
rect 12713 7355 12771 7361
rect 12820 7364 13185 7392
rect 12820 7336 12848 7364
rect 13173 7361 13185 7364
rect 13219 7361 13231 7395
rect 13173 7355 13231 7361
rect 13814 7352 13820 7404
rect 13872 7352 13878 7404
rect 14369 7395 14427 7401
rect 14369 7361 14381 7395
rect 14415 7361 14427 7395
rect 14369 7355 14427 7361
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7361 15255 7395
rect 15197 7355 15255 7361
rect 12069 7327 12127 7333
rect 12069 7324 12081 7327
rect 11808 7296 12081 7324
rect 10980 7265 11008 7296
rect 12069 7293 12081 7296
rect 12115 7293 12127 7327
rect 12069 7287 12127 7293
rect 12158 7284 12164 7336
rect 12216 7324 12222 7336
rect 12216 7296 12480 7324
rect 12216 7284 12222 7296
rect 10965 7259 11023 7265
rect 10965 7225 10977 7259
rect 11011 7225 11023 7259
rect 10965 7219 11023 7225
rect 11054 7216 11060 7268
rect 11112 7256 11118 7268
rect 11149 7259 11207 7265
rect 11149 7256 11161 7259
rect 11112 7228 11161 7256
rect 11112 7216 11118 7228
rect 11149 7225 11161 7228
rect 11195 7225 11207 7259
rect 12345 7259 12403 7265
rect 12345 7256 12357 7259
rect 11149 7219 11207 7225
rect 11440 7228 12357 7256
rect 11440 7200 11468 7228
rect 12345 7225 12357 7228
rect 12391 7225 12403 7259
rect 12452 7256 12480 7296
rect 12802 7284 12808 7336
rect 12860 7284 12866 7336
rect 12897 7327 12955 7333
rect 12897 7293 12909 7327
rect 12943 7293 12955 7327
rect 12897 7287 12955 7293
rect 12912 7256 12940 7287
rect 13262 7284 13268 7336
rect 13320 7324 13326 7336
rect 14090 7324 14096 7336
rect 13320 7296 14096 7324
rect 13320 7284 13326 7296
rect 14090 7284 14096 7296
rect 14148 7284 14154 7336
rect 12452 7228 12940 7256
rect 14384 7256 14412 7355
rect 14550 7284 14556 7336
rect 14608 7284 14614 7336
rect 15212 7324 15240 7355
rect 15470 7352 15476 7404
rect 15528 7352 15534 7404
rect 15562 7352 15568 7404
rect 15620 7392 15626 7404
rect 16025 7395 16083 7401
rect 16025 7392 16037 7395
rect 15620 7364 16037 7392
rect 15620 7352 15626 7364
rect 16025 7361 16037 7364
rect 16071 7361 16083 7395
rect 16025 7355 16083 7361
rect 16114 7352 16120 7404
rect 16172 7392 16178 7404
rect 16758 7392 16764 7404
rect 16172 7364 16764 7392
rect 16172 7352 16178 7364
rect 16758 7352 16764 7364
rect 16816 7352 16822 7404
rect 16960 7401 16988 7432
rect 17954 7420 17960 7472
rect 18012 7460 18018 7472
rect 18616 7460 18644 7491
rect 19518 7488 19524 7500
rect 19576 7488 19582 7540
rect 19628 7500 19840 7528
rect 18966 7460 18972 7472
rect 18012 7432 18644 7460
rect 18800 7432 18972 7460
rect 18012 7420 18018 7432
rect 16945 7395 17003 7401
rect 16945 7361 16957 7395
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 17218 7352 17224 7404
rect 17276 7352 17282 7404
rect 18141 7395 18199 7401
rect 18141 7361 18153 7395
rect 18187 7392 18199 7395
rect 18598 7392 18604 7404
rect 18187 7364 18604 7392
rect 18187 7361 18199 7364
rect 18141 7355 18199 7361
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 18800 7401 18828 7432
rect 18966 7420 18972 7432
rect 19024 7420 19030 7472
rect 19628 7460 19656 7500
rect 19076 7432 19656 7460
rect 19812 7460 19840 7500
rect 20438 7488 20444 7540
rect 20496 7488 20502 7540
rect 20530 7488 20536 7540
rect 20588 7528 20594 7540
rect 20993 7531 21051 7537
rect 20993 7528 21005 7531
rect 20588 7500 21005 7528
rect 20588 7488 20594 7500
rect 20993 7497 21005 7500
rect 21039 7497 21051 7531
rect 20993 7491 21051 7497
rect 22097 7531 22155 7537
rect 22097 7497 22109 7531
rect 22143 7528 22155 7531
rect 22738 7528 22744 7540
rect 22143 7500 22744 7528
rect 22143 7497 22155 7500
rect 22097 7491 22155 7497
rect 22738 7488 22744 7500
rect 22796 7488 22802 7540
rect 23201 7531 23259 7537
rect 23201 7497 23213 7531
rect 23247 7528 23259 7531
rect 23566 7528 23572 7540
rect 23247 7500 23572 7528
rect 23247 7497 23259 7500
rect 23201 7491 23259 7497
rect 23566 7488 23572 7500
rect 23624 7488 23630 7540
rect 24121 7531 24179 7537
rect 24121 7497 24133 7531
rect 24167 7528 24179 7531
rect 24578 7528 24584 7540
rect 24167 7500 24584 7528
rect 24167 7497 24179 7500
rect 24121 7491 24179 7497
rect 24578 7488 24584 7500
rect 24636 7488 24642 7540
rect 24670 7488 24676 7540
rect 24728 7528 24734 7540
rect 26786 7528 26792 7540
rect 24728 7500 26792 7528
rect 24728 7488 24734 7500
rect 26786 7488 26792 7500
rect 26844 7488 26850 7540
rect 27157 7531 27215 7537
rect 27157 7497 27169 7531
rect 27203 7528 27215 7531
rect 30466 7528 30472 7540
rect 27203 7500 30472 7528
rect 27203 7497 27215 7500
rect 27157 7491 27215 7497
rect 30466 7488 30472 7500
rect 30524 7488 30530 7540
rect 30558 7488 30564 7540
rect 30616 7488 30622 7540
rect 30834 7488 30840 7540
rect 30892 7528 30898 7540
rect 31110 7528 31116 7540
rect 30892 7500 31116 7528
rect 30892 7488 30898 7500
rect 31110 7488 31116 7500
rect 31168 7488 31174 7540
rect 31202 7488 31208 7540
rect 31260 7488 31266 7540
rect 31478 7488 31484 7540
rect 31536 7488 31542 7540
rect 31754 7488 31760 7540
rect 31812 7488 31818 7540
rect 32125 7531 32183 7537
rect 32125 7497 32137 7531
rect 32171 7528 32183 7531
rect 32398 7528 32404 7540
rect 32171 7500 32404 7528
rect 32171 7497 32183 7500
rect 32125 7491 32183 7497
rect 32398 7488 32404 7500
rect 32456 7488 32462 7540
rect 32493 7531 32551 7537
rect 32493 7497 32505 7531
rect 32539 7528 32551 7531
rect 32674 7528 32680 7540
rect 32539 7500 32680 7528
rect 32539 7497 32551 7500
rect 32493 7491 32551 7497
rect 32674 7488 32680 7500
rect 32732 7488 32738 7540
rect 35529 7531 35587 7537
rect 35529 7497 35541 7531
rect 35575 7528 35587 7531
rect 35802 7528 35808 7540
rect 35575 7500 35808 7528
rect 35575 7497 35587 7500
rect 35529 7491 35587 7497
rect 35802 7488 35808 7500
rect 35860 7488 35866 7540
rect 37090 7488 37096 7540
rect 37148 7528 37154 7540
rect 37461 7531 37519 7537
rect 37461 7528 37473 7531
rect 37148 7500 37473 7528
rect 37148 7488 37154 7500
rect 37461 7497 37473 7500
rect 37507 7497 37519 7531
rect 37461 7491 37519 7497
rect 38286 7488 38292 7540
rect 38344 7488 38350 7540
rect 38657 7531 38715 7537
rect 38657 7497 38669 7531
rect 38703 7528 38715 7531
rect 38746 7528 38752 7540
rect 38703 7500 38752 7528
rect 38703 7497 38715 7500
rect 38657 7491 38715 7497
rect 38746 7488 38752 7500
rect 38804 7488 38810 7540
rect 39025 7531 39083 7537
rect 39025 7497 39037 7531
rect 39071 7497 39083 7531
rect 39025 7491 39083 7497
rect 39393 7531 39451 7537
rect 39393 7497 39405 7531
rect 39439 7528 39451 7531
rect 39574 7528 39580 7540
rect 39439 7500 39580 7528
rect 39439 7497 39451 7500
rect 39393 7491 39451 7497
rect 22186 7460 22192 7472
rect 19812 7432 22192 7460
rect 18785 7395 18843 7401
rect 18785 7361 18797 7395
rect 18831 7361 18843 7395
rect 18785 7355 18843 7361
rect 18874 7352 18880 7404
rect 18932 7352 18938 7404
rect 19076 7392 19104 7432
rect 22186 7420 22192 7432
rect 22244 7420 22250 7472
rect 22370 7420 22376 7472
rect 22428 7460 22434 7472
rect 23753 7463 23811 7469
rect 23753 7460 23765 7463
rect 22428 7432 23765 7460
rect 22428 7420 22434 7432
rect 23753 7429 23765 7432
rect 23799 7429 23811 7463
rect 30576 7460 30604 7488
rect 31772 7460 31800 7488
rect 23753 7423 23811 7429
rect 24412 7432 29960 7460
rect 30576 7432 31340 7460
rect 31772 7432 32628 7460
rect 18984 7364 19104 7392
rect 16482 7324 16488 7336
rect 15212 7296 16488 7324
rect 16482 7284 16488 7296
rect 16540 7284 16546 7336
rect 16850 7284 16856 7336
rect 16908 7324 16914 7336
rect 17773 7327 17831 7333
rect 17773 7324 17785 7327
rect 16908 7296 17785 7324
rect 16908 7284 16914 7296
rect 17773 7293 17785 7296
rect 17819 7293 17831 7327
rect 17773 7287 17831 7293
rect 17862 7284 17868 7336
rect 17920 7284 17926 7336
rect 18984 7256 19012 7364
rect 19150 7352 19156 7404
rect 19208 7352 19214 7404
rect 19708 7396 19766 7401
rect 19794 7396 19800 7404
rect 19708 7395 19800 7396
rect 19708 7361 19720 7395
rect 19754 7368 19800 7395
rect 19754 7361 19766 7368
rect 19708 7355 19766 7361
rect 19794 7352 19800 7368
rect 19852 7352 19858 7404
rect 20714 7352 20720 7404
rect 20772 7352 20778 7404
rect 20806 7352 20812 7404
rect 20864 7392 20870 7404
rect 21177 7395 21235 7401
rect 21177 7392 21189 7395
rect 20864 7364 21189 7392
rect 20864 7352 20870 7364
rect 21177 7361 21189 7364
rect 21223 7361 21235 7395
rect 21177 7355 21235 7361
rect 21634 7352 21640 7404
rect 21692 7392 21698 7404
rect 21913 7395 21971 7401
rect 21913 7392 21925 7395
rect 21692 7364 21925 7392
rect 21692 7352 21698 7364
rect 21913 7361 21925 7364
rect 21959 7392 21971 7395
rect 22465 7395 22523 7401
rect 22465 7392 22477 7395
rect 21959 7364 22477 7392
rect 21959 7361 21971 7364
rect 21913 7355 21971 7361
rect 22465 7361 22477 7364
rect 22511 7361 22523 7395
rect 22465 7355 22523 7361
rect 23290 7352 23296 7404
rect 23348 7392 23354 7404
rect 23661 7395 23719 7401
rect 23661 7392 23673 7395
rect 23348 7364 23673 7392
rect 23348 7352 23354 7364
rect 23661 7361 23673 7364
rect 23707 7361 23719 7395
rect 23661 7355 23719 7361
rect 19058 7284 19064 7336
rect 19116 7324 19122 7336
rect 19242 7324 19248 7336
rect 19116 7296 19248 7324
rect 19116 7284 19122 7296
rect 19242 7284 19248 7296
rect 19300 7324 19306 7336
rect 19429 7327 19487 7333
rect 19429 7324 19441 7327
rect 19300 7296 19441 7324
rect 19300 7284 19306 7296
rect 19429 7293 19441 7296
rect 19475 7293 19487 7327
rect 19429 7287 19487 7293
rect 22186 7284 22192 7336
rect 22244 7284 22250 7336
rect 23566 7284 23572 7336
rect 23624 7284 23630 7336
rect 14384 7228 19012 7256
rect 20901 7259 20959 7265
rect 12345 7219 12403 7225
rect 20901 7225 20913 7259
rect 20947 7256 20959 7259
rect 20947 7228 22324 7256
rect 20947 7225 20959 7228
rect 20901 7219 20959 7225
rect 9364 7160 10640 7188
rect 9364 7148 9370 7160
rect 11422 7148 11428 7200
rect 11480 7148 11486 7200
rect 11514 7148 11520 7200
rect 11572 7148 11578 7200
rect 11606 7148 11612 7200
rect 11664 7188 11670 7200
rect 12894 7188 12900 7200
rect 11664 7160 12900 7188
rect 11664 7148 11670 7160
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 13354 7148 13360 7200
rect 13412 7188 13418 7200
rect 14550 7188 14556 7200
rect 13412 7160 14556 7188
rect 13412 7148 13418 7160
rect 14550 7148 14556 7160
rect 14608 7148 14614 7200
rect 15378 7148 15384 7200
rect 15436 7188 15442 7200
rect 16761 7191 16819 7197
rect 16761 7188 16773 7191
rect 15436 7160 16773 7188
rect 15436 7148 15442 7160
rect 16761 7157 16773 7160
rect 16807 7157 16819 7191
rect 16761 7151 16819 7157
rect 17402 7148 17408 7200
rect 17460 7188 17466 7200
rect 18230 7188 18236 7200
rect 17460 7160 18236 7188
rect 17460 7148 17466 7160
rect 18230 7148 18236 7160
rect 18288 7188 18294 7200
rect 18325 7191 18383 7197
rect 18325 7188 18337 7191
rect 18288 7160 18337 7188
rect 18288 7148 18294 7160
rect 18325 7157 18337 7160
rect 18371 7157 18383 7191
rect 18325 7151 18383 7157
rect 19337 7191 19395 7197
rect 19337 7157 19349 7191
rect 19383 7188 19395 7191
rect 22094 7188 22100 7200
rect 19383 7160 22100 7188
rect 19383 7157 19395 7160
rect 19337 7151 19395 7157
rect 22094 7148 22100 7160
rect 22152 7148 22158 7200
rect 22296 7188 22324 7228
rect 24412 7188 24440 7432
rect 25130 7352 25136 7404
rect 25188 7392 25194 7404
rect 25590 7392 25596 7404
rect 25188 7364 25596 7392
rect 25188 7352 25194 7364
rect 25590 7352 25596 7364
rect 25648 7352 25654 7404
rect 26786 7352 26792 7404
rect 26844 7392 26850 7404
rect 26973 7395 27031 7401
rect 26973 7392 26985 7395
rect 26844 7364 26985 7392
rect 26844 7352 26850 7364
rect 26973 7361 26985 7364
rect 27019 7392 27031 7395
rect 27525 7395 27583 7401
rect 27525 7392 27537 7395
rect 27019 7364 27537 7392
rect 27019 7361 27031 7364
rect 26973 7355 27031 7361
rect 27525 7361 27537 7364
rect 27571 7361 27583 7395
rect 27525 7355 27583 7361
rect 27614 7352 27620 7404
rect 27672 7392 27678 7404
rect 27672 7364 27844 7392
rect 27672 7352 27678 7364
rect 24486 7284 24492 7336
rect 24544 7324 24550 7336
rect 27249 7327 27307 7333
rect 27249 7324 27261 7327
rect 24544 7296 27261 7324
rect 24544 7284 24550 7296
rect 27249 7293 27261 7296
rect 27295 7293 27307 7327
rect 27816 7324 27844 7364
rect 28350 7352 28356 7404
rect 28408 7392 28414 7404
rect 28445 7395 28503 7401
rect 28445 7392 28457 7395
rect 28408 7364 28457 7392
rect 28408 7352 28414 7364
rect 28445 7361 28457 7364
rect 28491 7361 28503 7395
rect 28445 7355 28503 7361
rect 28994 7352 29000 7404
rect 29052 7392 29058 7404
rect 29089 7395 29147 7401
rect 29089 7392 29101 7395
rect 29052 7364 29101 7392
rect 29052 7352 29058 7364
rect 29089 7361 29101 7364
rect 29135 7361 29147 7395
rect 29089 7355 29147 7361
rect 29178 7352 29184 7404
rect 29236 7392 29242 7404
rect 29822 7392 29828 7404
rect 29236 7364 29828 7392
rect 29236 7352 29242 7364
rect 29822 7352 29828 7364
rect 29880 7352 29886 7404
rect 29932 7392 29960 7432
rect 30558 7392 30564 7404
rect 29932 7364 30564 7392
rect 30558 7352 30564 7364
rect 30616 7352 30622 7404
rect 31312 7401 31340 7432
rect 31021 7395 31079 7401
rect 31021 7361 31033 7395
rect 31067 7361 31079 7395
rect 31021 7355 31079 7361
rect 31297 7395 31355 7401
rect 31297 7361 31309 7395
rect 31343 7361 31355 7395
rect 31297 7355 31355 7361
rect 31757 7395 31815 7401
rect 31757 7361 31769 7395
rect 31803 7361 31815 7395
rect 32600 7392 32628 7432
rect 34146 7420 34152 7472
rect 34204 7460 34210 7472
rect 36630 7460 36636 7472
rect 34204 7432 36636 7460
rect 34204 7420 34210 7432
rect 36630 7420 36636 7432
rect 36688 7420 36694 7472
rect 39040 7460 39068 7491
rect 39574 7488 39580 7500
rect 39632 7488 39638 7540
rect 39482 7460 39488 7472
rect 36740 7432 38884 7460
rect 39040 7432 39488 7460
rect 32600 7364 32720 7392
rect 31757 7355 31815 7361
rect 29362 7324 29368 7336
rect 27816 7296 29368 7324
rect 27249 7287 27307 7293
rect 22296 7160 24440 7188
rect 25317 7191 25375 7197
rect 25317 7157 25329 7191
rect 25363 7188 25375 7191
rect 27154 7188 27160 7200
rect 25363 7160 27160 7188
rect 25363 7157 25375 7160
rect 25317 7151 25375 7157
rect 27154 7148 27160 7160
rect 27212 7148 27218 7200
rect 27264 7188 27292 7287
rect 28261 7259 28319 7265
rect 28261 7225 28273 7259
rect 28307 7256 28319 7259
rect 29178 7256 29184 7268
rect 28307 7228 29184 7256
rect 28307 7225 28319 7228
rect 28261 7219 28319 7225
rect 29178 7216 29184 7228
rect 29236 7216 29242 7268
rect 29288 7265 29316 7296
rect 29362 7284 29368 7296
rect 29420 7324 29426 7336
rect 29420 7296 30420 7324
rect 29420 7284 29426 7296
rect 29273 7259 29331 7265
rect 29273 7225 29285 7259
rect 29319 7225 29331 7259
rect 30098 7256 30104 7268
rect 29273 7219 29331 7225
rect 29380 7228 30104 7256
rect 29380 7200 29408 7228
rect 30098 7216 30104 7228
rect 30156 7216 30162 7268
rect 30392 7256 30420 7296
rect 30466 7284 30472 7336
rect 30524 7324 30530 7336
rect 30653 7327 30711 7333
rect 30653 7324 30665 7327
rect 30524 7296 30665 7324
rect 30524 7284 30530 7296
rect 30653 7293 30665 7296
rect 30699 7293 30711 7327
rect 30653 7287 30711 7293
rect 30742 7284 30748 7336
rect 30800 7284 30806 7336
rect 31036 7256 31064 7355
rect 31110 7284 31116 7336
rect 31168 7324 31174 7336
rect 31772 7324 31800 7355
rect 31168 7296 31800 7324
rect 31168 7284 31174 7296
rect 32490 7284 32496 7336
rect 32548 7324 32554 7336
rect 32692 7333 32720 7364
rect 34238 7352 34244 7404
rect 34296 7392 34302 7404
rect 35345 7395 35403 7401
rect 35345 7392 35357 7395
rect 34296 7364 35357 7392
rect 34296 7352 34302 7364
rect 35345 7361 35357 7364
rect 35391 7361 35403 7395
rect 35345 7355 35403 7361
rect 32585 7327 32643 7333
rect 32585 7324 32597 7327
rect 32548 7296 32597 7324
rect 32548 7284 32554 7296
rect 32585 7293 32597 7296
rect 32631 7293 32643 7327
rect 32585 7287 32643 7293
rect 32677 7327 32735 7333
rect 32677 7293 32689 7327
rect 32723 7293 32735 7327
rect 32677 7287 32735 7293
rect 34882 7284 34888 7336
rect 34940 7324 34946 7336
rect 36740 7324 36768 7432
rect 37642 7352 37648 7404
rect 37700 7352 37706 7404
rect 37737 7395 37795 7401
rect 37737 7361 37749 7395
rect 37783 7361 37795 7395
rect 37737 7355 37795 7361
rect 38105 7395 38163 7401
rect 38105 7361 38117 7395
rect 38151 7361 38163 7395
rect 38105 7355 38163 7361
rect 34940 7296 36768 7324
rect 34940 7284 34946 7296
rect 36906 7284 36912 7336
rect 36964 7324 36970 7336
rect 37752 7324 37780 7355
rect 38120 7324 38148 7355
rect 38378 7352 38384 7404
rect 38436 7392 38442 7404
rect 38856 7401 38884 7432
rect 39482 7420 39488 7432
rect 39540 7420 39546 7472
rect 38473 7395 38531 7401
rect 38473 7392 38485 7395
rect 38436 7364 38485 7392
rect 38436 7352 38442 7364
rect 38473 7361 38485 7364
rect 38519 7361 38531 7395
rect 38473 7355 38531 7361
rect 38841 7395 38899 7401
rect 38841 7361 38853 7395
rect 38887 7361 38899 7395
rect 38841 7355 38899 7361
rect 39209 7395 39267 7401
rect 39209 7361 39221 7395
rect 39255 7361 39267 7395
rect 39209 7355 39267 7361
rect 36964 7296 37780 7324
rect 37844 7296 38148 7324
rect 36964 7284 36970 7296
rect 30392 7228 31064 7256
rect 31386 7216 31392 7268
rect 31444 7256 31450 7268
rect 31573 7259 31631 7265
rect 31573 7256 31585 7259
rect 31444 7228 31585 7256
rect 31444 7216 31450 7228
rect 31573 7225 31585 7228
rect 31619 7225 31631 7259
rect 37458 7256 37464 7268
rect 31573 7219 31631 7225
rect 31726 7228 37464 7256
rect 28534 7188 28540 7200
rect 27264 7160 28540 7188
rect 28534 7148 28540 7160
rect 28592 7148 28598 7200
rect 28629 7191 28687 7197
rect 28629 7157 28641 7191
rect 28675 7188 28687 7191
rect 28902 7188 28908 7200
rect 28675 7160 28908 7188
rect 28675 7157 28687 7160
rect 28629 7151 28687 7157
rect 28902 7148 28908 7160
rect 28960 7148 28966 7200
rect 29362 7148 29368 7200
rect 29420 7148 29426 7200
rect 30006 7148 30012 7200
rect 30064 7148 30070 7200
rect 30190 7148 30196 7200
rect 30248 7148 30254 7200
rect 30282 7148 30288 7200
rect 30340 7188 30346 7200
rect 31726 7188 31754 7228
rect 37458 7216 37464 7228
rect 37516 7216 37522 7268
rect 37734 7216 37740 7268
rect 37792 7256 37798 7268
rect 37844 7256 37872 7296
rect 38194 7284 38200 7336
rect 38252 7324 38258 7336
rect 39224 7324 39252 7355
rect 38252 7296 39252 7324
rect 38252 7284 38258 7296
rect 37792 7228 37872 7256
rect 37921 7259 37979 7265
rect 37792 7216 37798 7228
rect 37921 7225 37933 7259
rect 37967 7256 37979 7259
rect 40034 7256 40040 7268
rect 37967 7228 40040 7256
rect 37967 7225 37979 7228
rect 37921 7219 37979 7225
rect 40034 7216 40040 7228
rect 40092 7216 40098 7268
rect 30340 7160 31754 7188
rect 30340 7148 30346 7160
rect 32674 7148 32680 7200
rect 32732 7188 32738 7200
rect 38838 7188 38844 7200
rect 32732 7160 38844 7188
rect 32732 7148 32738 7160
rect 38838 7148 38844 7160
rect 38896 7148 38902 7200
rect 1104 7098 39836 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 37950 7098
rect 38002 7046 38014 7098
rect 38066 7046 38078 7098
rect 38130 7046 38142 7098
rect 38194 7046 38206 7098
rect 38258 7046 39836 7098
rect 1104 7024 39836 7046
rect 2866 6944 2872 6996
rect 2924 6984 2930 6996
rect 2924 6956 4568 6984
rect 2924 6944 2930 6956
rect 4540 6916 4568 6956
rect 4890 6944 4896 6996
rect 4948 6944 4954 6996
rect 4982 6944 4988 6996
rect 5040 6984 5046 6996
rect 5040 6956 8616 6984
rect 5040 6944 5046 6956
rect 7558 6916 7564 6928
rect 4540 6888 7564 6916
rect 7558 6876 7564 6888
rect 7616 6876 7622 6928
rect 8588 6916 8616 6956
rect 8662 6944 8668 6996
rect 8720 6984 8726 6996
rect 8757 6987 8815 6993
rect 8757 6984 8769 6987
rect 8720 6956 8769 6984
rect 8720 6944 8726 6956
rect 8757 6953 8769 6956
rect 8803 6953 8815 6987
rect 9766 6984 9772 6996
rect 8757 6947 8815 6953
rect 9600 6956 9772 6984
rect 9600 6916 9628 6956
rect 9766 6944 9772 6956
rect 9824 6944 9830 6996
rect 9950 6944 9956 6996
rect 10008 6984 10014 6996
rect 10045 6987 10103 6993
rect 10045 6984 10057 6987
rect 10008 6956 10057 6984
rect 10008 6944 10014 6956
rect 10045 6953 10057 6956
rect 10091 6953 10103 6987
rect 10045 6947 10103 6953
rect 11241 6987 11299 6993
rect 11241 6953 11253 6987
rect 11287 6984 11299 6987
rect 11330 6984 11336 6996
rect 11287 6956 11336 6984
rect 11287 6953 11299 6956
rect 11241 6947 11299 6953
rect 11330 6944 11336 6956
rect 11388 6944 11394 6996
rect 12618 6944 12624 6996
rect 12676 6984 12682 6996
rect 15197 6987 15255 6993
rect 12676 6956 14412 6984
rect 12676 6944 12682 6956
rect 8588 6888 9628 6916
rect 9674 6876 9680 6928
rect 9732 6916 9738 6928
rect 13722 6916 13728 6928
rect 9732 6888 13728 6916
rect 9732 6876 9738 6888
rect 13722 6876 13728 6888
rect 13780 6876 13786 6928
rect 14384 6916 14412 6956
rect 15197 6953 15209 6987
rect 15243 6984 15255 6987
rect 15470 6984 15476 6996
rect 15243 6956 15476 6984
rect 15243 6953 15255 6956
rect 15197 6947 15255 6953
rect 15470 6944 15476 6956
rect 15528 6944 15534 6996
rect 16022 6944 16028 6996
rect 16080 6984 16086 6996
rect 16117 6987 16175 6993
rect 16117 6984 16129 6987
rect 16080 6956 16129 6984
rect 16080 6944 16086 6956
rect 16117 6953 16129 6956
rect 16163 6953 16175 6987
rect 16117 6947 16175 6953
rect 16206 6944 16212 6996
rect 16264 6984 16270 6996
rect 17402 6984 17408 6996
rect 16264 6956 17408 6984
rect 16264 6944 16270 6956
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 17862 6944 17868 6996
rect 17920 6984 17926 6996
rect 20714 6984 20720 6996
rect 17920 6956 20720 6984
rect 17920 6944 17926 6956
rect 20714 6944 20720 6956
rect 20772 6944 20778 6996
rect 27430 6984 27436 6996
rect 22066 6956 27436 6984
rect 16298 6916 16304 6928
rect 14384 6888 16304 6916
rect 16298 6876 16304 6888
rect 16356 6876 16362 6928
rect 16942 6876 16948 6928
rect 17000 6916 17006 6928
rect 20533 6919 20591 6925
rect 17000 6888 18000 6916
rect 17000 6876 17006 6888
rect 5994 6808 6000 6860
rect 6052 6848 6058 6860
rect 7006 6848 7012 6860
rect 6052 6820 7012 6848
rect 6052 6808 6058 6820
rect 7006 6808 7012 6820
rect 7064 6808 7070 6860
rect 8662 6848 8668 6860
rect 8312 6820 8668 6848
rect 198 6740 204 6792
rect 256 6780 262 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 256 6752 1409 6780
rect 256 6740 262 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6749 1731 6783
rect 1673 6743 1731 6749
rect 1688 6712 1716 6743
rect 3878 6740 3884 6792
rect 3936 6740 3942 6792
rect 4154 6740 4160 6792
rect 4212 6740 4218 6792
rect 5534 6740 5540 6792
rect 5592 6740 5598 6792
rect 6362 6740 6368 6792
rect 6420 6780 6426 6792
rect 6457 6783 6515 6789
rect 6457 6780 6469 6783
rect 6420 6752 6469 6780
rect 6420 6740 6426 6752
rect 6457 6749 6469 6752
rect 6503 6749 6515 6783
rect 6457 6743 6515 6749
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6780 7803 6783
rect 7926 6780 7932 6792
rect 7791 6752 7932 6780
rect 7791 6749 7803 6752
rect 7745 6743 7803 6749
rect 7926 6740 7932 6752
rect 7984 6740 7990 6792
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6780 8079 6783
rect 8312 6780 8340 6820
rect 8662 6808 8668 6820
rect 8720 6848 8726 6860
rect 9122 6848 9128 6860
rect 8720 6820 9128 6848
rect 8720 6808 8726 6820
rect 9122 6808 9128 6820
rect 9180 6808 9186 6860
rect 11330 6848 11336 6860
rect 9225 6820 11336 6848
rect 8067 6752 8340 6780
rect 8067 6749 8079 6752
rect 8021 6743 8079 6749
rect 8386 6740 8392 6792
rect 8444 6780 8450 6792
rect 9030 6780 9036 6792
rect 8444 6752 9036 6780
rect 8444 6740 8450 6752
rect 9030 6740 9036 6752
rect 9088 6740 9094 6792
rect 9225 6789 9253 6820
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 11974 6808 11980 6860
rect 12032 6848 12038 6860
rect 12253 6851 12311 6857
rect 12253 6848 12265 6851
rect 12032 6820 12265 6848
rect 12032 6808 12038 6820
rect 12253 6817 12265 6820
rect 12299 6817 12311 6851
rect 13262 6848 13268 6860
rect 12253 6811 12311 6817
rect 12544 6820 13268 6848
rect 9210 6783 9268 6789
rect 9210 6749 9222 6783
rect 9256 6749 9268 6783
rect 9210 6743 9268 6749
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 9401 6783 9459 6789
rect 9401 6780 9413 6783
rect 9364 6752 9413 6780
rect 9364 6740 9370 6752
rect 9401 6749 9413 6752
rect 9447 6749 9459 6783
rect 9401 6743 9459 6749
rect 9582 6740 9588 6792
rect 9640 6740 9646 6792
rect 10226 6740 10232 6792
rect 10284 6740 10290 6792
rect 10597 6783 10655 6789
rect 10597 6749 10609 6783
rect 10643 6749 10655 6783
rect 10597 6743 10655 6749
rect 5442 6712 5448 6724
rect 1688 6684 5448 6712
rect 5442 6672 5448 6684
rect 5500 6672 5506 6724
rect 9490 6712 9496 6724
rect 5552 6684 9496 6712
rect 1578 6604 1584 6656
rect 1636 6644 1642 6656
rect 5552 6644 5580 6684
rect 9490 6672 9496 6684
rect 9548 6672 9554 6724
rect 9600 6712 9628 6740
rect 10612 6712 10640 6743
rect 10686 6740 10692 6792
rect 10744 6740 10750 6792
rect 11422 6740 11428 6792
rect 11480 6740 11486 6792
rect 11514 6740 11520 6792
rect 11572 6740 11578 6792
rect 11698 6740 11704 6792
rect 11756 6780 11762 6792
rect 12544 6780 12572 6820
rect 13262 6808 13268 6820
rect 13320 6808 13326 6860
rect 14182 6808 14188 6860
rect 14240 6848 14246 6860
rect 14553 6851 14611 6857
rect 14553 6848 14565 6851
rect 14240 6820 14565 6848
rect 14240 6808 14246 6820
rect 14553 6817 14565 6820
rect 14599 6817 14611 6851
rect 14553 6811 14611 6817
rect 14734 6808 14740 6860
rect 14792 6848 14798 6860
rect 16850 6848 16856 6860
rect 14792 6820 16856 6848
rect 14792 6808 14798 6820
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 17037 6851 17095 6857
rect 17037 6817 17049 6851
rect 17083 6848 17095 6851
rect 17083 6820 17356 6848
rect 17083 6817 17095 6820
rect 17037 6811 17095 6817
rect 11756 6752 12572 6780
rect 11756 6740 11762 6752
rect 12618 6740 12624 6792
rect 12676 6780 12682 6792
rect 13173 6783 13231 6789
rect 13173 6780 13185 6783
rect 12676 6752 13185 6780
rect 12676 6740 12682 6752
rect 13173 6749 13185 6752
rect 13219 6749 13231 6783
rect 13173 6743 13231 6749
rect 13354 6740 13360 6792
rect 13412 6780 13418 6792
rect 15470 6780 15476 6792
rect 13412 6752 15476 6780
rect 13412 6740 13418 6752
rect 15470 6740 15476 6752
rect 15528 6740 15534 6792
rect 16301 6783 16359 6789
rect 16301 6749 16313 6783
rect 16347 6780 16359 6783
rect 16761 6783 16819 6789
rect 16347 6752 16436 6780
rect 16347 6749 16359 6752
rect 16301 6743 16359 6749
rect 11054 6712 11060 6724
rect 9600 6684 10456 6712
rect 10612 6684 11060 6712
rect 1636 6616 5580 6644
rect 5721 6647 5779 6653
rect 1636 6604 1642 6616
rect 5721 6613 5733 6647
rect 5767 6644 5779 6647
rect 5902 6644 5908 6656
rect 5767 6616 5908 6644
rect 5767 6613 5779 6616
rect 5721 6607 5779 6613
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 6270 6604 6276 6656
rect 6328 6644 6334 6656
rect 6641 6647 6699 6653
rect 6641 6644 6653 6647
rect 6328 6616 6653 6644
rect 6328 6604 6334 6616
rect 6641 6613 6653 6616
rect 6687 6644 6699 6647
rect 7190 6644 7196 6656
rect 6687 6616 7196 6644
rect 6687 6613 6699 6616
rect 6641 6607 6699 6613
rect 7190 6604 7196 6616
rect 7248 6644 7254 6656
rect 7558 6644 7564 6656
rect 7248 6616 7564 6644
rect 7248 6604 7254 6616
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 8754 6604 8760 6656
rect 8812 6644 8818 6656
rect 9033 6647 9091 6653
rect 9033 6644 9045 6647
rect 8812 6616 9045 6644
rect 8812 6604 8818 6616
rect 9033 6613 9045 6616
rect 9079 6613 9091 6647
rect 9033 6607 9091 6613
rect 9398 6604 9404 6656
rect 9456 6644 9462 6656
rect 10428 6653 10456 6684
rect 11054 6672 11060 6684
rect 11112 6672 11118 6724
rect 12250 6672 12256 6724
rect 12308 6712 12314 6724
rect 13262 6712 13268 6724
rect 12308 6684 13268 6712
rect 12308 6672 12314 6684
rect 13262 6672 13268 6684
rect 13320 6672 13326 6724
rect 13814 6672 13820 6724
rect 13872 6712 13878 6724
rect 14826 6712 14832 6724
rect 13872 6684 14832 6712
rect 13872 6672 13878 6684
rect 14826 6672 14832 6684
rect 14884 6672 14890 6724
rect 9585 6647 9643 6653
rect 9585 6644 9597 6647
rect 9456 6616 9597 6644
rect 9456 6604 9462 6616
rect 9585 6613 9597 6616
rect 9631 6613 9643 6647
rect 9585 6607 9643 6613
rect 10413 6647 10471 6653
rect 10413 6613 10425 6647
rect 10459 6613 10471 6647
rect 10413 6607 10471 6613
rect 10778 6604 10784 6656
rect 10836 6644 10842 6656
rect 10873 6647 10931 6653
rect 10873 6644 10885 6647
rect 10836 6616 10885 6644
rect 10836 6604 10842 6616
rect 10873 6613 10885 6616
rect 10919 6613 10931 6647
rect 10873 6607 10931 6613
rect 11701 6647 11759 6653
rect 11701 6613 11713 6647
rect 11747 6644 11759 6647
rect 11790 6644 11796 6656
rect 11747 6616 11796 6644
rect 11747 6613 11759 6616
rect 11701 6607 11759 6613
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 12434 6604 12440 6656
rect 12492 6604 12498 6656
rect 12526 6604 12532 6656
rect 12584 6604 12590 6656
rect 12618 6604 12624 6656
rect 12676 6644 12682 6656
rect 12897 6647 12955 6653
rect 12897 6644 12909 6647
rect 12676 6616 12909 6644
rect 12676 6604 12682 6616
rect 12897 6613 12909 6616
rect 12943 6613 12955 6647
rect 12897 6607 12955 6613
rect 12989 6647 13047 6653
rect 12989 6613 13001 6647
rect 13035 6644 13047 6647
rect 13078 6644 13084 6656
rect 13035 6616 13084 6644
rect 13035 6613 13047 6616
rect 12989 6607 13047 6613
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 13170 6604 13176 6656
rect 13228 6644 13234 6656
rect 15654 6644 15660 6656
rect 13228 6616 15660 6644
rect 13228 6604 13234 6616
rect 15654 6604 15660 6616
rect 15712 6604 15718 6656
rect 16408 6653 16436 6752
rect 16761 6749 16773 6783
rect 16807 6780 16819 6783
rect 16942 6780 16948 6792
rect 16807 6752 16948 6780
rect 16807 6749 16819 6752
rect 16761 6743 16819 6749
rect 16942 6740 16948 6752
rect 17000 6740 17006 6792
rect 17218 6740 17224 6792
rect 17276 6740 17282 6792
rect 16393 6647 16451 6653
rect 16393 6613 16405 6647
rect 16439 6613 16451 6647
rect 17328 6644 17356 6820
rect 17402 6808 17408 6860
rect 17460 6808 17466 6860
rect 17862 6808 17868 6860
rect 17920 6808 17926 6860
rect 17972 6848 18000 6888
rect 20533 6885 20545 6919
rect 20579 6885 20591 6919
rect 20533 6879 20591 6885
rect 18258 6851 18316 6857
rect 18258 6848 18270 6851
rect 17972 6820 18270 6848
rect 18258 6817 18270 6820
rect 18304 6817 18316 6851
rect 20548 6848 20576 6879
rect 20622 6876 20628 6928
rect 20680 6916 20686 6928
rect 22066 6916 22094 6956
rect 27430 6944 27436 6956
rect 27488 6944 27494 6996
rect 29822 6984 29828 6996
rect 28644 6956 29828 6984
rect 20680 6888 22094 6916
rect 22281 6919 22339 6925
rect 20680 6876 20686 6888
rect 22281 6885 22293 6919
rect 22327 6885 22339 6919
rect 22281 6879 22339 6885
rect 25133 6919 25191 6925
rect 25133 6885 25145 6919
rect 25179 6885 25191 6919
rect 25133 6879 25191 6885
rect 21177 6851 21235 6857
rect 21177 6848 21189 6851
rect 20548 6820 21189 6848
rect 18258 6811 18316 6817
rect 21177 6817 21189 6820
rect 21223 6817 21235 6851
rect 22296 6848 22324 6879
rect 21177 6811 21235 6817
rect 21284 6820 22324 6848
rect 18138 6740 18144 6792
rect 18196 6740 18202 6792
rect 18414 6740 18420 6792
rect 18472 6740 18478 6792
rect 19518 6740 19524 6792
rect 19576 6740 19582 6792
rect 19794 6740 19800 6792
rect 19852 6740 19858 6792
rect 20162 6740 20168 6792
rect 20220 6780 20226 6792
rect 21085 6783 21143 6789
rect 21085 6780 21097 6783
rect 20220 6752 21097 6780
rect 20220 6740 20226 6752
rect 21085 6749 21097 6752
rect 21131 6749 21143 6783
rect 21085 6743 21143 6749
rect 21284 6712 21312 6820
rect 25148 6792 25176 6879
rect 25406 6876 25412 6928
rect 25464 6916 25470 6928
rect 28644 6916 28672 6956
rect 29822 6944 29828 6956
rect 29880 6944 29886 6996
rect 30006 6944 30012 6996
rect 30064 6984 30070 6996
rect 30064 6956 33272 6984
rect 30064 6944 30070 6956
rect 25464 6888 28672 6916
rect 25464 6876 25470 6888
rect 28718 6876 28724 6928
rect 28776 6916 28782 6928
rect 30282 6916 30288 6928
rect 28776 6888 30288 6916
rect 28776 6876 28782 6888
rect 30282 6876 30288 6888
rect 30340 6876 30346 6928
rect 30558 6876 30564 6928
rect 30616 6916 30622 6928
rect 30616 6888 31708 6916
rect 30616 6876 30622 6888
rect 27154 6808 27160 6860
rect 27212 6848 27218 6860
rect 27212 6820 30052 6848
rect 27212 6808 27218 6820
rect 21634 6740 21640 6792
rect 21692 6780 21698 6792
rect 23017 6783 23075 6789
rect 23017 6780 23029 6783
rect 21692 6752 23029 6780
rect 21692 6740 21698 6752
rect 23017 6749 23029 6752
rect 23063 6749 23075 6783
rect 23017 6743 23075 6749
rect 23293 6783 23351 6789
rect 23293 6749 23305 6783
rect 23339 6780 23351 6783
rect 23750 6780 23756 6792
rect 23339 6752 23756 6780
rect 23339 6749 23351 6752
rect 23293 6743 23351 6749
rect 23750 6740 23756 6752
rect 23808 6740 23814 6792
rect 25130 6740 25136 6792
rect 25188 6740 25194 6792
rect 25317 6783 25375 6789
rect 25317 6749 25329 6783
rect 25363 6780 25375 6783
rect 25406 6780 25412 6792
rect 25363 6752 25412 6780
rect 25363 6749 25375 6752
rect 25317 6743 25375 6749
rect 25406 6740 25412 6752
rect 25464 6740 25470 6792
rect 28813 6783 28871 6789
rect 28813 6749 28825 6783
rect 28859 6780 28871 6783
rect 28859 6752 29592 6780
rect 28859 6749 28871 6752
rect 28813 6743 28871 6749
rect 18892 6684 21312 6712
rect 18892 6644 18920 6684
rect 21818 6672 21824 6724
rect 21876 6712 21882 6724
rect 28718 6712 28724 6724
rect 21876 6684 28724 6712
rect 21876 6672 21882 6684
rect 28718 6672 28724 6684
rect 28776 6672 28782 6724
rect 17328 6616 18920 6644
rect 16393 6607 16451 6613
rect 18966 6604 18972 6656
rect 19024 6644 19030 6656
rect 19061 6647 19119 6653
rect 19061 6644 19073 6647
rect 19024 6616 19073 6644
rect 19024 6604 19030 6616
rect 19061 6613 19073 6616
rect 19107 6613 19119 6647
rect 19061 6607 19119 6613
rect 19242 6604 19248 6656
rect 19300 6644 19306 6656
rect 20438 6644 20444 6656
rect 19300 6616 20444 6644
rect 19300 6604 19306 6616
rect 20438 6604 20444 6616
rect 20496 6604 20502 6656
rect 20625 6647 20683 6653
rect 20625 6613 20637 6647
rect 20671 6644 20683 6647
rect 20898 6644 20904 6656
rect 20671 6616 20904 6644
rect 20671 6613 20683 6616
rect 20625 6607 20683 6613
rect 20898 6604 20904 6616
rect 20956 6604 20962 6656
rect 20990 6604 20996 6656
rect 21048 6604 21054 6656
rect 21450 6604 21456 6656
rect 21508 6644 21514 6656
rect 25222 6644 25228 6656
rect 21508 6616 25228 6644
rect 21508 6604 21514 6616
rect 25222 6604 25228 6616
rect 25280 6604 25286 6656
rect 27522 6604 27528 6656
rect 27580 6644 27586 6656
rect 29564 6653 29592 6752
rect 29914 6740 29920 6792
rect 29972 6740 29978 6792
rect 30024 6712 30052 6820
rect 30098 6808 30104 6860
rect 30156 6808 30162 6860
rect 30374 6808 30380 6860
rect 30432 6848 30438 6860
rect 31680 6857 31708 6888
rect 31754 6876 31760 6928
rect 31812 6916 31818 6928
rect 32214 6916 32220 6928
rect 31812 6888 32220 6916
rect 31812 6876 31818 6888
rect 32214 6876 32220 6888
rect 32272 6876 32278 6928
rect 31665 6851 31723 6857
rect 30432 6820 31524 6848
rect 30432 6808 30438 6820
rect 30190 6740 30196 6792
rect 30248 6780 30254 6792
rect 30561 6783 30619 6789
rect 30561 6780 30573 6783
rect 30248 6752 30573 6780
rect 30248 6740 30254 6752
rect 30561 6749 30573 6752
rect 30607 6749 30619 6783
rect 30561 6743 30619 6749
rect 31110 6740 31116 6792
rect 31168 6780 31174 6792
rect 31389 6783 31447 6789
rect 31389 6780 31401 6783
rect 31168 6752 31401 6780
rect 31168 6740 31174 6752
rect 31389 6749 31401 6752
rect 31435 6749 31447 6783
rect 31496 6780 31524 6820
rect 31665 6817 31677 6851
rect 31711 6817 31723 6851
rect 32309 6851 32367 6857
rect 32309 6848 32321 6851
rect 31665 6811 31723 6817
rect 31772 6820 32321 6848
rect 31772 6780 31800 6820
rect 32309 6817 32321 6820
rect 32355 6817 32367 6851
rect 32309 6811 32367 6817
rect 32582 6808 32588 6860
rect 32640 6808 32646 6860
rect 33244 6848 33272 6956
rect 37826 6944 37832 6996
rect 37884 6944 37890 6996
rect 38930 6848 38936 6860
rect 33244 6820 38936 6848
rect 38930 6808 38936 6820
rect 38988 6808 38994 6860
rect 31496 6752 31800 6780
rect 31849 6783 31907 6789
rect 31389 6743 31447 6749
rect 31849 6749 31861 6783
rect 31895 6780 31907 6783
rect 32030 6780 32036 6792
rect 31895 6752 32036 6780
rect 31895 6749 31907 6752
rect 31849 6743 31907 6749
rect 32030 6740 32036 6752
rect 32088 6740 32094 6792
rect 32766 6789 32772 6792
rect 32723 6783 32772 6789
rect 32723 6749 32735 6783
rect 32769 6749 32772 6783
rect 32723 6743 32772 6749
rect 32766 6740 32772 6743
rect 32824 6740 32830 6792
rect 32858 6740 32864 6792
rect 32916 6740 32922 6792
rect 37645 6783 37703 6789
rect 37645 6749 37657 6783
rect 37691 6780 37703 6783
rect 38010 6780 38016 6792
rect 37691 6752 38016 6780
rect 37691 6749 37703 6752
rect 37645 6743 37703 6749
rect 38010 6740 38016 6752
rect 38068 6740 38074 6792
rect 38105 6783 38163 6789
rect 38105 6749 38117 6783
rect 38151 6780 38163 6783
rect 38381 6783 38439 6789
rect 38381 6780 38393 6783
rect 38151 6752 38393 6780
rect 38151 6749 38163 6752
rect 38105 6743 38163 6749
rect 38381 6749 38393 6752
rect 38427 6749 38439 6783
rect 38381 6743 38439 6749
rect 38473 6783 38531 6789
rect 38473 6749 38485 6783
rect 38519 6749 38531 6783
rect 38841 6783 38899 6789
rect 38841 6780 38853 6783
rect 38473 6743 38531 6749
rect 38580 6752 38853 6780
rect 35526 6712 35532 6724
rect 30024 6684 31754 6712
rect 28629 6647 28687 6653
rect 28629 6644 28641 6647
rect 27580 6616 28641 6644
rect 27580 6604 27586 6616
rect 28629 6613 28641 6616
rect 28675 6613 28687 6647
rect 28629 6607 28687 6613
rect 29549 6647 29607 6653
rect 29549 6613 29561 6647
rect 29595 6613 29607 6647
rect 29549 6607 29607 6613
rect 30009 6647 30067 6653
rect 30009 6613 30021 6647
rect 30055 6644 30067 6647
rect 30282 6644 30288 6656
rect 30055 6616 30288 6644
rect 30055 6613 30067 6616
rect 30009 6607 30067 6613
rect 30282 6604 30288 6616
rect 30340 6604 30346 6656
rect 30374 6604 30380 6656
rect 30432 6604 30438 6656
rect 30650 6604 30656 6656
rect 30708 6644 30714 6656
rect 31205 6647 31263 6653
rect 31205 6644 31217 6647
rect 30708 6616 31217 6644
rect 30708 6604 30714 6616
rect 31205 6613 31217 6616
rect 31251 6613 31263 6647
rect 31726 6644 31754 6684
rect 33428 6684 35532 6712
rect 33428 6644 33456 6684
rect 35526 6672 35532 6684
rect 35584 6672 35590 6724
rect 36998 6672 37004 6724
rect 37056 6712 37062 6724
rect 37056 6684 38240 6712
rect 37056 6672 37062 6684
rect 31726 6616 33456 6644
rect 31205 6607 31263 6613
rect 33502 6604 33508 6656
rect 33560 6604 33566 6656
rect 37826 6604 37832 6656
rect 37884 6644 37890 6656
rect 38212 6653 38240 6684
rect 38286 6672 38292 6724
rect 38344 6712 38350 6724
rect 38488 6712 38516 6743
rect 38344 6684 38516 6712
rect 38344 6672 38350 6684
rect 38013 6647 38071 6653
rect 38013 6644 38025 6647
rect 37884 6616 38025 6644
rect 37884 6604 37890 6616
rect 38013 6613 38025 6616
rect 38059 6613 38071 6647
rect 38013 6607 38071 6613
rect 38197 6647 38255 6653
rect 38197 6613 38209 6647
rect 38243 6613 38255 6647
rect 38197 6607 38255 6613
rect 38470 6604 38476 6656
rect 38528 6644 38534 6656
rect 38580 6644 38608 6752
rect 38841 6749 38853 6752
rect 38887 6749 38899 6783
rect 39209 6783 39267 6789
rect 39209 6780 39221 6783
rect 38841 6743 38899 6749
rect 38948 6752 39221 6780
rect 38746 6672 38752 6724
rect 38804 6712 38810 6724
rect 38948 6712 38976 6752
rect 39209 6749 39221 6752
rect 39255 6749 39267 6783
rect 39209 6743 39267 6749
rect 39666 6712 39672 6724
rect 38804 6684 38976 6712
rect 39040 6684 39672 6712
rect 38804 6672 38810 6684
rect 38528 6616 38608 6644
rect 38528 6604 38534 6616
rect 38654 6604 38660 6656
rect 38712 6604 38718 6656
rect 39040 6653 39068 6684
rect 39666 6672 39672 6684
rect 39724 6672 39730 6724
rect 39025 6647 39083 6653
rect 39025 6613 39037 6647
rect 39071 6613 39083 6647
rect 39025 6607 39083 6613
rect 39390 6604 39396 6656
rect 39448 6604 39454 6656
rect 1104 6554 39836 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 39010 6554
rect 39062 6502 39074 6554
rect 39126 6502 39138 6554
rect 39190 6502 39202 6554
rect 39254 6502 39266 6554
rect 39318 6502 39836 6554
rect 1104 6480 39836 6502
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 3878 6440 3884 6452
rect 2556 6412 3884 6440
rect 2556 6400 2562 6412
rect 3878 6400 3884 6412
rect 3936 6440 3942 6452
rect 5721 6443 5779 6449
rect 3936 6412 5120 6440
rect 3936 6400 3942 6412
rect 5092 6384 5120 6412
rect 5721 6409 5733 6443
rect 5767 6440 5779 6443
rect 6454 6440 6460 6452
rect 5767 6412 6460 6440
rect 5767 6409 5779 6412
rect 5721 6403 5779 6409
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 7745 6443 7803 6449
rect 7745 6409 7757 6443
rect 7791 6440 7803 6443
rect 7926 6440 7932 6452
rect 7791 6412 7932 6440
rect 7791 6409 7803 6412
rect 7745 6403 7803 6409
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 11698 6440 11704 6452
rect 8312 6412 11704 6440
rect 934 6332 940 6384
rect 992 6372 998 6384
rect 3697 6375 3755 6381
rect 992 6344 1808 6372
rect 992 6332 998 6344
rect 750 6264 756 6316
rect 808 6304 814 6316
rect 1780 6313 1808 6344
rect 3697 6341 3709 6375
rect 3743 6372 3755 6375
rect 4154 6372 4160 6384
rect 3743 6344 4160 6372
rect 3743 6341 3755 6344
rect 3697 6335 3755 6341
rect 1489 6307 1547 6313
rect 1489 6304 1501 6307
rect 808 6276 1501 6304
rect 808 6264 814 6276
rect 1489 6273 1501 6276
rect 1535 6273 1547 6307
rect 1489 6267 1547 6273
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6273 1823 6307
rect 1765 6267 1823 6273
rect 1854 6264 1860 6316
rect 1912 6304 1918 6316
rect 3712 6304 3740 6335
rect 4154 6332 4160 6344
rect 4212 6332 4218 6384
rect 4430 6332 4436 6384
rect 4488 6372 4494 6384
rect 4488 6344 5028 6372
rect 4488 6332 4494 6344
rect 1912 6276 3740 6304
rect 1912 6264 1918 6276
rect 4522 6264 4528 6316
rect 4580 6304 4586 6316
rect 4617 6307 4675 6313
rect 4617 6304 4629 6307
rect 4580 6276 4629 6304
rect 4580 6264 4586 6276
rect 4617 6273 4629 6276
rect 4663 6273 4675 6307
rect 4617 6267 4675 6273
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6304 4767 6307
rect 4890 6304 4896 6316
rect 4755 6276 4896 6304
rect 4755 6273 4767 6276
rect 4709 6267 4767 6273
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 5000 6313 5028 6344
rect 5074 6332 5080 6384
rect 5132 6372 5138 6384
rect 5132 6344 8064 6372
rect 5132 6332 5138 6344
rect 7852 6313 7880 6344
rect 8036 6334 8064 6344
rect 8312 6334 8340 6412
rect 11698 6400 11704 6412
rect 11756 6400 11762 6452
rect 11974 6400 11980 6452
rect 12032 6400 12038 6452
rect 17681 6443 17739 6449
rect 12820 6412 16988 6440
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6304 5043 6307
rect 7009 6307 7067 6313
rect 7009 6304 7021 6307
rect 5031 6276 6500 6304
rect 5031 6273 5043 6276
rect 4985 6267 5043 6273
rect 1670 6196 1676 6248
rect 1728 6196 1734 6248
rect 6472 6236 6500 6276
rect 6656 6276 7021 6304
rect 6546 6236 6552 6248
rect 6472 6208 6552 6236
rect 6546 6196 6552 6208
rect 6604 6236 6610 6248
rect 6656 6236 6684 6276
rect 7009 6273 7021 6276
rect 7055 6273 7067 6307
rect 7009 6267 7067 6273
rect 7837 6307 7895 6313
rect 7837 6273 7849 6307
rect 7883 6273 7895 6307
rect 8036 6306 8340 6334
rect 8754 6332 8760 6384
rect 8812 6372 8818 6384
rect 12342 6372 12348 6384
rect 8812 6344 12348 6372
rect 8812 6332 8818 6344
rect 12342 6332 12348 6344
rect 12400 6332 12406 6384
rect 8389 6307 8447 6313
rect 7837 6267 7895 6273
rect 8389 6273 8401 6307
rect 8435 6304 8447 6307
rect 8662 6304 8668 6316
rect 8435 6276 8668 6304
rect 8435 6273 8447 6276
rect 8389 6267 8447 6273
rect 8662 6264 8668 6276
rect 8720 6304 8726 6316
rect 9401 6307 9459 6313
rect 9401 6304 9413 6307
rect 8720 6276 9413 6304
rect 8720 6264 8726 6276
rect 9401 6273 9413 6276
rect 9447 6273 9459 6307
rect 9401 6267 9459 6273
rect 9490 6264 9496 6316
rect 9548 6304 9554 6316
rect 10502 6304 10508 6316
rect 9548 6276 10508 6304
rect 9548 6264 9554 6276
rect 10502 6264 10508 6276
rect 10560 6304 10566 6316
rect 12713 6307 12771 6313
rect 12713 6304 12725 6307
rect 10560 6276 12725 6304
rect 10560 6264 10566 6276
rect 12713 6273 12725 6276
rect 12759 6304 12771 6307
rect 12820 6304 12848 6412
rect 13262 6332 13268 6384
rect 13320 6372 13326 6384
rect 14366 6372 14372 6384
rect 13320 6344 14372 6372
rect 13320 6332 13326 6344
rect 14366 6332 14372 6344
rect 14424 6332 14430 6384
rect 12759 6276 12848 6304
rect 12989 6307 13047 6313
rect 12759 6273 12771 6276
rect 12713 6267 12771 6273
rect 12989 6273 13001 6307
rect 13035 6304 13047 6307
rect 13173 6307 13231 6313
rect 13173 6304 13185 6307
rect 13035 6276 13185 6304
rect 13035 6273 13047 6276
rect 12989 6267 13047 6273
rect 13173 6273 13185 6276
rect 13219 6304 13231 6307
rect 13354 6304 13360 6316
rect 13219 6276 13360 6304
rect 13219 6273 13231 6276
rect 13173 6267 13231 6273
rect 13354 6264 13360 6276
rect 13412 6264 13418 6316
rect 13446 6264 13452 6316
rect 13504 6264 13510 6316
rect 13538 6264 13544 6316
rect 13596 6304 13602 6316
rect 13596 6276 14596 6304
rect 13596 6264 13602 6276
rect 6604 6208 6684 6236
rect 6733 6239 6791 6245
rect 6604 6196 6610 6208
rect 6733 6205 6745 6239
rect 6779 6205 6791 6239
rect 6733 6199 6791 6205
rect 3878 6128 3884 6180
rect 3936 6128 3942 6180
rect 5442 6128 5448 6180
rect 5500 6168 5506 6180
rect 5500 6140 6408 6168
rect 5500 6128 5506 6140
rect 1949 6103 2007 6109
rect 1949 6069 1961 6103
rect 1995 6100 2007 6103
rect 6178 6100 6184 6112
rect 1995 6072 6184 6100
rect 1995 6069 2007 6072
rect 1949 6063 2007 6069
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 6380 6100 6408 6140
rect 6454 6128 6460 6180
rect 6512 6168 6518 6180
rect 6748 6168 6776 6199
rect 7650 6196 7656 6248
rect 7708 6236 7714 6248
rect 7708 6208 7972 6236
rect 7708 6196 7714 6208
rect 6512 6140 6776 6168
rect 6512 6128 6518 6140
rect 7558 6128 7564 6180
rect 7616 6168 7622 6180
rect 7834 6168 7840 6180
rect 7616 6140 7840 6168
rect 7616 6128 7622 6140
rect 7834 6128 7840 6140
rect 7892 6128 7898 6180
rect 7944 6168 7972 6208
rect 9122 6196 9128 6248
rect 9180 6196 9186 6248
rect 9766 6196 9772 6248
rect 9824 6236 9830 6248
rect 10134 6236 10140 6248
rect 9824 6208 10140 6236
rect 9824 6196 9830 6208
rect 10134 6196 10140 6208
rect 10192 6236 10198 6248
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 10192 6208 10241 6236
rect 10192 6196 10198 6208
rect 10229 6205 10241 6208
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 11606 6196 11612 6248
rect 11664 6236 11670 6248
rect 12066 6236 12072 6248
rect 11664 6208 12072 6236
rect 11664 6196 11670 6208
rect 12066 6196 12072 6208
rect 12124 6196 12130 6248
rect 12342 6196 12348 6248
rect 12400 6196 12406 6248
rect 14277 6239 14335 6245
rect 14277 6205 14289 6239
rect 14323 6205 14335 6239
rect 14277 6199 14335 6205
rect 9140 6168 9168 6196
rect 12250 6168 12256 6180
rect 7944 6140 9168 6168
rect 10060 6140 10364 6168
rect 7190 6100 7196 6112
rect 6380 6072 7196 6100
rect 7190 6060 7196 6072
rect 7248 6060 7254 6112
rect 8036 6109 8064 6140
rect 8021 6103 8079 6109
rect 8021 6069 8033 6103
rect 8067 6069 8079 6103
rect 8021 6063 8079 6069
rect 8481 6103 8539 6109
rect 8481 6069 8493 6103
rect 8527 6100 8539 6103
rect 8570 6100 8576 6112
rect 8527 6072 8576 6100
rect 8527 6069 8539 6072
rect 8481 6063 8539 6069
rect 8570 6060 8576 6072
rect 8628 6060 8634 6112
rect 9122 6060 9128 6112
rect 9180 6100 9186 6112
rect 10060 6100 10088 6140
rect 9180 6072 10088 6100
rect 9180 6060 9186 6072
rect 10134 6060 10140 6112
rect 10192 6060 10198 6112
rect 10336 6100 10364 6140
rect 11072 6140 12256 6168
rect 11072 6100 11100 6140
rect 12250 6128 12256 6140
rect 12308 6128 12314 6180
rect 10336 6072 11100 6100
rect 11241 6103 11299 6109
rect 11241 6069 11253 6103
rect 11287 6100 11299 6103
rect 11974 6100 11980 6112
rect 11287 6072 11980 6100
rect 11287 6069 11299 6072
rect 11241 6063 11299 6069
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 12360 6100 12388 6196
rect 14182 6128 14188 6180
rect 14240 6128 14246 6180
rect 14292 6168 14320 6199
rect 14366 6196 14372 6248
rect 14424 6236 14430 6248
rect 14461 6239 14519 6245
rect 14461 6236 14473 6239
rect 14424 6208 14473 6236
rect 14424 6196 14430 6208
rect 14461 6205 14473 6208
rect 14507 6205 14519 6239
rect 14568 6236 14596 6276
rect 15470 6264 15476 6316
rect 15528 6264 15534 6316
rect 16117 6307 16175 6313
rect 16117 6273 16129 6307
rect 16163 6304 16175 6307
rect 16850 6304 16856 6316
rect 16163 6276 16856 6304
rect 16163 6273 16175 6276
rect 16117 6267 16175 6273
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 16960 6313 16988 6412
rect 17681 6409 17693 6443
rect 17727 6440 17739 6443
rect 17862 6440 17868 6452
rect 17727 6412 17868 6440
rect 17727 6409 17739 6412
rect 17681 6403 17739 6409
rect 17862 6400 17868 6412
rect 17920 6400 17926 6452
rect 18141 6443 18199 6449
rect 18141 6409 18153 6443
rect 18187 6409 18199 6443
rect 18141 6403 18199 6409
rect 20257 6443 20315 6449
rect 20257 6409 20269 6443
rect 20303 6440 20315 6443
rect 20346 6440 20352 6452
rect 20303 6412 20352 6440
rect 20303 6409 20315 6412
rect 20257 6403 20315 6409
rect 16945 6307 17003 6313
rect 16945 6273 16957 6307
rect 16991 6273 17003 6307
rect 16945 6267 17003 6273
rect 17218 6264 17224 6316
rect 17276 6264 17282 6316
rect 18049 6307 18107 6313
rect 18049 6273 18061 6307
rect 18095 6304 18107 6307
rect 18156 6304 18184 6403
rect 20346 6400 20352 6412
rect 20404 6400 20410 6452
rect 20714 6400 20720 6452
rect 20772 6440 20778 6452
rect 22373 6443 22431 6449
rect 22373 6440 22385 6443
rect 20772 6412 22385 6440
rect 20772 6400 20778 6412
rect 22373 6409 22385 6412
rect 22419 6409 22431 6443
rect 22373 6403 22431 6409
rect 23474 6400 23480 6452
rect 23532 6400 23538 6452
rect 23934 6400 23940 6452
rect 23992 6440 23998 6452
rect 26418 6440 26424 6452
rect 23992 6412 26424 6440
rect 23992 6400 23998 6412
rect 26418 6400 26424 6412
rect 26476 6400 26482 6452
rect 26510 6400 26516 6452
rect 26568 6440 26574 6452
rect 27522 6440 27528 6452
rect 26568 6412 27528 6440
rect 26568 6400 26574 6412
rect 27522 6400 27528 6412
rect 27580 6400 27586 6452
rect 28442 6400 28448 6452
rect 28500 6440 28506 6452
rect 28721 6443 28779 6449
rect 28721 6440 28733 6443
rect 28500 6412 28733 6440
rect 28500 6400 28506 6412
rect 28721 6409 28733 6412
rect 28767 6409 28779 6443
rect 28721 6403 28779 6409
rect 31110 6400 31116 6452
rect 31168 6400 31174 6452
rect 31754 6400 31760 6452
rect 31812 6440 31818 6452
rect 32030 6440 32036 6452
rect 31812 6412 32036 6440
rect 31812 6400 31818 6412
rect 32030 6400 32036 6412
rect 32088 6400 32094 6452
rect 32125 6443 32183 6449
rect 32125 6409 32137 6443
rect 32171 6440 32183 6443
rect 32398 6440 32404 6452
rect 32171 6412 32404 6440
rect 32171 6409 32183 6412
rect 32125 6403 32183 6409
rect 32398 6400 32404 6412
rect 32456 6400 32462 6452
rect 32858 6400 32864 6452
rect 32916 6440 32922 6452
rect 33229 6443 33287 6449
rect 33229 6440 33241 6443
rect 32916 6412 33241 6440
rect 32916 6400 32922 6412
rect 33229 6409 33241 6412
rect 33275 6409 33287 6443
rect 33229 6403 33287 6409
rect 35434 6400 35440 6452
rect 35492 6440 35498 6452
rect 35713 6443 35771 6449
rect 35713 6440 35725 6443
rect 35492 6412 35725 6440
rect 35492 6400 35498 6412
rect 35713 6409 35725 6412
rect 35759 6409 35771 6443
rect 35713 6403 35771 6409
rect 36078 6400 36084 6452
rect 36136 6440 36142 6452
rect 38565 6443 38623 6449
rect 38565 6440 38577 6443
rect 36136 6412 38577 6440
rect 36136 6400 36142 6412
rect 38565 6409 38577 6412
rect 38611 6409 38623 6443
rect 38565 6403 38623 6409
rect 39393 6443 39451 6449
rect 39393 6409 39405 6443
rect 39439 6440 39451 6443
rect 39850 6440 39856 6452
rect 39439 6412 39856 6440
rect 39439 6409 39451 6412
rect 39393 6403 39451 6409
rect 39850 6400 39856 6412
rect 39908 6400 39914 6452
rect 18509 6375 18567 6381
rect 18509 6341 18521 6375
rect 18555 6372 18567 6375
rect 23842 6372 23848 6384
rect 18555 6344 23848 6372
rect 18555 6341 18567 6344
rect 18509 6335 18567 6341
rect 18095 6276 18184 6304
rect 18095 6273 18107 6276
rect 18049 6267 18107 6273
rect 15194 6236 15200 6248
rect 14568 6208 15200 6236
rect 14461 6199 14519 6205
rect 15194 6196 15200 6208
rect 15252 6196 15258 6248
rect 15335 6239 15393 6245
rect 15335 6205 15347 6239
rect 15381 6236 15393 6239
rect 16298 6236 16304 6248
rect 15381 6208 16304 6236
rect 15381 6205 15393 6208
rect 15335 6199 15393 6205
rect 16298 6196 16304 6208
rect 16356 6196 16362 6248
rect 16666 6196 16672 6248
rect 16724 6196 16730 6248
rect 17236 6236 17264 6264
rect 18524 6236 18552 6335
rect 23842 6332 23848 6344
rect 23900 6332 23906 6384
rect 24026 6332 24032 6384
rect 24084 6372 24090 6384
rect 29086 6372 29092 6384
rect 24084 6344 29092 6372
rect 24084 6332 24090 6344
rect 29086 6332 29092 6344
rect 29144 6332 29150 6384
rect 32766 6372 32772 6384
rect 32232 6344 32772 6372
rect 18601 6307 18659 6313
rect 18601 6273 18613 6307
rect 18647 6304 18659 6307
rect 18966 6304 18972 6316
rect 18647 6276 18972 6304
rect 18647 6273 18659 6276
rect 18601 6267 18659 6273
rect 18966 6264 18972 6276
rect 19024 6304 19030 6316
rect 20162 6304 20168 6316
rect 19024 6276 20168 6304
rect 19024 6264 19030 6276
rect 20162 6264 20168 6276
rect 20220 6264 20226 6316
rect 20898 6264 20904 6316
rect 20956 6264 20962 6316
rect 21177 6307 21235 6313
rect 21177 6273 21189 6307
rect 21223 6273 21235 6307
rect 21177 6267 21235 6273
rect 17236 6208 18552 6236
rect 18693 6239 18751 6245
rect 18693 6205 18705 6239
rect 18739 6205 18751 6239
rect 18693 6199 18751 6205
rect 20073 6239 20131 6245
rect 20073 6205 20085 6239
rect 20119 6205 20131 6239
rect 21192 6236 21220 6267
rect 22554 6264 22560 6316
rect 22612 6304 22618 6316
rect 23109 6307 23167 6313
rect 23109 6304 23121 6307
rect 22612 6276 23121 6304
rect 22612 6264 22618 6276
rect 23109 6273 23121 6276
rect 23155 6273 23167 6307
rect 24213 6307 24271 6313
rect 24213 6304 24225 6307
rect 23109 6267 23167 6273
rect 23952 6276 24225 6304
rect 20073 6199 20131 6205
rect 20640 6208 21220 6236
rect 14826 6168 14832 6180
rect 14292 6140 14832 6168
rect 14826 6128 14832 6140
rect 14884 6128 14890 6180
rect 14918 6128 14924 6180
rect 14976 6128 14982 6180
rect 18708 6168 18736 6199
rect 17328 6140 18736 6168
rect 20088 6168 20116 6199
rect 20346 6168 20352 6180
rect 20088 6140 20352 6168
rect 17328 6100 17356 6140
rect 20346 6128 20352 6140
rect 20404 6128 20410 6180
rect 20640 6177 20668 6208
rect 23382 6196 23388 6248
rect 23440 6196 23446 6248
rect 23658 6196 23664 6248
rect 23716 6236 23722 6248
rect 23952 6236 23980 6276
rect 24213 6273 24225 6276
rect 24259 6273 24271 6307
rect 24213 6267 24271 6273
rect 24486 6264 24492 6316
rect 24544 6264 24550 6316
rect 25038 6264 25044 6316
rect 25096 6264 25102 6316
rect 26237 6307 26295 6313
rect 26237 6304 26249 6307
rect 25424 6276 26249 6304
rect 23716 6208 23980 6236
rect 23716 6196 23722 6208
rect 24578 6196 24584 6248
rect 24636 6236 24642 6248
rect 24765 6239 24823 6245
rect 24765 6236 24777 6239
rect 24636 6208 24777 6236
rect 24636 6196 24642 6208
rect 24765 6205 24777 6208
rect 24811 6205 24823 6239
rect 24765 6199 24823 6205
rect 20625 6171 20683 6177
rect 20625 6137 20637 6171
rect 20671 6137 20683 6171
rect 20625 6131 20683 6137
rect 20806 6128 20812 6180
rect 20864 6168 20870 6180
rect 20993 6171 21051 6177
rect 20993 6168 21005 6171
rect 20864 6140 21005 6168
rect 20864 6128 20870 6140
rect 20993 6137 21005 6140
rect 21039 6137 21051 6171
rect 20993 6131 21051 6137
rect 23400 6140 23612 6168
rect 12360 6072 17356 6100
rect 17862 6060 17868 6112
rect 17920 6060 17926 6112
rect 19702 6060 19708 6112
rect 19760 6100 19766 6112
rect 20717 6103 20775 6109
rect 20717 6100 20729 6103
rect 19760 6072 20729 6100
rect 19760 6060 19766 6072
rect 20717 6069 20729 6072
rect 20763 6069 20775 6103
rect 20717 6063 20775 6069
rect 21082 6060 21088 6112
rect 21140 6100 21146 6112
rect 22278 6100 22284 6112
rect 21140 6072 22284 6100
rect 21140 6060 21146 6072
rect 22278 6060 22284 6072
rect 22336 6100 22342 6112
rect 23400 6100 23428 6140
rect 22336 6072 23428 6100
rect 23584 6100 23612 6140
rect 25424 6100 25452 6276
rect 26237 6273 26249 6276
rect 26283 6273 26295 6307
rect 26237 6267 26295 6273
rect 26786 6264 26792 6316
rect 26844 6304 26850 6316
rect 27249 6307 27307 6313
rect 27249 6304 27261 6307
rect 26844 6276 27261 6304
rect 26844 6264 26850 6276
rect 27249 6273 27261 6276
rect 27295 6273 27307 6307
rect 27249 6267 27307 6273
rect 27522 6264 27528 6316
rect 27580 6264 27586 6316
rect 28626 6264 28632 6316
rect 28684 6304 28690 6316
rect 28905 6307 28963 6313
rect 28905 6304 28917 6307
rect 28684 6276 28917 6304
rect 28684 6264 28690 6276
rect 28905 6273 28917 6276
rect 28951 6273 28963 6307
rect 28905 6267 28963 6273
rect 29638 6264 29644 6316
rect 29696 6264 29702 6316
rect 29914 6264 29920 6316
rect 29972 6264 29978 6316
rect 31294 6264 31300 6316
rect 31352 6304 31358 6316
rect 31481 6307 31539 6313
rect 31481 6304 31493 6307
rect 31352 6276 31493 6304
rect 31352 6264 31358 6276
rect 31481 6273 31493 6276
rect 31527 6304 31539 6307
rect 32232 6304 32260 6344
rect 32766 6332 32772 6344
rect 32824 6332 32830 6384
rect 33980 6344 34836 6372
rect 33980 6316 34008 6344
rect 31527 6276 32260 6304
rect 32309 6307 32367 6313
rect 31527 6273 31539 6276
rect 31481 6267 31539 6273
rect 32309 6273 32321 6307
rect 32355 6273 32367 6307
rect 32309 6267 32367 6273
rect 25866 6196 25872 6248
rect 25924 6236 25930 6248
rect 26329 6239 26387 6245
rect 26329 6236 26341 6239
rect 25924 6208 26341 6236
rect 25924 6196 25930 6208
rect 26329 6205 26341 6208
rect 26375 6205 26387 6239
rect 26329 6199 26387 6205
rect 26421 6239 26479 6245
rect 26421 6205 26433 6239
rect 26467 6205 26479 6239
rect 26973 6239 27031 6245
rect 26973 6236 26985 6239
rect 26421 6199 26479 6205
rect 26528 6208 26985 6236
rect 25777 6171 25835 6177
rect 25777 6137 25789 6171
rect 25823 6168 25835 6171
rect 26436 6168 26464 6199
rect 25823 6140 26464 6168
rect 25823 6137 25835 6140
rect 25777 6131 25835 6137
rect 23584 6072 25452 6100
rect 25869 6103 25927 6109
rect 22336 6060 22342 6072
rect 25869 6069 25881 6103
rect 25915 6100 25927 6103
rect 25958 6100 25964 6112
rect 25915 6072 25964 6100
rect 25915 6069 25927 6072
rect 25869 6063 25927 6069
rect 25958 6060 25964 6072
rect 26016 6060 26022 6112
rect 26326 6060 26332 6112
rect 26384 6100 26390 6112
rect 26528 6100 26556 6208
rect 26973 6205 26985 6208
rect 27019 6205 27031 6239
rect 27540 6236 27568 6264
rect 29779 6239 29837 6245
rect 29779 6236 29791 6239
rect 27540 6208 29791 6236
rect 26973 6199 27031 6205
rect 29779 6205 29791 6208
rect 29825 6205 29837 6239
rect 29779 6199 29837 6205
rect 30650 6196 30656 6248
rect 30708 6196 30714 6248
rect 30837 6239 30895 6245
rect 30837 6205 30849 6239
rect 30883 6236 30895 6239
rect 30926 6236 30932 6248
rect 30883 6208 30932 6236
rect 30883 6205 30895 6208
rect 30837 6199 30895 6205
rect 30926 6196 30932 6208
rect 30984 6236 30990 6248
rect 31110 6236 31116 6248
rect 30984 6208 31116 6236
rect 30984 6196 30990 6208
rect 31110 6196 31116 6208
rect 31168 6196 31174 6248
rect 31573 6239 31631 6245
rect 31573 6205 31585 6239
rect 31619 6205 31631 6239
rect 31573 6199 31631 6205
rect 31757 6239 31815 6245
rect 31757 6205 31769 6239
rect 31803 6236 31815 6239
rect 31846 6236 31852 6248
rect 31803 6208 31852 6236
rect 31803 6205 31815 6208
rect 31757 6199 31815 6205
rect 27985 6171 28043 6177
rect 27985 6137 27997 6171
rect 28031 6168 28043 6171
rect 28031 6140 29316 6168
rect 28031 6137 28043 6140
rect 27985 6131 28043 6137
rect 26384 6072 26556 6100
rect 26384 6060 26390 6072
rect 26602 6060 26608 6112
rect 26660 6100 26666 6112
rect 28718 6100 28724 6112
rect 26660 6072 28724 6100
rect 26660 6060 26666 6072
rect 28718 6060 28724 6072
rect 28776 6060 28782 6112
rect 28997 6103 29055 6109
rect 28997 6069 29009 6103
rect 29043 6100 29055 6103
rect 29086 6100 29092 6112
rect 29043 6072 29092 6100
rect 29043 6069 29055 6072
rect 28997 6063 29055 6069
rect 29086 6060 29092 6072
rect 29144 6060 29150 6112
rect 29288 6100 29316 6140
rect 30190 6128 30196 6180
rect 30248 6128 30254 6180
rect 31202 6128 31208 6180
rect 31260 6168 31266 6180
rect 31588 6168 31616 6199
rect 31846 6196 31852 6208
rect 31904 6196 31910 6248
rect 32324 6236 32352 6267
rect 32582 6264 32588 6316
rect 32640 6304 32646 6316
rect 33502 6304 33508 6316
rect 32640 6276 33508 6304
rect 32640 6264 32646 6276
rect 33502 6264 33508 6276
rect 33560 6264 33566 6316
rect 33962 6264 33968 6316
rect 34020 6264 34026 6316
rect 34517 6307 34575 6313
rect 34517 6273 34529 6307
rect 34563 6304 34575 6307
rect 34698 6304 34704 6316
rect 34563 6276 34704 6304
rect 34563 6273 34575 6276
rect 34517 6267 34575 6273
rect 34698 6264 34704 6276
rect 34756 6264 34762 6316
rect 34808 6313 34836 6344
rect 35526 6332 35532 6384
rect 35584 6372 35590 6384
rect 35584 6344 39252 6372
rect 35584 6332 35590 6344
rect 34793 6307 34851 6313
rect 34793 6273 34805 6307
rect 34839 6273 34851 6307
rect 34793 6267 34851 6273
rect 35805 6307 35863 6313
rect 35805 6273 35817 6307
rect 35851 6304 35863 6307
rect 35986 6304 35992 6316
rect 35851 6276 35992 6304
rect 35851 6273 35863 6276
rect 35805 6267 35863 6273
rect 35986 6264 35992 6276
rect 36044 6264 36050 6316
rect 38749 6307 38807 6313
rect 38749 6273 38761 6307
rect 38795 6273 38807 6307
rect 38749 6267 38807 6273
rect 38841 6307 38899 6313
rect 38841 6273 38853 6307
rect 38887 6304 38899 6307
rect 38930 6304 38936 6316
rect 38887 6276 38936 6304
rect 38887 6273 38899 6276
rect 38841 6267 38899 6273
rect 32766 6236 32772 6248
rect 32324 6208 32772 6236
rect 32766 6196 32772 6208
rect 32824 6196 32830 6248
rect 34241 6239 34299 6245
rect 34241 6205 34253 6239
rect 34287 6205 34299 6239
rect 38764 6236 38792 6267
rect 38930 6264 38936 6276
rect 38988 6264 38994 6316
rect 39224 6313 39252 6344
rect 39209 6307 39267 6313
rect 39209 6273 39221 6307
rect 39255 6273 39267 6307
rect 39209 6267 39267 6273
rect 39850 6236 39856 6248
rect 38764 6208 39856 6236
rect 34241 6199 34299 6205
rect 32490 6168 32496 6180
rect 31260 6140 32496 6168
rect 31260 6128 31266 6140
rect 32490 6128 32496 6140
rect 32548 6128 32554 6180
rect 31846 6100 31852 6112
rect 29288 6072 31852 6100
rect 31846 6060 31852 6072
rect 31904 6060 31910 6112
rect 32214 6060 32220 6112
rect 32272 6100 32278 6112
rect 34256 6100 34284 6199
rect 39850 6196 39856 6208
rect 39908 6196 39914 6248
rect 38010 6128 38016 6180
rect 38068 6168 38074 6180
rect 39574 6168 39580 6180
rect 38068 6140 39580 6168
rect 38068 6128 38074 6140
rect 39574 6128 39580 6140
rect 39632 6128 39638 6180
rect 32272 6072 34284 6100
rect 32272 6060 32278 6072
rect 35434 6060 35440 6112
rect 35492 6100 35498 6112
rect 35529 6103 35587 6109
rect 35529 6100 35541 6103
rect 35492 6072 35541 6100
rect 35492 6060 35498 6072
rect 35529 6069 35541 6072
rect 35575 6069 35587 6103
rect 35529 6063 35587 6069
rect 39022 6060 39028 6112
rect 39080 6060 39086 6112
rect 1104 6010 39836 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 37950 6010
rect 38002 5958 38014 6010
rect 38066 5958 38078 6010
rect 38130 5958 38142 6010
rect 38194 5958 38206 6010
rect 38258 5958 39836 6010
rect 1104 5936 39836 5958
rect 1578 5856 1584 5908
rect 1636 5856 1642 5908
rect 2133 5899 2191 5905
rect 2133 5865 2145 5899
rect 2179 5896 2191 5899
rect 6086 5896 6092 5908
rect 2179 5868 6092 5896
rect 2179 5865 2191 5868
rect 2133 5859 2191 5865
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 6196 5868 6960 5896
rect 5074 5788 5080 5840
rect 5132 5788 5138 5840
rect 1026 5720 1032 5772
rect 1084 5760 1090 5772
rect 1084 5732 1992 5760
rect 1084 5720 1090 5732
rect 750 5652 756 5704
rect 808 5692 814 5704
rect 1964 5701 1992 5732
rect 1397 5695 1455 5701
rect 1397 5692 1409 5695
rect 808 5664 1409 5692
rect 808 5652 814 5664
rect 1397 5661 1409 5664
rect 1443 5661 1455 5695
rect 1397 5655 1455 5661
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5661 1731 5695
rect 1673 5655 1731 5661
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5661 2007 5695
rect 1949 5655 2007 5661
rect 566 5584 572 5636
rect 624 5624 630 5636
rect 1688 5624 1716 5655
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 4525 5695 4583 5701
rect 4525 5692 4537 5695
rect 4212 5664 4537 5692
rect 4212 5652 4218 5664
rect 4525 5661 4537 5664
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 4798 5652 4804 5704
rect 4856 5652 4862 5704
rect 4890 5652 4896 5704
rect 4948 5692 4954 5704
rect 6196 5692 6224 5868
rect 6270 5720 6276 5772
rect 6328 5720 6334 5772
rect 6932 5760 6960 5868
rect 7006 5856 7012 5908
rect 7064 5896 7070 5908
rect 12250 5896 12256 5908
rect 7064 5868 12256 5896
rect 7064 5856 7070 5868
rect 12250 5856 12256 5868
rect 12308 5856 12314 5908
rect 12342 5856 12348 5908
rect 12400 5896 12406 5908
rect 12400 5868 14780 5896
rect 12400 5856 12406 5868
rect 8478 5788 8484 5840
rect 8536 5828 8542 5840
rect 9309 5831 9367 5837
rect 9309 5828 9321 5831
rect 8536 5800 9321 5828
rect 8536 5788 8542 5800
rect 9309 5797 9321 5800
rect 9355 5797 9367 5831
rect 9309 5791 9367 5797
rect 10134 5788 10140 5840
rect 10192 5828 10198 5840
rect 10192 5800 14044 5828
rect 10192 5788 10198 5800
rect 11790 5760 11796 5772
rect 6932 5732 11796 5760
rect 11790 5720 11796 5732
rect 11848 5720 11854 5772
rect 11974 5720 11980 5772
rect 12032 5720 12038 5772
rect 12710 5760 12716 5772
rect 12176 5732 12716 5760
rect 4948 5664 6224 5692
rect 4948 5652 4954 5664
rect 6546 5652 6552 5704
rect 6604 5652 6610 5704
rect 7190 5652 7196 5704
rect 7248 5692 7254 5704
rect 8478 5692 8484 5704
rect 7248 5664 8484 5692
rect 7248 5652 7254 5664
rect 8478 5652 8484 5664
rect 8536 5692 8542 5704
rect 9122 5692 9128 5704
rect 8536 5664 9128 5692
rect 8536 5652 8542 5664
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 10502 5652 10508 5704
rect 10560 5652 10566 5704
rect 11149 5695 11207 5701
rect 11149 5661 11161 5695
rect 11195 5692 11207 5695
rect 11885 5695 11943 5701
rect 11195 5664 11468 5692
rect 11195 5661 11207 5664
rect 11149 5655 11207 5661
rect 7006 5624 7012 5636
rect 624 5596 1716 5624
rect 1872 5596 7012 5624
rect 624 5584 630 5596
rect 1872 5565 1900 5596
rect 7006 5584 7012 5596
rect 7064 5584 7070 5636
rect 7116 5596 11192 5624
rect 1857 5559 1915 5565
rect 1857 5525 1869 5559
rect 1903 5525 1915 5559
rect 1857 5519 1915 5525
rect 3789 5559 3847 5565
rect 3789 5525 3801 5559
rect 3835 5556 3847 5559
rect 4154 5556 4160 5568
rect 3835 5528 4160 5556
rect 3835 5525 3847 5528
rect 3789 5519 3847 5525
rect 4154 5516 4160 5528
rect 4212 5516 4218 5568
rect 6086 5516 6092 5568
rect 6144 5556 6150 5568
rect 7116 5556 7144 5596
rect 11164 5568 11192 5596
rect 6144 5528 7144 5556
rect 7285 5559 7343 5565
rect 6144 5516 6150 5528
rect 7285 5525 7297 5559
rect 7331 5556 7343 5559
rect 7558 5556 7564 5568
rect 7331 5528 7564 5556
rect 7331 5525 7343 5528
rect 7285 5519 7343 5525
rect 7558 5516 7564 5528
rect 7616 5516 7622 5568
rect 7926 5516 7932 5568
rect 7984 5556 7990 5568
rect 8754 5556 8760 5568
rect 7984 5528 8760 5556
rect 7984 5516 7990 5528
rect 8754 5516 8760 5528
rect 8812 5516 8818 5568
rect 8846 5516 8852 5568
rect 8904 5556 8910 5568
rect 9398 5556 9404 5568
rect 8904 5528 9404 5556
rect 8904 5516 8910 5528
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 9950 5516 9956 5568
rect 10008 5556 10014 5568
rect 10597 5559 10655 5565
rect 10597 5556 10609 5559
rect 10008 5528 10609 5556
rect 10008 5516 10014 5528
rect 10597 5525 10609 5528
rect 10643 5525 10655 5559
rect 10597 5519 10655 5525
rect 11146 5516 11152 5568
rect 11204 5516 11210 5568
rect 11238 5516 11244 5568
rect 11296 5556 11302 5568
rect 11440 5565 11468 5664
rect 11885 5661 11897 5695
rect 11931 5692 11943 5695
rect 12176 5692 12204 5732
rect 12710 5720 12716 5732
rect 12768 5720 12774 5772
rect 12897 5763 12955 5769
rect 12897 5729 12909 5763
rect 12943 5760 12955 5763
rect 13814 5760 13820 5772
rect 12943 5732 13820 5760
rect 12943 5729 12955 5732
rect 12897 5723 12955 5729
rect 13814 5720 13820 5732
rect 13872 5720 13878 5772
rect 11931 5664 12204 5692
rect 11931 5661 11943 5664
rect 11885 5655 11943 5661
rect 12250 5652 12256 5704
rect 12308 5692 12314 5704
rect 13906 5692 13912 5704
rect 12308 5664 13912 5692
rect 12308 5652 12314 5664
rect 13906 5652 13912 5664
rect 13964 5652 13970 5704
rect 11793 5627 11851 5633
rect 11793 5593 11805 5627
rect 11839 5624 11851 5627
rect 12342 5624 12348 5636
rect 11839 5596 12348 5624
rect 11839 5593 11851 5596
rect 11793 5587 11851 5593
rect 12342 5584 12348 5596
rect 12400 5624 12406 5636
rect 13630 5624 13636 5636
rect 12400 5596 13636 5624
rect 12400 5584 12406 5596
rect 13630 5584 13636 5596
rect 13688 5584 13694 5636
rect 14016 5624 14044 5800
rect 14752 5760 14780 5868
rect 14918 5856 14924 5908
rect 14976 5896 14982 5908
rect 15105 5899 15163 5905
rect 15105 5896 15117 5899
rect 14976 5868 15117 5896
rect 14976 5856 14982 5868
rect 15105 5865 15117 5868
rect 15151 5865 15163 5899
rect 15105 5859 15163 5865
rect 16666 5856 16672 5908
rect 16724 5896 16730 5908
rect 18782 5896 18788 5908
rect 16724 5868 18788 5896
rect 16724 5856 16730 5868
rect 18782 5856 18788 5868
rect 18840 5856 18846 5908
rect 21821 5899 21879 5905
rect 20732 5868 21496 5896
rect 14826 5788 14832 5840
rect 14884 5828 14890 5840
rect 20622 5828 20628 5840
rect 14884 5800 20628 5828
rect 14884 5788 14890 5800
rect 20622 5788 20628 5800
rect 20680 5788 20686 5840
rect 19794 5760 19800 5772
rect 14752 5732 19800 5760
rect 19794 5720 19800 5732
rect 19852 5720 19858 5772
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5692 14151 5695
rect 14274 5692 14280 5704
rect 14139 5664 14280 5692
rect 14139 5661 14151 5664
rect 14093 5655 14151 5661
rect 14274 5652 14280 5664
rect 14332 5652 14338 5704
rect 14369 5695 14427 5701
rect 14369 5661 14381 5695
rect 14415 5692 14427 5695
rect 14734 5692 14740 5704
rect 14415 5664 14740 5692
rect 14415 5661 14427 5664
rect 14369 5655 14427 5661
rect 14734 5652 14740 5664
rect 14792 5652 14798 5704
rect 15194 5652 15200 5704
rect 15252 5692 15258 5704
rect 17034 5692 17040 5704
rect 15252 5664 17040 5692
rect 15252 5652 15258 5664
rect 17034 5652 17040 5664
rect 17092 5652 17098 5704
rect 20732 5692 20760 5868
rect 21468 5828 21496 5868
rect 21821 5865 21833 5899
rect 21867 5896 21879 5899
rect 21867 5868 23428 5896
rect 21867 5865 21879 5868
rect 21821 5859 21879 5865
rect 22646 5828 22652 5840
rect 21468 5800 22652 5828
rect 22646 5788 22652 5800
rect 22704 5788 22710 5840
rect 17328 5664 20760 5692
rect 17218 5624 17224 5636
rect 14016 5596 17224 5624
rect 17218 5584 17224 5596
rect 17276 5584 17282 5636
rect 11333 5559 11391 5565
rect 11333 5556 11345 5559
rect 11296 5528 11345 5556
rect 11296 5516 11302 5528
rect 11333 5525 11345 5528
rect 11379 5525 11391 5559
rect 11333 5519 11391 5525
rect 11425 5559 11483 5565
rect 11425 5525 11437 5559
rect 11471 5525 11483 5559
rect 11425 5519 11483 5525
rect 11974 5516 11980 5568
rect 12032 5556 12038 5568
rect 12253 5559 12311 5565
rect 12253 5556 12265 5559
rect 12032 5528 12265 5556
rect 12032 5516 12038 5528
rect 12253 5525 12265 5528
rect 12299 5525 12311 5559
rect 12253 5519 12311 5525
rect 12621 5559 12679 5565
rect 12621 5525 12633 5559
rect 12667 5556 12679 5559
rect 13170 5556 13176 5568
rect 12667 5528 13176 5556
rect 12667 5525 12679 5528
rect 12621 5519 12679 5525
rect 13170 5516 13176 5528
rect 13228 5516 13234 5568
rect 13722 5516 13728 5568
rect 13780 5556 13786 5568
rect 17328 5556 17356 5664
rect 20806 5652 20812 5704
rect 20864 5652 20870 5704
rect 21085 5695 21143 5701
rect 21085 5661 21097 5695
rect 21131 5692 21143 5695
rect 21542 5692 21548 5704
rect 21131 5664 21548 5692
rect 21131 5661 21143 5664
rect 21085 5655 21143 5661
rect 21542 5652 21548 5664
rect 21600 5652 21606 5704
rect 23400 5692 23428 5868
rect 23566 5856 23572 5908
rect 23624 5896 23630 5908
rect 24397 5899 24455 5905
rect 24397 5896 24409 5899
rect 23624 5868 24409 5896
rect 23624 5856 23630 5868
rect 24397 5865 24409 5868
rect 24443 5865 24455 5899
rect 26786 5896 26792 5908
rect 24397 5859 24455 5865
rect 24780 5868 26792 5896
rect 23658 5788 23664 5840
rect 23716 5828 23722 5840
rect 24780 5828 24808 5868
rect 26786 5856 26792 5868
rect 26844 5856 26850 5908
rect 27356 5868 28488 5896
rect 23716 5800 24808 5828
rect 23716 5788 23722 5800
rect 23474 5720 23480 5772
rect 23532 5760 23538 5772
rect 23750 5760 23756 5772
rect 23532 5732 23756 5760
rect 23532 5720 23538 5732
rect 23750 5720 23756 5732
rect 23808 5760 23814 5772
rect 24486 5760 24492 5772
rect 23808 5732 24492 5760
rect 23808 5720 23814 5732
rect 24486 5720 24492 5732
rect 24544 5720 24550 5772
rect 24026 5692 24032 5704
rect 23400 5664 24032 5692
rect 24026 5652 24032 5664
rect 24084 5652 24090 5704
rect 25133 5695 25191 5701
rect 25133 5661 25145 5695
rect 25179 5692 25191 5695
rect 25222 5692 25228 5704
rect 25179 5664 25228 5692
rect 25179 5661 25191 5664
rect 25133 5655 25191 5661
rect 25222 5652 25228 5664
rect 25280 5652 25286 5704
rect 25409 5695 25467 5701
rect 25409 5661 25421 5695
rect 25455 5692 25467 5695
rect 26326 5692 26332 5704
rect 25455 5664 26332 5692
rect 25455 5661 25467 5664
rect 25409 5655 25467 5661
rect 26326 5652 26332 5664
rect 26384 5692 26390 5704
rect 26421 5695 26479 5701
rect 26421 5692 26433 5695
rect 26384 5664 26433 5692
rect 26384 5652 26390 5664
rect 26421 5661 26433 5664
rect 26467 5661 26479 5695
rect 26421 5655 26479 5661
rect 26694 5652 26700 5704
rect 26752 5652 26758 5704
rect 18414 5584 18420 5636
rect 18472 5624 18478 5636
rect 21726 5624 21732 5636
rect 18472 5596 21732 5624
rect 18472 5584 18478 5596
rect 21726 5584 21732 5596
rect 21784 5584 21790 5636
rect 23106 5584 23112 5636
rect 23164 5624 23170 5636
rect 23934 5624 23940 5636
rect 23164 5596 23940 5624
rect 23164 5584 23170 5596
rect 23934 5584 23940 5596
rect 23992 5584 23998 5636
rect 13780 5528 17356 5556
rect 13780 5516 13786 5528
rect 18506 5516 18512 5568
rect 18564 5556 18570 5568
rect 27356 5556 27384 5868
rect 27430 5720 27436 5772
rect 27488 5760 27494 5772
rect 27525 5763 27583 5769
rect 27525 5760 27537 5763
rect 27488 5732 27537 5760
rect 27488 5720 27494 5732
rect 27525 5729 27537 5732
rect 27571 5729 27583 5763
rect 27525 5723 27583 5729
rect 27706 5652 27712 5704
rect 27764 5692 27770 5704
rect 27801 5695 27859 5701
rect 27801 5692 27813 5695
rect 27764 5664 27813 5692
rect 27764 5652 27770 5664
rect 27801 5661 27813 5664
rect 27847 5661 27859 5695
rect 28460 5692 28488 5868
rect 28626 5856 28632 5908
rect 28684 5856 28690 5908
rect 28718 5856 28724 5908
rect 28776 5896 28782 5908
rect 30834 5896 30840 5908
rect 28776 5868 30840 5896
rect 28776 5856 28782 5868
rect 30834 5856 30840 5868
rect 30892 5856 30898 5908
rect 31570 5856 31576 5908
rect 31628 5896 31634 5908
rect 32217 5899 32275 5905
rect 31628 5868 32168 5896
rect 31628 5856 31634 5868
rect 28537 5831 28595 5837
rect 28537 5797 28549 5831
rect 28583 5828 28595 5831
rect 30190 5828 30196 5840
rect 28583 5800 30196 5828
rect 28583 5797 28595 5800
rect 28537 5791 28595 5797
rect 30190 5788 30196 5800
rect 30248 5788 30254 5840
rect 32140 5828 32168 5868
rect 32217 5865 32229 5899
rect 32263 5896 32275 5899
rect 32766 5896 32772 5908
rect 32263 5868 32772 5896
rect 32263 5865 32275 5868
rect 32217 5859 32275 5865
rect 32766 5856 32772 5868
rect 32824 5856 32830 5908
rect 35986 5856 35992 5908
rect 36044 5856 36050 5908
rect 36446 5856 36452 5908
rect 36504 5896 36510 5908
rect 39393 5899 39451 5905
rect 36504 5868 38332 5896
rect 36504 5856 36510 5868
rect 30300 5800 31064 5828
rect 32140 5800 38240 5828
rect 28994 5720 29000 5772
rect 29052 5760 29058 5772
rect 29181 5763 29239 5769
rect 29181 5760 29193 5763
rect 29052 5732 29193 5760
rect 29052 5720 29058 5732
rect 29181 5729 29193 5732
rect 29227 5729 29239 5763
rect 29181 5723 29239 5729
rect 29362 5720 29368 5772
rect 29420 5760 29426 5772
rect 30300 5760 30328 5800
rect 29420 5732 30328 5760
rect 30469 5763 30527 5769
rect 29420 5720 29426 5732
rect 30469 5729 30481 5763
rect 30515 5760 30527 5763
rect 30650 5760 30656 5772
rect 30515 5732 30656 5760
rect 30515 5729 30527 5732
rect 30469 5723 30527 5729
rect 28460 5664 30236 5692
rect 27801 5655 27859 5661
rect 29362 5624 29368 5636
rect 27448 5596 29368 5624
rect 27448 5565 27476 5596
rect 29362 5584 29368 5596
rect 29420 5584 29426 5636
rect 30208 5624 30236 5664
rect 30282 5652 30288 5704
rect 30340 5652 30346 5704
rect 30484 5624 30512 5723
rect 30650 5720 30656 5732
rect 30708 5720 30714 5772
rect 30926 5720 30932 5772
rect 30984 5720 30990 5772
rect 31036 5760 31064 5800
rect 31481 5763 31539 5769
rect 31481 5760 31493 5763
rect 31036 5732 31493 5760
rect 31481 5729 31493 5732
rect 31527 5729 31539 5763
rect 31481 5723 31539 5729
rect 31846 5720 31852 5772
rect 31904 5760 31910 5772
rect 32769 5763 32827 5769
rect 32769 5760 32781 5763
rect 31904 5732 32781 5760
rect 31904 5720 31910 5732
rect 32769 5729 32781 5732
rect 32815 5729 32827 5763
rect 32769 5723 32827 5729
rect 35434 5720 35440 5772
rect 35492 5720 35498 5772
rect 31202 5652 31208 5704
rect 31260 5652 31266 5704
rect 31294 5652 31300 5704
rect 31352 5701 31358 5704
rect 31352 5695 31380 5701
rect 31368 5661 31380 5695
rect 31352 5655 31380 5661
rect 32125 5695 32183 5701
rect 32125 5661 32137 5695
rect 32171 5692 32183 5695
rect 32306 5692 32312 5704
rect 32171 5664 32312 5692
rect 32171 5661 32183 5664
rect 32125 5655 32183 5661
rect 31352 5652 31358 5655
rect 32306 5652 32312 5664
rect 32364 5652 32370 5704
rect 32490 5652 32496 5704
rect 32548 5692 32554 5704
rect 32677 5695 32735 5701
rect 32677 5692 32689 5695
rect 32548 5664 32689 5692
rect 32548 5652 32554 5664
rect 32677 5661 32689 5664
rect 32723 5661 32735 5695
rect 32677 5655 32735 5661
rect 33410 5652 33416 5704
rect 33468 5692 33474 5704
rect 38212 5701 38240 5800
rect 38304 5760 38332 5868
rect 39393 5865 39405 5899
rect 39439 5896 39451 5899
rect 39666 5896 39672 5908
rect 39439 5868 39672 5896
rect 39439 5865 39451 5868
rect 39393 5859 39451 5865
rect 39666 5856 39672 5868
rect 39724 5856 39730 5908
rect 39025 5831 39083 5837
rect 39025 5797 39037 5831
rect 39071 5828 39083 5831
rect 39942 5828 39948 5840
rect 39071 5800 39948 5828
rect 39071 5797 39083 5800
rect 39025 5791 39083 5797
rect 39942 5788 39948 5800
rect 40000 5788 40006 5840
rect 38304 5732 39252 5760
rect 38197 5695 38255 5701
rect 33468 5664 35756 5692
rect 33468 5652 33474 5664
rect 35621 5627 35679 5633
rect 35621 5624 35633 5627
rect 30208 5596 30512 5624
rect 32048 5596 35633 5624
rect 18564 5528 27384 5556
rect 27433 5559 27491 5565
rect 18564 5516 18570 5528
rect 27433 5525 27445 5559
rect 27479 5525 27491 5559
rect 27433 5519 27491 5525
rect 27522 5516 27528 5568
rect 27580 5556 27586 5568
rect 28997 5559 29055 5565
rect 28997 5556 29009 5559
rect 27580 5528 29009 5556
rect 27580 5516 27586 5528
rect 28997 5525 29009 5528
rect 29043 5525 29055 5559
rect 28997 5519 29055 5525
rect 29089 5559 29147 5565
rect 29089 5525 29101 5559
rect 29135 5556 29147 5559
rect 30466 5556 30472 5568
rect 29135 5528 30472 5556
rect 29135 5525 29147 5528
rect 29089 5519 29147 5525
rect 30466 5516 30472 5528
rect 30524 5516 30530 5568
rect 31110 5516 31116 5568
rect 31168 5556 31174 5568
rect 32048 5556 32076 5596
rect 35621 5593 35633 5596
rect 35667 5593 35679 5627
rect 35728 5624 35756 5664
rect 38197 5661 38209 5695
rect 38243 5661 38255 5695
rect 38197 5655 38255 5661
rect 38838 5652 38844 5704
rect 38896 5652 38902 5704
rect 39224 5701 39252 5732
rect 39209 5695 39267 5701
rect 39209 5661 39221 5695
rect 39255 5661 39267 5695
rect 39209 5655 39267 5661
rect 38470 5624 38476 5636
rect 35728 5596 38476 5624
rect 35621 5587 35679 5593
rect 38470 5584 38476 5596
rect 38528 5584 38534 5636
rect 31168 5528 32076 5556
rect 32585 5559 32643 5565
rect 31168 5516 31174 5528
rect 32585 5525 32597 5559
rect 32631 5556 32643 5559
rect 32674 5556 32680 5568
rect 32631 5528 32680 5556
rect 32631 5525 32643 5528
rect 32585 5519 32643 5525
rect 32674 5516 32680 5528
rect 32732 5516 32738 5568
rect 35526 5516 35532 5568
rect 35584 5516 35590 5568
rect 35710 5516 35716 5568
rect 35768 5556 35774 5568
rect 38013 5559 38071 5565
rect 38013 5556 38025 5559
rect 35768 5528 38025 5556
rect 35768 5516 35774 5528
rect 38013 5525 38025 5528
rect 38059 5525 38071 5559
rect 38013 5519 38071 5525
rect 1104 5466 39836 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 39010 5466
rect 39062 5414 39074 5466
rect 39126 5414 39138 5466
rect 39190 5414 39202 5466
rect 39254 5414 39266 5466
rect 39318 5414 39836 5466
rect 1104 5392 39836 5414
rect 2314 5312 2320 5364
rect 2372 5312 2378 5364
rect 4706 5312 4712 5364
rect 4764 5352 4770 5364
rect 6457 5355 6515 5361
rect 6457 5352 6469 5355
rect 4764 5324 6469 5352
rect 4764 5312 4770 5324
rect 6457 5321 6469 5324
rect 6503 5321 6515 5355
rect 6457 5315 6515 5321
rect 8404 5324 8708 5352
rect 934 5244 940 5296
rect 992 5284 998 5296
rect 1857 5287 1915 5293
rect 1857 5284 1869 5287
rect 992 5256 1869 5284
rect 992 5244 998 5256
rect 1857 5253 1869 5256
rect 1903 5253 1915 5287
rect 1857 5247 1915 5253
rect 2041 5287 2099 5293
rect 2041 5253 2053 5287
rect 2087 5284 2099 5287
rect 7926 5284 7932 5296
rect 2087 5256 7932 5284
rect 2087 5253 2099 5256
rect 2041 5247 2099 5253
rect 7926 5244 7932 5256
rect 7984 5244 7990 5296
rect 382 5176 388 5228
rect 440 5216 446 5228
rect 1489 5219 1547 5225
rect 1489 5216 1501 5219
rect 440 5188 1501 5216
rect 440 5176 446 5188
rect 1489 5185 1501 5188
rect 1535 5185 1547 5219
rect 1489 5179 1547 5185
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5216 2283 5219
rect 2682 5216 2688 5228
rect 2271 5188 2688 5216
rect 2271 5185 2283 5188
rect 2225 5179 2283 5185
rect 2682 5176 2688 5188
rect 2740 5176 2746 5228
rect 2777 5219 2835 5225
rect 2777 5185 2789 5219
rect 2823 5216 2835 5219
rect 2866 5216 2872 5228
rect 2823 5188 2872 5216
rect 2823 5185 2835 5188
rect 2777 5179 2835 5185
rect 2866 5176 2872 5188
rect 2924 5216 2930 5228
rect 4522 5216 4528 5228
rect 2924 5188 4528 5216
rect 2924 5176 2930 5188
rect 4522 5176 4528 5188
rect 4580 5176 4586 5228
rect 5445 5219 5503 5225
rect 5445 5216 5457 5219
rect 4632 5188 5457 5216
rect 2498 5108 2504 5160
rect 2556 5108 2562 5160
rect 3142 5108 3148 5160
rect 3200 5148 3206 5160
rect 3786 5148 3792 5160
rect 3200 5120 3792 5148
rect 3200 5108 3206 5120
rect 3786 5108 3792 5120
rect 3844 5148 3850 5160
rect 4632 5148 4660 5188
rect 5445 5185 5457 5188
rect 5491 5216 5503 5219
rect 6641 5219 6699 5225
rect 5491 5188 5764 5216
rect 5491 5185 5503 5188
rect 5445 5179 5503 5185
rect 3844 5120 4660 5148
rect 5169 5151 5227 5157
rect 3844 5108 3850 5120
rect 5169 5117 5181 5151
rect 5215 5117 5227 5151
rect 5736 5148 5764 5188
rect 6641 5185 6653 5219
rect 6687 5216 6699 5219
rect 7006 5216 7012 5228
rect 6687 5188 7012 5216
rect 6687 5185 6699 5188
rect 6641 5179 6699 5185
rect 7006 5176 7012 5188
rect 7064 5176 7070 5228
rect 7561 5219 7619 5225
rect 7561 5216 7573 5219
rect 7116 5188 7573 5216
rect 7116 5148 7144 5188
rect 7561 5185 7573 5188
rect 7607 5185 7619 5219
rect 7561 5179 7619 5185
rect 7650 5176 7656 5228
rect 7708 5216 7714 5228
rect 8404 5225 8432 5324
rect 8478 5244 8484 5296
rect 8536 5244 8542 5296
rect 8680 5284 8708 5324
rect 9490 5312 9496 5364
rect 9548 5352 9554 5364
rect 9548 5324 10640 5352
rect 9548 5312 9554 5324
rect 8680 5256 8800 5284
rect 8389 5219 8447 5225
rect 8389 5216 8401 5219
rect 7708 5188 8401 5216
rect 7708 5176 7714 5188
rect 8389 5185 8401 5188
rect 8435 5185 8447 5219
rect 8496 5216 8524 5244
rect 8652 5219 8710 5225
rect 8652 5216 8664 5219
rect 8496 5188 8664 5216
rect 8389 5179 8447 5185
rect 8652 5185 8664 5188
rect 8698 5185 8710 5219
rect 8772 5216 8800 5256
rect 8846 5244 8852 5296
rect 8904 5284 8910 5296
rect 10502 5284 10508 5296
rect 8904 5256 10508 5284
rect 8904 5244 8910 5256
rect 10502 5244 10508 5256
rect 10560 5244 10566 5296
rect 8772 5188 9674 5216
rect 8652 5179 8710 5185
rect 5736 5120 7144 5148
rect 5169 5111 5227 5117
rect 1578 4972 1584 5024
rect 1636 4972 1642 5024
rect 3510 4972 3516 5024
rect 3568 4972 3574 5024
rect 5184 5012 5212 5111
rect 7282 5108 7288 5160
rect 7340 5108 7346 5160
rect 9646 5148 9674 5188
rect 9766 5176 9772 5228
rect 9824 5216 9830 5228
rect 9953 5219 10011 5225
rect 9953 5216 9965 5219
rect 9824 5188 9965 5216
rect 9824 5176 9830 5188
rect 9953 5185 9965 5188
rect 9999 5216 10011 5219
rect 10042 5216 10048 5228
rect 9999 5188 10048 5216
rect 9999 5185 10011 5188
rect 9953 5179 10011 5185
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 10612 5225 10640 5324
rect 11330 5312 11336 5364
rect 11388 5352 11394 5364
rect 11609 5355 11667 5361
rect 11609 5352 11621 5355
rect 11388 5324 11621 5352
rect 11388 5312 11394 5324
rect 11609 5321 11621 5324
rect 11655 5321 11667 5355
rect 12526 5352 12532 5364
rect 11609 5315 11667 5321
rect 11992 5324 12532 5352
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5216 10655 5219
rect 10686 5216 10692 5228
rect 10643 5188 10692 5216
rect 10643 5185 10655 5188
rect 10597 5179 10655 5185
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 11793 5219 11851 5225
rect 11793 5185 11805 5219
rect 11839 5216 11851 5219
rect 11882 5216 11888 5228
rect 11839 5188 11888 5216
rect 11839 5185 11851 5188
rect 11793 5179 11851 5185
rect 11882 5176 11888 5188
rect 11940 5176 11946 5228
rect 11992 5225 12020 5324
rect 12526 5312 12532 5324
rect 12584 5352 12590 5364
rect 13722 5352 13728 5364
rect 12584 5324 13728 5352
rect 12584 5312 12590 5324
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 14366 5312 14372 5364
rect 14424 5352 14430 5364
rect 16853 5355 16911 5361
rect 14424 5324 16804 5352
rect 14424 5312 14430 5324
rect 16776 5284 16804 5324
rect 16853 5321 16865 5355
rect 16899 5352 16911 5355
rect 16942 5352 16948 5364
rect 16899 5324 16948 5352
rect 16899 5321 16911 5324
rect 16853 5315 16911 5321
rect 16942 5312 16948 5324
rect 17000 5312 17006 5364
rect 17052 5324 19840 5352
rect 17052 5284 17080 5324
rect 14660 5256 16712 5284
rect 16776 5256 17080 5284
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5185 12035 5219
rect 11977 5179 12035 5185
rect 12158 5176 12164 5228
rect 12216 5176 12222 5228
rect 13906 5176 13912 5228
rect 13964 5216 13970 5228
rect 14660 5225 14688 5256
rect 14645 5219 14703 5225
rect 14645 5216 14657 5219
rect 13964 5188 14657 5216
rect 13964 5176 13970 5188
rect 14645 5185 14657 5188
rect 14691 5185 14703 5219
rect 14645 5179 14703 5185
rect 14734 5176 14740 5228
rect 14792 5216 14798 5228
rect 16684 5225 16712 5256
rect 15749 5219 15807 5225
rect 15749 5216 15761 5219
rect 14792 5188 15761 5216
rect 14792 5176 14798 5188
rect 15749 5185 15761 5188
rect 15795 5185 15807 5219
rect 15749 5179 15807 5185
rect 16669 5219 16727 5225
rect 16669 5185 16681 5219
rect 16715 5216 16727 5219
rect 17221 5219 17279 5225
rect 17221 5216 17233 5219
rect 16715 5188 17233 5216
rect 16715 5185 16727 5188
rect 16669 5179 16727 5185
rect 17221 5185 17233 5188
rect 17267 5216 17279 5219
rect 17678 5216 17684 5228
rect 17267 5188 17684 5216
rect 17267 5185 17279 5188
rect 17221 5179 17279 5185
rect 17678 5176 17684 5188
rect 17736 5176 17742 5228
rect 18230 5176 18236 5228
rect 18288 5176 18294 5228
rect 18966 5176 18972 5228
rect 19024 5176 19030 5228
rect 19242 5176 19248 5228
rect 19300 5176 19306 5228
rect 10321 5151 10379 5157
rect 10321 5148 10333 5151
rect 9646 5120 10333 5148
rect 10321 5117 10333 5120
rect 10367 5117 10379 5151
rect 10321 5111 10379 5117
rect 6181 5083 6239 5089
rect 6181 5049 6193 5083
rect 6227 5080 6239 5083
rect 6546 5080 6552 5092
rect 6227 5052 6552 5080
rect 6227 5049 6239 5052
rect 6181 5043 6239 5049
rect 6546 5040 6552 5052
rect 6604 5040 6610 5092
rect 6362 5012 6368 5024
rect 5184 4984 6368 5012
rect 6362 4972 6368 4984
rect 6420 5012 6426 5024
rect 7650 5012 7656 5024
rect 6420 4984 7656 5012
rect 6420 4972 6426 4984
rect 7650 4972 7656 4984
rect 7708 4972 7714 5024
rect 8297 5015 8355 5021
rect 8297 4981 8309 5015
rect 8343 5012 8355 5015
rect 8846 5012 8852 5024
rect 8343 4984 8852 5012
rect 8343 4981 8355 4984
rect 8297 4975 8355 4981
rect 8846 4972 8852 4984
rect 8904 4972 8910 5024
rect 9401 5015 9459 5021
rect 9401 4981 9413 5015
rect 9447 5012 9459 5015
rect 10042 5012 10048 5024
rect 9447 4984 10048 5012
rect 9447 4981 9459 4984
rect 9401 4975 9459 4981
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 10137 5015 10195 5021
rect 10137 4981 10149 5015
rect 10183 5012 10195 5015
rect 10336 5012 10364 5111
rect 12342 5108 12348 5160
rect 12400 5148 12406 5160
rect 13078 5157 13084 5160
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 12400 5120 12909 5148
rect 12400 5108 12406 5120
rect 12897 5117 12909 5120
rect 12943 5117 12955 5151
rect 12897 5111 12955 5117
rect 13035 5151 13084 5157
rect 13035 5117 13047 5151
rect 13081 5117 13084 5151
rect 13035 5111 13084 5117
rect 13078 5108 13084 5111
rect 13136 5108 13142 5160
rect 13173 5151 13231 5157
rect 13173 5117 13185 5151
rect 13219 5148 13231 5151
rect 13219 5120 13584 5148
rect 13219 5117 13231 5120
rect 13173 5111 13231 5117
rect 11333 5083 11391 5089
rect 11333 5049 11345 5083
rect 11379 5080 11391 5083
rect 11379 5052 12204 5080
rect 11379 5049 11391 5052
rect 11333 5043 11391 5049
rect 11422 5012 11428 5024
rect 10183 4984 11428 5012
rect 10183 4981 10195 4984
rect 10137 4975 10195 4981
rect 11422 4972 11428 4984
rect 11480 4972 11486 5024
rect 12176 5012 12204 5052
rect 12250 5040 12256 5092
rect 12308 5080 12314 5092
rect 12621 5083 12679 5089
rect 12621 5080 12633 5083
rect 12308 5052 12633 5080
rect 12308 5040 12314 5052
rect 12621 5049 12633 5052
rect 12667 5049 12679 5083
rect 12621 5043 12679 5049
rect 13556 5012 13584 5120
rect 14366 5108 14372 5160
rect 14424 5108 14430 5160
rect 15010 5108 15016 5160
rect 15068 5148 15074 5160
rect 15473 5151 15531 5157
rect 15473 5148 15485 5151
rect 15068 5120 15485 5148
rect 15068 5108 15074 5120
rect 15473 5117 15485 5120
rect 15519 5117 15531 5151
rect 16942 5148 16948 5160
rect 15473 5111 15531 5117
rect 16408 5120 16948 5148
rect 15286 5040 15292 5092
rect 15344 5080 15350 5092
rect 15381 5083 15439 5089
rect 15381 5080 15393 5083
rect 15344 5052 15393 5080
rect 15344 5040 15350 5052
rect 15381 5049 15393 5052
rect 15427 5049 15439 5083
rect 15381 5043 15439 5049
rect 12176 4984 13584 5012
rect 13817 5015 13875 5021
rect 13817 4981 13829 5015
rect 13863 5012 13875 5015
rect 14826 5012 14832 5024
rect 13863 4984 14832 5012
rect 13863 4981 13875 4984
rect 13817 4975 13875 4981
rect 14826 4972 14832 4984
rect 14884 4972 14890 5024
rect 15488 5012 15516 5111
rect 16408 5012 16436 5120
rect 16942 5108 16948 5120
rect 17000 5108 17006 5160
rect 18046 5108 18052 5160
rect 18104 5108 18110 5160
rect 19107 5151 19165 5157
rect 19107 5117 19119 5151
rect 19153 5148 19165 5151
rect 19426 5148 19432 5160
rect 19153 5120 19432 5148
rect 19153 5117 19165 5120
rect 19107 5111 19165 5117
rect 19426 5108 19432 5120
rect 19484 5108 19490 5160
rect 19812 5148 19840 5324
rect 20622 5312 20628 5364
rect 20680 5352 20686 5364
rect 24578 5352 24584 5364
rect 20680 5324 24584 5352
rect 20680 5312 20686 5324
rect 24578 5312 24584 5324
rect 24636 5352 24642 5364
rect 27706 5352 27712 5364
rect 24636 5324 27712 5352
rect 24636 5312 24642 5324
rect 27706 5312 27712 5324
rect 27764 5312 27770 5364
rect 27985 5355 28043 5361
rect 27985 5321 27997 5355
rect 28031 5352 28043 5355
rect 30926 5352 30932 5364
rect 28031 5324 30932 5352
rect 28031 5321 28043 5324
rect 27985 5315 28043 5321
rect 30926 5312 30932 5324
rect 30984 5312 30990 5364
rect 31018 5312 31024 5364
rect 31076 5352 31082 5364
rect 31076 5324 31800 5352
rect 31076 5312 31082 5324
rect 20438 5244 20444 5296
rect 20496 5284 20502 5296
rect 26145 5287 26203 5293
rect 26145 5284 26157 5287
rect 20496 5256 26157 5284
rect 20496 5244 20502 5256
rect 26145 5253 26157 5256
rect 26191 5253 26203 5287
rect 26145 5247 26203 5253
rect 19889 5219 19947 5225
rect 19889 5185 19901 5219
rect 19935 5216 19947 5219
rect 20165 5219 20223 5225
rect 20165 5216 20177 5219
rect 19935 5188 20177 5216
rect 19935 5185 19947 5188
rect 19889 5179 19947 5185
rect 20165 5185 20177 5188
rect 20211 5185 20223 5219
rect 20165 5179 20223 5185
rect 21085 5219 21143 5225
rect 21085 5185 21097 5219
rect 21131 5216 21143 5219
rect 21542 5216 21548 5228
rect 21131 5188 21548 5216
rect 21131 5185 21143 5188
rect 21085 5179 21143 5185
rect 21542 5176 21548 5188
rect 21600 5176 21606 5228
rect 22097 5219 22155 5225
rect 22097 5185 22109 5219
rect 22143 5216 22155 5219
rect 22554 5216 22560 5228
rect 22143 5188 22560 5216
rect 22143 5185 22155 5188
rect 22097 5179 22155 5185
rect 22554 5176 22560 5188
rect 22612 5216 22618 5228
rect 22649 5219 22707 5225
rect 22649 5216 22661 5219
rect 22612 5188 22661 5216
rect 22612 5176 22618 5188
rect 22649 5185 22661 5188
rect 22695 5185 22707 5219
rect 22649 5179 22707 5185
rect 24946 5176 24952 5228
rect 25004 5176 25010 5228
rect 25133 5219 25191 5225
rect 25133 5185 25145 5219
rect 25179 5216 25191 5219
rect 25590 5216 25596 5228
rect 25179 5188 25596 5216
rect 25179 5185 25191 5188
rect 25133 5179 25191 5185
rect 25590 5176 25596 5188
rect 25648 5176 25654 5228
rect 22370 5148 22376 5160
rect 19812 5120 22376 5148
rect 22370 5108 22376 5120
rect 22428 5108 22434 5160
rect 24964 5148 24992 5176
rect 26050 5148 26056 5160
rect 24964 5120 26056 5148
rect 26050 5108 26056 5120
rect 26108 5108 26114 5160
rect 16485 5083 16543 5089
rect 16485 5049 16497 5083
rect 16531 5080 16543 5083
rect 18693 5083 18751 5089
rect 18693 5080 18705 5083
rect 16531 5052 17080 5080
rect 16531 5049 16543 5052
rect 16485 5043 16543 5049
rect 15488 4984 16436 5012
rect 17052 5012 17080 5052
rect 17604 5052 18705 5080
rect 17604 5012 17632 5052
rect 18693 5049 18705 5052
rect 18739 5049 18751 5083
rect 18693 5043 18751 5049
rect 19978 5040 19984 5092
rect 20036 5040 20042 5092
rect 24854 5080 24860 5092
rect 23308 5052 24860 5080
rect 17052 4984 17632 5012
rect 17957 5015 18015 5021
rect 17957 4981 17969 5015
rect 18003 5012 18015 5015
rect 18598 5012 18604 5024
rect 18003 4984 18604 5012
rect 18003 4981 18015 4984
rect 17957 4975 18015 4981
rect 18598 4972 18604 4984
rect 18656 4972 18662 5024
rect 19150 4972 19156 5024
rect 19208 5012 19214 5024
rect 20898 5012 20904 5024
rect 19208 4984 20904 5012
rect 19208 4972 19214 4984
rect 20898 4972 20904 4984
rect 20956 4972 20962 5024
rect 21269 5015 21327 5021
rect 21269 4981 21281 5015
rect 21315 5012 21327 5015
rect 21726 5012 21732 5024
rect 21315 4984 21732 5012
rect 21315 4981 21327 4984
rect 21269 4975 21327 4981
rect 21726 4972 21732 4984
rect 21784 4972 21790 5024
rect 22281 5015 22339 5021
rect 22281 4981 22293 5015
rect 22327 5012 22339 5015
rect 23308 5012 23336 5052
rect 24854 5040 24860 5052
rect 24912 5040 24918 5092
rect 22327 4984 23336 5012
rect 23385 5015 23443 5021
rect 22327 4981 22339 4984
rect 22281 4975 22339 4981
rect 23385 4981 23397 5015
rect 23431 5012 23443 5015
rect 23566 5012 23572 5024
rect 23431 4984 23572 5012
rect 23431 4981 23443 4984
rect 23385 4975 23443 4981
rect 23566 4972 23572 4984
rect 23624 4972 23630 5024
rect 24118 4972 24124 5024
rect 24176 5012 24182 5024
rect 24949 5015 25007 5021
rect 24949 5012 24961 5015
rect 24176 4984 24961 5012
rect 24176 4972 24182 4984
rect 24949 4981 24961 4984
rect 24995 4981 25007 5015
rect 26160 5012 26188 5247
rect 26418 5244 26424 5296
rect 26476 5284 26482 5296
rect 31386 5284 31392 5296
rect 26476 5256 31392 5284
rect 26476 5244 26482 5256
rect 31386 5244 31392 5256
rect 31444 5244 31450 5296
rect 31772 5284 31800 5324
rect 31846 5312 31852 5364
rect 31904 5352 31910 5364
rect 32674 5352 32680 5364
rect 31904 5324 32680 5352
rect 31904 5312 31910 5324
rect 32674 5312 32680 5324
rect 32732 5312 32738 5364
rect 38562 5312 38568 5364
rect 38620 5312 38626 5364
rect 39390 5312 39396 5364
rect 39448 5312 39454 5364
rect 32766 5284 32772 5296
rect 31772 5256 32772 5284
rect 32766 5244 32772 5256
rect 32824 5284 32830 5296
rect 35250 5284 35256 5296
rect 32824 5256 35256 5284
rect 32824 5244 32830 5256
rect 35250 5244 35256 5256
rect 35308 5244 35314 5296
rect 27154 5176 27160 5228
rect 27212 5216 27218 5228
rect 27249 5219 27307 5225
rect 27249 5216 27261 5219
rect 27212 5188 27261 5216
rect 27212 5176 27218 5188
rect 27249 5185 27261 5188
rect 27295 5185 27307 5219
rect 27249 5179 27307 5185
rect 27706 5176 27712 5228
rect 27764 5216 27770 5228
rect 28169 5219 28227 5225
rect 28169 5216 28181 5219
rect 27764 5188 28181 5216
rect 27764 5176 27770 5188
rect 28169 5185 28181 5188
rect 28215 5216 28227 5219
rect 28258 5216 28264 5228
rect 28215 5188 28264 5216
rect 28215 5185 28227 5188
rect 28169 5179 28227 5185
rect 28258 5176 28264 5188
rect 28316 5176 28322 5228
rect 28813 5219 28871 5225
rect 28813 5185 28825 5219
rect 28859 5216 28871 5219
rect 28859 5188 29132 5216
rect 28859 5185 28871 5188
rect 28813 5179 28871 5185
rect 26973 5151 27031 5157
rect 26973 5148 26985 5151
rect 26344 5120 26985 5148
rect 26344 5092 26372 5120
rect 26973 5117 26985 5120
rect 27019 5117 27031 5151
rect 26973 5111 27031 5117
rect 28074 5108 28080 5160
rect 28132 5148 28138 5160
rect 28537 5151 28595 5157
rect 28537 5148 28549 5151
rect 28132 5120 28549 5148
rect 28132 5108 28138 5120
rect 28537 5117 28549 5120
rect 28583 5117 28595 5151
rect 29104 5148 29132 5188
rect 30558 5176 30564 5228
rect 30616 5216 30622 5228
rect 32125 5219 32183 5225
rect 32125 5216 32137 5219
rect 30616 5188 32137 5216
rect 30616 5176 30622 5188
rect 32125 5185 32137 5188
rect 32171 5185 32183 5219
rect 32125 5179 32183 5185
rect 32306 5176 32312 5228
rect 32364 5176 32370 5228
rect 35713 5219 35771 5225
rect 35713 5185 35725 5219
rect 35759 5216 35771 5219
rect 35894 5216 35900 5228
rect 35759 5188 35900 5216
rect 35759 5185 35771 5188
rect 35713 5179 35771 5185
rect 35894 5176 35900 5188
rect 35952 5176 35958 5228
rect 38746 5176 38752 5228
rect 38804 5176 38810 5228
rect 38841 5219 38899 5225
rect 38841 5185 38853 5219
rect 38887 5185 38899 5219
rect 38841 5179 38899 5185
rect 39209 5219 39267 5225
rect 39209 5185 39221 5219
rect 39255 5216 39267 5219
rect 39666 5216 39672 5228
rect 39255 5188 39672 5216
rect 39255 5185 39267 5188
rect 39209 5179 39267 5185
rect 29270 5148 29276 5160
rect 29104 5120 29276 5148
rect 28537 5111 28595 5117
rect 29270 5108 29276 5120
rect 29328 5108 29334 5160
rect 31478 5108 31484 5160
rect 31536 5148 31542 5160
rect 32674 5148 32680 5160
rect 31536 5120 32680 5148
rect 31536 5108 31542 5120
rect 32674 5108 32680 5120
rect 32732 5108 32738 5160
rect 38856 5148 38884 5179
rect 39666 5176 39672 5188
rect 39724 5176 39730 5228
rect 32784 5120 38884 5148
rect 26326 5040 26332 5092
rect 26384 5040 26390 5092
rect 28353 5015 28411 5021
rect 28353 5012 28365 5015
rect 26160 4984 28365 5012
rect 24949 4975 25007 4981
rect 28353 4981 28365 4984
rect 28399 5012 28411 5015
rect 29454 5012 29460 5024
rect 28399 4984 29460 5012
rect 28399 4981 28411 4984
rect 28353 4975 28411 4981
rect 29454 4972 29460 4984
rect 29512 4972 29518 5024
rect 29549 5015 29607 5021
rect 29549 4981 29561 5015
rect 29595 5012 29607 5015
rect 31846 5012 31852 5024
rect 29595 4984 31852 5012
rect 29595 4981 29607 4984
rect 29549 4975 29607 4981
rect 31846 4972 31852 4984
rect 31904 4972 31910 5024
rect 32306 4972 32312 5024
rect 32364 5012 32370 5024
rect 32784 5012 32812 5120
rect 33962 5040 33968 5092
rect 34020 5080 34026 5092
rect 38654 5080 38660 5092
rect 34020 5052 38660 5080
rect 34020 5040 34026 5052
rect 38654 5040 38660 5052
rect 38712 5040 38718 5092
rect 32364 4984 32812 5012
rect 32364 4972 32370 4984
rect 35066 4972 35072 5024
rect 35124 5012 35130 5024
rect 35529 5015 35587 5021
rect 35529 5012 35541 5015
rect 35124 4984 35541 5012
rect 35124 4972 35130 4984
rect 35529 4981 35541 4984
rect 35575 4981 35587 5015
rect 35529 4975 35587 4981
rect 39022 4972 39028 5024
rect 39080 4972 39086 5024
rect 1104 4922 39836 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 37950 4922
rect 38002 4870 38014 4922
rect 38066 4870 38078 4922
rect 38130 4870 38142 4922
rect 38194 4870 38206 4922
rect 38258 4870 39836 4922
rect 1104 4848 39836 4870
rect 1578 4768 1584 4820
rect 1636 4808 1642 4820
rect 1636 4780 6868 4808
rect 1636 4768 1642 4780
rect 1673 4743 1731 4749
rect 1673 4709 1685 4743
rect 1719 4740 1731 4743
rect 1854 4740 1860 4752
rect 1719 4712 1860 4740
rect 1719 4709 1731 4712
rect 1673 4703 1731 4709
rect 1854 4700 1860 4712
rect 1912 4700 1918 4752
rect 3053 4743 3111 4749
rect 3053 4709 3065 4743
rect 3099 4740 3111 4743
rect 3418 4740 3424 4752
rect 3099 4712 3424 4740
rect 3099 4709 3111 4712
rect 3053 4703 3111 4709
rect 3418 4700 3424 4712
rect 3476 4700 3482 4752
rect 5902 4632 5908 4684
rect 5960 4632 5966 4684
rect 566 4564 572 4616
rect 624 4604 630 4616
rect 1765 4607 1823 4613
rect 1765 4604 1777 4607
rect 624 4576 1777 4604
rect 624 4564 630 4576
rect 1765 4573 1777 4576
rect 1811 4573 1823 4607
rect 1765 4567 1823 4573
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4573 2099 4607
rect 2041 4567 2099 4573
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4604 2375 4607
rect 2774 4604 2780 4616
rect 2363 4576 2780 4604
rect 2363 4573 2375 4576
rect 2317 4567 2375 4573
rect 750 4496 756 4548
rect 808 4536 814 4548
rect 1489 4539 1547 4545
rect 1489 4536 1501 4539
rect 808 4508 1501 4536
rect 808 4496 814 4508
rect 1489 4505 1501 4508
rect 1535 4505 1547 4539
rect 2056 4536 2084 4567
rect 2774 4564 2780 4576
rect 2832 4564 2838 4616
rect 4522 4564 4528 4616
rect 4580 4564 4586 4616
rect 4798 4564 4804 4616
rect 4856 4604 4862 4616
rect 4856 4576 6132 4604
rect 4856 4564 4862 4576
rect 2498 4536 2504 4548
rect 2056 4508 2504 4536
rect 1489 4499 1547 4505
rect 2498 4496 2504 4508
rect 2556 4496 2562 4548
rect 5994 4536 6000 4548
rect 3712 4508 6000 4536
rect 1949 4471 2007 4477
rect 1949 4437 1961 4471
rect 1995 4468 2007 4471
rect 3712 4468 3740 4508
rect 5994 4496 6000 4508
rect 6052 4496 6058 4548
rect 1995 4440 3740 4468
rect 3789 4471 3847 4477
rect 1995 4437 2007 4440
rect 1949 4431 2007 4437
rect 3789 4437 3801 4471
rect 3835 4468 3847 4471
rect 4706 4468 4712 4480
rect 3835 4440 4712 4468
rect 3835 4437 3847 4440
rect 3789 4431 3847 4437
rect 4706 4428 4712 4440
rect 4764 4428 4770 4480
rect 6104 4468 6132 4576
rect 6178 4564 6184 4616
rect 6236 4564 6242 4616
rect 6840 4604 6868 4780
rect 7006 4768 7012 4820
rect 7064 4768 7070 4820
rect 7466 4768 7472 4820
rect 7524 4808 7530 4820
rect 8113 4811 8171 4817
rect 8113 4808 8125 4811
rect 7524 4780 8125 4808
rect 7524 4768 7530 4780
rect 8113 4777 8125 4780
rect 8159 4777 8171 4811
rect 9766 4808 9772 4820
rect 8113 4771 8171 4777
rect 8220 4780 9772 4808
rect 6917 4743 6975 4749
rect 6917 4709 6929 4743
rect 6963 4740 6975 4743
rect 6963 4712 7604 4740
rect 6963 4709 6975 4712
rect 6917 4703 6975 4709
rect 7576 4681 7604 4712
rect 7834 4700 7840 4752
rect 7892 4740 7898 4752
rect 8220 4740 8248 4780
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 10594 4768 10600 4820
rect 10652 4808 10658 4820
rect 10781 4811 10839 4817
rect 10781 4808 10793 4811
rect 10652 4780 10793 4808
rect 10652 4768 10658 4780
rect 10781 4777 10793 4780
rect 10827 4777 10839 4811
rect 10781 4771 10839 4777
rect 10962 4768 10968 4820
rect 11020 4768 11026 4820
rect 12161 4811 12219 4817
rect 12161 4777 12173 4811
rect 12207 4808 12219 4811
rect 12250 4808 12256 4820
rect 12207 4780 12256 4808
rect 12207 4777 12219 4780
rect 12161 4771 12219 4777
rect 12250 4768 12256 4780
rect 12308 4768 12314 4820
rect 12360 4780 13492 4808
rect 7892 4712 8248 4740
rect 7892 4700 7898 4712
rect 8294 4700 8300 4752
rect 8352 4740 8358 4752
rect 8754 4740 8760 4752
rect 8352 4712 8760 4740
rect 8352 4700 8358 4712
rect 8754 4700 8760 4712
rect 8812 4700 8818 4752
rect 7561 4675 7619 4681
rect 7561 4641 7573 4675
rect 7607 4641 7619 4675
rect 7561 4635 7619 4641
rect 7650 4632 7656 4684
rect 7708 4672 7714 4684
rect 12360 4672 12388 4780
rect 13464 4752 13492 4780
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 14737 4811 14795 4817
rect 14737 4808 14749 4811
rect 13872 4780 14749 4808
rect 13872 4768 13878 4780
rect 14737 4777 14749 4780
rect 14783 4777 14795 4811
rect 16853 4811 16911 4817
rect 14737 4771 14795 4777
rect 14844 4780 15884 4808
rect 13446 4700 13452 4752
rect 13504 4740 13510 4752
rect 14182 4740 14188 4752
rect 13504 4712 14188 4740
rect 13504 4700 13510 4712
rect 14182 4700 14188 4712
rect 14240 4700 14246 4752
rect 14274 4700 14280 4752
rect 14332 4740 14338 4752
rect 14844 4740 14872 4780
rect 14332 4712 14872 4740
rect 14332 4700 14338 4712
rect 15856 4684 15884 4780
rect 16853 4777 16865 4811
rect 16899 4808 16911 4811
rect 19334 4808 19340 4820
rect 16899 4780 19340 4808
rect 16899 4777 16911 4780
rect 16853 4771 16911 4777
rect 19334 4768 19340 4780
rect 19392 4768 19398 4820
rect 19426 4768 19432 4820
rect 19484 4808 19490 4820
rect 19978 4808 19984 4820
rect 19484 4780 19984 4808
rect 19484 4768 19490 4780
rect 19978 4768 19984 4780
rect 20036 4768 20042 4820
rect 21450 4808 21456 4820
rect 20088 4780 21456 4808
rect 18322 4700 18328 4752
rect 18380 4740 18386 4752
rect 19150 4740 19156 4752
rect 18380 4712 19156 4740
rect 18380 4700 18386 4712
rect 19150 4700 19156 4712
rect 19208 4700 19214 4752
rect 19242 4700 19248 4752
rect 19300 4740 19306 4752
rect 19300 4712 19564 4740
rect 19300 4700 19306 4712
rect 7708 4644 10640 4672
rect 7708 4632 7714 4644
rect 6840 4576 7788 4604
rect 6730 4496 6736 4548
rect 6788 4536 6794 4548
rect 7377 4539 7435 4545
rect 7377 4536 7389 4539
rect 6788 4508 7389 4536
rect 6788 4496 6794 4508
rect 7377 4505 7389 4508
rect 7423 4536 7435 4539
rect 7650 4536 7656 4548
rect 7423 4508 7656 4536
rect 7423 4505 7435 4508
rect 7377 4499 7435 4505
rect 7650 4496 7656 4508
rect 7708 4496 7714 4548
rect 7760 4536 7788 4576
rect 8294 4564 8300 4616
rect 8352 4564 8358 4616
rect 9766 4536 9772 4548
rect 7760 4508 9772 4536
rect 9766 4496 9772 4508
rect 9824 4496 9830 4548
rect 10612 4536 10640 4644
rect 11072 4644 12388 4672
rect 10686 4564 10692 4616
rect 10744 4604 10750 4616
rect 11072 4604 11100 4644
rect 13630 4632 13636 4684
rect 13688 4672 13694 4684
rect 14366 4672 14372 4684
rect 13688 4644 14372 4672
rect 13688 4632 13694 4644
rect 14366 4632 14372 4644
rect 14424 4632 14430 4684
rect 15838 4632 15844 4684
rect 15896 4632 15902 4684
rect 19536 4681 19564 4712
rect 20088 4684 20116 4780
rect 21450 4768 21456 4780
rect 21508 4768 21514 4820
rect 23124 4780 25176 4808
rect 21269 4743 21327 4749
rect 21269 4709 21281 4743
rect 21315 4709 21327 4743
rect 22830 4740 22836 4752
rect 21269 4703 21327 4709
rect 22388 4712 22836 4740
rect 19521 4675 19579 4681
rect 19521 4641 19533 4675
rect 19567 4641 19579 4675
rect 19521 4635 19579 4641
rect 19886 4632 19892 4684
rect 19944 4672 19950 4684
rect 19981 4675 20039 4681
rect 19981 4672 19993 4675
rect 19944 4644 19993 4672
rect 19944 4632 19950 4644
rect 19981 4641 19993 4644
rect 20027 4641 20039 4675
rect 19981 4635 20039 4641
rect 20070 4632 20076 4684
rect 20128 4672 20134 4684
rect 20374 4675 20432 4681
rect 20374 4672 20386 4675
rect 20128 4644 20386 4672
rect 20128 4632 20134 4644
rect 20374 4641 20386 4644
rect 20420 4641 20432 4675
rect 20374 4635 20432 4641
rect 20533 4675 20591 4681
rect 20533 4641 20545 4675
rect 20579 4672 20591 4675
rect 21284 4672 21312 4703
rect 20579 4644 21312 4672
rect 20579 4641 20591 4644
rect 20533 4635 20591 4641
rect 22278 4632 22284 4684
rect 22336 4632 22342 4684
rect 22388 4681 22416 4712
rect 22830 4700 22836 4712
rect 22888 4700 22894 4752
rect 22373 4675 22431 4681
rect 22373 4641 22385 4675
rect 22419 4641 22431 4675
rect 22373 4635 22431 4641
rect 22462 4632 22468 4684
rect 22520 4672 22526 4684
rect 22557 4675 22615 4681
rect 22557 4672 22569 4675
rect 22520 4644 22569 4672
rect 22520 4632 22526 4644
rect 22557 4641 22569 4644
rect 22603 4641 22615 4675
rect 22557 4635 22615 4641
rect 23014 4632 23020 4684
rect 23072 4632 23078 4684
rect 23124 4672 23152 4780
rect 23293 4675 23351 4681
rect 23293 4672 23305 4675
rect 23124 4644 23305 4672
rect 23293 4641 23305 4644
rect 23339 4641 23351 4675
rect 23293 4635 23351 4641
rect 23431 4675 23489 4681
rect 23431 4641 23443 4675
rect 23477 4672 23489 4675
rect 25148 4672 25176 4780
rect 25590 4768 25596 4820
rect 25648 4768 25654 4820
rect 27249 4811 27307 4817
rect 27249 4777 27261 4811
rect 27295 4808 27307 4811
rect 28905 4811 28963 4817
rect 27295 4780 28856 4808
rect 27295 4777 27307 4780
rect 27249 4771 27307 4777
rect 25501 4743 25559 4749
rect 25501 4709 25513 4743
rect 25547 4740 25559 4743
rect 28828 4740 28856 4780
rect 28905 4777 28917 4811
rect 28951 4808 28963 4811
rect 29638 4808 29644 4820
rect 28951 4780 29644 4808
rect 28951 4777 28963 4780
rect 28905 4771 28963 4777
rect 29638 4768 29644 4780
rect 29696 4768 29702 4820
rect 31478 4808 31484 4820
rect 30024 4780 31484 4808
rect 30024 4740 30052 4780
rect 31478 4768 31484 4780
rect 31536 4768 31542 4820
rect 31588 4780 31892 4808
rect 25547 4712 26188 4740
rect 28828 4712 30052 4740
rect 25547 4709 25559 4712
rect 25501 4703 25559 4709
rect 23477 4644 24440 4672
rect 25148 4644 25820 4672
rect 23477 4641 23489 4644
rect 23431 4635 23489 4641
rect 10744 4576 11100 4604
rect 10744 4564 10750 4576
rect 11146 4564 11152 4616
rect 11204 4564 11210 4616
rect 12894 4564 12900 4616
rect 12952 4564 12958 4616
rect 13173 4607 13231 4613
rect 13173 4573 13185 4607
rect 13219 4573 13231 4607
rect 13173 4567 13231 4573
rect 13188 4536 13216 4567
rect 13722 4564 13728 4616
rect 13780 4604 13786 4616
rect 13780 4576 14872 4604
rect 13780 4564 13786 4576
rect 10612 4508 13216 4536
rect 7190 4468 7196 4480
rect 6104 4440 7196 4468
rect 7190 4428 7196 4440
rect 7248 4428 7254 4480
rect 7466 4428 7472 4480
rect 7524 4468 7530 4480
rect 10410 4468 10416 4480
rect 7524 4440 10416 4468
rect 7524 4428 7530 4440
rect 10410 4428 10416 4440
rect 10468 4428 10474 4480
rect 10502 4428 10508 4480
rect 10560 4468 10566 4480
rect 13078 4468 13084 4480
rect 10560 4440 13084 4468
rect 10560 4428 10566 4440
rect 13078 4428 13084 4440
rect 13136 4428 13142 4480
rect 13188 4468 13216 4508
rect 13814 4496 13820 4548
rect 13872 4536 13878 4548
rect 14734 4536 14740 4548
rect 13872 4508 14740 4536
rect 13872 4496 13878 4508
rect 14734 4496 14740 4508
rect 14792 4496 14798 4548
rect 14844 4536 14872 4576
rect 15470 4564 15476 4616
rect 15528 4564 15534 4616
rect 15749 4607 15807 4613
rect 15749 4573 15761 4607
rect 15795 4604 15807 4607
rect 16022 4604 16028 4616
rect 15795 4576 16028 4604
rect 15795 4573 15807 4576
rect 15749 4567 15807 4573
rect 16022 4564 16028 4576
rect 16080 4564 16086 4616
rect 16117 4607 16175 4613
rect 16117 4573 16129 4607
rect 16163 4600 16175 4607
rect 17405 4607 17463 4613
rect 16163 4573 16252 4600
rect 16117 4572 16252 4573
rect 16117 4567 16175 4572
rect 15194 4536 15200 4548
rect 14844 4508 15200 4536
rect 15194 4496 15200 4508
rect 15252 4496 15258 4548
rect 15488 4536 15516 4564
rect 16224 4536 16252 4572
rect 17405 4573 17417 4607
rect 17451 4604 17463 4607
rect 17586 4604 17592 4616
rect 17451 4576 17592 4604
rect 17451 4573 17463 4576
rect 17405 4567 17463 4573
rect 17586 4564 17592 4576
rect 17644 4564 17650 4616
rect 17678 4564 17684 4616
rect 17736 4564 17742 4616
rect 18230 4564 18236 4616
rect 18288 4604 18294 4616
rect 19242 4604 19248 4616
rect 18288 4576 19248 4604
rect 18288 4564 18294 4576
rect 19242 4564 19248 4576
rect 19300 4564 19306 4616
rect 19337 4607 19395 4613
rect 19337 4573 19349 4607
rect 19383 4594 19395 4607
rect 19426 4594 19432 4616
rect 19383 4573 19432 4594
rect 19337 4567 19432 4573
rect 19352 4566 19432 4567
rect 19426 4564 19432 4566
rect 19484 4564 19490 4616
rect 20254 4564 20260 4616
rect 20312 4564 20318 4616
rect 21542 4564 21548 4616
rect 21600 4604 21606 4616
rect 22005 4607 22063 4613
rect 22005 4604 22017 4607
rect 21600 4576 22017 4604
rect 21600 4564 21606 4576
rect 22005 4573 22017 4576
rect 22051 4573 22063 4607
rect 22005 4567 22063 4573
rect 23566 4564 23572 4616
rect 23624 4564 23630 4616
rect 15488 4508 16252 4536
rect 16942 4496 16948 4548
rect 17000 4536 17006 4548
rect 24412 4536 24440 4644
rect 24486 4564 24492 4616
rect 24544 4564 24550 4616
rect 24765 4607 24823 4613
rect 24765 4573 24777 4607
rect 24811 4604 24823 4607
rect 25314 4604 25320 4616
rect 24811 4576 25320 4604
rect 24811 4573 24823 4576
rect 24765 4567 24823 4573
rect 25314 4564 25320 4576
rect 25372 4564 25378 4616
rect 25792 4604 25820 4644
rect 25866 4632 25872 4684
rect 25924 4672 25930 4684
rect 26160 4681 26188 4712
rect 26053 4675 26111 4681
rect 26053 4672 26065 4675
rect 25924 4644 26065 4672
rect 25924 4632 25930 4644
rect 26053 4641 26065 4644
rect 26099 4641 26111 4675
rect 26053 4635 26111 4641
rect 26145 4675 26203 4681
rect 26145 4641 26157 4675
rect 26191 4641 26203 4675
rect 26145 4635 26203 4641
rect 26786 4632 26792 4684
rect 26844 4672 26850 4684
rect 27522 4672 27528 4684
rect 26844 4644 27528 4672
rect 26844 4632 26850 4644
rect 25961 4607 26019 4613
rect 25961 4604 25973 4607
rect 25792 4576 25973 4604
rect 25961 4573 25973 4576
rect 26007 4604 26019 4607
rect 26418 4604 26424 4616
rect 26007 4576 26424 4604
rect 26007 4573 26019 4576
rect 25961 4567 26019 4573
rect 26418 4564 26424 4576
rect 26476 4564 26482 4616
rect 27062 4564 27068 4616
rect 27120 4564 27126 4616
rect 27356 4613 27384 4644
rect 27522 4632 27528 4644
rect 27580 4632 27586 4684
rect 29454 4632 29460 4684
rect 29512 4672 29518 4684
rect 29917 4675 29975 4681
rect 29917 4672 29929 4675
rect 29512 4644 29929 4672
rect 29512 4632 29518 4644
rect 29917 4641 29929 4644
rect 29963 4641 29975 4675
rect 29917 4635 29975 4641
rect 27341 4607 27399 4613
rect 27341 4573 27353 4607
rect 27387 4573 27399 4607
rect 27341 4567 27399 4573
rect 27430 4564 27436 4616
rect 27488 4604 27494 4616
rect 27893 4607 27951 4613
rect 27893 4604 27905 4607
rect 27488 4576 27905 4604
rect 27488 4564 27494 4576
rect 27893 4573 27905 4576
rect 27939 4604 27951 4607
rect 28074 4604 28080 4616
rect 27939 4576 28080 4604
rect 27939 4573 27951 4576
rect 27893 4567 27951 4573
rect 28074 4564 28080 4576
rect 28132 4564 28138 4616
rect 28166 4564 28172 4616
rect 28224 4564 28230 4616
rect 28994 4564 29000 4616
rect 29052 4604 29058 4616
rect 29270 4604 29276 4616
rect 29052 4576 29276 4604
rect 29052 4564 29058 4576
rect 29270 4564 29276 4576
rect 29328 4564 29334 4616
rect 29546 4564 29552 4616
rect 29604 4604 29610 4616
rect 30193 4607 30251 4613
rect 30193 4604 30205 4607
rect 29604 4576 30205 4604
rect 29604 4564 29610 4576
rect 30193 4573 30205 4576
rect 30239 4604 30251 4607
rect 30466 4604 30472 4616
rect 30239 4576 30472 4604
rect 30239 4573 30251 4576
rect 30193 4567 30251 4573
rect 30466 4564 30472 4576
rect 30524 4564 30530 4616
rect 31588 4604 31616 4780
rect 31864 4740 31892 4780
rect 32674 4768 32680 4820
rect 32732 4808 32738 4820
rect 32732 4780 35480 4808
rect 32732 4768 32738 4780
rect 32306 4740 32312 4752
rect 31864 4712 32312 4740
rect 32306 4700 32312 4712
rect 32364 4700 32370 4752
rect 33873 4743 33931 4749
rect 33873 4709 33885 4743
rect 33919 4740 33931 4743
rect 33962 4740 33968 4752
rect 33919 4712 33968 4740
rect 33919 4709 33931 4712
rect 33873 4703 33931 4709
rect 33962 4700 33968 4712
rect 34020 4700 34026 4752
rect 34790 4700 34796 4752
rect 34848 4700 34854 4752
rect 34974 4700 34980 4752
rect 35032 4740 35038 4752
rect 35069 4743 35127 4749
rect 35069 4740 35081 4743
rect 35032 4712 35081 4740
rect 35032 4700 35038 4712
rect 35069 4709 35081 4712
rect 35115 4709 35127 4743
rect 35069 4703 35127 4709
rect 31754 4632 31760 4684
rect 31812 4632 31818 4684
rect 31846 4632 31852 4684
rect 31904 4672 31910 4684
rect 32401 4675 32459 4681
rect 32401 4672 32413 4675
rect 31904 4644 32413 4672
rect 31904 4632 31910 4644
rect 32401 4641 32413 4644
rect 32447 4641 32459 4675
rect 32401 4635 32459 4641
rect 32674 4632 32680 4684
rect 32732 4632 32738 4684
rect 32766 4632 32772 4684
rect 32824 4681 32830 4684
rect 32824 4675 32852 4681
rect 32840 4641 32852 4675
rect 32824 4635 32852 4641
rect 32824 4632 32830 4635
rect 30944 4576 31616 4604
rect 31941 4607 31999 4613
rect 17000 4508 19472 4536
rect 24412 4508 24808 4536
rect 17000 4496 17006 4508
rect 18322 4468 18328 4480
rect 13188 4440 18328 4468
rect 18322 4428 18328 4440
rect 18380 4428 18386 4480
rect 18417 4471 18475 4477
rect 18417 4437 18429 4471
rect 18463 4468 18475 4471
rect 19242 4468 19248 4480
rect 18463 4440 19248 4468
rect 18463 4437 18475 4440
rect 18417 4431 18475 4437
rect 19242 4428 19248 4440
rect 19300 4428 19306 4480
rect 19444 4468 19472 4508
rect 24780 4480 24808 4508
rect 27706 4496 27712 4548
rect 27764 4536 27770 4548
rect 30944 4536 30972 4576
rect 31941 4573 31953 4607
rect 31987 4573 31999 4607
rect 31941 4567 31999 4573
rect 27764 4508 30972 4536
rect 27764 4496 27770 4508
rect 31018 4496 31024 4548
rect 31076 4496 31082 4548
rect 31202 4496 31208 4548
rect 31260 4496 31266 4548
rect 31846 4496 31852 4548
rect 31904 4536 31910 4548
rect 31956 4536 31984 4567
rect 32950 4564 32956 4616
rect 33008 4564 33014 4616
rect 33686 4564 33692 4616
rect 33744 4564 33750 4616
rect 34974 4564 34980 4616
rect 35032 4564 35038 4616
rect 35452 4613 35480 4780
rect 35894 4768 35900 4820
rect 35952 4768 35958 4820
rect 36814 4768 36820 4820
rect 36872 4808 36878 4820
rect 38289 4811 38347 4817
rect 38289 4808 38301 4811
rect 36872 4780 38301 4808
rect 36872 4768 36878 4780
rect 38289 4777 38301 4780
rect 38335 4777 38347 4811
rect 38289 4771 38347 4777
rect 39390 4768 39396 4820
rect 39448 4768 39454 4820
rect 36722 4700 36728 4752
rect 36780 4740 36786 4752
rect 38565 4743 38623 4749
rect 38565 4740 38577 4743
rect 36780 4712 38577 4740
rect 36780 4700 36786 4712
rect 38565 4709 38577 4712
rect 38611 4709 38623 4743
rect 38565 4703 38623 4709
rect 39025 4743 39083 4749
rect 39025 4709 39037 4743
rect 39071 4740 39083 4743
rect 39942 4740 39948 4752
rect 39071 4712 39948 4740
rect 39071 4709 39083 4712
rect 39025 4703 39083 4709
rect 39942 4700 39948 4712
rect 40000 4700 40006 4752
rect 35618 4632 35624 4684
rect 35676 4632 35682 4684
rect 36446 4632 36452 4684
rect 36504 4632 36510 4684
rect 37182 4632 37188 4684
rect 37240 4672 37246 4684
rect 37240 4644 39252 4672
rect 37240 4632 37246 4644
rect 35437 4607 35495 4613
rect 35437 4573 35449 4607
rect 35483 4573 35495 4607
rect 35437 4567 35495 4573
rect 38470 4564 38476 4616
rect 38528 4564 38534 4616
rect 38562 4564 38568 4616
rect 38620 4604 38626 4616
rect 39224 4613 39252 4644
rect 38749 4607 38807 4613
rect 38749 4604 38761 4607
rect 38620 4576 38761 4604
rect 38620 4564 38626 4576
rect 38749 4573 38761 4576
rect 38795 4573 38807 4607
rect 38749 4567 38807 4573
rect 38841 4607 38899 4613
rect 38841 4573 38853 4607
rect 38887 4573 38899 4607
rect 38841 4567 38899 4573
rect 39209 4607 39267 4613
rect 39209 4573 39221 4607
rect 39255 4573 39267 4607
rect 39209 4567 39267 4573
rect 31904 4508 31984 4536
rect 33520 4508 34928 4536
rect 31904 4496 31910 4508
rect 20622 4468 20628 4480
rect 19444 4440 20628 4468
rect 20622 4428 20628 4440
rect 20680 4428 20686 4480
rect 20806 4428 20812 4480
rect 20864 4468 20870 4480
rect 21177 4471 21235 4477
rect 21177 4468 21189 4471
rect 20864 4440 21189 4468
rect 20864 4428 20870 4440
rect 21177 4437 21189 4440
rect 21223 4437 21235 4471
rect 21177 4431 21235 4437
rect 21450 4428 21456 4480
rect 21508 4468 21514 4480
rect 24213 4471 24271 4477
rect 24213 4468 24225 4471
rect 21508 4440 24225 4468
rect 21508 4428 21514 4440
rect 24213 4437 24225 4440
rect 24259 4437 24271 4471
rect 24213 4431 24271 4437
rect 24762 4428 24768 4480
rect 24820 4428 24826 4480
rect 25314 4428 25320 4480
rect 25372 4468 25378 4480
rect 26050 4468 26056 4480
rect 25372 4440 26056 4468
rect 25372 4428 25378 4440
rect 26050 4428 26056 4440
rect 26108 4428 26114 4480
rect 26234 4428 26240 4480
rect 26292 4468 26298 4480
rect 27430 4468 27436 4480
rect 26292 4440 27436 4468
rect 26292 4428 26298 4440
rect 27430 4428 27436 4440
rect 27488 4428 27494 4480
rect 27522 4428 27528 4480
rect 27580 4428 27586 4480
rect 29178 4428 29184 4480
rect 29236 4428 29242 4480
rect 30558 4428 30564 4480
rect 30616 4468 30622 4480
rect 30929 4471 30987 4477
rect 30929 4468 30941 4471
rect 30616 4440 30941 4468
rect 30616 4428 30622 4440
rect 30929 4437 30941 4440
rect 30975 4437 30987 4471
rect 30929 4431 30987 4437
rect 31938 4428 31944 4480
rect 31996 4468 32002 4480
rect 33520 4468 33548 4508
rect 31996 4440 33548 4468
rect 31996 4428 32002 4440
rect 33594 4428 33600 4480
rect 33652 4428 33658 4480
rect 34900 4468 34928 4508
rect 35250 4496 35256 4548
rect 35308 4536 35314 4548
rect 36265 4539 36323 4545
rect 36265 4536 36277 4539
rect 35308 4508 36277 4536
rect 35308 4496 35314 4508
rect 36265 4505 36277 4508
rect 36311 4505 36323 4539
rect 36265 4499 36323 4505
rect 37274 4496 37280 4548
rect 37332 4536 37338 4548
rect 38856 4536 38884 4567
rect 37332 4508 38884 4536
rect 37332 4496 37338 4508
rect 35526 4468 35532 4480
rect 34900 4440 35532 4468
rect 35526 4428 35532 4440
rect 35584 4468 35590 4480
rect 36357 4471 36415 4477
rect 36357 4468 36369 4471
rect 35584 4440 36369 4468
rect 35584 4428 35590 4440
rect 36357 4437 36369 4440
rect 36403 4437 36415 4471
rect 36357 4431 36415 4437
rect 1104 4378 39836 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 39010 4378
rect 39062 4326 39074 4378
rect 39126 4326 39138 4378
rect 39190 4326 39202 4378
rect 39254 4326 39266 4378
rect 39318 4326 39836 4378
rect 1104 4304 39836 4326
rect 1946 4224 1952 4276
rect 2004 4224 2010 4276
rect 3053 4267 3111 4273
rect 3053 4233 3065 4267
rect 3099 4264 3111 4267
rect 4338 4264 4344 4276
rect 3099 4236 4344 4264
rect 3099 4233 3111 4236
rect 3053 4227 3111 4233
rect 4338 4224 4344 4236
rect 4396 4224 4402 4276
rect 6546 4224 6552 4276
rect 6604 4264 6610 4276
rect 7006 4264 7012 4276
rect 6604 4236 7012 4264
rect 6604 4224 6610 4236
rect 7006 4224 7012 4236
rect 7064 4224 7070 4276
rect 7282 4224 7288 4276
rect 7340 4264 7346 4276
rect 7340 4236 8156 4264
rect 7340 4224 7346 4236
rect 750 4156 756 4208
rect 808 4196 814 4208
rect 1489 4199 1547 4205
rect 1489 4196 1501 4199
rect 808 4168 1501 4196
rect 808 4156 814 4168
rect 1489 4165 1501 4168
rect 1535 4165 1547 4199
rect 1489 4159 1547 4165
rect 934 4088 940 4140
rect 992 4128 998 4140
rect 1765 4131 1823 4137
rect 1765 4128 1777 4131
rect 992 4100 1777 4128
rect 992 4088 998 4100
rect 1765 4097 1777 4100
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4097 2191 4131
rect 2133 4091 2191 4097
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4128 2467 4131
rect 2455 4100 2728 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 2148 4060 2176 4091
rect 2498 4060 2504 4072
rect 2148 4032 2504 4060
rect 2498 4020 2504 4032
rect 2556 4020 2562 4072
rect 1673 3995 1731 4001
rect 1673 3961 1685 3995
rect 1719 3992 1731 3995
rect 1719 3964 2268 3992
rect 1719 3961 1731 3964
rect 1673 3955 1731 3961
rect 2240 3924 2268 3964
rect 2314 3952 2320 4004
rect 2372 3952 2378 4004
rect 2590 3952 2596 4004
rect 2648 3952 2654 4004
rect 2700 4001 2728 4100
rect 4154 4088 4160 4140
rect 4212 4088 4218 4140
rect 4338 4137 4344 4140
rect 4316 4131 4344 4137
rect 4316 4097 4328 4131
rect 4316 4091 4344 4097
rect 4338 4088 4344 4091
rect 4396 4088 4402 4140
rect 4430 4088 4436 4140
rect 4488 4088 4494 4140
rect 5169 4131 5227 4137
rect 5169 4097 5181 4131
rect 5215 4128 5227 4131
rect 6365 4131 6423 4137
rect 5215 4100 6316 4128
rect 5215 4097 5227 4100
rect 5169 4091 5227 4097
rect 3142 4020 3148 4072
rect 3200 4020 3206 4072
rect 3329 4063 3387 4069
rect 3329 4029 3341 4063
rect 3375 4060 3387 4063
rect 3510 4060 3516 4072
rect 3375 4032 3516 4060
rect 3375 4029 3387 4032
rect 3329 4023 3387 4029
rect 3510 4020 3516 4032
rect 3568 4020 3574 4072
rect 4706 4020 4712 4072
rect 4764 4020 4770 4072
rect 5353 4063 5411 4069
rect 5353 4029 5365 4063
rect 5399 4060 5411 4063
rect 5442 4060 5448 4072
rect 5399 4032 5448 4060
rect 5399 4029 5411 4032
rect 5353 4023 5411 4029
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 6288 4060 6316 4100
rect 6365 4097 6377 4131
rect 6411 4128 6423 4131
rect 6730 4128 6736 4140
rect 6411 4100 6736 4128
rect 6411 4097 6423 4100
rect 6365 4091 6423 4097
rect 6730 4088 6736 4100
rect 6788 4088 6794 4140
rect 7558 4088 7564 4140
rect 7616 4088 7622 4140
rect 8128 4128 8156 4236
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 8481 4267 8539 4273
rect 8481 4264 8493 4267
rect 8352 4236 8493 4264
rect 8352 4224 8358 4236
rect 8481 4233 8493 4236
rect 8527 4233 8539 4267
rect 8481 4227 8539 4233
rect 8772 4236 11100 4264
rect 8772 4128 8800 4236
rect 10410 4137 10416 4140
rect 8128 4100 8800 4128
rect 8849 4131 8907 4137
rect 8849 4097 8861 4131
rect 8895 4097 8907 4131
rect 8849 4091 8907 4097
rect 8941 4131 8999 4137
rect 8941 4097 8953 4131
rect 8987 4128 8999 4131
rect 10367 4131 10416 4137
rect 8987 4100 9720 4128
rect 8987 4097 8999 4100
rect 8941 4091 8999 4097
rect 6546 4060 6552 4072
rect 6288 4032 6552 4060
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 7006 4020 7012 4072
rect 7064 4020 7070 4072
rect 7285 4063 7343 4069
rect 7285 4060 7297 4063
rect 7116 4032 7297 4060
rect 2685 3995 2743 4001
rect 2685 3961 2697 3995
rect 2731 3961 2743 3995
rect 2685 3955 2743 3961
rect 6914 3952 6920 4004
rect 6972 3992 6978 4004
rect 7116 3992 7144 4032
rect 7285 4029 7297 4032
rect 7331 4029 7343 4063
rect 7285 4023 7343 4029
rect 7423 4063 7481 4069
rect 7423 4029 7435 4063
rect 7469 4060 7481 4063
rect 7469 4032 7972 4060
rect 7469 4029 7481 4032
rect 7423 4023 7481 4029
rect 6972 3964 7144 3992
rect 6972 3952 6978 3964
rect 2866 3924 2872 3936
rect 2240 3896 2872 3924
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 3513 3927 3571 3933
rect 3513 3893 3525 3927
rect 3559 3924 3571 3927
rect 3786 3924 3792 3936
rect 3559 3896 3792 3924
rect 3559 3893 3571 3896
rect 3513 3887 3571 3893
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 7282 3924 7288 3936
rect 4028 3896 7288 3924
rect 4028 3884 4034 3896
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 7650 3884 7656 3936
rect 7708 3924 7714 3936
rect 7944 3924 7972 4032
rect 8754 4020 8760 4072
rect 8812 4060 8818 4072
rect 8864 4060 8892 4091
rect 9692 4072 9720 4100
rect 10367 4097 10379 4131
rect 10413 4097 10416 4131
rect 10367 4091 10416 4097
rect 10410 4088 10416 4091
rect 10468 4088 10474 4140
rect 8812 4032 8892 4060
rect 9033 4063 9091 4069
rect 8812 4020 8818 4032
rect 9033 4029 9045 4063
rect 9079 4029 9091 4063
rect 9033 4023 9091 4029
rect 8018 3952 8024 4004
rect 8076 3992 8082 4004
rect 8205 3995 8263 4001
rect 8205 3992 8217 3995
rect 8076 3964 8217 3992
rect 8076 3952 8082 3964
rect 8205 3961 8217 3964
rect 8251 3961 8263 3995
rect 8205 3955 8263 3961
rect 8846 3952 8852 4004
rect 8904 3992 8910 4004
rect 9048 3992 9076 4023
rect 9306 4020 9312 4072
rect 9364 4020 9370 4072
rect 9490 4020 9496 4072
rect 9548 4020 9554 4072
rect 9674 4020 9680 4072
rect 9732 4060 9738 4072
rect 10229 4063 10287 4069
rect 10229 4060 10241 4063
rect 9732 4032 10241 4060
rect 9732 4020 9738 4032
rect 10229 4029 10241 4032
rect 10275 4029 10287 4063
rect 10229 4023 10287 4029
rect 10502 4020 10508 4072
rect 10560 4020 10566 4072
rect 11072 4060 11100 4236
rect 11146 4224 11152 4276
rect 11204 4224 11210 4276
rect 11422 4224 11428 4276
rect 11480 4264 11486 4276
rect 11480 4236 13032 4264
rect 11480 4224 11486 4236
rect 13004 4196 13032 4236
rect 13078 4224 13084 4276
rect 13136 4264 13142 4276
rect 17218 4264 17224 4276
rect 13136 4236 17224 4264
rect 13136 4224 13142 4236
rect 17218 4224 17224 4236
rect 17276 4224 17282 4276
rect 18046 4224 18052 4276
rect 18104 4264 18110 4276
rect 19153 4267 19211 4273
rect 19153 4264 19165 4267
rect 18104 4236 19165 4264
rect 18104 4224 18110 4236
rect 19153 4233 19165 4236
rect 19199 4233 19211 4267
rect 19426 4264 19432 4276
rect 19153 4227 19211 4233
rect 19260 4236 19432 4264
rect 13630 4196 13636 4208
rect 13004 4168 13636 4196
rect 13630 4156 13636 4168
rect 13688 4156 13694 4208
rect 13814 4196 13820 4208
rect 13740 4168 13820 4196
rect 11238 4088 11244 4140
rect 11296 4128 11302 4140
rect 13170 4128 13176 4140
rect 11296 4100 13176 4128
rect 11296 4088 11302 4100
rect 13170 4088 13176 4100
rect 13228 4128 13234 4140
rect 13740 4128 13768 4168
rect 13814 4156 13820 4168
rect 13872 4156 13878 4208
rect 14108 4168 14320 4196
rect 14108 4128 14136 4168
rect 13228 4100 13768 4128
rect 13832 4100 14136 4128
rect 13228 4088 13234 4100
rect 13832 4060 13860 4100
rect 14182 4088 14188 4140
rect 14240 4088 14246 4140
rect 14292 4128 14320 4168
rect 14366 4156 14372 4208
rect 14424 4196 14430 4208
rect 15562 4196 15568 4208
rect 14424 4168 15568 4196
rect 14424 4156 14430 4168
rect 15562 4156 15568 4168
rect 15620 4156 15626 4208
rect 16850 4156 16856 4208
rect 16908 4196 16914 4208
rect 18966 4196 18972 4208
rect 16908 4168 18972 4196
rect 16908 4156 16914 4168
rect 18966 4156 18972 4168
rect 19024 4156 19030 4208
rect 19061 4199 19119 4205
rect 19061 4165 19073 4199
rect 19107 4196 19119 4199
rect 19260 4196 19288 4236
rect 19426 4224 19432 4236
rect 19484 4224 19490 4276
rect 19702 4224 19708 4276
rect 19760 4264 19766 4276
rect 20254 4264 20260 4276
rect 19760 4236 20260 4264
rect 19760 4224 19766 4236
rect 20254 4224 20260 4236
rect 20312 4264 20318 4276
rect 21818 4264 21824 4276
rect 20312 4236 21824 4264
rect 20312 4224 20318 4236
rect 21818 4224 21824 4236
rect 21876 4224 21882 4276
rect 22925 4267 22983 4273
rect 22925 4233 22937 4267
rect 22971 4264 22983 4267
rect 23014 4264 23020 4276
rect 22971 4236 23020 4264
rect 22971 4233 22983 4236
rect 22925 4227 22983 4233
rect 23014 4224 23020 4236
rect 23072 4224 23078 4276
rect 24949 4267 25007 4273
rect 24949 4233 24961 4267
rect 24995 4233 25007 4267
rect 24949 4227 25007 4233
rect 19107 4168 19288 4196
rect 19107 4165 19119 4168
rect 19061 4159 19119 4165
rect 19978 4156 19984 4208
rect 20036 4196 20042 4208
rect 20165 4199 20223 4205
rect 20165 4196 20177 4199
rect 20036 4168 20177 4196
rect 20036 4156 20042 4168
rect 20165 4165 20177 4168
rect 20211 4165 20223 4199
rect 20165 4159 20223 4165
rect 20456 4168 21864 4196
rect 15470 4128 15476 4140
rect 14292 4100 15476 4128
rect 15470 4088 15476 4100
rect 15528 4128 15534 4140
rect 15657 4131 15715 4137
rect 15657 4128 15669 4131
rect 15528 4100 15669 4128
rect 15528 4088 15534 4100
rect 15657 4097 15669 4100
rect 15703 4097 15715 4131
rect 15657 4091 15715 4097
rect 15746 4088 15752 4140
rect 15804 4128 15810 4140
rect 17954 4128 17960 4140
rect 15804 4100 17960 4128
rect 15804 4088 15810 4100
rect 17954 4088 17960 4100
rect 18012 4088 18018 4140
rect 18601 4131 18659 4137
rect 18601 4097 18613 4131
rect 18647 4128 18659 4131
rect 18647 4100 18736 4128
rect 18647 4097 18659 4100
rect 18601 4091 18659 4097
rect 11072 4032 13860 4060
rect 13909 4063 13967 4069
rect 13909 4029 13921 4063
rect 13955 4029 13967 4063
rect 17218 4060 17224 4072
rect 13909 4023 13967 4029
rect 14568 4032 17224 4060
rect 8904 3964 9076 3992
rect 9953 3995 10011 4001
rect 8904 3952 8910 3964
rect 9953 3961 9965 3995
rect 9999 3961 10011 3995
rect 9953 3955 10011 3961
rect 7708 3896 7972 3924
rect 7708 3884 7714 3896
rect 9306 3884 9312 3936
rect 9364 3924 9370 3936
rect 9766 3924 9772 3936
rect 9364 3896 9772 3924
rect 9364 3884 9370 3896
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 9968 3924 9996 3955
rect 10962 3952 10968 4004
rect 11020 3992 11026 4004
rect 12618 3992 12624 4004
rect 11020 3964 12624 3992
rect 11020 3952 11026 3964
rect 12618 3952 12624 3964
rect 12676 3952 12682 4004
rect 12986 3952 12992 4004
rect 13044 3992 13050 4004
rect 13722 3992 13728 4004
rect 13044 3964 13728 3992
rect 13044 3952 13050 3964
rect 13722 3952 13728 3964
rect 13780 3992 13786 4004
rect 13924 3992 13952 4023
rect 13780 3964 13952 3992
rect 13780 3952 13786 3964
rect 13262 3924 13268 3936
rect 9968 3896 13268 3924
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 13354 3884 13360 3936
rect 13412 3884 13418 3936
rect 13446 3884 13452 3936
rect 13504 3924 13510 3936
rect 14568 3924 14596 4032
rect 17218 4020 17224 4032
rect 17276 4020 17282 4072
rect 14921 3995 14979 4001
rect 14921 3961 14933 3995
rect 14967 3992 14979 3995
rect 18598 3992 18604 4004
rect 14967 3964 18604 3992
rect 14967 3961 14979 3964
rect 14921 3955 14979 3961
rect 18598 3952 18604 3964
rect 18656 3952 18662 4004
rect 18708 4001 18736 4100
rect 19150 4088 19156 4140
rect 19208 4128 19214 4140
rect 20073 4131 20131 4137
rect 20073 4128 20085 4131
rect 19208 4100 20085 4128
rect 19208 4088 19214 4100
rect 20073 4097 20085 4100
rect 20119 4097 20131 4131
rect 20073 4091 20131 4097
rect 19242 4020 19248 4072
rect 19300 4020 19306 4072
rect 19334 4020 19340 4072
rect 19392 4060 19398 4072
rect 19886 4060 19892 4072
rect 19392 4032 19892 4060
rect 19392 4020 19398 4032
rect 19886 4020 19892 4032
rect 19944 4020 19950 4072
rect 19981 4063 20039 4069
rect 19981 4029 19993 4063
rect 20027 4060 20039 4063
rect 20456 4060 20484 4168
rect 20809 4131 20867 4137
rect 20809 4128 20821 4131
rect 20027 4032 20484 4060
rect 20548 4100 20821 4128
rect 20027 4029 20039 4032
rect 19981 4023 20039 4029
rect 20548 4001 20576 4100
rect 20809 4097 20821 4100
rect 20855 4097 20867 4131
rect 20809 4091 20867 4097
rect 18693 3995 18751 4001
rect 18693 3961 18705 3995
rect 18739 3961 18751 3995
rect 18693 3955 18751 3961
rect 20533 3995 20591 4001
rect 20533 3961 20545 3995
rect 20579 3961 20591 3995
rect 20533 3955 20591 3961
rect 20622 3952 20628 4004
rect 20680 3952 20686 4004
rect 21836 4001 21864 4168
rect 22554 4088 22560 4140
rect 22612 4088 22618 4140
rect 23658 4088 23664 4140
rect 23716 4088 23722 4140
rect 24857 4131 24915 4137
rect 24857 4097 24869 4131
rect 24903 4128 24915 4131
rect 24964 4128 24992 4227
rect 25406 4224 25412 4276
rect 25464 4264 25470 4276
rect 25866 4264 25872 4276
rect 25464 4236 25872 4264
rect 25464 4224 25470 4236
rect 25866 4224 25872 4236
rect 25924 4224 25930 4276
rect 26050 4224 26056 4276
rect 26108 4264 26114 4276
rect 28994 4264 29000 4276
rect 26108 4236 29000 4264
rect 26108 4224 26114 4236
rect 28994 4224 29000 4236
rect 29052 4224 29058 4276
rect 30837 4267 30895 4273
rect 30837 4233 30849 4267
rect 30883 4264 30895 4267
rect 31202 4264 31208 4276
rect 30883 4236 31208 4264
rect 30883 4233 30895 4236
rect 30837 4227 30895 4233
rect 31202 4224 31208 4236
rect 31260 4224 31266 4276
rect 31941 4267 31999 4273
rect 31941 4233 31953 4267
rect 31987 4264 31999 4267
rect 32858 4264 32864 4276
rect 31987 4236 32864 4264
rect 31987 4233 31999 4236
rect 31941 4227 31999 4233
rect 32858 4224 32864 4236
rect 32916 4224 32922 4276
rect 33686 4264 33692 4276
rect 33428 4236 33692 4264
rect 25038 4156 25044 4208
rect 25096 4196 25102 4208
rect 25317 4199 25375 4205
rect 25317 4196 25329 4199
rect 25096 4168 25329 4196
rect 25096 4156 25102 4168
rect 25317 4165 25329 4168
rect 25363 4196 25375 4199
rect 27890 4196 27896 4208
rect 25363 4168 27896 4196
rect 25363 4165 25375 4168
rect 25317 4159 25375 4165
rect 27890 4156 27896 4168
rect 27948 4156 27954 4208
rect 30374 4156 30380 4208
rect 30432 4156 30438 4208
rect 30469 4199 30527 4205
rect 30469 4165 30481 4199
rect 30515 4196 30527 4199
rect 31754 4196 31760 4208
rect 30515 4168 31760 4196
rect 30515 4165 30527 4168
rect 30469 4159 30527 4165
rect 31754 4156 31760 4168
rect 31812 4196 31818 4208
rect 32214 4196 32220 4208
rect 31812 4168 32220 4196
rect 31812 4156 31818 4168
rect 32214 4156 32220 4168
rect 32272 4156 32278 4208
rect 26234 4128 26240 4140
rect 24903 4100 24992 4128
rect 25516 4100 26240 4128
rect 24903 4097 24915 4100
rect 24857 4091 24915 4097
rect 22830 4020 22836 4072
rect 22888 4020 22894 4072
rect 23937 4063 23995 4069
rect 23937 4029 23949 4063
rect 23983 4060 23995 4063
rect 25516 4060 25544 4100
rect 26234 4088 26240 4100
rect 26292 4088 26298 4140
rect 27430 4088 27436 4140
rect 27488 4128 27494 4140
rect 27709 4131 27767 4137
rect 27709 4128 27721 4131
rect 27488 4100 27721 4128
rect 27488 4088 27494 4100
rect 27709 4097 27721 4100
rect 27755 4128 27767 4131
rect 28166 4128 28172 4140
rect 27755 4100 28172 4128
rect 27755 4097 27767 4100
rect 27709 4091 27767 4097
rect 28166 4088 28172 4100
rect 28224 4088 28230 4140
rect 30558 4128 30564 4140
rect 30392 4100 30564 4128
rect 23983 4032 25544 4060
rect 23983 4029 23995 4032
rect 23937 4023 23995 4029
rect 25590 4020 25596 4072
rect 25648 4020 25654 4072
rect 27985 4063 28043 4069
rect 27985 4029 27997 4063
rect 28031 4029 28043 4063
rect 27985 4023 28043 4029
rect 30285 4063 30343 4069
rect 30285 4029 30297 4063
rect 30331 4060 30343 4063
rect 30392 4060 30420 4100
rect 30558 4088 30564 4100
rect 30616 4088 30622 4140
rect 31205 4132 31263 4137
rect 31205 4131 31340 4132
rect 31205 4128 31217 4131
rect 30668 4100 31217 4128
rect 30331 4032 30420 4060
rect 30331 4029 30343 4032
rect 30285 4023 30343 4029
rect 21821 3995 21879 4001
rect 21821 3961 21833 3995
rect 21867 3961 21879 3995
rect 21821 3955 21879 3961
rect 26326 3952 26332 4004
rect 26384 3992 26390 4004
rect 26384 3964 27384 3992
rect 26384 3952 26390 3964
rect 13504 3896 14596 3924
rect 15841 3927 15899 3933
rect 13504 3884 13510 3896
rect 15841 3893 15853 3927
rect 15887 3924 15899 3927
rect 16390 3924 16396 3936
rect 15887 3896 16396 3924
rect 15887 3893 15899 3896
rect 15841 3887 15899 3893
rect 16390 3884 16396 3896
rect 16448 3884 16454 3936
rect 16574 3884 16580 3936
rect 16632 3924 16638 3936
rect 18417 3927 18475 3933
rect 18417 3924 18429 3927
rect 16632 3896 18429 3924
rect 16632 3884 16638 3896
rect 18417 3893 18429 3896
rect 18463 3893 18475 3927
rect 18417 3887 18475 3893
rect 19058 3884 19064 3936
rect 19116 3924 19122 3936
rect 22186 3924 22192 3936
rect 19116 3896 22192 3924
rect 19116 3884 19122 3896
rect 22186 3884 22192 3896
rect 22244 3884 22250 3936
rect 24670 3884 24676 3936
rect 24728 3884 24734 3936
rect 26602 3884 26608 3936
rect 26660 3924 26666 3936
rect 26973 3927 27031 3933
rect 26973 3924 26985 3927
rect 26660 3896 26985 3924
rect 26660 3884 26666 3896
rect 26973 3893 26985 3896
rect 27019 3893 27031 3927
rect 27356 3924 27384 3964
rect 28000 3924 28028 4023
rect 30466 4020 30472 4072
rect 30524 4060 30530 4072
rect 30668 4060 30696 4100
rect 31205 4097 31217 4100
rect 31251 4128 31340 4131
rect 33428 4128 33456 4236
rect 33686 4224 33692 4236
rect 33744 4264 33750 4276
rect 34054 4264 34060 4276
rect 33744 4236 34060 4264
rect 33744 4224 33750 4236
rect 34054 4224 34060 4236
rect 34112 4224 34118 4276
rect 34793 4267 34851 4273
rect 34793 4233 34805 4267
rect 34839 4264 34851 4267
rect 35618 4264 35624 4276
rect 34839 4236 35624 4264
rect 34839 4233 34851 4236
rect 34793 4227 34851 4233
rect 35618 4224 35624 4236
rect 35676 4224 35682 4276
rect 35897 4267 35955 4273
rect 35897 4233 35909 4267
rect 35943 4264 35955 4267
rect 36446 4264 36452 4276
rect 35943 4236 36452 4264
rect 35943 4233 35955 4236
rect 35897 4227 35955 4233
rect 36446 4224 36452 4236
rect 36504 4224 36510 4276
rect 33980 4168 34192 4196
rect 31251 4104 33456 4128
rect 31251 4097 31263 4104
rect 31312 4100 33456 4104
rect 31205 4091 31263 4097
rect 33502 4088 33508 4140
rect 33560 4128 33566 4140
rect 33980 4128 34008 4168
rect 33560 4100 34008 4128
rect 33560 4088 33566 4100
rect 34054 4088 34060 4140
rect 34112 4088 34118 4140
rect 34164 4128 34192 4168
rect 34330 4156 34336 4208
rect 34388 4196 34394 4208
rect 38470 4196 38476 4208
rect 34388 4168 38476 4196
rect 34388 4156 34394 4168
rect 38470 4156 38476 4168
rect 38528 4156 38534 4208
rect 35161 4131 35219 4137
rect 35161 4128 35173 4131
rect 34164 4100 35173 4128
rect 35161 4097 35173 4100
rect 35207 4097 35219 4131
rect 35161 4091 35219 4097
rect 35250 4088 35256 4140
rect 35308 4128 35314 4140
rect 35308 4100 35480 4128
rect 35308 4088 35314 4100
rect 30524 4032 30696 4060
rect 30929 4063 30987 4069
rect 30524 4020 30530 4032
rect 30929 4029 30941 4063
rect 30975 4029 30987 4063
rect 30929 4023 30987 4029
rect 28074 3952 28080 4004
rect 28132 3992 28138 4004
rect 30944 3992 30972 4023
rect 33410 4020 33416 4072
rect 33468 4060 33474 4072
rect 33781 4063 33839 4069
rect 33781 4060 33793 4063
rect 33468 4032 33793 4060
rect 33468 4020 33474 4032
rect 33781 4029 33793 4032
rect 33827 4029 33839 4063
rect 33781 4023 33839 4029
rect 34422 4020 34428 4072
rect 34480 4060 34486 4072
rect 34885 4063 34943 4069
rect 34885 4060 34897 4063
rect 34480 4032 34897 4060
rect 34480 4020 34486 4032
rect 34885 4029 34897 4032
rect 34931 4029 34943 4063
rect 35452 4060 35480 4100
rect 37550 4088 37556 4140
rect 37608 4088 37614 4140
rect 38841 4131 38899 4137
rect 38841 4097 38853 4131
rect 38887 4097 38899 4131
rect 38841 4091 38899 4097
rect 38856 4060 38884 4091
rect 38930 4088 38936 4140
rect 38988 4128 38994 4140
rect 39209 4131 39267 4137
rect 39209 4128 39221 4131
rect 38988 4100 39221 4128
rect 38988 4088 38994 4100
rect 39209 4097 39221 4100
rect 39255 4097 39267 4131
rect 39209 4091 39267 4097
rect 35452 4032 38884 4060
rect 34885 4023 34943 4029
rect 37737 3995 37795 4001
rect 37737 3992 37749 3995
rect 28132 3964 30972 3992
rect 34716 3964 35020 3992
rect 28132 3952 28138 3964
rect 27356 3896 28028 3924
rect 26973 3887 27031 3893
rect 28902 3884 28908 3936
rect 28960 3924 28966 3936
rect 31202 3924 31208 3936
rect 28960 3896 31208 3924
rect 28960 3884 28966 3896
rect 31202 3884 31208 3896
rect 31260 3884 31266 3936
rect 32766 3884 32772 3936
rect 32824 3924 32830 3936
rect 33318 3924 33324 3936
rect 32824 3896 33324 3924
rect 32824 3884 32830 3896
rect 33318 3884 33324 3896
rect 33376 3884 33382 3936
rect 33686 3884 33692 3936
rect 33744 3884 33750 3936
rect 33870 3884 33876 3936
rect 33928 3924 33934 3936
rect 34716 3924 34744 3964
rect 33928 3896 34744 3924
rect 34992 3924 35020 3964
rect 35636 3964 37749 3992
rect 35636 3924 35664 3964
rect 37737 3961 37749 3964
rect 37783 3961 37795 3995
rect 37737 3955 37795 3961
rect 39393 3995 39451 4001
rect 39393 3961 39405 3995
rect 39439 3992 39451 3995
rect 39482 3992 39488 4004
rect 39439 3964 39488 3992
rect 39439 3961 39451 3964
rect 39393 3955 39451 3961
rect 39482 3952 39488 3964
rect 39540 3952 39546 4004
rect 34992 3896 35664 3924
rect 33928 3884 33934 3896
rect 39022 3884 39028 3936
rect 39080 3884 39086 3936
rect 1104 3834 39836 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 37950 3834
rect 38002 3782 38014 3834
rect 38066 3782 38078 3834
rect 38130 3782 38142 3834
rect 38194 3782 38206 3834
rect 38258 3782 39836 3834
rect 1104 3760 39836 3782
rect 2498 3680 2504 3732
rect 2556 3720 2562 3732
rect 2869 3723 2927 3729
rect 2869 3720 2881 3723
rect 2556 3692 2881 3720
rect 2556 3680 2562 3692
rect 2869 3689 2881 3692
rect 2915 3689 2927 3723
rect 5626 3720 5632 3732
rect 2869 3683 2927 3689
rect 4908 3692 5632 3720
rect 2777 3655 2835 3661
rect 2777 3621 2789 3655
rect 2823 3652 2835 3655
rect 4908 3652 4936 3692
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 6546 3680 6552 3732
rect 6604 3720 6610 3732
rect 9490 3720 9496 3732
rect 6604 3692 9496 3720
rect 6604 3680 6610 3692
rect 9490 3680 9496 3692
rect 9548 3720 9554 3732
rect 10962 3720 10968 3732
rect 9548 3692 10968 3720
rect 9548 3680 9554 3692
rect 2823 3624 4936 3652
rect 8205 3655 8263 3661
rect 2823 3621 2835 3624
rect 2777 3615 2835 3621
rect 8205 3621 8217 3655
rect 8251 3652 8263 3655
rect 9585 3655 9643 3661
rect 9585 3652 9597 3655
rect 8251 3624 9597 3652
rect 8251 3621 8263 3624
rect 8205 3615 8263 3621
rect 9585 3621 9597 3624
rect 9631 3621 9643 3655
rect 9585 3615 9643 3621
rect 1673 3587 1731 3593
rect 1673 3553 1685 3587
rect 1719 3584 1731 3587
rect 2866 3584 2872 3596
rect 1719 3556 2872 3584
rect 1719 3553 1731 3556
rect 1673 3547 1731 3553
rect 2866 3544 2872 3556
rect 2924 3544 2930 3596
rect 3142 3544 3148 3596
rect 3200 3584 3206 3596
rect 3329 3587 3387 3593
rect 3329 3584 3341 3587
rect 3200 3556 3341 3584
rect 3200 3544 3206 3556
rect 3329 3553 3341 3556
rect 3375 3553 3387 3587
rect 3329 3547 3387 3553
rect 3418 3544 3424 3596
rect 3476 3544 3482 3596
rect 5902 3544 5908 3596
rect 5960 3544 5966 3596
rect 6730 3544 6736 3596
rect 6788 3544 6794 3596
rect 7190 3544 7196 3596
rect 7248 3544 7254 3596
rect 8754 3544 8760 3596
rect 8812 3584 8818 3596
rect 8941 3587 8999 3593
rect 8941 3584 8953 3587
rect 8812 3556 8953 3584
rect 8812 3544 8818 3556
rect 8941 3553 8953 3556
rect 8987 3553 8999 3587
rect 8941 3547 8999 3553
rect 9125 3587 9183 3593
rect 9125 3553 9137 3587
rect 9171 3584 9183 3587
rect 9692 3584 9720 3692
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 12529 3723 12587 3729
rect 12529 3720 12541 3723
rect 11072 3692 12541 3720
rect 9171 3556 9720 3584
rect 9171 3553 9183 3556
rect 9125 3547 9183 3553
rect 9858 3544 9864 3596
rect 9916 3544 9922 3596
rect 10134 3544 10140 3596
rect 10192 3544 10198 3596
rect 10318 3544 10324 3596
rect 10376 3584 10382 3596
rect 11072 3593 11100 3692
rect 12529 3689 12541 3692
rect 12575 3689 12587 3723
rect 12529 3683 12587 3689
rect 13538 3680 13544 3732
rect 13596 3720 13602 3732
rect 17221 3723 17279 3729
rect 17221 3720 17233 3723
rect 13596 3692 17233 3720
rect 13596 3680 13602 3692
rect 17221 3689 17233 3692
rect 17267 3689 17279 3723
rect 17221 3683 17279 3689
rect 17770 3680 17776 3732
rect 17828 3720 17834 3732
rect 20165 3723 20223 3729
rect 20165 3720 20177 3723
rect 17828 3692 20177 3720
rect 17828 3680 17834 3692
rect 20165 3689 20177 3692
rect 20211 3689 20223 3723
rect 20165 3683 20223 3689
rect 20254 3680 20260 3732
rect 20312 3720 20318 3732
rect 22830 3720 22836 3732
rect 20312 3692 22836 3720
rect 20312 3680 20318 3692
rect 22830 3680 22836 3692
rect 22888 3720 22894 3732
rect 26326 3720 26332 3732
rect 22888 3692 26332 3720
rect 22888 3680 22894 3692
rect 11514 3612 11520 3664
rect 11572 3652 11578 3664
rect 11701 3655 11759 3661
rect 11701 3652 11713 3655
rect 11572 3624 11713 3652
rect 11572 3612 11578 3624
rect 11701 3621 11713 3624
rect 11747 3621 11759 3655
rect 11701 3615 11759 3621
rect 12161 3655 12219 3661
rect 12161 3621 12173 3655
rect 12207 3652 12219 3655
rect 12802 3652 12808 3664
rect 12207 3624 12808 3652
rect 12207 3621 12219 3624
rect 12161 3615 12219 3621
rect 12802 3612 12808 3624
rect 12860 3612 12866 3664
rect 14550 3612 14556 3664
rect 14608 3652 14614 3664
rect 15197 3655 15255 3661
rect 15197 3652 15209 3655
rect 14608 3624 15209 3652
rect 14608 3612 14614 3624
rect 15197 3621 15209 3624
rect 15243 3621 15255 3655
rect 15197 3615 15255 3621
rect 18138 3612 18144 3664
rect 18196 3652 18202 3664
rect 20622 3652 20628 3664
rect 18196 3624 20628 3652
rect 18196 3612 18202 3624
rect 20622 3612 20628 3624
rect 20680 3612 20686 3664
rect 22186 3612 22192 3664
rect 22244 3652 22250 3664
rect 23014 3652 23020 3664
rect 22244 3624 23020 3652
rect 22244 3612 22250 3624
rect 23014 3612 23020 3624
rect 23072 3612 23078 3664
rect 11057 3587 11115 3593
rect 10376 3556 10732 3584
rect 10376 3544 10382 3556
rect 198 3476 204 3528
rect 256 3516 262 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 256 3488 1409 3516
rect 256 3476 262 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 2314 3476 2320 3528
rect 2372 3476 2378 3528
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3485 2651 3519
rect 2593 3479 2651 3485
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 4430 3516 4436 3528
rect 3283 3488 4436 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 1302 3408 1308 3460
rect 1360 3448 1366 3460
rect 2608 3448 2636 3479
rect 4430 3476 4436 3488
rect 4488 3476 4494 3528
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3516 5043 3519
rect 5031 3488 5580 3516
rect 5031 3485 5043 3488
rect 4985 3479 5043 3485
rect 1360 3420 2636 3448
rect 1360 3408 1366 3420
rect 2498 3340 2504 3392
rect 2556 3340 2562 3392
rect 3329 3383 3387 3389
rect 3329 3349 3341 3383
rect 3375 3380 3387 3383
rect 4338 3380 4344 3392
rect 3375 3352 4344 3380
rect 3375 3349 3387 3352
rect 3329 3343 3387 3349
rect 4338 3340 4344 3352
rect 4396 3340 4402 3392
rect 5166 3340 5172 3392
rect 5224 3340 5230 3392
rect 5350 3340 5356 3392
rect 5408 3340 5414 3392
rect 5552 3380 5580 3488
rect 5718 3476 5724 3528
rect 5776 3476 5782 3528
rect 6549 3519 6607 3525
rect 6549 3485 6561 3519
rect 6595 3516 6607 3519
rect 6914 3516 6920 3528
rect 6595 3488 6920 3516
rect 6595 3485 6607 3488
rect 6549 3479 6607 3485
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 7469 3519 7527 3525
rect 7469 3485 7481 3519
rect 7515 3516 7527 3519
rect 7558 3516 7564 3528
rect 7515 3488 7564 3516
rect 7515 3485 7527 3488
rect 7469 3479 7527 3485
rect 7558 3476 7564 3488
rect 7616 3476 7622 3528
rect 10042 3525 10048 3528
rect 9999 3519 10048 3525
rect 9999 3485 10011 3519
rect 10045 3485 10048 3519
rect 9999 3479 10048 3485
rect 10042 3476 10048 3479
rect 10100 3476 10106 3528
rect 10704 3516 10732 3556
rect 11057 3553 11069 3587
rect 11103 3553 11115 3587
rect 11057 3547 11115 3553
rect 11256 3556 12434 3584
rect 11256 3525 11284 3556
rect 11149 3519 11207 3525
rect 11149 3516 11161 3519
rect 10704 3488 11161 3516
rect 11149 3485 11161 3488
rect 11195 3485 11207 3519
rect 11149 3479 11207 3485
rect 11241 3519 11299 3525
rect 11241 3485 11253 3519
rect 11287 3485 11299 3519
rect 11241 3479 11299 3485
rect 5813 3451 5871 3457
rect 5813 3417 5825 3451
rect 5859 3448 5871 3451
rect 11256 3448 11284 3479
rect 11882 3476 11888 3528
rect 11940 3476 11946 3528
rect 11977 3519 12035 3525
rect 11977 3485 11989 3519
rect 12023 3485 12035 3519
rect 11977 3479 12035 3485
rect 11992 3448 12020 3479
rect 5859 3420 6684 3448
rect 5859 3417 5871 3420
rect 5813 3411 5871 3417
rect 6656 3389 6684 3420
rect 10612 3420 11284 3448
rect 11624 3420 12020 3448
rect 12406 3448 12434 3556
rect 13538 3544 13544 3596
rect 13596 3584 13602 3596
rect 13722 3584 13728 3596
rect 13596 3556 13728 3584
rect 13596 3544 13602 3556
rect 13722 3544 13728 3556
rect 13780 3584 13786 3596
rect 17129 3587 17187 3593
rect 13780 3556 16620 3584
rect 13780 3544 13786 3556
rect 16592 3528 16620 3556
rect 17129 3553 17141 3587
rect 17175 3584 17187 3587
rect 17218 3584 17224 3596
rect 17175 3556 17224 3584
rect 17175 3553 17187 3556
rect 17129 3547 17187 3553
rect 17218 3544 17224 3556
rect 17276 3584 17282 3596
rect 18230 3584 18236 3596
rect 17276 3556 18236 3584
rect 17276 3544 17282 3556
rect 18230 3544 18236 3556
rect 18288 3544 18294 3596
rect 18598 3544 18604 3596
rect 18656 3584 18662 3596
rect 19429 3587 19487 3593
rect 19429 3584 19441 3587
rect 18656 3556 19441 3584
rect 18656 3544 18662 3556
rect 19429 3553 19441 3556
rect 19475 3553 19487 3587
rect 22830 3584 22836 3596
rect 19429 3547 19487 3553
rect 19628 3556 22836 3584
rect 13170 3476 13176 3528
rect 13228 3516 13234 3528
rect 13265 3519 13323 3525
rect 13265 3516 13277 3519
rect 13228 3488 13277 3516
rect 13228 3476 13234 3488
rect 13265 3485 13277 3488
rect 13311 3485 13323 3519
rect 13265 3479 13323 3485
rect 15378 3476 15384 3528
rect 15436 3476 15442 3528
rect 16574 3476 16580 3528
rect 16632 3476 16638 3528
rect 16853 3519 16911 3525
rect 16853 3485 16865 3519
rect 16899 3516 16911 3519
rect 16942 3516 16948 3528
rect 16899 3488 16948 3516
rect 16899 3485 16911 3488
rect 16853 3479 16911 3485
rect 16942 3476 16948 3488
rect 17000 3476 17006 3528
rect 17402 3476 17408 3528
rect 17460 3476 17466 3528
rect 17770 3476 17776 3528
rect 17828 3476 17834 3528
rect 17862 3476 17868 3528
rect 17920 3516 17926 3528
rect 19628 3516 19656 3556
rect 22830 3544 22836 3556
rect 22888 3544 22894 3596
rect 23768 3593 23796 3692
rect 26326 3680 26332 3692
rect 26384 3680 26390 3732
rect 26973 3723 27031 3729
rect 26973 3689 26985 3723
rect 27019 3720 27031 3723
rect 27019 3692 31524 3720
rect 27019 3689 27031 3692
rect 26973 3683 27031 3689
rect 28258 3612 28264 3664
rect 28316 3652 28322 3664
rect 29181 3655 29239 3661
rect 29181 3652 29193 3655
rect 28316 3624 29193 3652
rect 28316 3612 28322 3624
rect 29181 3621 29193 3624
rect 29227 3652 29239 3655
rect 30466 3652 30472 3664
rect 29227 3624 30472 3652
rect 29227 3621 29239 3624
rect 29181 3615 29239 3621
rect 30466 3612 30472 3624
rect 30524 3612 30530 3664
rect 31496 3661 31524 3692
rect 31662 3680 31668 3732
rect 31720 3720 31726 3732
rect 33318 3720 33324 3732
rect 31720 3692 33324 3720
rect 31720 3680 31726 3692
rect 33318 3680 33324 3692
rect 33376 3680 33382 3732
rect 33410 3680 33416 3732
rect 33468 3720 33474 3732
rect 34422 3720 34428 3732
rect 33468 3692 34428 3720
rect 33468 3680 33474 3692
rect 34422 3680 34428 3692
rect 34480 3680 34486 3732
rect 34514 3680 34520 3732
rect 34572 3720 34578 3732
rect 34701 3723 34759 3729
rect 34701 3720 34713 3723
rect 34572 3692 34713 3720
rect 34572 3680 34578 3692
rect 34701 3689 34713 3692
rect 34747 3689 34759 3723
rect 34701 3683 34759 3689
rect 35986 3680 35992 3732
rect 36044 3680 36050 3732
rect 39390 3680 39396 3732
rect 39448 3680 39454 3732
rect 31481 3655 31539 3661
rect 31481 3621 31493 3655
rect 31527 3621 31539 3655
rect 31481 3615 31539 3621
rect 32030 3612 32036 3664
rect 32088 3652 32094 3664
rect 38930 3652 38936 3664
rect 32088 3624 38936 3652
rect 32088 3612 32094 3624
rect 38930 3612 38936 3624
rect 38988 3612 38994 3664
rect 39025 3655 39083 3661
rect 39025 3621 39037 3655
rect 39071 3652 39083 3655
rect 39942 3652 39948 3664
rect 39071 3624 39948 3652
rect 39071 3621 39083 3624
rect 39025 3615 39083 3621
rect 39942 3612 39948 3624
rect 40000 3612 40006 3664
rect 23753 3587 23811 3593
rect 23753 3553 23765 3587
rect 23799 3553 23811 3587
rect 23753 3547 23811 3553
rect 29822 3544 29828 3596
rect 29880 3584 29886 3596
rect 30742 3584 30748 3596
rect 29880 3556 30748 3584
rect 29880 3544 29886 3556
rect 30742 3544 30748 3556
rect 30800 3584 30806 3596
rect 31067 3587 31125 3593
rect 31067 3584 31079 3587
rect 30800 3556 31079 3584
rect 30800 3544 30806 3556
rect 31067 3553 31079 3556
rect 31113 3553 31125 3587
rect 31067 3547 31125 3553
rect 31846 3544 31852 3596
rect 31904 3584 31910 3596
rect 31941 3587 31999 3593
rect 31941 3584 31953 3587
rect 31904 3556 31953 3584
rect 31904 3544 31910 3556
rect 31941 3553 31953 3556
rect 31987 3553 31999 3587
rect 31941 3547 31999 3553
rect 33686 3544 33692 3596
rect 33744 3584 33750 3596
rect 38654 3584 38660 3596
rect 33744 3556 38660 3584
rect 33744 3544 33750 3556
rect 38654 3544 38660 3556
rect 38712 3544 38718 3596
rect 17920 3488 19656 3516
rect 17920 3476 17926 3488
rect 19702 3476 19708 3528
rect 19760 3476 19766 3528
rect 20349 3519 20407 3525
rect 20349 3485 20361 3519
rect 20395 3512 20407 3519
rect 22097 3519 22155 3525
rect 20395 3485 20417 3512
rect 20349 3479 20417 3485
rect 22097 3485 22109 3519
rect 22143 3516 22155 3519
rect 22554 3516 22560 3528
rect 22143 3488 22560 3516
rect 22143 3485 22155 3488
rect 22097 3479 22155 3485
rect 19288 3448 19294 3460
rect 12406 3420 19294 3448
rect 10612 3392 10640 3420
rect 6181 3383 6239 3389
rect 6181 3380 6193 3383
rect 5552 3352 6193 3380
rect 6181 3349 6193 3352
rect 6227 3349 6239 3383
rect 6181 3343 6239 3349
rect 6641 3383 6699 3389
rect 6641 3349 6653 3383
rect 6687 3380 6699 3383
rect 9674 3380 9680 3392
rect 6687 3352 9680 3380
rect 6687 3349 6699 3352
rect 6641 3343 6699 3349
rect 9674 3340 9680 3352
rect 9732 3380 9738 3392
rect 10226 3380 10232 3392
rect 9732 3352 10232 3380
rect 9732 3340 9738 3352
rect 10226 3340 10232 3352
rect 10284 3340 10290 3392
rect 10594 3340 10600 3392
rect 10652 3340 10658 3392
rect 10781 3383 10839 3389
rect 10781 3349 10793 3383
rect 10827 3380 10839 3383
rect 10962 3380 10968 3392
rect 10827 3352 10968 3380
rect 10827 3349 10839 3352
rect 10781 3343 10839 3349
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 11149 3383 11207 3389
rect 11149 3349 11161 3383
rect 11195 3380 11207 3383
rect 11422 3380 11428 3392
rect 11195 3352 11428 3380
rect 11195 3349 11207 3352
rect 11149 3343 11207 3349
rect 11422 3340 11428 3352
rect 11480 3340 11486 3392
rect 11624 3389 11652 3420
rect 19288 3408 19294 3420
rect 19346 3408 19352 3460
rect 20389 3448 20417 3479
rect 22554 3476 22560 3488
rect 22612 3476 22618 3528
rect 23477 3519 23535 3525
rect 23477 3485 23489 3519
rect 23523 3516 23535 3519
rect 23566 3516 23572 3528
rect 23523 3488 23572 3516
rect 23523 3485 23535 3488
rect 23477 3479 23535 3485
rect 23566 3476 23572 3488
rect 23624 3476 23630 3528
rect 25961 3519 26019 3525
rect 25961 3516 25973 3519
rect 23676 3488 25973 3516
rect 20088 3420 20417 3448
rect 11609 3383 11667 3389
rect 11609 3349 11621 3383
rect 11655 3349 11667 3383
rect 11609 3343 11667 3349
rect 11698 3340 11704 3392
rect 11756 3380 11762 3392
rect 15746 3380 15752 3392
rect 11756 3352 15752 3380
rect 11756 3340 11762 3352
rect 15746 3340 15752 3352
rect 15804 3340 15810 3392
rect 16114 3340 16120 3392
rect 16172 3340 16178 3392
rect 16482 3340 16488 3392
rect 16540 3380 16546 3392
rect 17589 3383 17647 3389
rect 17589 3380 17601 3383
rect 16540 3352 17601 3380
rect 16540 3340 16546 3352
rect 17589 3349 17601 3352
rect 17635 3349 17647 3383
rect 17589 3343 17647 3349
rect 19150 3340 19156 3392
rect 19208 3380 19214 3392
rect 20088 3389 20116 3420
rect 20622 3408 20628 3460
rect 20680 3448 20686 3460
rect 22186 3448 22192 3460
rect 20680 3420 22192 3448
rect 20680 3408 20686 3420
rect 22186 3408 22192 3420
rect 22244 3408 22250 3460
rect 22370 3408 22376 3460
rect 22428 3448 22434 3460
rect 23676 3448 23704 3488
rect 25961 3485 25973 3488
rect 26007 3516 26019 3519
rect 26142 3516 26148 3528
rect 26007 3488 26148 3516
rect 26007 3485 26019 3488
rect 25961 3479 26019 3485
rect 26142 3476 26148 3488
rect 26200 3476 26206 3528
rect 26237 3519 26295 3525
rect 26237 3485 26249 3519
rect 26283 3485 26295 3519
rect 26237 3479 26295 3485
rect 22428 3420 23704 3448
rect 22428 3408 22434 3420
rect 25866 3408 25872 3460
rect 25924 3448 25930 3460
rect 26252 3448 26280 3479
rect 26326 3476 26332 3528
rect 26384 3516 26390 3528
rect 27249 3519 27307 3525
rect 27249 3516 27261 3519
rect 26384 3488 27261 3516
rect 26384 3476 26390 3488
rect 27249 3485 27261 3488
rect 27295 3485 27307 3519
rect 27249 3479 27307 3485
rect 27430 3476 27436 3528
rect 27488 3516 27494 3528
rect 27525 3519 27583 3525
rect 27525 3516 27537 3519
rect 27488 3488 27537 3516
rect 27488 3476 27494 3488
rect 27525 3485 27537 3488
rect 27571 3485 27583 3519
rect 27525 3479 27583 3485
rect 27614 3476 27620 3528
rect 27672 3516 27678 3528
rect 30282 3516 30288 3528
rect 27672 3488 30288 3516
rect 27672 3476 27678 3488
rect 30282 3476 30288 3488
rect 30340 3476 30346 3528
rect 30926 3476 30932 3528
rect 30984 3476 30990 3528
rect 31202 3476 31208 3528
rect 31260 3476 31266 3528
rect 31754 3476 31760 3528
rect 31812 3516 31818 3528
rect 32125 3519 32183 3525
rect 32125 3516 32137 3519
rect 31812 3488 32137 3516
rect 31812 3476 31818 3488
rect 32125 3485 32137 3488
rect 32171 3485 32183 3519
rect 32125 3479 32183 3485
rect 33318 3476 33324 3528
rect 33376 3516 33382 3528
rect 34698 3516 34704 3528
rect 33376 3488 34704 3516
rect 33376 3476 33382 3488
rect 34698 3476 34704 3488
rect 34756 3516 34762 3528
rect 34885 3519 34943 3525
rect 34885 3516 34897 3519
rect 34756 3488 34897 3516
rect 34756 3476 34762 3488
rect 34885 3485 34897 3488
rect 34931 3485 34943 3519
rect 34885 3479 34943 3485
rect 34974 3476 34980 3528
rect 35032 3476 35038 3528
rect 36173 3519 36231 3525
rect 36173 3485 36185 3519
rect 36219 3485 36231 3519
rect 36173 3479 36231 3485
rect 25924 3420 26280 3448
rect 25924 3408 25930 3420
rect 28994 3408 29000 3460
rect 29052 3408 29058 3460
rect 29270 3408 29276 3460
rect 29328 3448 29334 3460
rect 29328 3420 30420 3448
rect 29328 3408 29334 3420
rect 19613 3383 19671 3389
rect 19613 3380 19625 3383
rect 19208 3352 19625 3380
rect 19208 3340 19214 3352
rect 19613 3349 19625 3352
rect 19659 3349 19671 3383
rect 19613 3343 19671 3349
rect 20073 3383 20131 3389
rect 20073 3349 20085 3383
rect 20119 3349 20131 3383
rect 20073 3343 20131 3349
rect 22281 3383 22339 3389
rect 22281 3349 22293 3383
rect 22327 3380 22339 3383
rect 22646 3380 22652 3392
rect 22327 3352 22652 3380
rect 22327 3349 22339 3352
rect 22281 3343 22339 3349
rect 22646 3340 22652 3352
rect 22704 3340 22710 3392
rect 22738 3340 22744 3392
rect 22796 3340 22802 3392
rect 23014 3340 23020 3392
rect 23072 3380 23078 3392
rect 27338 3380 27344 3392
rect 23072 3352 27344 3380
rect 23072 3340 23078 3352
rect 27338 3340 27344 3352
rect 27396 3340 27402 3392
rect 28258 3340 28264 3392
rect 28316 3340 28322 3392
rect 29178 3340 29184 3392
rect 29236 3380 29242 3392
rect 30285 3383 30343 3389
rect 30285 3380 30297 3383
rect 29236 3352 30297 3380
rect 29236 3340 29242 3352
rect 30285 3349 30297 3352
rect 30331 3349 30343 3383
rect 30392 3380 30420 3420
rect 33686 3408 33692 3460
rect 33744 3448 33750 3460
rect 36188 3448 36216 3479
rect 38838 3476 38844 3528
rect 38896 3476 38902 3528
rect 39209 3519 39267 3525
rect 39209 3485 39221 3519
rect 39255 3485 39267 3519
rect 39209 3479 39267 3485
rect 33744 3420 36216 3448
rect 33744 3408 33750 3420
rect 36262 3408 36268 3460
rect 36320 3448 36326 3460
rect 39224 3448 39252 3479
rect 36320 3420 39252 3448
rect 36320 3408 36326 3420
rect 33410 3380 33416 3392
rect 30392 3352 33416 3380
rect 30285 3343 30343 3349
rect 33410 3340 33416 3352
rect 33468 3340 33474 3392
rect 33870 3340 33876 3392
rect 33928 3380 33934 3392
rect 34146 3380 34152 3392
rect 33928 3352 34152 3380
rect 33928 3340 33934 3352
rect 34146 3340 34152 3352
rect 34204 3380 34210 3392
rect 34974 3380 34980 3392
rect 34204 3352 34980 3380
rect 34204 3340 34210 3352
rect 34974 3340 34980 3352
rect 35032 3340 35038 3392
rect 35161 3383 35219 3389
rect 35161 3349 35173 3383
rect 35207 3380 35219 3383
rect 38378 3380 38384 3392
rect 35207 3352 38384 3380
rect 35207 3349 35219 3352
rect 35161 3343 35219 3349
rect 38378 3340 38384 3352
rect 38436 3340 38442 3392
rect 1104 3290 39836 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 39010 3290
rect 39062 3238 39074 3290
rect 39126 3238 39138 3290
rect 39190 3238 39202 3290
rect 39254 3238 39266 3290
rect 39318 3238 39836 3290
rect 1104 3216 39836 3238
rect 3697 3179 3755 3185
rect 3697 3145 3709 3179
rect 3743 3176 3755 3179
rect 3970 3176 3976 3188
rect 3743 3148 3976 3176
rect 3743 3145 3755 3148
rect 3697 3139 3755 3145
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 4338 3136 4344 3188
rect 4396 3136 4402 3188
rect 4801 3179 4859 3185
rect 4801 3145 4813 3179
rect 4847 3176 4859 3179
rect 5905 3179 5963 3185
rect 4847 3148 5856 3176
rect 4847 3145 4859 3148
rect 4801 3139 4859 3145
rect 1854 3068 1860 3120
rect 1912 3108 1918 3120
rect 5350 3108 5356 3120
rect 1912 3080 3832 3108
rect 1912 3068 1918 3080
rect 1210 3000 1216 3052
rect 1268 3040 1274 3052
rect 2409 3043 2467 3049
rect 2409 3040 2421 3043
rect 1268 3012 2421 3040
rect 1268 3000 1274 3012
rect 2409 3009 2421 3012
rect 2455 3009 2467 3043
rect 2409 3003 2467 3009
rect 2774 3000 2780 3052
rect 2832 3040 2838 3052
rect 3804 3049 3832 3080
rect 4632 3080 5356 3108
rect 4632 3049 4660 3080
rect 5350 3068 5356 3080
rect 5408 3068 5414 3120
rect 5828 3108 5856 3148
rect 5905 3145 5917 3179
rect 5951 3176 5963 3179
rect 6730 3176 6736 3188
rect 5951 3148 6736 3176
rect 5951 3145 5963 3148
rect 5905 3139 5963 3145
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 11517 3179 11575 3185
rect 11517 3176 11529 3179
rect 9232 3148 11529 3176
rect 8386 3108 8392 3120
rect 5828 3080 8392 3108
rect 8386 3068 8392 3080
rect 8444 3068 8450 3120
rect 2961 3043 3019 3049
rect 2961 3040 2973 3043
rect 2832 3012 2973 3040
rect 2832 3000 2838 3012
rect 2961 3009 2973 3012
rect 3007 3009 3019 3043
rect 2961 3003 3019 3009
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3009 3571 3043
rect 3513 3003 3571 3009
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3009 3847 3043
rect 3789 3003 3847 3009
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3009 4583 3043
rect 4525 3003 4583 3009
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3009 4675 3043
rect 5074 3040 5080 3052
rect 4617 3003 4675 3009
rect 4908 3012 5080 3040
rect 382 2932 388 2984
rect 440 2972 446 2984
rect 1397 2975 1455 2981
rect 1397 2972 1409 2975
rect 440 2944 1409 2972
rect 440 2932 446 2944
rect 1397 2941 1409 2944
rect 1443 2941 1455 2975
rect 1397 2935 1455 2941
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2972 1731 2975
rect 2682 2972 2688 2984
rect 1719 2944 2688 2972
rect 1719 2941 1731 2944
rect 1673 2935 1731 2941
rect 2682 2932 2688 2944
rect 2740 2932 2746 2984
rect 3142 2932 3148 2984
rect 3200 2932 3206 2984
rect 1118 2864 1124 2916
rect 1176 2904 1182 2916
rect 3252 2904 3280 3003
rect 1176 2876 3280 2904
rect 1176 2864 1182 2876
rect 3418 2864 3424 2916
rect 3476 2864 3482 2916
rect 2498 2796 2504 2848
rect 2556 2796 2562 2848
rect 2590 2796 2596 2848
rect 2648 2836 2654 2848
rect 3528 2836 3556 3003
rect 4540 2972 4568 3003
rect 4908 2984 4936 3012
rect 5074 3000 5080 3012
rect 5132 3000 5138 3052
rect 5169 3043 5227 3049
rect 5169 3009 5181 3043
rect 5215 3040 5227 3043
rect 6086 3040 6092 3052
rect 5215 3012 6092 3040
rect 5215 3009 5227 3012
rect 5169 3003 5227 3009
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 6270 3000 6276 3052
rect 6328 3040 6334 3052
rect 9232 3049 9260 3148
rect 11517 3145 11529 3148
rect 11563 3145 11575 3179
rect 11517 3139 11575 3145
rect 11790 3136 11796 3188
rect 11848 3176 11854 3188
rect 11885 3179 11943 3185
rect 11885 3176 11897 3179
rect 11848 3148 11897 3176
rect 11848 3136 11854 3148
rect 11885 3145 11897 3148
rect 11931 3145 11943 3179
rect 11885 3139 11943 3145
rect 12618 3136 12624 3188
rect 12676 3176 12682 3188
rect 17494 3176 17500 3188
rect 12676 3148 17500 3176
rect 12676 3136 12682 3148
rect 17494 3136 17500 3148
rect 17552 3136 17558 3188
rect 17770 3136 17776 3188
rect 17828 3136 17834 3188
rect 18138 3136 18144 3188
rect 18196 3136 18202 3188
rect 18230 3136 18236 3188
rect 18288 3176 18294 3188
rect 20254 3176 20260 3188
rect 18288 3148 20260 3176
rect 18288 3136 18294 3148
rect 20254 3136 20260 3148
rect 20312 3136 20318 3188
rect 20346 3136 20352 3188
rect 20404 3176 20410 3188
rect 20717 3179 20775 3185
rect 20717 3176 20729 3179
rect 20404 3148 20729 3176
rect 20404 3136 20410 3148
rect 20717 3145 20729 3148
rect 20763 3145 20775 3179
rect 20717 3139 20775 3145
rect 23106 3136 23112 3188
rect 23164 3136 23170 3188
rect 25590 3136 25596 3188
rect 25648 3176 25654 3188
rect 25777 3179 25835 3185
rect 25777 3176 25789 3179
rect 25648 3148 25789 3176
rect 25648 3136 25654 3148
rect 25777 3145 25789 3148
rect 25823 3145 25835 3179
rect 25777 3139 25835 3145
rect 26326 3136 26332 3188
rect 26384 3136 26390 3188
rect 27617 3179 27675 3185
rect 27617 3145 27629 3179
rect 27663 3176 27675 3179
rect 27706 3176 27712 3188
rect 27663 3148 27712 3176
rect 27663 3145 27675 3148
rect 27617 3139 27675 3145
rect 27706 3136 27712 3148
rect 27764 3136 27770 3188
rect 29270 3176 29276 3188
rect 27816 3148 29276 3176
rect 11422 3068 11428 3120
rect 11480 3108 11486 3120
rect 11977 3111 12035 3117
rect 11977 3108 11989 3111
rect 11480 3080 11989 3108
rect 11480 3068 11486 3080
rect 11977 3077 11989 3080
rect 12023 3077 12035 3111
rect 11977 3071 12035 3077
rect 13262 3068 13268 3120
rect 13320 3108 13326 3120
rect 21818 3108 21824 3120
rect 13320 3080 21824 3108
rect 13320 3068 13326 3080
rect 21818 3068 21824 3080
rect 21876 3068 21882 3120
rect 26344 3108 26372 3136
rect 27816 3108 27844 3148
rect 29270 3136 29276 3148
rect 29328 3136 29334 3188
rect 30377 3179 30435 3185
rect 30377 3145 30389 3179
rect 30423 3176 30435 3179
rect 30926 3176 30932 3188
rect 30423 3148 30932 3176
rect 30423 3145 30435 3148
rect 30377 3139 30435 3145
rect 30926 3136 30932 3148
rect 30984 3136 30990 3188
rect 31294 3136 31300 3188
rect 31352 3136 31358 3188
rect 33778 3136 33784 3188
rect 33836 3176 33842 3188
rect 34057 3179 34115 3185
rect 34057 3176 34069 3179
rect 33836 3148 34069 3176
rect 33836 3136 33842 3148
rect 34057 3145 34069 3148
rect 34103 3145 34115 3179
rect 34057 3139 34115 3145
rect 36538 3136 36544 3188
rect 36596 3176 36602 3188
rect 38197 3179 38255 3185
rect 38197 3176 38209 3179
rect 36596 3148 38209 3176
rect 36596 3136 36602 3148
rect 38197 3145 38209 3148
rect 38243 3145 38255 3179
rect 38197 3139 38255 3145
rect 39390 3136 39396 3188
rect 39448 3136 39454 3188
rect 22848 3080 26372 3108
rect 26436 3080 27844 3108
rect 22848 3052 22876 3080
rect 6917 3043 6975 3049
rect 6917 3040 6929 3043
rect 6328 3012 6929 3040
rect 6328 3000 6334 3012
rect 6917 3009 6929 3012
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 9217 3043 9275 3049
rect 9217 3009 9229 3043
rect 9263 3009 9275 3043
rect 9217 3003 9275 3009
rect 9493 3043 9551 3049
rect 9493 3009 9505 3043
rect 9539 3040 9551 3043
rect 9858 3040 9864 3052
rect 9539 3012 9864 3040
rect 9539 3009 9551 3012
rect 9493 3003 9551 3009
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 10594 3049 10600 3052
rect 10551 3043 10600 3049
rect 10551 3009 10563 3043
rect 10597 3009 10600 3043
rect 10551 3003 10600 3009
rect 10594 3000 10600 3003
rect 10652 3000 10658 3052
rect 10686 3000 10692 3052
rect 10744 3000 10750 3052
rect 12894 3000 12900 3052
rect 12952 3040 12958 3052
rect 13173 3043 13231 3049
rect 13173 3040 13185 3043
rect 12952 3012 13185 3040
rect 12952 3000 12958 3012
rect 13173 3009 13185 3012
rect 13219 3040 13231 3043
rect 13633 3043 13691 3049
rect 13633 3040 13645 3043
rect 13219 3012 13645 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 13633 3009 13645 3012
rect 13679 3040 13691 3043
rect 14829 3043 14887 3049
rect 14829 3040 14841 3043
rect 13679 3012 14841 3040
rect 13679 3009 13691 3012
rect 13633 3003 13691 3009
rect 14829 3009 14841 3012
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 15304 3012 15976 3040
rect 4798 2972 4804 2984
rect 4540 2944 4804 2972
rect 4798 2932 4804 2944
rect 4856 2932 4862 2984
rect 4890 2932 4896 2984
rect 4948 2932 4954 2984
rect 6362 2932 6368 2984
rect 6420 2972 6426 2984
rect 6641 2975 6699 2981
rect 6641 2972 6653 2975
rect 6420 2944 6653 2972
rect 6420 2932 6426 2944
rect 6641 2941 6653 2944
rect 6687 2941 6699 2975
rect 6641 2935 6699 2941
rect 9582 2932 9588 2984
rect 9640 2972 9646 2984
rect 9677 2975 9735 2981
rect 9677 2972 9689 2975
rect 9640 2944 9689 2972
rect 9640 2932 9646 2944
rect 9677 2941 9689 2944
rect 9723 2941 9735 2975
rect 9677 2935 9735 2941
rect 10413 2975 10471 2981
rect 10413 2941 10425 2975
rect 10459 2972 10471 2975
rect 11790 2972 11796 2984
rect 10459 2944 11796 2972
rect 10459 2941 10471 2944
rect 10413 2935 10471 2941
rect 11790 2932 11796 2944
rect 11848 2932 11854 2984
rect 12161 2975 12219 2981
rect 12161 2941 12173 2975
rect 12207 2941 12219 2975
rect 12161 2935 12219 2941
rect 13449 2975 13507 2981
rect 13449 2941 13461 2975
rect 13495 2972 13507 2975
rect 13538 2972 13544 2984
rect 13495 2944 13544 2972
rect 13495 2941 13507 2944
rect 13449 2935 13507 2941
rect 7653 2907 7711 2913
rect 7653 2873 7665 2907
rect 7699 2904 7711 2907
rect 10137 2907 10195 2913
rect 10137 2904 10149 2907
rect 7699 2876 10149 2904
rect 7699 2873 7711 2876
rect 7653 2867 7711 2873
rect 10137 2873 10149 2876
rect 10183 2873 10195 2907
rect 12176 2904 12204 2935
rect 13538 2932 13544 2944
rect 13596 2932 13602 2984
rect 14553 2975 14611 2981
rect 14553 2941 14565 2975
rect 14599 2941 14611 2975
rect 14553 2935 14611 2941
rect 12437 2907 12495 2913
rect 12437 2904 12449 2907
rect 10137 2867 10195 2873
rect 11256 2876 11468 2904
rect 12176 2876 12449 2904
rect 2648 2808 3556 2836
rect 3973 2839 4031 2845
rect 2648 2796 2654 2808
rect 3973 2805 3985 2839
rect 4019 2836 4031 2839
rect 4154 2836 4160 2848
rect 4019 2808 4160 2836
rect 4019 2805 4031 2808
rect 3973 2799 4031 2805
rect 4154 2796 4160 2808
rect 4212 2796 4218 2848
rect 4341 2839 4399 2845
rect 4341 2805 4353 2839
rect 4387 2836 4399 2839
rect 4706 2836 4712 2848
rect 4387 2808 4712 2836
rect 4387 2805 4399 2808
rect 4341 2799 4399 2805
rect 4706 2796 4712 2808
rect 4764 2796 4770 2848
rect 6546 2796 6552 2848
rect 6604 2836 6610 2848
rect 7466 2836 7472 2848
rect 6604 2808 7472 2836
rect 6604 2796 6610 2808
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 9401 2839 9459 2845
rect 9401 2805 9413 2839
rect 9447 2836 9459 2839
rect 9766 2836 9772 2848
rect 9447 2808 9772 2836
rect 9447 2805 9459 2808
rect 9401 2799 9459 2805
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 10042 2796 10048 2848
rect 10100 2836 10106 2848
rect 11256 2836 11284 2876
rect 10100 2808 11284 2836
rect 10100 2796 10106 2808
rect 11330 2796 11336 2848
rect 11388 2796 11394 2848
rect 11440 2836 11468 2876
rect 12437 2873 12449 2876
rect 12483 2873 12495 2907
rect 12437 2867 12495 2873
rect 13817 2907 13875 2913
rect 13817 2873 13829 2907
rect 13863 2904 13875 2907
rect 14458 2904 14464 2916
rect 13863 2876 14464 2904
rect 13863 2873 13875 2876
rect 13817 2867 13875 2873
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
rect 13722 2836 13728 2848
rect 11440 2808 13728 2836
rect 13722 2796 13728 2808
rect 13780 2796 13786 2848
rect 14568 2836 14596 2935
rect 15304 2904 15332 3012
rect 15378 2932 15384 2984
rect 15436 2972 15442 2984
rect 15948 2972 15976 3012
rect 16022 3000 16028 3052
rect 16080 3000 16086 3052
rect 16117 3043 16175 3049
rect 16117 3009 16129 3043
rect 16163 3040 16175 3043
rect 16574 3040 16580 3052
rect 16163 3012 16580 3040
rect 16163 3009 16175 3012
rect 16117 3003 16175 3009
rect 16574 3000 16580 3012
rect 16632 3000 16638 3052
rect 16942 3000 16948 3052
rect 17000 3040 17006 3052
rect 17000 3012 18460 3040
rect 17000 3000 17006 3012
rect 16209 2975 16267 2981
rect 16209 2972 16221 2975
rect 15436 2944 15700 2972
rect 15948 2944 16221 2972
rect 15436 2932 15442 2944
rect 15672 2913 15700 2944
rect 16209 2941 16221 2944
rect 16255 2941 16267 2975
rect 16209 2935 16267 2941
rect 16666 2932 16672 2984
rect 16724 2932 16730 2984
rect 17494 2932 17500 2984
rect 17552 2972 17558 2984
rect 18233 2975 18291 2981
rect 18233 2972 18245 2975
rect 17552 2944 18245 2972
rect 17552 2932 17558 2944
rect 18233 2941 18245 2944
rect 18279 2941 18291 2975
rect 18233 2935 18291 2941
rect 18325 2975 18383 2981
rect 18325 2941 18337 2975
rect 18371 2941 18383 2975
rect 18325 2935 18383 2941
rect 15565 2907 15623 2913
rect 15565 2904 15577 2907
rect 15304 2876 15577 2904
rect 15565 2873 15577 2876
rect 15611 2873 15623 2907
rect 15565 2867 15623 2873
rect 15657 2907 15715 2913
rect 15657 2873 15669 2907
rect 15703 2873 15715 2907
rect 15657 2867 15715 2873
rect 14918 2836 14924 2848
rect 14568 2808 14924 2836
rect 14918 2796 14924 2808
rect 14976 2796 14982 2848
rect 16684 2836 16712 2932
rect 17681 2907 17739 2913
rect 17681 2873 17693 2907
rect 17727 2904 17739 2907
rect 18340 2904 18368 2935
rect 17727 2876 18368 2904
rect 18432 2904 18460 3012
rect 19426 3000 19432 3052
rect 19484 3040 19490 3052
rect 19981 3043 20039 3049
rect 19981 3040 19993 3043
rect 19484 3012 19993 3040
rect 19484 3000 19490 3012
rect 19981 3009 19993 3012
rect 20027 3009 20039 3043
rect 19981 3003 20039 3009
rect 22554 3000 22560 3052
rect 22612 3000 22618 3052
rect 22830 3000 22836 3052
rect 22888 3000 22894 3052
rect 22925 3043 22983 3049
rect 22925 3009 22937 3043
rect 22971 3040 22983 3043
rect 23658 3040 23664 3052
rect 22971 3012 23664 3040
rect 22971 3009 22983 3012
rect 22925 3003 22983 3009
rect 19518 2932 19524 2984
rect 19576 2972 19582 2984
rect 19705 2975 19763 2981
rect 19705 2972 19717 2975
rect 19576 2944 19717 2972
rect 19576 2932 19582 2944
rect 19705 2941 19717 2944
rect 19751 2941 19763 2975
rect 19705 2935 19763 2941
rect 18432 2876 19748 2904
rect 17727 2873 17739 2876
rect 17681 2867 17739 2873
rect 17586 2836 17592 2848
rect 16684 2808 17592 2836
rect 17586 2796 17592 2808
rect 17644 2796 17650 2848
rect 19610 2796 19616 2848
rect 19668 2796 19674 2848
rect 19720 2836 19748 2876
rect 20364 2876 22094 2904
rect 20364 2836 20392 2876
rect 19720 2808 20392 2836
rect 21818 2796 21824 2848
rect 21876 2796 21882 2848
rect 22066 2836 22094 2876
rect 22940 2836 22968 3003
rect 23658 3000 23664 3012
rect 23716 3000 23722 3052
rect 25038 3000 25044 3052
rect 25096 3040 25102 3052
rect 25866 3040 25872 3052
rect 25096 3012 25872 3040
rect 25096 3000 25102 3012
rect 25866 3000 25872 3012
rect 25924 3000 25930 3052
rect 26145 3043 26203 3049
rect 26145 3009 26157 3043
rect 26191 3040 26203 3043
rect 26436 3040 26464 3080
rect 28258 3068 28264 3120
rect 28316 3108 28322 3120
rect 28316 3080 31064 3108
rect 28316 3068 28322 3080
rect 26191 3012 26464 3040
rect 26191 3009 26203 3012
rect 26145 3003 26203 3009
rect 24486 2932 24492 2984
rect 24544 2972 24550 2984
rect 24765 2975 24823 2981
rect 24765 2972 24777 2975
rect 24544 2944 24777 2972
rect 24544 2932 24550 2944
rect 24765 2941 24777 2944
rect 24811 2941 24823 2975
rect 26160 2972 26188 3003
rect 27430 3000 27436 3052
rect 27488 3000 27494 3052
rect 29546 3000 29552 3052
rect 29604 3040 29610 3052
rect 29641 3043 29699 3049
rect 29641 3040 29653 3043
rect 29604 3012 29653 3040
rect 29604 3000 29610 3012
rect 29641 3009 29653 3012
rect 29687 3009 29699 3043
rect 29641 3003 29699 3009
rect 30834 3000 30840 3052
rect 30892 3000 30898 3052
rect 24765 2935 24823 2941
rect 25424 2944 26188 2972
rect 22066 2808 22968 2836
rect 24780 2836 24808 2935
rect 25424 2836 25452 2944
rect 26234 2932 26240 2984
rect 26292 2972 26298 2984
rect 29365 2975 29423 2981
rect 29365 2972 29377 2975
rect 26292 2944 29377 2972
rect 26292 2932 26298 2944
rect 29365 2941 29377 2944
rect 29411 2941 29423 2975
rect 29365 2935 29423 2941
rect 30742 2932 30748 2984
rect 30800 2972 30806 2984
rect 31036 2981 31064 3080
rect 31726 3080 38516 3108
rect 31478 3000 31484 3052
rect 31536 3000 31542 3052
rect 30929 2975 30987 2981
rect 30929 2972 30941 2975
rect 30800 2944 30941 2972
rect 30800 2932 30806 2944
rect 30929 2941 30941 2944
rect 30975 2941 30987 2975
rect 30929 2935 30987 2941
rect 31021 2975 31079 2981
rect 31021 2941 31033 2975
rect 31067 2941 31079 2975
rect 31021 2935 31079 2941
rect 26053 2907 26111 2913
rect 26053 2873 26065 2907
rect 26099 2904 26111 2907
rect 31726 2904 31754 3080
rect 33689 3043 33747 3049
rect 33689 3009 33701 3043
rect 33735 3040 33747 3043
rect 33778 3040 33784 3052
rect 33735 3012 33784 3040
rect 33735 3009 33747 3012
rect 33689 3003 33747 3009
rect 33778 3000 33784 3012
rect 33836 3000 33842 3052
rect 33965 3043 34023 3049
rect 33965 3009 33977 3043
rect 34011 3040 34023 3043
rect 34241 3043 34299 3049
rect 34241 3040 34253 3043
rect 34011 3012 34253 3040
rect 34011 3009 34023 3012
rect 33965 3003 34023 3009
rect 34241 3009 34253 3012
rect 34287 3040 34299 3043
rect 34422 3040 34428 3052
rect 34287 3012 34428 3040
rect 34287 3009 34299 3012
rect 34241 3003 34299 3009
rect 34422 3000 34428 3012
rect 34480 3000 34486 3052
rect 38378 3000 38384 3052
rect 38436 3000 38442 3052
rect 38488 3049 38516 3080
rect 38473 3043 38531 3049
rect 38473 3009 38485 3043
rect 38519 3009 38531 3043
rect 38473 3003 38531 3009
rect 38654 3000 38660 3052
rect 38712 3040 38718 3052
rect 38841 3043 38899 3049
rect 38841 3040 38853 3043
rect 38712 3012 38853 3040
rect 38712 3000 38718 3012
rect 38841 3009 38853 3012
rect 38887 3009 38899 3043
rect 38841 3003 38899 3009
rect 38930 3000 38936 3052
rect 38988 3040 38994 3052
rect 39209 3043 39267 3049
rect 39209 3040 39221 3043
rect 38988 3012 39221 3040
rect 38988 3000 38994 3012
rect 39209 3009 39221 3012
rect 39255 3009 39267 3043
rect 39209 3003 39267 3009
rect 26099 2876 29500 2904
rect 26099 2873 26111 2876
rect 26053 2867 26111 2873
rect 24780 2808 25452 2836
rect 29472 2836 29500 2876
rect 30392 2876 31754 2904
rect 30392 2836 30420 2876
rect 29472 2808 30420 2836
rect 30466 2796 30472 2848
rect 30524 2796 30530 2848
rect 32950 2796 32956 2848
rect 33008 2796 33014 2848
rect 38654 2796 38660 2848
rect 38712 2796 38718 2848
rect 39022 2796 39028 2848
rect 39080 2796 39086 2848
rect 1104 2746 39836 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 37950 2746
rect 38002 2694 38014 2746
rect 38066 2694 38078 2746
rect 38130 2694 38142 2746
rect 38194 2694 38206 2746
rect 38258 2694 39836 2746
rect 1104 2672 39836 2694
rect 4798 2632 4804 2644
rect 2608 2604 4804 2632
rect 1210 2456 1216 2508
rect 1268 2496 1274 2508
rect 2608 2505 2636 2604
rect 4798 2592 4804 2604
rect 4856 2592 4862 2644
rect 5902 2592 5908 2644
rect 5960 2592 5966 2644
rect 10226 2592 10232 2644
rect 10284 2632 10290 2644
rect 10321 2635 10379 2641
rect 10321 2632 10333 2635
rect 10284 2604 10333 2632
rect 10284 2592 10290 2604
rect 10321 2601 10333 2604
rect 10367 2601 10379 2635
rect 10321 2595 10379 2601
rect 11333 2635 11391 2641
rect 11333 2601 11345 2635
rect 11379 2632 11391 2635
rect 11882 2632 11888 2644
rect 11379 2604 11888 2632
rect 11379 2601 11391 2604
rect 11333 2595 11391 2601
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 12621 2635 12679 2641
rect 12621 2601 12633 2635
rect 12667 2632 12679 2635
rect 12802 2632 12808 2644
rect 12667 2604 12808 2632
rect 12667 2601 12679 2604
rect 12621 2595 12679 2601
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 12986 2592 12992 2644
rect 13044 2632 13050 2644
rect 16850 2632 16856 2644
rect 13044 2604 16856 2632
rect 13044 2592 13050 2604
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 17037 2635 17095 2641
rect 17037 2601 17049 2635
rect 17083 2632 17095 2635
rect 17402 2632 17408 2644
rect 17083 2604 17408 2632
rect 17083 2601 17095 2604
rect 17037 2595 17095 2601
rect 17402 2592 17408 2604
rect 17460 2592 17466 2644
rect 21818 2632 21824 2644
rect 17696 2604 21824 2632
rect 4154 2524 4160 2576
rect 4212 2564 4218 2576
rect 4706 2564 4712 2576
rect 4212 2536 4712 2564
rect 4212 2524 4218 2536
rect 4706 2524 4712 2536
rect 4764 2524 4770 2576
rect 5718 2524 5724 2576
rect 5776 2564 5782 2576
rect 5776 2536 7236 2564
rect 5776 2524 5782 2536
rect 2317 2499 2375 2505
rect 2317 2496 2329 2499
rect 1268 2468 2329 2496
rect 1268 2456 1274 2468
rect 2317 2465 2329 2468
rect 2363 2465 2375 2499
rect 2317 2459 2375 2465
rect 2593 2499 2651 2505
rect 2593 2465 2605 2499
rect 2639 2465 2651 2499
rect 2593 2459 2651 2465
rect 4246 2456 4252 2508
rect 4304 2496 4310 2508
rect 4801 2499 4859 2505
rect 4801 2496 4813 2499
rect 4304 2468 4813 2496
rect 4304 2456 4310 2468
rect 4801 2465 4813 2468
rect 4847 2465 4859 2499
rect 4801 2459 4859 2465
rect 4890 2456 4896 2508
rect 4948 2456 4954 2508
rect 6178 2456 6184 2508
rect 6236 2496 6242 2508
rect 6236 2468 6868 2496
rect 6236 2456 6242 2468
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 1360 2400 1409 2428
rect 1360 2388 1366 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2428 3479 2431
rect 3510 2428 3516 2440
rect 3467 2400 3516 2428
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 3510 2388 3516 2400
rect 3568 2388 3574 2440
rect 4525 2431 4583 2437
rect 4525 2397 4537 2431
rect 4571 2397 4583 2431
rect 4525 2391 4583 2397
rect 4540 2360 4568 2391
rect 4706 2388 4712 2440
rect 4764 2428 4770 2440
rect 5169 2431 5227 2437
rect 5169 2428 5181 2431
rect 4764 2400 5181 2428
rect 4764 2388 4770 2400
rect 5169 2397 5181 2400
rect 5215 2428 5227 2431
rect 5997 2431 6055 2437
rect 5215 2400 5948 2428
rect 5215 2397 5227 2400
rect 5169 2391 5227 2397
rect 5810 2360 5816 2372
rect 4540 2332 5816 2360
rect 5810 2320 5816 2332
rect 5868 2320 5874 2372
rect 5920 2360 5948 2400
rect 5997 2397 6009 2431
rect 6043 2428 6055 2431
rect 6362 2428 6368 2440
rect 6043 2400 6368 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 6362 2388 6368 2400
rect 6420 2388 6426 2440
rect 6840 2437 6868 2468
rect 7208 2437 7236 2536
rect 9858 2524 9864 2576
rect 9916 2564 9922 2576
rect 11054 2564 11060 2576
rect 9916 2536 11060 2564
rect 9916 2524 9922 2536
rect 11054 2524 11060 2536
rect 11112 2524 11118 2576
rect 16114 2564 16120 2576
rect 11256 2536 16120 2564
rect 7377 2499 7435 2505
rect 7377 2465 7389 2499
rect 7423 2496 7435 2499
rect 9766 2496 9772 2508
rect 7423 2468 9772 2496
rect 7423 2465 7435 2468
rect 7377 2459 7435 2465
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 10781 2499 10839 2505
rect 10781 2465 10793 2499
rect 10827 2496 10839 2499
rect 11256 2496 11284 2536
rect 16114 2524 16120 2536
rect 16172 2524 16178 2576
rect 16574 2524 16580 2576
rect 16632 2564 16638 2576
rect 16632 2536 17540 2564
rect 16632 2524 16638 2536
rect 17512 2508 17540 2536
rect 10827 2468 11284 2496
rect 10827 2465 10839 2468
rect 10781 2459 10839 2465
rect 11330 2456 11336 2508
rect 11388 2496 11394 2508
rect 11388 2468 14136 2496
rect 11388 2456 11394 2468
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2428 6883 2431
rect 7193 2431 7251 2437
rect 6871 2400 7144 2428
rect 6871 2397 6883 2400
rect 6825 2391 6883 2397
rect 6270 2360 6276 2372
rect 5920 2332 6276 2360
rect 6270 2320 6276 2332
rect 6328 2360 6334 2372
rect 6457 2363 6515 2369
rect 6457 2360 6469 2363
rect 6328 2332 6469 2360
rect 6328 2320 6334 2332
rect 6457 2329 6469 2332
rect 6503 2329 6515 2363
rect 6457 2323 6515 2329
rect 6638 2320 6644 2372
rect 6696 2320 6702 2372
rect 7006 2320 7012 2372
rect 7064 2320 7070 2372
rect 7116 2360 7144 2400
rect 7193 2397 7205 2431
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 7282 2388 7288 2440
rect 7340 2428 7346 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 7340 2400 7481 2428
rect 7340 2388 7346 2400
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 7926 2388 7932 2440
rect 7984 2428 7990 2440
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7984 2400 8033 2428
rect 7984 2388 7990 2400
rect 8021 2397 8033 2400
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 9398 2388 9404 2440
rect 9456 2428 9462 2440
rect 9493 2431 9551 2437
rect 9493 2428 9505 2431
rect 9456 2400 9505 2428
rect 9456 2388 9462 2400
rect 9493 2397 9505 2400
rect 9539 2397 9551 2431
rect 9493 2391 9551 2397
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 10134 2428 10140 2440
rect 10091 2400 10140 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2428 10563 2431
rect 10870 2428 10876 2440
rect 10551 2400 10876 2428
rect 10551 2397 10563 2400
rect 10505 2391 10563 2397
rect 10870 2388 10876 2400
rect 10928 2388 10934 2440
rect 10965 2431 11023 2437
rect 10965 2397 10977 2431
rect 11011 2428 11023 2431
rect 11054 2428 11060 2440
rect 11011 2400 11060 2428
rect 11011 2397 11023 2400
rect 10965 2391 11023 2397
rect 11054 2388 11060 2400
rect 11112 2428 11118 2440
rect 11698 2428 11704 2440
rect 11112 2400 11704 2428
rect 11112 2388 11118 2400
rect 11698 2388 11704 2400
rect 11756 2388 11762 2440
rect 12342 2388 12348 2440
rect 12400 2428 12406 2440
rect 14108 2437 14136 2468
rect 17494 2456 17500 2508
rect 17552 2456 17558 2508
rect 17696 2505 17724 2604
rect 21818 2592 21824 2604
rect 21876 2592 21882 2644
rect 22278 2632 22284 2644
rect 22020 2604 22284 2632
rect 22020 2505 22048 2604
rect 22278 2592 22284 2604
rect 22336 2592 22342 2644
rect 22646 2592 22652 2644
rect 22704 2632 22710 2644
rect 23661 2635 23719 2641
rect 23661 2632 23673 2635
rect 22704 2604 23673 2632
rect 22704 2592 22710 2604
rect 23661 2601 23673 2604
rect 23707 2601 23719 2635
rect 23661 2595 23719 2601
rect 24044 2604 31064 2632
rect 22922 2524 22928 2576
rect 22980 2564 22986 2576
rect 23017 2567 23075 2573
rect 23017 2564 23029 2567
rect 22980 2536 23029 2564
rect 22980 2524 22986 2536
rect 23017 2533 23029 2536
rect 23063 2533 23075 2567
rect 23017 2527 23075 2533
rect 23290 2524 23296 2576
rect 23348 2524 23354 2576
rect 23382 2524 23388 2576
rect 23440 2564 23446 2576
rect 23937 2567 23995 2573
rect 23937 2564 23949 2567
rect 23440 2536 23949 2564
rect 23440 2524 23446 2536
rect 23937 2533 23949 2536
rect 23983 2533 23995 2567
rect 23937 2527 23995 2533
rect 17681 2499 17739 2505
rect 17681 2465 17693 2499
rect 17727 2465 17739 2499
rect 20349 2499 20407 2505
rect 17681 2459 17739 2465
rect 17788 2468 18460 2496
rect 12437 2431 12495 2437
rect 12437 2428 12449 2431
rect 12400 2400 12449 2428
rect 12400 2388 12406 2400
rect 12437 2397 12449 2400
rect 12483 2397 12495 2431
rect 12437 2391 12495 2397
rect 13449 2431 13507 2437
rect 13449 2397 13461 2431
rect 13495 2397 13507 2431
rect 13449 2391 13507 2397
rect 14093 2431 14151 2437
rect 14093 2397 14105 2431
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 7558 2360 7564 2372
rect 7116 2332 7564 2360
rect 7558 2320 7564 2332
rect 7616 2320 7622 2372
rect 8662 2320 8668 2372
rect 8720 2360 8726 2372
rect 9033 2363 9091 2369
rect 9033 2360 9045 2363
rect 8720 2332 9045 2360
rect 8720 2320 8726 2332
rect 9033 2329 9045 2332
rect 9079 2329 9091 2363
rect 9033 2323 9091 2329
rect 9214 2320 9220 2372
rect 9272 2320 9278 2372
rect 10244 2332 11560 2360
rect 3513 2295 3571 2301
rect 3513 2261 3525 2295
rect 3559 2292 3571 2295
rect 3694 2292 3700 2304
rect 3559 2264 3700 2292
rect 3559 2261 3571 2264
rect 3513 2255 3571 2261
rect 3694 2252 3700 2264
rect 3752 2252 3758 2304
rect 6178 2252 6184 2304
rect 6236 2252 6242 2304
rect 7650 2252 7656 2304
rect 7708 2252 7714 2304
rect 8202 2252 8208 2304
rect 8260 2252 8266 2304
rect 9674 2252 9680 2304
rect 9732 2252 9738 2304
rect 10244 2301 10272 2332
rect 10229 2295 10287 2301
rect 10229 2261 10241 2295
rect 10275 2261 10287 2295
rect 10229 2255 10287 2261
rect 10318 2252 10324 2304
rect 10376 2292 10382 2304
rect 10873 2295 10931 2301
rect 10873 2292 10885 2295
rect 10376 2264 10885 2292
rect 10376 2252 10382 2264
rect 10873 2261 10885 2264
rect 10919 2261 10931 2295
rect 11532 2292 11560 2332
rect 11606 2320 11612 2372
rect 11664 2360 11670 2372
rect 11793 2363 11851 2369
rect 11793 2360 11805 2363
rect 11664 2332 11805 2360
rect 11664 2320 11670 2332
rect 11793 2329 11805 2332
rect 11839 2329 11851 2363
rect 11793 2323 11851 2329
rect 11974 2320 11980 2372
rect 12032 2320 12038 2372
rect 13464 2360 13492 2391
rect 14918 2388 14924 2440
rect 14976 2388 14982 2440
rect 15654 2388 15660 2440
rect 15712 2388 15718 2440
rect 15746 2388 15752 2440
rect 15804 2428 15810 2440
rect 16117 2431 16175 2437
rect 16117 2428 16129 2431
rect 15804 2400 16129 2428
rect 15804 2388 15810 2400
rect 16117 2397 16129 2400
rect 16163 2397 16175 2431
rect 16117 2391 16175 2397
rect 16206 2388 16212 2440
rect 16264 2428 16270 2440
rect 16669 2431 16727 2437
rect 16264 2418 16574 2428
rect 16669 2418 16681 2431
rect 16264 2400 16681 2418
rect 16264 2388 16270 2400
rect 16546 2397 16681 2400
rect 16715 2397 16727 2431
rect 17788 2428 17816 2468
rect 16546 2391 16727 2397
rect 16776 2400 17816 2428
rect 16546 2390 16712 2391
rect 16776 2360 16804 2400
rect 18138 2388 18144 2440
rect 18196 2388 18202 2440
rect 18325 2431 18383 2437
rect 18325 2397 18337 2431
rect 18371 2397 18383 2431
rect 18325 2391 18383 2397
rect 13464 2332 16804 2360
rect 17126 2320 17132 2372
rect 17184 2360 17190 2372
rect 18340 2360 18368 2391
rect 17184 2332 18368 2360
rect 18432 2360 18460 2468
rect 20349 2465 20361 2499
rect 20395 2496 20407 2499
rect 22005 2499 22063 2505
rect 22005 2496 22017 2499
rect 20395 2468 22017 2496
rect 20395 2465 20407 2468
rect 20349 2459 20407 2465
rect 22005 2465 22017 2468
rect 22051 2465 22063 2499
rect 22005 2459 22063 2465
rect 22738 2456 22744 2508
rect 22796 2496 22802 2508
rect 24044 2496 24072 2604
rect 29822 2564 29828 2576
rect 22796 2468 24072 2496
rect 24136 2536 29828 2564
rect 22796 2456 22802 2468
rect 18782 2388 18788 2440
rect 18840 2428 18846 2440
rect 19061 2431 19119 2437
rect 19061 2428 19073 2431
rect 18840 2400 19073 2428
rect 18840 2388 18846 2400
rect 19061 2397 19073 2400
rect 19107 2397 19119 2431
rect 19061 2391 19119 2397
rect 19426 2388 19432 2440
rect 19484 2428 19490 2440
rect 20073 2431 20131 2437
rect 20073 2428 20085 2431
rect 19484 2400 20085 2428
rect 19484 2388 19490 2400
rect 20073 2397 20085 2400
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 20714 2388 20720 2440
rect 20772 2388 20778 2440
rect 20809 2431 20867 2437
rect 20809 2397 20821 2431
rect 20855 2397 20867 2431
rect 20809 2391 20867 2397
rect 20732 2360 20760 2388
rect 18432 2332 20760 2360
rect 20824 2360 20852 2391
rect 20898 2388 20904 2440
rect 20956 2388 20962 2440
rect 21450 2388 21456 2440
rect 21508 2428 21514 2440
rect 21545 2431 21603 2437
rect 21545 2428 21557 2431
rect 21508 2400 21557 2428
rect 21508 2388 21514 2400
rect 21545 2397 21557 2400
rect 21591 2397 21603 2431
rect 21545 2391 21603 2397
rect 21818 2388 21824 2440
rect 21876 2428 21882 2440
rect 22281 2431 22339 2437
rect 22281 2428 22293 2431
rect 21876 2400 22293 2428
rect 21876 2388 21882 2400
rect 22281 2397 22293 2400
rect 22327 2397 22339 2431
rect 22281 2391 22339 2397
rect 22296 2360 22324 2391
rect 22370 2388 22376 2440
rect 22428 2428 22434 2440
rect 23109 2431 23167 2437
rect 23109 2428 23121 2431
rect 22428 2400 23121 2428
rect 22428 2388 22434 2400
rect 23109 2397 23121 2400
rect 23155 2397 23167 2431
rect 23109 2391 23167 2397
rect 23474 2388 23480 2440
rect 23532 2388 23538 2440
rect 24136 2437 24164 2536
rect 29822 2524 29828 2536
rect 29880 2524 29886 2576
rect 31036 2564 31064 2604
rect 31478 2592 31484 2644
rect 31536 2632 31542 2644
rect 31665 2635 31723 2641
rect 31665 2632 31677 2635
rect 31536 2604 31677 2632
rect 31536 2592 31542 2604
rect 31665 2601 31677 2604
rect 31711 2601 31723 2635
rect 31665 2595 31723 2601
rect 33321 2635 33379 2641
rect 33321 2601 33333 2635
rect 33367 2632 33379 2635
rect 33410 2632 33416 2644
rect 33367 2604 33416 2632
rect 33367 2601 33379 2604
rect 33321 2595 33379 2601
rect 33410 2592 33416 2604
rect 33468 2592 33474 2644
rect 39390 2592 39396 2644
rect 39448 2592 39454 2644
rect 39025 2567 39083 2573
rect 31036 2536 35894 2564
rect 31113 2499 31171 2505
rect 26206 2468 30604 2496
rect 24121 2431 24179 2437
rect 24121 2397 24133 2431
rect 24167 2397 24179 2431
rect 24121 2391 24179 2397
rect 24394 2388 24400 2440
rect 24452 2388 24458 2440
rect 22554 2360 22560 2372
rect 20824 2332 22232 2360
rect 22296 2332 22560 2360
rect 17184 2320 17190 2332
rect 12986 2292 12992 2304
rect 11532 2264 12992 2292
rect 10873 2255 10931 2261
rect 12986 2252 12992 2264
rect 13044 2252 13050 2304
rect 13078 2252 13084 2304
rect 13136 2292 13142 2304
rect 13265 2295 13323 2301
rect 13265 2292 13277 2295
rect 13136 2264 13277 2292
rect 13136 2252 13142 2264
rect 13265 2261 13277 2264
rect 13311 2261 13323 2295
rect 13265 2255 13323 2261
rect 13814 2252 13820 2304
rect 13872 2292 13878 2304
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 13872 2264 14289 2292
rect 13872 2252 13878 2264
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 14277 2255 14335 2261
rect 14550 2252 14556 2304
rect 14608 2292 14614 2304
rect 14737 2295 14795 2301
rect 14737 2292 14749 2295
rect 14608 2264 14749 2292
rect 14608 2252 14614 2264
rect 14737 2261 14749 2264
rect 14783 2261 14795 2295
rect 14737 2255 14795 2261
rect 15378 2252 15384 2304
rect 15436 2292 15442 2304
rect 15473 2295 15531 2301
rect 15473 2292 15485 2295
rect 15436 2264 15485 2292
rect 15436 2252 15442 2264
rect 15473 2261 15485 2264
rect 15519 2261 15531 2295
rect 15473 2255 15531 2261
rect 16022 2252 16028 2304
rect 16080 2292 16086 2304
rect 16301 2295 16359 2301
rect 16301 2292 16313 2295
rect 16080 2264 16313 2292
rect 16080 2252 16086 2264
rect 16301 2261 16313 2264
rect 16347 2261 16359 2295
rect 16301 2255 16359 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 16853 2295 16911 2301
rect 16853 2292 16865 2295
rect 16816 2264 16865 2292
rect 16816 2252 16822 2264
rect 16853 2261 16865 2264
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 17405 2295 17463 2301
rect 17405 2261 17417 2295
rect 17451 2292 17463 2295
rect 17678 2292 17684 2304
rect 17451 2264 17684 2292
rect 17451 2261 17463 2264
rect 17405 2255 17463 2261
rect 17678 2252 17684 2264
rect 17736 2252 17742 2304
rect 17770 2252 17776 2304
rect 17828 2292 17834 2304
rect 17957 2295 18015 2301
rect 17957 2292 17969 2295
rect 17828 2264 17969 2292
rect 17828 2252 17834 2264
rect 17957 2261 17969 2264
rect 18003 2261 18015 2295
rect 17957 2255 18015 2261
rect 18230 2252 18236 2304
rect 18288 2292 18294 2304
rect 18509 2295 18567 2301
rect 18509 2292 18521 2295
rect 18288 2264 18521 2292
rect 18288 2252 18294 2264
rect 18509 2261 18521 2264
rect 18555 2261 18567 2295
rect 18509 2255 18567 2261
rect 18877 2295 18935 2301
rect 18877 2261 18889 2295
rect 18923 2292 18935 2295
rect 18966 2292 18972 2304
rect 18923 2264 18972 2292
rect 18923 2261 18935 2264
rect 18877 2255 18935 2261
rect 18966 2252 18972 2264
rect 19024 2252 19030 2304
rect 19334 2252 19340 2304
rect 19392 2252 19398 2304
rect 20438 2252 20444 2304
rect 20496 2292 20502 2304
rect 20625 2295 20683 2301
rect 20625 2292 20637 2295
rect 20496 2264 20637 2292
rect 20496 2252 20502 2264
rect 20625 2261 20637 2264
rect 20671 2261 20683 2295
rect 20625 2255 20683 2261
rect 20714 2252 20720 2304
rect 20772 2292 20778 2304
rect 21085 2295 21143 2301
rect 21085 2292 21097 2295
rect 20772 2264 21097 2292
rect 20772 2252 20778 2264
rect 21085 2261 21097 2264
rect 21131 2261 21143 2295
rect 21085 2255 21143 2261
rect 21358 2252 21364 2304
rect 21416 2252 21422 2304
rect 22204 2292 22232 2332
rect 22554 2320 22560 2332
rect 22612 2320 22618 2372
rect 26206 2360 26234 2468
rect 30466 2388 30472 2440
rect 30524 2388 30530 2440
rect 30576 2428 30604 2468
rect 31113 2465 31125 2499
rect 31159 2496 31171 2499
rect 32950 2496 32956 2508
rect 31159 2468 32956 2496
rect 31159 2465 31171 2468
rect 31113 2459 31171 2465
rect 32950 2456 32956 2468
rect 33008 2456 33014 2508
rect 33594 2496 33600 2508
rect 33060 2468 33600 2496
rect 33060 2428 33088 2468
rect 33594 2456 33600 2468
rect 33652 2456 33658 2508
rect 35866 2496 35894 2536
rect 39025 2533 39037 2567
rect 39071 2564 39083 2567
rect 39942 2564 39948 2576
rect 39071 2536 39948 2564
rect 39071 2533 39083 2536
rect 39025 2527 39083 2533
rect 39942 2524 39948 2536
rect 40000 2524 40006 2576
rect 35866 2468 39252 2496
rect 30576 2400 33088 2428
rect 33410 2388 33416 2440
rect 33468 2428 33474 2440
rect 37737 2431 37795 2437
rect 37737 2428 37749 2431
rect 33468 2400 37749 2428
rect 33468 2388 33474 2400
rect 37737 2397 37749 2400
rect 37783 2397 37795 2431
rect 37737 2391 37795 2397
rect 38102 2388 38108 2440
rect 38160 2388 38166 2440
rect 38470 2388 38476 2440
rect 38528 2388 38534 2440
rect 38562 2388 38568 2440
rect 38620 2428 38626 2440
rect 39224 2437 39252 2468
rect 38841 2431 38899 2437
rect 38841 2428 38853 2431
rect 38620 2400 38853 2428
rect 38620 2388 38626 2400
rect 38841 2397 38853 2400
rect 38887 2397 38899 2431
rect 38841 2391 38899 2397
rect 39209 2431 39267 2437
rect 39209 2397 39221 2431
rect 39255 2397 39267 2431
rect 39209 2391 39267 2397
rect 23492 2332 26234 2360
rect 23492 2292 23520 2332
rect 26326 2320 26332 2372
rect 26384 2360 26390 2372
rect 33229 2363 33287 2369
rect 33229 2360 33241 2363
rect 26384 2332 33241 2360
rect 26384 2320 26390 2332
rect 33229 2329 33241 2332
rect 33275 2329 33287 2363
rect 33229 2323 33287 2329
rect 22204 2264 23520 2292
rect 24118 2252 24124 2304
rect 24176 2292 24182 2304
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 24176 2264 24593 2292
rect 24176 2252 24182 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 30282 2252 30288 2304
rect 30340 2252 30346 2304
rect 30742 2252 30748 2304
rect 30800 2292 30806 2304
rect 31205 2295 31263 2301
rect 31205 2292 31217 2295
rect 30800 2264 31217 2292
rect 30800 2252 30806 2264
rect 31205 2261 31217 2264
rect 31251 2261 31263 2295
rect 31205 2255 31263 2261
rect 31294 2252 31300 2304
rect 31352 2252 31358 2304
rect 37918 2252 37924 2304
rect 37976 2252 37982 2304
rect 38286 2252 38292 2304
rect 38344 2252 38350 2304
rect 38654 2252 38660 2304
rect 38712 2252 38718 2304
rect 1104 2202 39836 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 39010 2202
rect 39062 2150 39074 2202
rect 39126 2150 39138 2202
rect 39190 2150 39202 2202
rect 39254 2150 39266 2202
rect 39318 2150 39836 2202
rect 1104 2128 39836 2150
rect 4798 2048 4804 2100
rect 4856 2088 4862 2100
rect 7558 2088 7564 2100
rect 4856 2060 7564 2088
rect 4856 2048 4862 2060
rect 7558 2048 7564 2060
rect 7616 2048 7622 2100
rect 10962 2048 10968 2100
rect 11020 2088 11026 2100
rect 20898 2088 20904 2100
rect 11020 2060 20904 2088
rect 11020 2048 11026 2060
rect 20898 2048 20904 2060
rect 20956 2048 20962 2100
rect 29822 2048 29828 2100
rect 29880 2088 29886 2100
rect 32306 2088 32312 2100
rect 29880 2060 32312 2088
rect 29880 2048 29886 2060
rect 32306 2048 32312 2060
rect 32364 2048 32370 2100
rect 32950 2048 32956 2100
rect 33008 2088 33014 2100
rect 38378 2088 38384 2100
rect 33008 2060 38384 2088
rect 33008 2048 33014 2060
rect 38378 2048 38384 2060
rect 38436 2048 38442 2100
rect 9674 1980 9680 2032
rect 9732 2020 9738 2032
rect 25406 2020 25412 2032
rect 9732 1992 25412 2020
rect 9732 1980 9738 1992
rect 25406 1980 25412 1992
rect 25464 1980 25470 2032
rect 1670 1912 1676 1964
rect 1728 1952 1734 1964
rect 19242 1952 19248 1964
rect 1728 1924 19248 1952
rect 1728 1912 1734 1924
rect 19242 1912 19248 1924
rect 19300 1912 19306 1964
rect 19610 1912 19616 1964
rect 19668 1952 19674 1964
rect 38562 1952 38568 1964
rect 19668 1924 38568 1952
rect 19668 1912 19674 1924
rect 38562 1912 38568 1924
rect 38620 1912 38626 1964
rect 3694 1844 3700 1896
rect 3752 1884 3758 1896
rect 11514 1884 11520 1896
rect 3752 1856 11520 1884
rect 3752 1844 3758 1856
rect 11514 1844 11520 1856
rect 11572 1844 11578 1896
rect 15654 1844 15660 1896
rect 15712 1884 15718 1896
rect 24302 1884 24308 1896
rect 15712 1856 24308 1884
rect 15712 1844 15718 1856
rect 24302 1844 24308 1856
rect 24360 1844 24366 1896
rect 2866 1776 2872 1828
rect 2924 1816 2930 1828
rect 21634 1816 21640 1828
rect 2924 1788 21640 1816
rect 2924 1776 2930 1788
rect 21634 1776 21640 1788
rect 21692 1776 21698 1828
rect 21910 1776 21916 1828
rect 21968 1816 21974 1828
rect 23290 1816 23296 1828
rect 21968 1788 23296 1816
rect 21968 1776 21974 1788
rect 23290 1776 23296 1788
rect 23348 1776 23354 1828
rect 25590 1776 25596 1828
rect 25648 1816 25654 1828
rect 27798 1816 27804 1828
rect 25648 1788 27804 1816
rect 25648 1776 25654 1788
rect 27798 1776 27804 1788
rect 27856 1776 27862 1828
rect 6178 1708 6184 1760
rect 6236 1748 6242 1760
rect 12434 1748 12440 1760
rect 6236 1720 12440 1748
rect 6236 1708 6242 1720
rect 12434 1708 12440 1720
rect 12492 1708 12498 1760
rect 14826 1708 14832 1760
rect 14884 1748 14890 1760
rect 24394 1748 24400 1760
rect 14884 1720 24400 1748
rect 14884 1708 14890 1720
rect 24394 1708 24400 1720
rect 24452 1708 24458 1760
rect 7650 1640 7656 1692
rect 7708 1680 7714 1692
rect 14734 1680 14740 1692
rect 7708 1652 14740 1680
rect 7708 1640 7714 1652
rect 14734 1640 14740 1652
rect 14792 1640 14798 1692
rect 14918 1640 14924 1692
rect 14976 1680 14982 1692
rect 29178 1680 29184 1692
rect 14976 1652 29184 1680
rect 14976 1640 14982 1652
rect 29178 1640 29184 1652
rect 29236 1640 29242 1692
rect 18138 1572 18144 1624
rect 18196 1612 18202 1624
rect 29086 1612 29092 1624
rect 18196 1584 29092 1612
rect 18196 1572 18202 1584
rect 29086 1572 29092 1584
rect 29144 1572 29150 1624
rect 8202 1504 8208 1556
rect 8260 1544 8266 1556
rect 16574 1544 16580 1556
rect 8260 1516 16580 1544
rect 8260 1504 8266 1516
rect 16574 1504 16580 1516
rect 16632 1504 16638 1556
rect 21726 1504 21732 1556
rect 21784 1544 21790 1556
rect 38102 1544 38108 1556
rect 21784 1516 38108 1544
rect 21784 1504 21790 1516
rect 38102 1504 38108 1516
rect 38160 1504 38166 1556
rect 10778 1436 10784 1488
rect 10836 1476 10842 1488
rect 19334 1476 19340 1488
rect 10836 1448 19340 1476
rect 10836 1436 10842 1448
rect 19334 1436 19340 1448
rect 19392 1436 19398 1488
rect 27062 1368 27068 1420
rect 27120 1408 27126 1420
rect 28994 1408 29000 1420
rect 27120 1380 29000 1408
rect 27120 1368 27126 1380
rect 28994 1368 29000 1380
rect 29052 1368 29058 1420
rect 35710 1368 35716 1420
rect 35768 1408 35774 1420
rect 38102 1408 38108 1420
rect 35768 1380 38108 1408
rect 35768 1368 35774 1380
rect 38102 1368 38108 1380
rect 38160 1368 38166 1420
rect 14458 1300 14464 1352
rect 14516 1340 14522 1352
rect 32766 1340 32772 1352
rect 14516 1312 32772 1340
rect 14516 1300 14522 1312
rect 32766 1300 32772 1312
rect 32824 1300 32830 1352
rect 9950 1232 9956 1284
rect 10008 1272 10014 1284
rect 39666 1272 39672 1284
rect 10008 1244 39672 1272
rect 10008 1232 10014 1244
rect 39666 1232 39672 1244
rect 39724 1232 39730 1284
rect 7558 1164 7564 1216
rect 7616 1204 7622 1216
rect 21542 1204 21548 1216
rect 7616 1176 21548 1204
rect 7616 1164 7622 1176
rect 21542 1164 21548 1176
rect 21600 1164 21606 1216
rect 2498 1096 2504 1148
rect 2556 1136 2562 1148
rect 29454 1136 29460 1148
rect 2556 1108 29460 1136
rect 2556 1096 2562 1108
rect 29454 1096 29460 1108
rect 29512 1096 29518 1148
rect 8570 1028 8576 1080
rect 8628 1068 8634 1080
rect 35066 1068 35072 1080
rect 8628 1040 35072 1068
rect 8628 1028 8634 1040
rect 35066 1028 35072 1040
rect 35124 1028 35130 1080
rect 2682 960 2688 1012
rect 2740 1000 2746 1012
rect 25038 1000 25044 1012
rect 2740 972 25044 1000
rect 2740 960 2746 972
rect 25038 960 25044 972
rect 25096 960 25102 1012
rect 32214 960 32220 1012
rect 32272 1000 32278 1012
rect 34238 1000 34244 1012
rect 32272 972 34244 1000
rect 32272 960 32278 972
rect 34238 960 34244 972
rect 34296 960 34302 1012
rect 13354 892 13360 944
rect 13412 932 13418 944
rect 37182 932 37188 944
rect 13412 904 37188 932
rect 13412 892 13418 904
rect 37182 892 37188 904
rect 37240 892 37246 944
rect 10502 824 10508 876
rect 10560 864 10566 876
rect 26602 864 26608 876
rect 10560 836 26608 864
rect 10560 824 10566 836
rect 26602 824 26608 836
rect 26660 824 26666 876
rect 7006 756 7012 808
rect 7064 796 7070 808
rect 38194 796 38200 808
rect 7064 768 38200 796
rect 7064 756 7070 768
rect 38194 756 38200 768
rect 38252 756 38258 808
rect 6638 688 6644 740
rect 6696 728 6702 740
rect 33410 728 33416 740
rect 6696 700 33416 728
rect 6696 688 6702 700
rect 33410 688 33416 700
rect 33468 688 33474 740
rect 7834 620 7840 672
rect 7892 660 7898 672
rect 23474 660 23480 672
rect 7892 632 23480 660
rect 7892 620 7898 632
rect 23474 620 23480 632
rect 23532 620 23538 672
rect 28626 8 28632 60
rect 28684 48 28690 60
rect 39850 48 39856 60
rect 28684 20 39856 48
rect 28684 8 28690 20
rect 39850 8 39856 20
rect 39908 8 39914 60
<< via1 >>
rect 10600 10820 10652 10872
rect 17224 10820 17276 10872
rect 10784 10684 10836 10736
rect 17408 10684 17460 10736
rect 8576 10412 8628 10464
rect 36452 10412 36504 10464
rect 4252 10344 4304 10396
rect 29828 10344 29880 10396
rect 17224 10276 17276 10328
rect 4160 10208 4212 10260
rect 25228 10208 25280 10260
rect 25596 10208 25648 10260
rect 26516 10208 26568 10260
rect 37648 10208 37700 10260
rect 11888 10140 11940 10192
rect 29000 10140 29052 10192
rect 6920 10072 6972 10124
rect 17224 10072 17276 10124
rect 17408 10072 17460 10124
rect 30380 10072 30432 10124
rect 8668 10004 8720 10056
rect 30748 10004 30800 10056
rect 2596 9936 2648 9988
rect 24584 9936 24636 9988
rect 14740 9868 14792 9920
rect 15108 9868 15160 9920
rect 17224 9868 17276 9920
rect 31484 9868 31536 9920
rect 9956 9800 10008 9852
rect 29552 9800 29604 9852
rect 10876 9732 10928 9784
rect 11796 9732 11848 9784
rect 12164 9732 12216 9784
rect 13084 9732 13136 9784
rect 14464 9732 14516 9784
rect 21548 9732 21600 9784
rect 25872 9732 25924 9784
rect 27436 9732 27488 9784
rect 10048 9664 10100 9716
rect 11244 9664 11296 9716
rect 11704 9664 11756 9716
rect 12900 9664 12952 9716
rect 19432 9664 19484 9716
rect 20352 9664 20404 9716
rect 20812 9664 20864 9716
rect 31760 9664 31812 9716
rect 4528 9596 4580 9648
rect 12440 9596 12492 9648
rect 12992 9596 13044 9648
rect 15568 9596 15620 9648
rect 5264 9528 5316 9580
rect 12256 9528 12308 9580
rect 13084 9528 13136 9580
rect 16580 9528 16632 9580
rect 17040 9528 17092 9580
rect 19708 9528 19760 9580
rect 28080 9596 28132 9648
rect 28908 9596 28960 9648
rect 30012 9596 30064 9648
rect 31576 9596 31628 9648
rect 28724 9528 28776 9580
rect 31852 9596 31904 9648
rect 32680 9596 32732 9648
rect 7288 9460 7340 9512
rect 7932 9460 7984 9512
rect 6368 9392 6420 9444
rect 14096 9392 14148 9444
rect 5632 9324 5684 9376
rect 11612 9324 11664 9376
rect 12716 9324 12768 9376
rect 28448 9460 28500 9512
rect 31760 9460 31812 9512
rect 18052 9392 18104 9444
rect 16948 9324 17000 9376
rect 26700 9324 26752 9376
rect 31944 9324 31996 9376
rect 2688 9256 2740 9308
rect 10324 9256 10376 9308
rect 11336 9256 11388 9308
rect 22192 9256 22244 9308
rect 24860 9256 24912 9308
rect 32864 9256 32916 9308
rect 1676 9188 1728 9240
rect 9680 9188 9732 9240
rect 11428 9188 11480 9240
rect 3608 9120 3660 9172
rect 8484 9120 8536 9172
rect 13360 9188 13412 9240
rect 19616 9188 19668 9240
rect 19708 9188 19760 9240
rect 31024 9188 31076 9240
rect 5356 9052 5408 9104
rect 9772 9052 9824 9104
rect 10140 9052 10192 9104
rect 11244 9052 11296 9104
rect 25780 9120 25832 9172
rect 25872 9120 25924 9172
rect 28080 9120 28132 9172
rect 10232 8984 10284 9036
rect 12716 8984 12768 9036
rect 14648 9052 14700 9104
rect 17868 9052 17920 9104
rect 18512 9052 18564 9104
rect 18788 9052 18840 9104
rect 22652 9052 22704 9104
rect 16028 8984 16080 9036
rect 16304 8984 16356 9036
rect 21916 8984 21968 9036
rect 22100 8984 22152 9036
rect 30288 9052 30340 9104
rect 23204 8984 23256 9036
rect 30472 8984 30524 9036
rect 7012 8916 7064 8968
rect 15476 8916 15528 8968
rect 19524 8916 19576 8968
rect 32404 9120 32456 9172
rect 5908 8848 5960 8900
rect 10508 8848 10560 8900
rect 11796 8848 11848 8900
rect 13544 8848 13596 8900
rect 13820 8848 13872 8900
rect 35348 8916 35400 8968
rect 36544 8916 36596 8968
rect 30380 8848 30432 8900
rect 38936 8848 38988 8900
rect 5816 8780 5868 8832
rect 12992 8780 13044 8832
rect 13268 8780 13320 8832
rect 19340 8780 19392 8832
rect 21916 8780 21968 8832
rect 26608 8780 26660 8832
rect 26976 8780 27028 8832
rect 28264 8780 28316 8832
rect 28632 8780 28684 8832
rect 30656 8780 30708 8832
rect 33048 8780 33100 8832
rect 33784 8780 33836 8832
rect 33876 8780 33928 8832
rect 34336 8780 34388 8832
rect 34520 8780 34572 8832
rect 37004 8780 37056 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 39010 8678 39062 8730
rect 39074 8678 39126 8730
rect 39138 8678 39190 8730
rect 39202 8678 39254 8730
rect 39266 8678 39318 8730
rect 3792 8576 3844 8628
rect 4344 8576 4396 8628
rect 4896 8576 4948 8628
rect 1308 8508 1360 8560
rect 6276 8576 6328 8628
rect 480 8440 532 8492
rect 3608 8483 3660 8492
rect 3608 8449 3617 8483
rect 3617 8449 3651 8483
rect 3651 8449 3660 8483
rect 3608 8440 3660 8449
rect 6000 8508 6052 8560
rect 6644 8576 6696 8628
rect 8852 8576 8904 8628
rect 9680 8576 9732 8628
rect 7288 8508 7340 8560
rect 8484 8508 8536 8560
rect 4528 8440 4580 8492
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 5632 8440 5684 8492
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 6184 8483 6236 8492
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 6184 8440 6236 8449
rect 6644 8483 6696 8492
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 6644 8440 6696 8449
rect 7012 8483 7064 8492
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 7380 8483 7432 8492
rect 7380 8449 7389 8483
rect 7389 8449 7423 8483
rect 7423 8449 7432 8483
rect 7380 8440 7432 8449
rect 7840 8440 7892 8492
rect 9220 8440 9272 8492
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 9680 8440 9732 8492
rect 756 8372 808 8424
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 4804 8372 4856 8424
rect 3792 8304 3844 8356
rect 5448 8304 5500 8356
rect 6828 8372 6880 8424
rect 7196 8372 7248 8424
rect 9956 8576 10008 8628
rect 10048 8619 10100 8628
rect 10048 8585 10057 8619
rect 10057 8585 10091 8619
rect 10091 8585 10100 8619
rect 10048 8576 10100 8585
rect 10876 8619 10928 8628
rect 10876 8585 10885 8619
rect 10885 8585 10919 8619
rect 10919 8585 10928 8619
rect 10876 8576 10928 8585
rect 12072 8576 12124 8628
rect 12164 8619 12216 8628
rect 12164 8585 12173 8619
rect 12173 8585 12207 8619
rect 12207 8585 12216 8619
rect 12164 8576 12216 8585
rect 12808 8619 12860 8628
rect 12808 8585 12817 8619
rect 12817 8585 12851 8619
rect 12851 8585 12860 8619
rect 12808 8576 12860 8585
rect 13176 8619 13228 8628
rect 13176 8585 13185 8619
rect 13185 8585 13219 8619
rect 13219 8585 13228 8619
rect 13176 8576 13228 8585
rect 14556 8576 14608 8628
rect 14648 8576 14700 8628
rect 11244 8508 11296 8560
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 10324 8483 10376 8492
rect 10324 8449 10333 8483
rect 10333 8449 10367 8483
rect 10367 8449 10376 8483
rect 10324 8440 10376 8449
rect 10508 8440 10560 8492
rect 11336 8483 11388 8492
rect 11336 8449 11345 8483
rect 11345 8449 11379 8483
rect 11379 8449 11388 8483
rect 11336 8440 11388 8449
rect 13084 8508 13136 8560
rect 13544 8508 13596 8560
rect 14924 8619 14976 8628
rect 14924 8585 14933 8619
rect 14933 8585 14967 8619
rect 14967 8585 14976 8619
rect 14924 8576 14976 8585
rect 16212 8576 16264 8628
rect 16396 8619 16448 8628
rect 16396 8585 16405 8619
rect 16405 8585 16439 8619
rect 16439 8585 16448 8619
rect 16396 8576 16448 8585
rect 17316 8576 17368 8628
rect 17684 8576 17736 8628
rect 7472 8236 7524 8288
rect 8208 8236 8260 8288
rect 8484 8279 8536 8288
rect 8484 8245 8493 8279
rect 8493 8245 8527 8279
rect 8527 8245 8536 8279
rect 8484 8236 8536 8245
rect 8944 8236 8996 8288
rect 11244 8372 11296 8424
rect 12256 8440 12308 8492
rect 13268 8440 13320 8492
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13360 8440 13412 8449
rect 13636 8483 13688 8492
rect 13636 8449 13645 8483
rect 13645 8449 13679 8483
rect 13679 8449 13688 8483
rect 13636 8440 13688 8449
rect 14280 8483 14332 8492
rect 14280 8449 14289 8483
rect 14289 8449 14323 8483
rect 14323 8449 14332 8483
rect 14280 8440 14332 8449
rect 15844 8508 15896 8560
rect 12440 8372 12492 8424
rect 13176 8372 13228 8424
rect 13544 8372 13596 8424
rect 14372 8372 14424 8424
rect 15752 8483 15804 8492
rect 15752 8449 15761 8483
rect 15761 8449 15795 8483
rect 15795 8449 15804 8483
rect 15752 8440 15804 8449
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 17500 8508 17552 8560
rect 19708 8576 19760 8628
rect 21180 8576 21232 8628
rect 21548 8576 21600 8628
rect 22008 8576 22060 8628
rect 17776 8440 17828 8492
rect 21640 8508 21692 8560
rect 21732 8508 21784 8560
rect 18144 8483 18196 8492
rect 18144 8449 18153 8483
rect 18153 8449 18187 8483
rect 18187 8449 18196 8483
rect 18144 8440 18196 8449
rect 18696 8440 18748 8492
rect 15384 8372 15436 8424
rect 11520 8304 11572 8356
rect 11704 8347 11756 8356
rect 11704 8313 11713 8347
rect 11713 8313 11747 8347
rect 11747 8313 11756 8347
rect 11704 8304 11756 8313
rect 13728 8304 13780 8356
rect 14096 8347 14148 8356
rect 14096 8313 14105 8347
rect 14105 8313 14139 8347
rect 14139 8313 14148 8347
rect 14096 8304 14148 8313
rect 14740 8304 14792 8356
rect 14924 8304 14976 8356
rect 10692 8236 10744 8288
rect 11336 8236 11388 8288
rect 13544 8236 13596 8288
rect 13636 8236 13688 8288
rect 15292 8236 15344 8288
rect 16488 8372 16540 8424
rect 17592 8372 17644 8424
rect 16764 8304 16816 8356
rect 20536 8440 20588 8492
rect 21364 8440 21416 8492
rect 21548 8440 21600 8492
rect 22560 8576 22612 8628
rect 22468 8508 22520 8560
rect 18788 8236 18840 8288
rect 20076 8372 20128 8424
rect 20628 8304 20680 8356
rect 20352 8279 20404 8288
rect 20352 8245 20361 8279
rect 20361 8245 20395 8279
rect 20395 8245 20404 8279
rect 20352 8236 20404 8245
rect 20444 8236 20496 8288
rect 20996 8372 21048 8424
rect 23112 8440 23164 8492
rect 24400 8619 24452 8628
rect 24400 8585 24409 8619
rect 24409 8585 24443 8619
rect 24443 8585 24452 8619
rect 24400 8576 24452 8585
rect 24860 8619 24912 8628
rect 24860 8585 24869 8619
rect 24869 8585 24903 8619
rect 24903 8585 24912 8619
rect 24860 8576 24912 8585
rect 25780 8619 25832 8628
rect 25780 8585 25789 8619
rect 25789 8585 25823 8619
rect 25823 8585 25832 8619
rect 25780 8576 25832 8585
rect 26516 8576 26568 8628
rect 27160 8576 27212 8628
rect 27528 8576 27580 8628
rect 24492 8508 24544 8560
rect 24676 8483 24728 8492
rect 24676 8449 24685 8483
rect 24685 8449 24719 8483
rect 24719 8449 24728 8483
rect 24676 8440 24728 8449
rect 25136 8483 25188 8492
rect 25136 8449 25145 8483
rect 25145 8449 25179 8483
rect 25179 8449 25188 8483
rect 25136 8440 25188 8449
rect 25412 8483 25464 8492
rect 25412 8449 25421 8483
rect 25421 8449 25455 8483
rect 25455 8449 25464 8483
rect 25412 8440 25464 8449
rect 26148 8508 26200 8560
rect 23296 8372 23348 8424
rect 23572 8415 23624 8424
rect 23572 8381 23581 8415
rect 23581 8381 23615 8415
rect 23615 8381 23624 8415
rect 23572 8372 23624 8381
rect 23664 8372 23716 8424
rect 26240 8483 26292 8492
rect 26240 8449 26249 8483
rect 26249 8449 26283 8483
rect 26283 8449 26292 8483
rect 26240 8440 26292 8449
rect 26332 8483 26384 8492
rect 26332 8449 26341 8483
rect 26341 8449 26375 8483
rect 26375 8449 26384 8483
rect 26332 8440 26384 8449
rect 26792 8483 26844 8492
rect 26792 8449 26801 8483
rect 26801 8449 26835 8483
rect 26835 8449 26844 8483
rect 26792 8440 26844 8449
rect 25780 8372 25832 8424
rect 27068 8440 27120 8492
rect 27160 8483 27212 8492
rect 27160 8449 27169 8483
rect 27169 8449 27203 8483
rect 27203 8449 27212 8483
rect 27160 8440 27212 8449
rect 27344 8508 27396 8560
rect 27436 8483 27488 8492
rect 27436 8449 27445 8483
rect 27445 8449 27479 8483
rect 27479 8449 27488 8483
rect 27436 8440 27488 8449
rect 21916 8304 21968 8356
rect 22100 8304 22152 8356
rect 22376 8304 22428 8356
rect 22652 8347 22704 8356
rect 22652 8313 22661 8347
rect 22661 8313 22695 8347
rect 22695 8313 22704 8347
rect 22652 8304 22704 8313
rect 22836 8304 22888 8356
rect 22008 8236 22060 8288
rect 23848 8279 23900 8288
rect 23848 8245 23857 8279
rect 23857 8245 23891 8279
rect 23891 8245 23900 8279
rect 23848 8236 23900 8245
rect 24768 8236 24820 8288
rect 26424 8304 26476 8356
rect 28264 8483 28316 8492
rect 28264 8449 28273 8483
rect 28273 8449 28307 8483
rect 28307 8449 28316 8483
rect 28264 8440 28316 8449
rect 29000 8576 29052 8628
rect 29736 8576 29788 8628
rect 28908 8508 28960 8560
rect 29460 8508 29512 8560
rect 27804 8372 27856 8424
rect 29828 8483 29880 8492
rect 29828 8449 29837 8483
rect 29837 8449 29871 8483
rect 29871 8449 29880 8483
rect 29828 8440 29880 8449
rect 30656 8483 30708 8492
rect 30656 8449 30665 8483
rect 30665 8449 30699 8483
rect 30699 8449 30708 8483
rect 30656 8440 30708 8449
rect 30932 8483 30984 8492
rect 30932 8449 30941 8483
rect 30941 8449 30975 8483
rect 30975 8449 30984 8483
rect 30932 8440 30984 8449
rect 31944 8576 31996 8628
rect 32496 8576 32548 8628
rect 33784 8576 33836 8628
rect 34152 8576 34204 8628
rect 31668 8508 31720 8560
rect 31576 8440 31628 8492
rect 29184 8372 29236 8424
rect 27712 8347 27764 8356
rect 27712 8313 27721 8347
rect 27721 8313 27755 8347
rect 27755 8313 27764 8347
rect 27712 8304 27764 8313
rect 28080 8347 28132 8356
rect 28080 8313 28089 8347
rect 28089 8313 28123 8347
rect 28123 8313 28132 8347
rect 28080 8304 28132 8313
rect 31300 8372 31352 8424
rect 31392 8372 31444 8424
rect 33784 8440 33836 8492
rect 34520 8508 34572 8560
rect 29920 8304 29972 8356
rect 31208 8304 31260 8356
rect 33416 8372 33468 8424
rect 32772 8304 32824 8356
rect 34520 8372 34572 8424
rect 34704 8576 34756 8628
rect 35808 8576 35860 8628
rect 36912 8576 36964 8628
rect 37096 8508 37148 8560
rect 37464 8508 37516 8560
rect 38936 8576 38988 8628
rect 35348 8483 35400 8492
rect 35348 8449 35357 8483
rect 35357 8449 35391 8483
rect 35391 8449 35400 8483
rect 35348 8440 35400 8449
rect 35716 8483 35768 8492
rect 35716 8449 35725 8483
rect 35725 8449 35759 8483
rect 35759 8449 35768 8483
rect 35716 8440 35768 8449
rect 35808 8483 35860 8492
rect 35808 8449 35817 8483
rect 35817 8449 35851 8483
rect 35851 8449 35860 8483
rect 35808 8440 35860 8449
rect 36728 8440 36780 8492
rect 36820 8483 36872 8492
rect 36820 8449 36829 8483
rect 36829 8449 36863 8483
rect 36863 8449 36872 8483
rect 36820 8440 36872 8449
rect 37280 8483 37332 8492
rect 37280 8449 37289 8483
rect 37289 8449 37323 8483
rect 37323 8449 37332 8483
rect 37280 8440 37332 8449
rect 37832 8440 37884 8492
rect 34336 8304 34388 8356
rect 34980 8304 35032 8356
rect 35624 8372 35676 8424
rect 38568 8440 38620 8492
rect 25228 8279 25280 8288
rect 25228 8245 25237 8279
rect 25237 8245 25271 8279
rect 25271 8245 25280 8279
rect 25228 8236 25280 8245
rect 25504 8279 25556 8288
rect 25504 8245 25513 8279
rect 25513 8245 25547 8279
rect 25547 8245 25556 8279
rect 25504 8236 25556 8245
rect 26516 8279 26568 8288
rect 26516 8245 26525 8279
rect 26525 8245 26559 8279
rect 26559 8245 26568 8279
rect 26516 8236 26568 8245
rect 26608 8279 26660 8288
rect 26608 8245 26617 8279
rect 26617 8245 26651 8279
rect 26651 8245 26660 8279
rect 26608 8236 26660 8245
rect 26700 8236 26752 8288
rect 27068 8236 27120 8288
rect 27896 8236 27948 8288
rect 28724 8236 28776 8288
rect 28816 8236 28868 8288
rect 30472 8279 30524 8288
rect 30472 8245 30481 8279
rect 30481 8245 30515 8279
rect 30515 8245 30524 8279
rect 30472 8236 30524 8245
rect 30748 8279 30800 8288
rect 30748 8245 30757 8279
rect 30757 8245 30791 8279
rect 30791 8245 30800 8279
rect 30748 8236 30800 8245
rect 30932 8236 30984 8288
rect 31668 8236 31720 8288
rect 34888 8236 34940 8288
rect 35256 8304 35308 8356
rect 36360 8304 36412 8356
rect 37188 8304 37240 8356
rect 39396 8347 39448 8356
rect 39396 8313 39405 8347
rect 39405 8313 39439 8347
rect 39439 8313 39448 8347
rect 39396 8304 39448 8313
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 37950 8134 38002 8186
rect 38014 8134 38066 8186
rect 38078 8134 38130 8186
rect 38142 8134 38194 8186
rect 38206 8134 38258 8186
rect 3424 8075 3476 8084
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 3516 8032 3568 8084
rect 4068 8032 4120 8084
rect 4620 8032 4672 8084
rect 5172 8032 5224 8084
rect 5724 8032 5776 8084
rect 6552 8032 6604 8084
rect 6736 8032 6788 8084
rect 7472 8075 7524 8084
rect 7472 8041 7481 8075
rect 7481 8041 7515 8075
rect 7515 8041 7524 8075
rect 7472 8032 7524 8041
rect 2596 8007 2648 8016
rect 2596 7973 2605 8007
rect 2605 7973 2639 8007
rect 2639 7973 2648 8007
rect 2596 7964 2648 7973
rect 5080 7964 5132 8016
rect 664 7896 716 7948
rect 6828 7896 6880 7948
rect 7656 7964 7708 8016
rect 8944 8032 8996 8084
rect 10416 8032 10468 8084
rect 12348 7964 12400 8016
rect 12808 8032 12860 8084
rect 13268 8032 13320 8084
rect 13360 8032 13412 8084
rect 14096 8032 14148 8084
rect 14372 7964 14424 8016
rect 8668 7896 8720 7948
rect 8852 7896 8904 7948
rect 10232 7896 10284 7948
rect 11520 7896 11572 7948
rect 15108 7939 15160 7948
rect 15108 7905 15117 7939
rect 15117 7905 15151 7939
rect 15151 7905 15160 7939
rect 15108 7896 15160 7905
rect 15660 8032 15712 8084
rect 15660 7896 15712 7948
rect 388 7760 440 7812
rect 2780 7871 2832 7880
rect 2780 7837 2789 7871
rect 2789 7837 2823 7871
rect 2823 7837 2832 7871
rect 2780 7828 2832 7837
rect 2872 7828 2924 7880
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 3976 7828 4028 7880
rect 4896 7828 4948 7880
rect 4988 7871 5040 7880
rect 4988 7837 4997 7871
rect 4997 7837 5031 7871
rect 5031 7837 5040 7871
rect 4988 7828 5040 7837
rect 5540 7871 5592 7880
rect 5540 7837 5549 7871
rect 5549 7837 5583 7871
rect 5583 7837 5592 7871
rect 5540 7828 5592 7837
rect 6000 7871 6052 7880
rect 6000 7837 6009 7871
rect 6009 7837 6043 7871
rect 6043 7837 6052 7871
rect 6000 7828 6052 7837
rect 6368 7871 6420 7880
rect 6368 7837 6377 7871
rect 6377 7837 6411 7871
rect 6411 7837 6420 7871
rect 6368 7828 6420 7837
rect 7288 7871 7340 7880
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7288 7828 7340 7837
rect 7380 7828 7432 7880
rect 7748 7871 7800 7880
rect 7748 7837 7757 7871
rect 7757 7837 7791 7871
rect 7791 7837 7800 7871
rect 7748 7828 7800 7837
rect 8024 7871 8076 7880
rect 8024 7837 8033 7871
rect 8033 7837 8067 7871
rect 8067 7837 8076 7871
rect 8024 7828 8076 7837
rect 7564 7760 7616 7812
rect 8392 7760 8444 7812
rect 9220 7871 9272 7880
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 10692 7871 10744 7880
rect 10692 7837 10701 7871
rect 10701 7837 10735 7871
rect 10735 7837 10744 7871
rect 10692 7828 10744 7837
rect 11152 7828 11204 7880
rect 1216 7692 1268 7744
rect 1952 7692 2004 7744
rect 4436 7692 4488 7744
rect 6644 7692 6696 7744
rect 6736 7692 6788 7744
rect 8668 7692 8720 7744
rect 9956 7760 10008 7812
rect 10416 7760 10468 7812
rect 9036 7692 9088 7744
rect 11152 7692 11204 7744
rect 11428 7735 11480 7744
rect 11428 7701 11437 7735
rect 11437 7701 11471 7735
rect 11471 7701 11480 7735
rect 11428 7692 11480 7701
rect 11980 7871 12032 7880
rect 11980 7837 11989 7871
rect 11989 7837 12023 7871
rect 12023 7837 12032 7871
rect 11980 7828 12032 7837
rect 12072 7871 12124 7880
rect 12072 7837 12081 7871
rect 12081 7837 12115 7871
rect 12115 7837 12124 7871
rect 12072 7828 12124 7837
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 12256 7828 12308 7837
rect 12992 7871 13044 7880
rect 12992 7837 13001 7871
rect 13001 7837 13035 7871
rect 13035 7837 13044 7871
rect 12992 7828 13044 7837
rect 13084 7871 13136 7880
rect 13084 7837 13118 7871
rect 13118 7837 13136 7871
rect 13084 7828 13136 7837
rect 14924 7828 14976 7880
rect 16212 7828 16264 7880
rect 19432 8032 19484 8084
rect 19708 8075 19760 8084
rect 19708 8041 19717 8075
rect 19717 8041 19751 8075
rect 19751 8041 19760 8075
rect 19708 8032 19760 8041
rect 19892 8032 19944 8084
rect 20352 8032 20404 8084
rect 23112 8032 23164 8084
rect 18972 7964 19024 8016
rect 18420 7896 18472 7948
rect 18512 7871 18564 7880
rect 18512 7837 18521 7871
rect 18521 7837 18555 7871
rect 18555 7837 18564 7871
rect 18512 7828 18564 7837
rect 18972 7828 19024 7880
rect 19248 7828 19300 7880
rect 14188 7692 14240 7744
rect 14372 7692 14424 7744
rect 15200 7735 15252 7744
rect 15200 7701 15209 7735
rect 15209 7701 15243 7735
rect 15243 7701 15252 7735
rect 15200 7692 15252 7701
rect 17408 7760 17460 7812
rect 18328 7760 18380 7812
rect 19800 7828 19852 7880
rect 19892 7867 19944 7880
rect 19892 7833 19901 7867
rect 19901 7833 19935 7867
rect 19935 7833 19944 7867
rect 20536 7964 20588 8016
rect 20628 8007 20680 8016
rect 20628 7973 20637 8007
rect 20637 7973 20671 8007
rect 20671 7973 20680 8007
rect 20628 7964 20680 7973
rect 21640 7964 21692 8016
rect 22192 7964 22244 8016
rect 21548 7896 21600 7948
rect 19892 7828 19944 7833
rect 16212 7692 16264 7744
rect 16396 7692 16448 7744
rect 17224 7692 17276 7744
rect 17592 7735 17644 7744
rect 17592 7701 17601 7735
rect 17601 7701 17635 7735
rect 17635 7701 17644 7735
rect 17592 7692 17644 7701
rect 19340 7692 19392 7744
rect 20352 7828 20404 7880
rect 20904 7871 20956 7880
rect 20904 7837 20913 7871
rect 20913 7837 20947 7871
rect 20947 7837 20956 7871
rect 20904 7828 20956 7837
rect 22008 7828 22060 7880
rect 22100 7760 22152 7812
rect 22376 7760 22428 7812
rect 22560 7939 22612 7948
rect 22560 7905 22569 7939
rect 22569 7905 22603 7939
rect 22603 7905 22612 7939
rect 22560 7896 22612 7905
rect 22928 7896 22980 7948
rect 23112 7896 23164 7948
rect 30380 8032 30432 8084
rect 30472 8032 30524 8084
rect 31668 8032 31720 8084
rect 32312 8032 32364 8084
rect 33600 8032 33652 8084
rect 34428 8032 34480 8084
rect 35532 8032 35584 8084
rect 36084 8032 36136 8084
rect 36636 8032 36688 8084
rect 37280 8075 37332 8084
rect 37280 8041 37289 8075
rect 37289 8041 37323 8075
rect 37323 8041 37332 8075
rect 37280 8032 37332 8041
rect 37832 8032 37884 8084
rect 38660 8075 38712 8084
rect 38660 8041 38669 8075
rect 38669 8041 38703 8075
rect 38703 8041 38712 8075
rect 38660 8032 38712 8041
rect 24032 7964 24084 8016
rect 27436 8007 27488 8016
rect 27436 7973 27445 8007
rect 27445 7973 27479 8007
rect 27479 7973 27488 8007
rect 27436 7964 27488 7973
rect 23572 7871 23624 7880
rect 23572 7837 23581 7871
rect 23581 7837 23615 7871
rect 23615 7837 23624 7871
rect 23572 7828 23624 7837
rect 24400 7828 24452 7880
rect 24584 7871 24636 7880
rect 24584 7837 24593 7871
rect 24593 7837 24627 7871
rect 24627 7837 24636 7871
rect 24584 7828 24636 7837
rect 24860 7896 24912 7948
rect 32404 8007 32456 8016
rect 32404 7973 32413 8007
rect 32413 7973 32447 8007
rect 32447 7973 32456 8007
rect 32404 7964 32456 7973
rect 25596 7828 25648 7880
rect 26792 7828 26844 7880
rect 27160 7828 27212 7880
rect 27344 7871 27396 7880
rect 27344 7837 27353 7871
rect 27353 7837 27387 7871
rect 27387 7837 27396 7871
rect 27344 7828 27396 7837
rect 22008 7692 22060 7744
rect 22192 7692 22244 7744
rect 22836 7692 22888 7744
rect 24216 7692 24268 7744
rect 24308 7692 24360 7744
rect 25412 7692 25464 7744
rect 26332 7735 26384 7744
rect 26332 7701 26341 7735
rect 26341 7701 26375 7735
rect 26375 7701 26384 7735
rect 26332 7692 26384 7701
rect 26608 7760 26660 7812
rect 27620 7871 27672 7880
rect 27620 7837 27629 7871
rect 27629 7837 27663 7871
rect 27663 7837 27672 7871
rect 27620 7828 27672 7837
rect 29092 7871 29144 7880
rect 29092 7837 29101 7871
rect 29101 7837 29135 7871
rect 29135 7837 29144 7871
rect 29092 7828 29144 7837
rect 29368 7871 29420 7880
rect 29368 7837 29377 7871
rect 29377 7837 29411 7871
rect 29411 7837 29420 7871
rect 29368 7828 29420 7837
rect 29460 7828 29512 7880
rect 29828 7828 29880 7880
rect 31852 7896 31904 7948
rect 27804 7760 27856 7812
rect 28540 7760 28592 7812
rect 31392 7828 31444 7880
rect 31760 7828 31812 7880
rect 29000 7692 29052 7744
rect 30748 7692 30800 7744
rect 31116 7760 31168 7812
rect 32404 7828 32456 7880
rect 32680 7828 32732 7880
rect 33876 7828 33928 7880
rect 34152 7871 34204 7880
rect 34152 7837 34161 7871
rect 34161 7837 34195 7871
rect 34195 7837 34204 7871
rect 34152 7828 34204 7837
rect 35348 7964 35400 8016
rect 36084 7896 36136 7948
rect 36176 7896 36228 7948
rect 35164 7828 35216 7880
rect 35532 7828 35584 7880
rect 35900 7871 35952 7880
rect 35900 7837 35909 7871
rect 35909 7837 35943 7871
rect 35943 7837 35952 7871
rect 35900 7828 35952 7837
rect 36360 7828 36412 7880
rect 36636 7828 36688 7880
rect 37740 7964 37792 8016
rect 37372 7896 37424 7948
rect 37832 7871 37884 7880
rect 37832 7837 37841 7871
rect 37841 7837 37875 7871
rect 37875 7837 37884 7871
rect 37832 7828 37884 7837
rect 38476 7871 38528 7880
rect 38476 7837 38485 7871
rect 38485 7837 38519 7871
rect 38519 7837 38528 7871
rect 38476 7828 38528 7837
rect 38844 7871 38896 7880
rect 38844 7837 38853 7871
rect 38853 7837 38887 7871
rect 38887 7837 38896 7871
rect 38844 7828 38896 7837
rect 37464 7760 37516 7812
rect 31668 7692 31720 7744
rect 31760 7735 31812 7744
rect 31760 7701 31769 7735
rect 31769 7701 31803 7735
rect 31803 7701 31812 7735
rect 31760 7692 31812 7701
rect 31852 7735 31904 7744
rect 31852 7701 31861 7735
rect 31861 7701 31895 7735
rect 31895 7701 31904 7735
rect 31852 7692 31904 7701
rect 32128 7735 32180 7744
rect 32128 7701 32137 7735
rect 32137 7701 32171 7735
rect 32171 7701 32180 7735
rect 32128 7692 32180 7701
rect 32680 7735 32732 7744
rect 32680 7701 32689 7735
rect 32689 7701 32723 7735
rect 32723 7701 32732 7735
rect 32680 7692 32732 7701
rect 32956 7735 33008 7744
rect 32956 7701 32965 7735
rect 32965 7701 32999 7735
rect 32999 7701 33008 7735
rect 32956 7692 33008 7701
rect 34336 7735 34388 7744
rect 34336 7701 34345 7735
rect 34345 7701 34379 7735
rect 34379 7701 34388 7735
rect 34336 7692 34388 7701
rect 35624 7692 35676 7744
rect 36360 7692 36412 7744
rect 37556 7692 37608 7744
rect 38200 7692 38252 7744
rect 38936 7692 38988 7744
rect 39396 7735 39448 7744
rect 39396 7701 39405 7735
rect 39405 7701 39439 7735
rect 39439 7701 39448 7735
rect 39396 7692 39448 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 39010 7590 39062 7642
rect 39074 7590 39126 7642
rect 39138 7590 39190 7642
rect 39202 7590 39254 7642
rect 39266 7590 39318 7642
rect 5264 7488 5316 7540
rect 5356 7531 5408 7540
rect 5356 7497 5365 7531
rect 5365 7497 5399 7531
rect 5399 7497 5408 7531
rect 5356 7488 5408 7497
rect 940 7420 992 7472
rect 1952 7420 2004 7472
rect 4160 7420 4212 7472
rect 4896 7420 4948 7472
rect 6092 7420 6144 7472
rect 6736 7463 6788 7472
rect 6736 7429 6745 7463
rect 6745 7429 6779 7463
rect 6779 7429 6788 7463
rect 6736 7420 6788 7429
rect 7104 7488 7156 7540
rect 7564 7488 7616 7540
rect 9956 7488 10008 7540
rect 11336 7488 11388 7540
rect 11428 7488 11480 7540
rect 756 7352 808 7404
rect 1124 7284 1176 7336
rect 2964 7395 3016 7404
rect 2964 7361 2973 7395
rect 2973 7361 3007 7395
rect 3007 7361 3016 7395
rect 2964 7352 3016 7361
rect 5080 7284 5132 7336
rect 3608 7216 3660 7268
rect 5816 7284 5868 7336
rect 7104 7352 7156 7404
rect 6092 7327 6144 7336
rect 6092 7293 6101 7327
rect 6101 7293 6135 7327
rect 6135 7293 6144 7327
rect 6092 7284 6144 7293
rect 6460 7216 6512 7268
rect 7012 7284 7064 7336
rect 8024 7352 8076 7404
rect 11612 7420 11664 7472
rect 8668 7395 8720 7404
rect 8668 7361 8677 7395
rect 8677 7361 8711 7395
rect 8711 7361 8720 7395
rect 8668 7352 8720 7361
rect 8944 7395 8996 7404
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 9772 7352 9824 7404
rect 10140 7352 10192 7404
rect 9680 7327 9732 7336
rect 9680 7293 9689 7327
rect 9689 7293 9723 7327
rect 9723 7293 9732 7327
rect 9680 7284 9732 7293
rect 9956 7327 10008 7336
rect 9956 7293 9965 7327
rect 9965 7293 9999 7327
rect 9999 7293 10008 7327
rect 9956 7284 10008 7293
rect 7748 7216 7800 7268
rect 2872 7148 2924 7200
rect 5540 7148 5592 7200
rect 6000 7148 6052 7200
rect 7104 7148 7156 7200
rect 7380 7148 7432 7200
rect 8484 7148 8536 7200
rect 9496 7216 9548 7268
rect 9312 7148 9364 7200
rect 11336 7395 11388 7404
rect 11336 7361 11345 7395
rect 11345 7361 11379 7395
rect 11379 7361 11388 7395
rect 11336 7352 11388 7361
rect 11520 7352 11572 7404
rect 12532 7488 12584 7540
rect 12624 7488 12676 7540
rect 13452 7488 13504 7540
rect 14280 7488 14332 7540
rect 14832 7488 14884 7540
rect 15476 7488 15528 7540
rect 15936 7488 15988 7540
rect 13084 7420 13136 7472
rect 13268 7420 13320 7472
rect 15752 7420 15804 7472
rect 18052 7488 18104 7540
rect 18328 7531 18380 7540
rect 18328 7497 18337 7531
rect 18337 7497 18371 7531
rect 18371 7497 18380 7531
rect 18328 7488 18380 7497
rect 12440 7352 12492 7404
rect 12624 7352 12676 7404
rect 13820 7395 13872 7404
rect 13820 7361 13829 7395
rect 13829 7361 13863 7395
rect 13863 7361 13872 7395
rect 13820 7352 13872 7361
rect 12164 7284 12216 7336
rect 11060 7216 11112 7268
rect 12808 7284 12860 7336
rect 13268 7284 13320 7336
rect 14096 7284 14148 7336
rect 14556 7327 14608 7336
rect 14556 7293 14565 7327
rect 14565 7293 14599 7327
rect 14599 7293 14608 7327
rect 14556 7284 14608 7293
rect 15476 7395 15528 7404
rect 15476 7361 15485 7395
rect 15485 7361 15519 7395
rect 15519 7361 15528 7395
rect 15476 7352 15528 7361
rect 15568 7352 15620 7404
rect 16120 7352 16172 7404
rect 16764 7352 16816 7404
rect 17960 7420 18012 7472
rect 19524 7488 19576 7540
rect 17224 7395 17276 7404
rect 17224 7361 17233 7395
rect 17233 7361 17267 7395
rect 17267 7361 17276 7395
rect 17224 7352 17276 7361
rect 18604 7352 18656 7404
rect 18972 7420 19024 7472
rect 20444 7531 20496 7540
rect 20444 7497 20453 7531
rect 20453 7497 20487 7531
rect 20487 7497 20496 7531
rect 20444 7488 20496 7497
rect 20536 7488 20588 7540
rect 22744 7488 22796 7540
rect 23572 7488 23624 7540
rect 24584 7488 24636 7540
rect 24676 7488 24728 7540
rect 26792 7488 26844 7540
rect 30472 7488 30524 7540
rect 30564 7488 30616 7540
rect 30840 7488 30892 7540
rect 31116 7488 31168 7540
rect 31208 7531 31260 7540
rect 31208 7497 31217 7531
rect 31217 7497 31251 7531
rect 31251 7497 31260 7531
rect 31208 7488 31260 7497
rect 31484 7531 31536 7540
rect 31484 7497 31493 7531
rect 31493 7497 31527 7531
rect 31527 7497 31536 7531
rect 31484 7488 31536 7497
rect 31760 7488 31812 7540
rect 32404 7488 32456 7540
rect 32680 7488 32732 7540
rect 35808 7488 35860 7540
rect 37096 7488 37148 7540
rect 38292 7531 38344 7540
rect 38292 7497 38301 7531
rect 38301 7497 38335 7531
rect 38335 7497 38344 7531
rect 38292 7488 38344 7497
rect 38752 7488 38804 7540
rect 18880 7395 18932 7404
rect 18880 7361 18889 7395
rect 18889 7361 18923 7395
rect 18923 7361 18932 7395
rect 18880 7352 18932 7361
rect 22192 7420 22244 7472
rect 22376 7420 22428 7472
rect 16488 7284 16540 7336
rect 16856 7284 16908 7336
rect 17868 7327 17920 7336
rect 17868 7293 17877 7327
rect 17877 7293 17911 7327
rect 17911 7293 17920 7327
rect 17868 7284 17920 7293
rect 19156 7395 19208 7404
rect 19156 7361 19165 7395
rect 19165 7361 19199 7395
rect 19199 7361 19208 7395
rect 19156 7352 19208 7361
rect 19800 7352 19852 7404
rect 20720 7395 20772 7404
rect 20720 7361 20729 7395
rect 20729 7361 20763 7395
rect 20763 7361 20772 7395
rect 20720 7352 20772 7361
rect 20812 7352 20864 7404
rect 21640 7352 21692 7404
rect 23296 7352 23348 7404
rect 19064 7284 19116 7336
rect 19248 7284 19300 7336
rect 22192 7327 22244 7336
rect 22192 7293 22201 7327
rect 22201 7293 22235 7327
rect 22235 7293 22244 7327
rect 22192 7284 22244 7293
rect 23572 7327 23624 7336
rect 23572 7293 23581 7327
rect 23581 7293 23615 7327
rect 23615 7293 23624 7327
rect 23572 7284 23624 7293
rect 11428 7148 11480 7200
rect 11520 7191 11572 7200
rect 11520 7157 11529 7191
rect 11529 7157 11563 7191
rect 11563 7157 11572 7191
rect 11520 7148 11572 7157
rect 11612 7148 11664 7200
rect 12900 7148 12952 7200
rect 13360 7148 13412 7200
rect 14556 7148 14608 7200
rect 15384 7148 15436 7200
rect 17408 7148 17460 7200
rect 18236 7148 18288 7200
rect 22100 7148 22152 7200
rect 25136 7395 25188 7404
rect 25136 7361 25145 7395
rect 25145 7361 25179 7395
rect 25179 7361 25188 7395
rect 25136 7352 25188 7361
rect 25596 7352 25648 7404
rect 26792 7352 26844 7404
rect 27620 7352 27672 7404
rect 24492 7284 24544 7336
rect 28356 7352 28408 7404
rect 29000 7352 29052 7404
rect 29184 7352 29236 7404
rect 29828 7395 29880 7404
rect 29828 7361 29837 7395
rect 29837 7361 29871 7395
rect 29871 7361 29880 7395
rect 29828 7352 29880 7361
rect 30564 7395 30616 7404
rect 30564 7361 30573 7395
rect 30573 7361 30607 7395
rect 30607 7361 30616 7395
rect 30564 7352 30616 7361
rect 34152 7420 34204 7472
rect 36636 7420 36688 7472
rect 39580 7488 39632 7540
rect 27160 7148 27212 7200
rect 29184 7216 29236 7268
rect 29368 7284 29420 7336
rect 30104 7216 30156 7268
rect 30472 7284 30524 7336
rect 30748 7327 30800 7336
rect 30748 7293 30757 7327
rect 30757 7293 30791 7327
rect 30791 7293 30800 7327
rect 30748 7284 30800 7293
rect 31116 7284 31168 7336
rect 32496 7284 32548 7336
rect 34244 7352 34296 7404
rect 34888 7284 34940 7336
rect 37648 7395 37700 7404
rect 37648 7361 37657 7395
rect 37657 7361 37691 7395
rect 37691 7361 37700 7395
rect 37648 7352 37700 7361
rect 36912 7284 36964 7336
rect 38384 7352 38436 7404
rect 39488 7420 39540 7472
rect 31392 7216 31444 7268
rect 28540 7148 28592 7200
rect 28908 7148 28960 7200
rect 29368 7148 29420 7200
rect 30012 7191 30064 7200
rect 30012 7157 30021 7191
rect 30021 7157 30055 7191
rect 30055 7157 30064 7191
rect 30012 7148 30064 7157
rect 30196 7191 30248 7200
rect 30196 7157 30205 7191
rect 30205 7157 30239 7191
rect 30239 7157 30248 7191
rect 30196 7148 30248 7157
rect 30288 7148 30340 7200
rect 37464 7216 37516 7268
rect 37740 7216 37792 7268
rect 38200 7284 38252 7336
rect 40040 7216 40092 7268
rect 32680 7148 32732 7200
rect 38844 7148 38896 7200
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 37950 7046 38002 7098
rect 38014 7046 38066 7098
rect 38078 7046 38130 7098
rect 38142 7046 38194 7098
rect 38206 7046 38258 7098
rect 2872 6944 2924 6996
rect 4896 6987 4948 6996
rect 4896 6953 4905 6987
rect 4905 6953 4939 6987
rect 4939 6953 4948 6987
rect 4896 6944 4948 6953
rect 4988 6944 5040 6996
rect 7564 6876 7616 6928
rect 8668 6944 8720 6996
rect 9772 6944 9824 6996
rect 9956 6944 10008 6996
rect 11336 6944 11388 6996
rect 12624 6944 12676 6996
rect 9680 6876 9732 6928
rect 13728 6876 13780 6928
rect 15476 6944 15528 6996
rect 16028 6944 16080 6996
rect 16212 6944 16264 6996
rect 17408 6944 17460 6996
rect 17868 6944 17920 6996
rect 20720 6944 20772 6996
rect 16304 6876 16356 6928
rect 16948 6876 17000 6928
rect 6000 6808 6052 6860
rect 7012 6808 7064 6860
rect 204 6740 256 6792
rect 3884 6783 3936 6792
rect 3884 6749 3893 6783
rect 3893 6749 3927 6783
rect 3927 6749 3936 6783
rect 3884 6740 3936 6749
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 5540 6783 5592 6792
rect 5540 6749 5549 6783
rect 5549 6749 5583 6783
rect 5583 6749 5592 6783
rect 5540 6740 5592 6749
rect 6368 6740 6420 6792
rect 7932 6740 7984 6792
rect 8668 6808 8720 6860
rect 9128 6808 9180 6860
rect 8392 6740 8444 6792
rect 9036 6740 9088 6792
rect 11336 6808 11388 6860
rect 11980 6808 12032 6860
rect 9312 6740 9364 6792
rect 9588 6740 9640 6792
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 5448 6672 5500 6724
rect 1584 6604 1636 6656
rect 9496 6672 9548 6724
rect 10692 6783 10744 6792
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 11428 6783 11480 6792
rect 11428 6749 11437 6783
rect 11437 6749 11471 6783
rect 11471 6749 11480 6783
rect 11428 6740 11480 6749
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 11704 6740 11756 6792
rect 13268 6808 13320 6860
rect 14188 6808 14240 6860
rect 14740 6851 14792 6860
rect 14740 6817 14749 6851
rect 14749 6817 14783 6851
rect 14783 6817 14792 6851
rect 16856 6851 16908 6860
rect 14740 6808 14792 6817
rect 16856 6817 16865 6851
rect 16865 6817 16899 6851
rect 16899 6817 16908 6851
rect 16856 6808 16908 6817
rect 12624 6740 12676 6792
rect 13360 6740 13412 6792
rect 15476 6740 15528 6792
rect 5908 6604 5960 6656
rect 6276 6604 6328 6656
rect 7196 6604 7248 6656
rect 7564 6604 7616 6656
rect 8760 6604 8812 6656
rect 9404 6604 9456 6656
rect 11060 6672 11112 6724
rect 12256 6672 12308 6724
rect 13268 6672 13320 6724
rect 13820 6672 13872 6724
rect 14832 6715 14884 6724
rect 14832 6681 14841 6715
rect 14841 6681 14875 6715
rect 14875 6681 14884 6715
rect 14832 6672 14884 6681
rect 10784 6604 10836 6656
rect 11796 6604 11848 6656
rect 12440 6647 12492 6656
rect 12440 6613 12449 6647
rect 12449 6613 12483 6647
rect 12483 6613 12492 6647
rect 12440 6604 12492 6613
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 12532 6604 12584 6613
rect 12624 6604 12676 6656
rect 13084 6604 13136 6656
rect 13176 6604 13228 6656
rect 15660 6604 15712 6656
rect 16948 6740 17000 6792
rect 17224 6783 17276 6792
rect 17224 6749 17233 6783
rect 17233 6749 17267 6783
rect 17267 6749 17276 6783
rect 17224 6740 17276 6749
rect 17408 6851 17460 6860
rect 17408 6817 17417 6851
rect 17417 6817 17451 6851
rect 17451 6817 17460 6851
rect 17408 6808 17460 6817
rect 17868 6851 17920 6860
rect 17868 6817 17877 6851
rect 17877 6817 17911 6851
rect 17911 6817 17920 6851
rect 17868 6808 17920 6817
rect 20628 6876 20680 6928
rect 27436 6944 27488 6996
rect 18144 6783 18196 6792
rect 18144 6749 18153 6783
rect 18153 6749 18187 6783
rect 18187 6749 18196 6783
rect 18144 6740 18196 6749
rect 18420 6783 18472 6792
rect 18420 6749 18429 6783
rect 18429 6749 18463 6783
rect 18463 6749 18472 6783
rect 18420 6740 18472 6749
rect 19524 6783 19576 6792
rect 19524 6749 19533 6783
rect 19533 6749 19567 6783
rect 19567 6749 19576 6783
rect 19524 6740 19576 6749
rect 19800 6783 19852 6792
rect 19800 6749 19809 6783
rect 19809 6749 19843 6783
rect 19843 6749 19852 6783
rect 19800 6740 19852 6749
rect 20168 6740 20220 6792
rect 25412 6876 25464 6928
rect 29828 6944 29880 6996
rect 30012 6944 30064 6996
rect 28724 6876 28776 6928
rect 30288 6876 30340 6928
rect 30564 6876 30616 6928
rect 27160 6808 27212 6860
rect 21640 6740 21692 6792
rect 23756 6740 23808 6792
rect 25136 6740 25188 6792
rect 25412 6740 25464 6792
rect 21824 6672 21876 6724
rect 28724 6672 28776 6724
rect 18972 6604 19024 6656
rect 19248 6604 19300 6656
rect 20444 6604 20496 6656
rect 20904 6604 20956 6656
rect 20996 6647 21048 6656
rect 20996 6613 21005 6647
rect 21005 6613 21039 6647
rect 21039 6613 21048 6647
rect 20996 6604 21048 6613
rect 21456 6604 21508 6656
rect 25228 6604 25280 6656
rect 27528 6604 27580 6656
rect 29920 6783 29972 6792
rect 29920 6749 29929 6783
rect 29929 6749 29963 6783
rect 29963 6749 29972 6783
rect 29920 6740 29972 6749
rect 30104 6851 30156 6860
rect 30104 6817 30113 6851
rect 30113 6817 30147 6851
rect 30147 6817 30156 6851
rect 30104 6808 30156 6817
rect 30380 6808 30432 6860
rect 31760 6876 31812 6928
rect 32220 6876 32272 6928
rect 30196 6740 30248 6792
rect 31116 6740 31168 6792
rect 32588 6851 32640 6860
rect 32588 6817 32597 6851
rect 32597 6817 32631 6851
rect 32631 6817 32640 6851
rect 32588 6808 32640 6817
rect 37832 6987 37884 6996
rect 37832 6953 37841 6987
rect 37841 6953 37875 6987
rect 37875 6953 37884 6987
rect 37832 6944 37884 6953
rect 38936 6808 38988 6860
rect 32036 6740 32088 6792
rect 32772 6740 32824 6792
rect 32864 6783 32916 6792
rect 32864 6749 32873 6783
rect 32873 6749 32907 6783
rect 32907 6749 32916 6783
rect 32864 6740 32916 6749
rect 38016 6740 38068 6792
rect 30288 6604 30340 6656
rect 30380 6647 30432 6656
rect 30380 6613 30389 6647
rect 30389 6613 30423 6647
rect 30423 6613 30432 6647
rect 30380 6604 30432 6613
rect 30656 6604 30708 6656
rect 35532 6672 35584 6724
rect 37004 6672 37056 6724
rect 33508 6647 33560 6656
rect 33508 6613 33517 6647
rect 33517 6613 33551 6647
rect 33551 6613 33560 6647
rect 33508 6604 33560 6613
rect 37832 6604 37884 6656
rect 38292 6672 38344 6724
rect 38476 6604 38528 6656
rect 38752 6672 38804 6724
rect 38660 6647 38712 6656
rect 38660 6613 38669 6647
rect 38669 6613 38703 6647
rect 38703 6613 38712 6647
rect 38660 6604 38712 6613
rect 39672 6672 39724 6724
rect 39396 6647 39448 6656
rect 39396 6613 39405 6647
rect 39405 6613 39439 6647
rect 39439 6613 39448 6647
rect 39396 6604 39448 6613
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 39010 6502 39062 6554
rect 39074 6502 39126 6554
rect 39138 6502 39190 6554
rect 39202 6502 39254 6554
rect 39266 6502 39318 6554
rect 2504 6400 2556 6452
rect 3884 6400 3936 6452
rect 6460 6400 6512 6452
rect 7932 6400 7984 6452
rect 940 6332 992 6384
rect 756 6264 808 6316
rect 1860 6264 1912 6316
rect 4160 6332 4212 6384
rect 4436 6375 4488 6384
rect 4436 6341 4445 6375
rect 4445 6341 4479 6375
rect 4479 6341 4488 6375
rect 4436 6332 4488 6341
rect 4528 6264 4580 6316
rect 4896 6264 4948 6316
rect 5080 6332 5132 6384
rect 11704 6400 11756 6452
rect 11980 6443 12032 6452
rect 11980 6409 11989 6443
rect 11989 6409 12023 6443
rect 12023 6409 12032 6443
rect 11980 6400 12032 6409
rect 1676 6239 1728 6248
rect 1676 6205 1685 6239
rect 1685 6205 1719 6239
rect 1719 6205 1728 6239
rect 1676 6196 1728 6205
rect 6552 6196 6604 6248
rect 8760 6332 8812 6384
rect 12348 6332 12400 6384
rect 8668 6264 8720 6316
rect 9496 6264 9548 6316
rect 10508 6307 10560 6316
rect 10508 6273 10517 6307
rect 10517 6273 10551 6307
rect 10551 6273 10560 6307
rect 10508 6264 10560 6273
rect 13268 6332 13320 6384
rect 14372 6332 14424 6384
rect 13360 6264 13412 6316
rect 13452 6307 13504 6316
rect 13452 6273 13461 6307
rect 13461 6273 13495 6307
rect 13495 6273 13504 6307
rect 13452 6264 13504 6273
rect 13544 6264 13596 6316
rect 3884 6171 3936 6180
rect 3884 6137 3893 6171
rect 3893 6137 3927 6171
rect 3927 6137 3936 6171
rect 3884 6128 3936 6137
rect 5448 6128 5500 6180
rect 6184 6060 6236 6112
rect 6460 6128 6512 6180
rect 7656 6196 7708 6248
rect 7564 6128 7616 6180
rect 7840 6128 7892 6180
rect 9128 6239 9180 6248
rect 9128 6205 9137 6239
rect 9137 6205 9171 6239
rect 9171 6205 9180 6239
rect 9128 6196 9180 6205
rect 9772 6196 9824 6248
rect 10140 6196 10192 6248
rect 11612 6196 11664 6248
rect 12072 6196 12124 6248
rect 12348 6196 12400 6248
rect 7196 6060 7248 6112
rect 8576 6060 8628 6112
rect 9128 6060 9180 6112
rect 10140 6103 10192 6112
rect 10140 6069 10149 6103
rect 10149 6069 10183 6103
rect 10183 6069 10192 6103
rect 10140 6060 10192 6069
rect 12256 6128 12308 6180
rect 11980 6060 12032 6112
rect 14188 6171 14240 6180
rect 14188 6137 14197 6171
rect 14197 6137 14231 6171
rect 14231 6137 14240 6171
rect 14188 6128 14240 6137
rect 14372 6196 14424 6248
rect 15476 6307 15528 6316
rect 15476 6273 15485 6307
rect 15485 6273 15519 6307
rect 15519 6273 15528 6307
rect 15476 6264 15528 6273
rect 16856 6264 16908 6316
rect 17868 6400 17920 6452
rect 17224 6264 17276 6316
rect 20352 6400 20404 6452
rect 20720 6400 20772 6452
rect 23480 6443 23532 6452
rect 23480 6409 23489 6443
rect 23489 6409 23523 6443
rect 23523 6409 23532 6443
rect 23480 6400 23532 6409
rect 23940 6400 23992 6452
rect 26424 6400 26476 6452
rect 26516 6400 26568 6452
rect 27528 6400 27580 6452
rect 28448 6400 28500 6452
rect 31116 6443 31168 6452
rect 31116 6409 31125 6443
rect 31125 6409 31159 6443
rect 31159 6409 31168 6443
rect 31116 6400 31168 6409
rect 31760 6400 31812 6452
rect 32036 6400 32088 6452
rect 32404 6400 32456 6452
rect 32864 6400 32916 6452
rect 35440 6400 35492 6452
rect 36084 6400 36136 6452
rect 39856 6400 39908 6452
rect 15200 6239 15252 6248
rect 15200 6205 15209 6239
rect 15209 6205 15243 6239
rect 15243 6205 15252 6239
rect 15200 6196 15252 6205
rect 16304 6196 16356 6248
rect 16672 6239 16724 6248
rect 16672 6205 16681 6239
rect 16681 6205 16715 6239
rect 16715 6205 16724 6239
rect 16672 6196 16724 6205
rect 23848 6332 23900 6384
rect 24032 6332 24084 6384
rect 29092 6332 29144 6384
rect 18972 6264 19024 6316
rect 20168 6307 20220 6316
rect 20168 6273 20177 6307
rect 20177 6273 20211 6307
rect 20211 6273 20220 6307
rect 20168 6264 20220 6273
rect 20904 6307 20956 6316
rect 20904 6273 20913 6307
rect 20913 6273 20947 6307
rect 20947 6273 20956 6307
rect 20904 6264 20956 6273
rect 22560 6264 22612 6316
rect 14832 6128 14884 6180
rect 14924 6171 14976 6180
rect 14924 6137 14933 6171
rect 14933 6137 14967 6171
rect 14967 6137 14976 6171
rect 14924 6128 14976 6137
rect 20352 6128 20404 6180
rect 23388 6239 23440 6248
rect 23388 6205 23397 6239
rect 23397 6205 23431 6239
rect 23431 6205 23440 6239
rect 23388 6196 23440 6205
rect 23664 6196 23716 6248
rect 24492 6307 24544 6316
rect 24492 6273 24501 6307
rect 24501 6273 24535 6307
rect 24535 6273 24544 6307
rect 24492 6264 24544 6273
rect 25044 6307 25096 6316
rect 25044 6273 25053 6307
rect 25053 6273 25087 6307
rect 25087 6273 25096 6307
rect 25044 6264 25096 6273
rect 24584 6196 24636 6248
rect 20812 6128 20864 6180
rect 17868 6103 17920 6112
rect 17868 6069 17877 6103
rect 17877 6069 17911 6103
rect 17911 6069 17920 6103
rect 17868 6060 17920 6069
rect 19708 6060 19760 6112
rect 21088 6060 21140 6112
rect 22284 6060 22336 6112
rect 26792 6264 26844 6316
rect 27528 6264 27580 6316
rect 28632 6264 28684 6316
rect 29644 6307 29696 6316
rect 29644 6273 29653 6307
rect 29653 6273 29687 6307
rect 29687 6273 29696 6307
rect 29644 6264 29696 6273
rect 29920 6307 29972 6316
rect 29920 6273 29929 6307
rect 29929 6273 29963 6307
rect 29963 6273 29972 6307
rect 29920 6264 29972 6273
rect 31300 6264 31352 6316
rect 32772 6332 32824 6384
rect 25872 6196 25924 6248
rect 25964 6060 26016 6112
rect 26332 6060 26384 6112
rect 30656 6239 30708 6248
rect 30656 6205 30665 6239
rect 30665 6205 30699 6239
rect 30699 6205 30708 6239
rect 30656 6196 30708 6205
rect 30932 6196 30984 6248
rect 31116 6196 31168 6248
rect 26608 6060 26660 6112
rect 28724 6060 28776 6112
rect 29092 6060 29144 6112
rect 30196 6171 30248 6180
rect 30196 6137 30205 6171
rect 30205 6137 30239 6171
rect 30239 6137 30248 6171
rect 30196 6128 30248 6137
rect 31208 6128 31260 6180
rect 31852 6196 31904 6248
rect 32588 6264 32640 6316
rect 33508 6264 33560 6316
rect 33968 6307 34020 6316
rect 33968 6273 33977 6307
rect 33977 6273 34011 6307
rect 34011 6273 34020 6307
rect 33968 6264 34020 6273
rect 34704 6264 34756 6316
rect 35532 6332 35584 6384
rect 35992 6264 36044 6316
rect 32772 6196 32824 6248
rect 38936 6264 38988 6316
rect 32496 6128 32548 6180
rect 31852 6060 31904 6112
rect 32220 6060 32272 6112
rect 39856 6196 39908 6248
rect 38016 6128 38068 6180
rect 39580 6128 39632 6180
rect 35440 6060 35492 6112
rect 39028 6103 39080 6112
rect 39028 6069 39037 6103
rect 39037 6069 39071 6103
rect 39071 6069 39080 6103
rect 39028 6060 39080 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 37950 5958 38002 6010
rect 38014 5958 38066 6010
rect 38078 5958 38130 6010
rect 38142 5958 38194 6010
rect 38206 5958 38258 6010
rect 1584 5899 1636 5908
rect 1584 5865 1593 5899
rect 1593 5865 1627 5899
rect 1627 5865 1636 5899
rect 1584 5856 1636 5865
rect 6092 5856 6144 5908
rect 5080 5831 5132 5840
rect 5080 5797 5089 5831
rect 5089 5797 5123 5831
rect 5123 5797 5132 5831
rect 5080 5788 5132 5797
rect 1032 5720 1084 5772
rect 756 5652 808 5704
rect 572 5584 624 5636
rect 4160 5652 4212 5704
rect 4804 5695 4856 5704
rect 4804 5661 4813 5695
rect 4813 5661 4847 5695
rect 4847 5661 4856 5695
rect 4804 5652 4856 5661
rect 4896 5695 4948 5704
rect 4896 5661 4905 5695
rect 4905 5661 4939 5695
rect 4939 5661 4948 5695
rect 6276 5763 6328 5772
rect 6276 5729 6285 5763
rect 6285 5729 6319 5763
rect 6319 5729 6328 5763
rect 6276 5720 6328 5729
rect 7012 5856 7064 5908
rect 12256 5856 12308 5908
rect 12348 5856 12400 5908
rect 8484 5788 8536 5840
rect 10140 5788 10192 5840
rect 11796 5720 11848 5772
rect 11980 5763 12032 5772
rect 11980 5729 11989 5763
rect 11989 5729 12023 5763
rect 12023 5729 12032 5763
rect 11980 5720 12032 5729
rect 12716 5763 12768 5772
rect 4896 5652 4948 5661
rect 6552 5695 6604 5704
rect 6552 5661 6561 5695
rect 6561 5661 6595 5695
rect 6595 5661 6604 5695
rect 6552 5652 6604 5661
rect 7196 5652 7248 5704
rect 8484 5652 8536 5704
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 10508 5695 10560 5704
rect 10508 5661 10517 5695
rect 10517 5661 10551 5695
rect 10551 5661 10560 5695
rect 10508 5652 10560 5661
rect 7012 5584 7064 5636
rect 4160 5516 4212 5568
rect 6092 5516 6144 5568
rect 7564 5516 7616 5568
rect 7932 5516 7984 5568
rect 8760 5516 8812 5568
rect 8852 5516 8904 5568
rect 9404 5516 9456 5568
rect 9956 5516 10008 5568
rect 11152 5516 11204 5568
rect 11244 5516 11296 5568
rect 12716 5729 12725 5763
rect 12725 5729 12759 5763
rect 12759 5729 12768 5763
rect 12716 5720 12768 5729
rect 13820 5720 13872 5772
rect 12256 5652 12308 5704
rect 13912 5652 13964 5704
rect 12348 5584 12400 5636
rect 13636 5584 13688 5636
rect 14924 5856 14976 5908
rect 16672 5856 16724 5908
rect 18788 5856 18840 5908
rect 14832 5788 14884 5840
rect 20628 5788 20680 5840
rect 19800 5720 19852 5772
rect 14280 5652 14332 5704
rect 14740 5652 14792 5704
rect 15200 5652 15252 5704
rect 17040 5652 17092 5704
rect 22652 5788 22704 5840
rect 17224 5584 17276 5636
rect 11980 5516 12032 5568
rect 13176 5516 13228 5568
rect 13728 5516 13780 5568
rect 20812 5695 20864 5704
rect 20812 5661 20821 5695
rect 20821 5661 20855 5695
rect 20855 5661 20864 5695
rect 20812 5652 20864 5661
rect 21548 5652 21600 5704
rect 23572 5856 23624 5908
rect 23664 5788 23716 5840
rect 26792 5856 26844 5908
rect 23480 5720 23532 5772
rect 23756 5720 23808 5772
rect 24492 5720 24544 5772
rect 24032 5652 24084 5704
rect 25228 5652 25280 5704
rect 26332 5652 26384 5704
rect 26700 5695 26752 5704
rect 26700 5661 26709 5695
rect 26709 5661 26743 5695
rect 26743 5661 26752 5695
rect 26700 5652 26752 5661
rect 18420 5584 18472 5636
rect 21732 5584 21784 5636
rect 23112 5584 23164 5636
rect 23940 5584 23992 5636
rect 18512 5516 18564 5568
rect 27436 5720 27488 5772
rect 27712 5652 27764 5704
rect 28632 5899 28684 5908
rect 28632 5865 28641 5899
rect 28641 5865 28675 5899
rect 28675 5865 28684 5899
rect 28632 5856 28684 5865
rect 28724 5856 28776 5908
rect 30840 5856 30892 5908
rect 31576 5856 31628 5908
rect 30196 5788 30248 5840
rect 32772 5856 32824 5908
rect 35992 5899 36044 5908
rect 35992 5865 36001 5899
rect 36001 5865 36035 5899
rect 36035 5865 36044 5899
rect 35992 5856 36044 5865
rect 36452 5856 36504 5908
rect 29000 5720 29052 5772
rect 29368 5720 29420 5772
rect 29368 5584 29420 5636
rect 30288 5695 30340 5704
rect 30288 5661 30297 5695
rect 30297 5661 30331 5695
rect 30331 5661 30340 5695
rect 30288 5652 30340 5661
rect 30656 5720 30708 5772
rect 30932 5763 30984 5772
rect 30932 5729 30941 5763
rect 30941 5729 30975 5763
rect 30975 5729 30984 5763
rect 30932 5720 30984 5729
rect 31852 5720 31904 5772
rect 35440 5763 35492 5772
rect 35440 5729 35449 5763
rect 35449 5729 35483 5763
rect 35483 5729 35492 5763
rect 35440 5720 35492 5729
rect 31208 5695 31260 5704
rect 31208 5661 31217 5695
rect 31217 5661 31251 5695
rect 31251 5661 31260 5695
rect 31208 5652 31260 5661
rect 31300 5695 31352 5704
rect 31300 5661 31334 5695
rect 31334 5661 31352 5695
rect 31300 5652 31352 5661
rect 32312 5652 32364 5704
rect 32496 5652 32548 5704
rect 33416 5652 33468 5704
rect 39672 5856 39724 5908
rect 39948 5788 40000 5840
rect 27528 5516 27580 5568
rect 30472 5516 30524 5568
rect 31116 5516 31168 5568
rect 38844 5695 38896 5704
rect 38844 5661 38853 5695
rect 38853 5661 38887 5695
rect 38887 5661 38896 5695
rect 38844 5652 38896 5661
rect 38476 5584 38528 5636
rect 32680 5516 32732 5568
rect 35532 5559 35584 5568
rect 35532 5525 35541 5559
rect 35541 5525 35575 5559
rect 35575 5525 35584 5559
rect 35532 5516 35584 5525
rect 35716 5516 35768 5568
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 39010 5414 39062 5466
rect 39074 5414 39126 5466
rect 39138 5414 39190 5466
rect 39202 5414 39254 5466
rect 39266 5414 39318 5466
rect 2320 5355 2372 5364
rect 2320 5321 2329 5355
rect 2329 5321 2363 5355
rect 2363 5321 2372 5355
rect 2320 5312 2372 5321
rect 4712 5312 4764 5364
rect 940 5244 992 5296
rect 7932 5244 7984 5296
rect 388 5176 440 5228
rect 2688 5176 2740 5228
rect 2872 5176 2924 5228
rect 4528 5176 4580 5228
rect 2504 5151 2556 5160
rect 2504 5117 2513 5151
rect 2513 5117 2547 5151
rect 2547 5117 2556 5151
rect 2504 5108 2556 5117
rect 3148 5108 3200 5160
rect 3792 5108 3844 5160
rect 7012 5176 7064 5228
rect 7656 5176 7708 5228
rect 8484 5244 8536 5296
rect 9496 5312 9548 5364
rect 8852 5244 8904 5296
rect 10508 5244 10560 5296
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 3516 5015 3568 5024
rect 3516 4981 3525 5015
rect 3525 4981 3559 5015
rect 3559 4981 3568 5015
rect 3516 4972 3568 4981
rect 7288 5151 7340 5160
rect 7288 5117 7297 5151
rect 7297 5117 7331 5151
rect 7331 5117 7340 5151
rect 7288 5108 7340 5117
rect 9772 5176 9824 5228
rect 10048 5176 10100 5228
rect 11336 5312 11388 5364
rect 10692 5176 10744 5228
rect 11888 5176 11940 5228
rect 12532 5312 12584 5364
rect 13728 5312 13780 5364
rect 14372 5312 14424 5364
rect 16948 5312 17000 5364
rect 12164 5219 12216 5228
rect 12164 5185 12173 5219
rect 12173 5185 12207 5219
rect 12207 5185 12216 5219
rect 12164 5176 12216 5185
rect 13912 5176 13964 5228
rect 14740 5176 14792 5228
rect 17684 5176 17736 5228
rect 18236 5219 18288 5228
rect 18236 5185 18245 5219
rect 18245 5185 18279 5219
rect 18279 5185 18288 5219
rect 18236 5176 18288 5185
rect 18972 5219 19024 5228
rect 18972 5185 18981 5219
rect 18981 5185 19015 5219
rect 19015 5185 19024 5219
rect 18972 5176 19024 5185
rect 19248 5219 19300 5228
rect 19248 5185 19257 5219
rect 19257 5185 19291 5219
rect 19291 5185 19300 5219
rect 19248 5176 19300 5185
rect 6552 5040 6604 5092
rect 6368 4972 6420 5024
rect 7656 4972 7708 5024
rect 8852 4972 8904 5024
rect 10048 4972 10100 5024
rect 12348 5108 12400 5160
rect 13084 5108 13136 5160
rect 11428 4972 11480 5024
rect 12256 5040 12308 5092
rect 14372 5151 14424 5160
rect 14372 5117 14381 5151
rect 14381 5117 14415 5151
rect 14415 5117 14424 5151
rect 14372 5108 14424 5117
rect 15016 5108 15068 5160
rect 16948 5151 17000 5160
rect 15292 5040 15344 5092
rect 14832 4972 14884 5024
rect 16948 5117 16957 5151
rect 16957 5117 16991 5151
rect 16991 5117 17000 5151
rect 16948 5108 17000 5117
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 19432 5108 19484 5160
rect 20628 5312 20680 5364
rect 24584 5312 24636 5364
rect 27712 5312 27764 5364
rect 30932 5312 30984 5364
rect 31024 5312 31076 5364
rect 20444 5244 20496 5296
rect 21548 5176 21600 5228
rect 22560 5176 22612 5228
rect 24952 5176 25004 5228
rect 25596 5176 25648 5228
rect 22376 5151 22428 5160
rect 22376 5117 22385 5151
rect 22385 5117 22419 5151
rect 22419 5117 22428 5151
rect 22376 5108 22428 5117
rect 26056 5108 26108 5160
rect 19984 5083 20036 5092
rect 19984 5049 19993 5083
rect 19993 5049 20027 5083
rect 20027 5049 20036 5083
rect 19984 5040 20036 5049
rect 18604 4972 18656 5024
rect 19156 4972 19208 5024
rect 20904 4972 20956 5024
rect 21732 4972 21784 5024
rect 24860 5040 24912 5092
rect 23572 4972 23624 5024
rect 24124 4972 24176 5024
rect 26424 5244 26476 5296
rect 31392 5244 31444 5296
rect 31852 5312 31904 5364
rect 32680 5312 32732 5364
rect 38568 5355 38620 5364
rect 38568 5321 38577 5355
rect 38577 5321 38611 5355
rect 38611 5321 38620 5355
rect 38568 5312 38620 5321
rect 39396 5355 39448 5364
rect 39396 5321 39405 5355
rect 39405 5321 39439 5355
rect 39439 5321 39448 5355
rect 39396 5312 39448 5321
rect 32772 5244 32824 5296
rect 35256 5244 35308 5296
rect 27160 5176 27212 5228
rect 27712 5176 27764 5228
rect 28264 5176 28316 5228
rect 28080 5108 28132 5160
rect 30564 5176 30616 5228
rect 32312 5219 32364 5228
rect 32312 5185 32321 5219
rect 32321 5185 32355 5219
rect 32355 5185 32364 5219
rect 32312 5176 32364 5185
rect 35900 5176 35952 5228
rect 38752 5219 38804 5228
rect 38752 5185 38761 5219
rect 38761 5185 38795 5219
rect 38795 5185 38804 5219
rect 38752 5176 38804 5185
rect 29276 5108 29328 5160
rect 31484 5108 31536 5160
rect 32680 5108 32732 5160
rect 39672 5176 39724 5228
rect 26332 5083 26384 5092
rect 26332 5049 26341 5083
rect 26341 5049 26375 5083
rect 26375 5049 26384 5083
rect 26332 5040 26384 5049
rect 29460 4972 29512 5024
rect 31852 4972 31904 5024
rect 32312 4972 32364 5024
rect 33968 5040 34020 5092
rect 38660 5040 38712 5092
rect 35072 4972 35124 5024
rect 39028 5015 39080 5024
rect 39028 4981 39037 5015
rect 39037 4981 39071 5015
rect 39071 4981 39080 5015
rect 39028 4972 39080 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 37950 4870 38002 4922
rect 38014 4870 38066 4922
rect 38078 4870 38130 4922
rect 38142 4870 38194 4922
rect 38206 4870 38258 4922
rect 1584 4768 1636 4820
rect 1860 4700 1912 4752
rect 3424 4700 3476 4752
rect 5908 4675 5960 4684
rect 5908 4641 5917 4675
rect 5917 4641 5951 4675
rect 5951 4641 5960 4675
rect 5908 4632 5960 4641
rect 572 4564 624 4616
rect 756 4496 808 4548
rect 2780 4564 2832 4616
rect 4528 4607 4580 4616
rect 4528 4573 4537 4607
rect 4537 4573 4571 4607
rect 4571 4573 4580 4607
rect 4528 4564 4580 4573
rect 4804 4607 4856 4616
rect 4804 4573 4813 4607
rect 4813 4573 4847 4607
rect 4847 4573 4856 4607
rect 4804 4564 4856 4573
rect 2504 4496 2556 4548
rect 6000 4496 6052 4548
rect 4712 4428 4764 4480
rect 6184 4607 6236 4616
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 7012 4811 7064 4820
rect 7012 4777 7021 4811
rect 7021 4777 7055 4811
rect 7055 4777 7064 4811
rect 7012 4768 7064 4777
rect 7472 4768 7524 4820
rect 7840 4700 7892 4752
rect 9772 4768 9824 4820
rect 10600 4768 10652 4820
rect 10968 4811 11020 4820
rect 10968 4777 10977 4811
rect 10977 4777 11011 4811
rect 11011 4777 11020 4811
rect 10968 4768 11020 4777
rect 12256 4768 12308 4820
rect 8300 4700 8352 4752
rect 8760 4700 8812 4752
rect 7656 4632 7708 4684
rect 13820 4768 13872 4820
rect 13452 4700 13504 4752
rect 14188 4700 14240 4752
rect 14280 4700 14332 4752
rect 19340 4768 19392 4820
rect 19432 4768 19484 4820
rect 19984 4768 20036 4820
rect 18328 4700 18380 4752
rect 19156 4700 19208 4752
rect 19248 4700 19300 4752
rect 6736 4496 6788 4548
rect 7656 4496 7708 4548
rect 8300 4607 8352 4616
rect 8300 4573 8309 4607
rect 8309 4573 8343 4607
rect 8343 4573 8352 4607
rect 8300 4564 8352 4573
rect 9772 4496 9824 4548
rect 10692 4607 10744 4616
rect 10692 4573 10703 4607
rect 10703 4573 10737 4607
rect 10737 4573 10744 4607
rect 13636 4632 13688 4684
rect 14372 4632 14424 4684
rect 15844 4675 15896 4684
rect 15844 4641 15853 4675
rect 15853 4641 15887 4675
rect 15887 4641 15896 4675
rect 15844 4632 15896 4641
rect 21456 4768 21508 4820
rect 19892 4632 19944 4684
rect 20076 4632 20128 4684
rect 22284 4675 22336 4684
rect 22284 4641 22293 4675
rect 22293 4641 22327 4675
rect 22327 4641 22336 4675
rect 22284 4632 22336 4641
rect 22836 4700 22888 4752
rect 22468 4632 22520 4684
rect 23020 4675 23072 4684
rect 23020 4641 23029 4675
rect 23029 4641 23063 4675
rect 23063 4641 23072 4675
rect 23020 4632 23072 4641
rect 25596 4811 25648 4820
rect 25596 4777 25605 4811
rect 25605 4777 25639 4811
rect 25639 4777 25648 4811
rect 25596 4768 25648 4777
rect 29644 4768 29696 4820
rect 31484 4768 31536 4820
rect 10692 4564 10744 4573
rect 11152 4607 11204 4616
rect 11152 4573 11161 4607
rect 11161 4573 11195 4607
rect 11195 4573 11204 4607
rect 11152 4564 11204 4573
rect 12900 4607 12952 4616
rect 12900 4573 12909 4607
rect 12909 4573 12943 4607
rect 12943 4573 12952 4607
rect 12900 4564 12952 4573
rect 13728 4564 13780 4616
rect 7196 4428 7248 4480
rect 7472 4471 7524 4480
rect 7472 4437 7481 4471
rect 7481 4437 7515 4471
rect 7515 4437 7524 4471
rect 7472 4428 7524 4437
rect 10416 4428 10468 4480
rect 10508 4428 10560 4480
rect 13084 4428 13136 4480
rect 13820 4496 13872 4548
rect 14740 4496 14792 4548
rect 15476 4607 15528 4616
rect 15476 4573 15485 4607
rect 15485 4573 15519 4607
rect 15519 4573 15528 4607
rect 15476 4564 15528 4573
rect 16028 4564 16080 4616
rect 15200 4496 15252 4548
rect 17592 4564 17644 4616
rect 17684 4607 17736 4616
rect 17684 4573 17693 4607
rect 17693 4573 17727 4607
rect 17727 4573 17736 4607
rect 17684 4564 17736 4573
rect 18236 4564 18288 4616
rect 19248 4564 19300 4616
rect 19432 4564 19484 4616
rect 20260 4607 20312 4616
rect 20260 4573 20269 4607
rect 20269 4573 20303 4607
rect 20303 4573 20312 4607
rect 20260 4564 20312 4573
rect 21548 4564 21600 4616
rect 23572 4607 23624 4616
rect 23572 4573 23581 4607
rect 23581 4573 23615 4607
rect 23615 4573 23624 4607
rect 23572 4564 23624 4573
rect 16948 4496 17000 4548
rect 24492 4607 24544 4616
rect 24492 4573 24501 4607
rect 24501 4573 24535 4607
rect 24535 4573 24544 4607
rect 24492 4564 24544 4573
rect 25320 4564 25372 4616
rect 25872 4632 25924 4684
rect 26792 4632 26844 4684
rect 26424 4564 26476 4616
rect 27068 4607 27120 4616
rect 27068 4573 27077 4607
rect 27077 4573 27111 4607
rect 27111 4573 27120 4607
rect 27068 4564 27120 4573
rect 27528 4632 27580 4684
rect 29460 4632 29512 4684
rect 27436 4564 27488 4616
rect 28080 4564 28132 4616
rect 28172 4607 28224 4616
rect 28172 4573 28181 4607
rect 28181 4573 28215 4607
rect 28215 4573 28224 4607
rect 28172 4564 28224 4573
rect 29000 4607 29052 4616
rect 29000 4573 29009 4607
rect 29009 4573 29043 4607
rect 29043 4573 29052 4607
rect 29000 4564 29052 4573
rect 29276 4564 29328 4616
rect 29552 4564 29604 4616
rect 30472 4564 30524 4616
rect 32680 4768 32732 4820
rect 32312 4700 32364 4752
rect 33968 4700 34020 4752
rect 34796 4743 34848 4752
rect 34796 4709 34805 4743
rect 34805 4709 34839 4743
rect 34839 4709 34848 4743
rect 34796 4700 34848 4709
rect 34980 4700 35032 4752
rect 31760 4675 31812 4684
rect 31760 4641 31769 4675
rect 31769 4641 31803 4675
rect 31803 4641 31812 4675
rect 31760 4632 31812 4641
rect 31852 4632 31904 4684
rect 32680 4675 32732 4684
rect 32680 4641 32689 4675
rect 32689 4641 32723 4675
rect 32723 4641 32732 4675
rect 32680 4632 32732 4641
rect 32772 4675 32824 4684
rect 32772 4641 32806 4675
rect 32806 4641 32824 4675
rect 32772 4632 32824 4641
rect 18328 4428 18380 4480
rect 19248 4428 19300 4480
rect 27712 4496 27764 4548
rect 31024 4539 31076 4548
rect 31024 4505 31033 4539
rect 31033 4505 31067 4539
rect 31067 4505 31076 4539
rect 31024 4496 31076 4505
rect 31208 4539 31260 4548
rect 31208 4505 31217 4539
rect 31217 4505 31251 4539
rect 31251 4505 31260 4539
rect 31208 4496 31260 4505
rect 31852 4496 31904 4548
rect 32956 4607 33008 4616
rect 32956 4573 32965 4607
rect 32965 4573 32999 4607
rect 32999 4573 33008 4607
rect 32956 4564 33008 4573
rect 33692 4607 33744 4616
rect 33692 4573 33701 4607
rect 33701 4573 33735 4607
rect 33735 4573 33744 4607
rect 33692 4564 33744 4573
rect 34980 4607 35032 4616
rect 34980 4573 34989 4607
rect 34989 4573 35023 4607
rect 35023 4573 35032 4607
rect 34980 4564 35032 4573
rect 35900 4811 35952 4820
rect 35900 4777 35909 4811
rect 35909 4777 35943 4811
rect 35943 4777 35952 4811
rect 35900 4768 35952 4777
rect 36820 4768 36872 4820
rect 39396 4811 39448 4820
rect 39396 4777 39405 4811
rect 39405 4777 39439 4811
rect 39439 4777 39448 4811
rect 39396 4768 39448 4777
rect 36728 4700 36780 4752
rect 39948 4700 40000 4752
rect 35624 4675 35676 4684
rect 35624 4641 35633 4675
rect 35633 4641 35667 4675
rect 35667 4641 35676 4675
rect 35624 4632 35676 4641
rect 36452 4675 36504 4684
rect 36452 4641 36461 4675
rect 36461 4641 36495 4675
rect 36495 4641 36504 4675
rect 36452 4632 36504 4641
rect 37188 4632 37240 4684
rect 38476 4607 38528 4616
rect 38476 4573 38485 4607
rect 38485 4573 38519 4607
rect 38519 4573 38528 4607
rect 38476 4564 38528 4573
rect 38568 4564 38620 4616
rect 20628 4428 20680 4480
rect 20812 4428 20864 4480
rect 21456 4428 21508 4480
rect 24768 4428 24820 4480
rect 25320 4428 25372 4480
rect 26056 4428 26108 4480
rect 26240 4428 26292 4480
rect 27436 4428 27488 4480
rect 27528 4471 27580 4480
rect 27528 4437 27537 4471
rect 27537 4437 27571 4471
rect 27571 4437 27580 4471
rect 27528 4428 27580 4437
rect 29184 4471 29236 4480
rect 29184 4437 29193 4471
rect 29193 4437 29227 4471
rect 29227 4437 29236 4471
rect 29184 4428 29236 4437
rect 30564 4428 30616 4480
rect 31944 4428 31996 4480
rect 33600 4471 33652 4480
rect 33600 4437 33609 4471
rect 33609 4437 33643 4471
rect 33643 4437 33652 4471
rect 33600 4428 33652 4437
rect 35256 4496 35308 4548
rect 37280 4496 37332 4548
rect 35532 4471 35584 4480
rect 35532 4437 35541 4471
rect 35541 4437 35575 4471
rect 35575 4437 35584 4471
rect 35532 4428 35584 4437
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 39010 4326 39062 4378
rect 39074 4326 39126 4378
rect 39138 4326 39190 4378
rect 39202 4326 39254 4378
rect 39266 4326 39318 4378
rect 1952 4267 2004 4276
rect 1952 4233 1961 4267
rect 1961 4233 1995 4267
rect 1995 4233 2004 4267
rect 1952 4224 2004 4233
rect 4344 4224 4396 4276
rect 6552 4224 6604 4276
rect 7012 4224 7064 4276
rect 7288 4224 7340 4276
rect 756 4156 808 4208
rect 940 4088 992 4140
rect 2504 4020 2556 4072
rect 2320 3995 2372 4004
rect 2320 3961 2329 3995
rect 2329 3961 2363 3995
rect 2363 3961 2372 3995
rect 2320 3952 2372 3961
rect 2596 3995 2648 4004
rect 2596 3961 2605 3995
rect 2605 3961 2639 3995
rect 2639 3961 2648 3995
rect 2596 3952 2648 3961
rect 4160 4131 4212 4140
rect 4160 4097 4169 4131
rect 4169 4097 4203 4131
rect 4203 4097 4212 4131
rect 4160 4088 4212 4097
rect 4344 4131 4396 4140
rect 4344 4097 4362 4131
rect 4362 4097 4396 4131
rect 4344 4088 4396 4097
rect 4436 4131 4488 4140
rect 4436 4097 4445 4131
rect 4445 4097 4479 4131
rect 4479 4097 4488 4131
rect 4436 4088 4488 4097
rect 3148 4063 3200 4072
rect 3148 4029 3157 4063
rect 3157 4029 3191 4063
rect 3191 4029 3200 4063
rect 3148 4020 3200 4029
rect 3516 4020 3568 4072
rect 4712 4063 4764 4072
rect 4712 4029 4721 4063
rect 4721 4029 4755 4063
rect 4755 4029 4764 4063
rect 4712 4020 4764 4029
rect 5448 4020 5500 4072
rect 6736 4088 6788 4140
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 8300 4224 8352 4276
rect 6552 4063 6604 4072
rect 6552 4029 6561 4063
rect 6561 4029 6595 4063
rect 6595 4029 6604 4063
rect 6552 4020 6604 4029
rect 7012 4063 7064 4072
rect 7012 4029 7021 4063
rect 7021 4029 7055 4063
rect 7055 4029 7064 4063
rect 7012 4020 7064 4029
rect 6920 3952 6972 4004
rect 2872 3884 2924 3936
rect 3792 3884 3844 3936
rect 3976 3884 4028 3936
rect 7288 3884 7340 3936
rect 7656 3884 7708 3936
rect 8760 4020 8812 4072
rect 10416 4088 10468 4140
rect 8024 3952 8076 4004
rect 8852 3952 8904 4004
rect 9312 4063 9364 4072
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 9312 4020 9364 4029
rect 9496 4063 9548 4072
rect 9496 4029 9505 4063
rect 9505 4029 9539 4063
rect 9539 4029 9548 4063
rect 9496 4020 9548 4029
rect 9680 4020 9732 4072
rect 10508 4063 10560 4072
rect 10508 4029 10517 4063
rect 10517 4029 10551 4063
rect 10551 4029 10560 4063
rect 10508 4020 10560 4029
rect 11152 4267 11204 4276
rect 11152 4233 11161 4267
rect 11161 4233 11195 4267
rect 11195 4233 11204 4267
rect 11152 4224 11204 4233
rect 11428 4224 11480 4276
rect 13084 4224 13136 4276
rect 17224 4224 17276 4276
rect 18052 4224 18104 4276
rect 13636 4156 13688 4208
rect 11244 4088 11296 4140
rect 13176 4131 13228 4140
rect 13176 4097 13185 4131
rect 13185 4097 13219 4131
rect 13219 4097 13228 4131
rect 13820 4156 13872 4208
rect 13176 4088 13228 4097
rect 14188 4131 14240 4140
rect 14188 4097 14197 4131
rect 14197 4097 14231 4131
rect 14231 4097 14240 4131
rect 14188 4088 14240 4097
rect 14372 4156 14424 4208
rect 15568 4156 15620 4208
rect 16856 4156 16908 4208
rect 18972 4156 19024 4208
rect 19432 4224 19484 4276
rect 19708 4224 19760 4276
rect 20260 4224 20312 4276
rect 21824 4224 21876 4276
rect 23020 4224 23072 4276
rect 19984 4156 20036 4208
rect 15476 4088 15528 4140
rect 15752 4088 15804 4140
rect 17960 4088 18012 4140
rect 9312 3884 9364 3936
rect 9772 3884 9824 3936
rect 10968 3952 11020 4004
rect 12624 3952 12676 4004
rect 12992 3952 13044 4004
rect 13728 3952 13780 4004
rect 13268 3884 13320 3936
rect 13360 3927 13412 3936
rect 13360 3893 13369 3927
rect 13369 3893 13403 3927
rect 13403 3893 13412 3927
rect 13360 3884 13412 3893
rect 13452 3884 13504 3936
rect 17224 4020 17276 4072
rect 18604 3952 18656 4004
rect 19156 4131 19208 4140
rect 19156 4097 19165 4131
rect 19165 4097 19199 4131
rect 19199 4097 19208 4131
rect 19156 4088 19208 4097
rect 19248 4063 19300 4072
rect 19248 4029 19257 4063
rect 19257 4029 19291 4063
rect 19291 4029 19300 4063
rect 19248 4020 19300 4029
rect 19340 4020 19392 4072
rect 19892 4020 19944 4072
rect 20628 3995 20680 4004
rect 20628 3961 20637 3995
rect 20637 3961 20671 3995
rect 20671 3961 20680 3995
rect 20628 3952 20680 3961
rect 22560 4131 22612 4140
rect 22560 4097 22569 4131
rect 22569 4097 22603 4131
rect 22603 4097 22612 4131
rect 22560 4088 22612 4097
rect 23664 4131 23716 4140
rect 23664 4097 23673 4131
rect 23673 4097 23707 4131
rect 23707 4097 23716 4131
rect 23664 4088 23716 4097
rect 25412 4267 25464 4276
rect 25412 4233 25421 4267
rect 25421 4233 25455 4267
rect 25455 4233 25464 4267
rect 25412 4224 25464 4233
rect 25872 4224 25924 4276
rect 26056 4224 26108 4276
rect 29000 4224 29052 4276
rect 31208 4224 31260 4276
rect 32864 4224 32916 4276
rect 25044 4156 25096 4208
rect 27896 4156 27948 4208
rect 30380 4199 30432 4208
rect 30380 4165 30389 4199
rect 30389 4165 30423 4199
rect 30423 4165 30432 4199
rect 30380 4156 30432 4165
rect 31760 4156 31812 4208
rect 32220 4156 32272 4208
rect 22836 4063 22888 4072
rect 22836 4029 22845 4063
rect 22845 4029 22879 4063
rect 22879 4029 22888 4063
rect 22836 4020 22888 4029
rect 26240 4088 26292 4140
rect 27436 4088 27488 4140
rect 28172 4088 28224 4140
rect 25596 4063 25648 4072
rect 25596 4029 25605 4063
rect 25605 4029 25639 4063
rect 25639 4029 25648 4063
rect 25596 4020 25648 4029
rect 30564 4088 30616 4140
rect 26332 3952 26384 4004
rect 16396 3884 16448 3936
rect 16580 3884 16632 3936
rect 19064 3884 19116 3936
rect 22192 3884 22244 3936
rect 24676 3927 24728 3936
rect 24676 3893 24685 3927
rect 24685 3893 24719 3927
rect 24719 3893 24728 3927
rect 24676 3884 24728 3893
rect 26608 3884 26660 3936
rect 30472 4020 30524 4072
rect 33692 4224 33744 4276
rect 34060 4224 34112 4276
rect 35624 4224 35676 4276
rect 36452 4224 36504 4276
rect 33508 4131 33560 4140
rect 33508 4097 33517 4131
rect 33517 4097 33551 4131
rect 33551 4097 33560 4131
rect 33508 4088 33560 4097
rect 34060 4131 34112 4140
rect 34060 4097 34069 4131
rect 34069 4097 34103 4131
rect 34103 4097 34112 4131
rect 34060 4088 34112 4097
rect 34336 4156 34388 4208
rect 38476 4156 38528 4208
rect 35256 4088 35308 4140
rect 28080 3952 28132 4004
rect 33416 4020 33468 4072
rect 34428 4020 34480 4072
rect 37556 4131 37608 4140
rect 37556 4097 37565 4131
rect 37565 4097 37599 4131
rect 37599 4097 37608 4131
rect 37556 4088 37608 4097
rect 38936 4088 38988 4140
rect 28908 3884 28960 3936
rect 31208 3884 31260 3936
rect 32772 3884 32824 3936
rect 33324 3884 33376 3936
rect 33692 3927 33744 3936
rect 33692 3893 33701 3927
rect 33701 3893 33735 3927
rect 33735 3893 33744 3927
rect 33692 3884 33744 3893
rect 33876 3884 33928 3936
rect 39488 3952 39540 4004
rect 39028 3927 39080 3936
rect 39028 3893 39037 3927
rect 39037 3893 39071 3927
rect 39071 3893 39080 3927
rect 39028 3884 39080 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 37950 3782 38002 3834
rect 38014 3782 38066 3834
rect 38078 3782 38130 3834
rect 38142 3782 38194 3834
rect 38206 3782 38258 3834
rect 2504 3680 2556 3732
rect 5632 3680 5684 3732
rect 6552 3680 6604 3732
rect 9496 3680 9548 3732
rect 2872 3544 2924 3596
rect 3148 3544 3200 3596
rect 3424 3587 3476 3596
rect 3424 3553 3433 3587
rect 3433 3553 3467 3587
rect 3467 3553 3476 3587
rect 3424 3544 3476 3553
rect 5908 3587 5960 3596
rect 5908 3553 5917 3587
rect 5917 3553 5951 3587
rect 5951 3553 5960 3587
rect 5908 3544 5960 3553
rect 6736 3587 6788 3596
rect 6736 3553 6745 3587
rect 6745 3553 6779 3587
rect 6779 3553 6788 3587
rect 6736 3544 6788 3553
rect 7196 3587 7248 3596
rect 7196 3553 7205 3587
rect 7205 3553 7239 3587
rect 7239 3553 7248 3587
rect 7196 3544 7248 3553
rect 8760 3544 8812 3596
rect 10968 3680 11020 3732
rect 9864 3587 9916 3596
rect 9864 3553 9873 3587
rect 9873 3553 9907 3587
rect 9907 3553 9916 3587
rect 9864 3544 9916 3553
rect 10140 3587 10192 3596
rect 10140 3553 10149 3587
rect 10149 3553 10183 3587
rect 10183 3553 10192 3587
rect 10140 3544 10192 3553
rect 10324 3544 10376 3596
rect 13544 3680 13596 3732
rect 17776 3680 17828 3732
rect 20260 3680 20312 3732
rect 22836 3680 22888 3732
rect 11520 3612 11572 3664
rect 12808 3612 12860 3664
rect 14556 3612 14608 3664
rect 18144 3612 18196 3664
rect 20628 3612 20680 3664
rect 22192 3612 22244 3664
rect 23020 3612 23072 3664
rect 204 3476 256 3528
rect 2320 3519 2372 3528
rect 2320 3485 2329 3519
rect 2329 3485 2363 3519
rect 2363 3485 2372 3519
rect 2320 3476 2372 3485
rect 1308 3408 1360 3460
rect 4436 3476 4488 3528
rect 2504 3383 2556 3392
rect 2504 3349 2513 3383
rect 2513 3349 2547 3383
rect 2547 3349 2556 3383
rect 2504 3340 2556 3349
rect 4344 3340 4396 3392
rect 5172 3383 5224 3392
rect 5172 3349 5181 3383
rect 5181 3349 5215 3383
rect 5215 3349 5224 3383
rect 5172 3340 5224 3349
rect 5356 3383 5408 3392
rect 5356 3349 5365 3383
rect 5365 3349 5399 3383
rect 5399 3349 5408 3383
rect 5356 3340 5408 3349
rect 5724 3519 5776 3528
rect 5724 3485 5733 3519
rect 5733 3485 5767 3519
rect 5767 3485 5776 3519
rect 5724 3476 5776 3485
rect 6920 3476 6972 3528
rect 7564 3476 7616 3528
rect 10048 3476 10100 3528
rect 11888 3519 11940 3528
rect 11888 3485 11897 3519
rect 11897 3485 11931 3519
rect 11931 3485 11940 3519
rect 11888 3476 11940 3485
rect 13544 3587 13596 3596
rect 13544 3553 13553 3587
rect 13553 3553 13587 3587
rect 13587 3553 13596 3587
rect 13544 3544 13596 3553
rect 13728 3544 13780 3596
rect 17224 3544 17276 3596
rect 18236 3544 18288 3596
rect 18604 3544 18656 3596
rect 13176 3476 13228 3528
rect 15384 3519 15436 3528
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 16580 3476 16632 3528
rect 16948 3476 17000 3528
rect 17408 3519 17460 3528
rect 17408 3485 17417 3519
rect 17417 3485 17451 3519
rect 17451 3485 17460 3519
rect 17408 3476 17460 3485
rect 17776 3519 17828 3528
rect 17776 3485 17785 3519
rect 17785 3485 17819 3519
rect 17819 3485 17828 3519
rect 17776 3476 17828 3485
rect 17868 3476 17920 3528
rect 22836 3544 22888 3596
rect 26332 3680 26384 3732
rect 28264 3612 28316 3664
rect 30472 3612 30524 3664
rect 31668 3680 31720 3732
rect 33324 3680 33376 3732
rect 33416 3680 33468 3732
rect 34428 3680 34480 3732
rect 34520 3680 34572 3732
rect 35992 3723 36044 3732
rect 35992 3689 36001 3723
rect 36001 3689 36035 3723
rect 36035 3689 36044 3723
rect 35992 3680 36044 3689
rect 39396 3723 39448 3732
rect 39396 3689 39405 3723
rect 39405 3689 39439 3723
rect 39439 3689 39448 3723
rect 39396 3680 39448 3689
rect 32036 3612 32088 3664
rect 38936 3612 38988 3664
rect 39948 3612 40000 3664
rect 29828 3544 29880 3596
rect 30748 3544 30800 3596
rect 31852 3544 31904 3596
rect 33692 3544 33744 3596
rect 38660 3544 38712 3596
rect 19708 3519 19760 3528
rect 19708 3485 19717 3519
rect 19717 3485 19751 3519
rect 19751 3485 19760 3519
rect 19708 3476 19760 3485
rect 9680 3340 9732 3392
rect 10232 3340 10284 3392
rect 10600 3340 10652 3392
rect 10968 3340 11020 3392
rect 11428 3340 11480 3392
rect 19294 3408 19346 3460
rect 22560 3476 22612 3528
rect 23572 3476 23624 3528
rect 11704 3340 11756 3392
rect 15752 3340 15804 3392
rect 16120 3383 16172 3392
rect 16120 3349 16129 3383
rect 16129 3349 16163 3383
rect 16163 3349 16172 3383
rect 16120 3340 16172 3349
rect 16488 3340 16540 3392
rect 19156 3340 19208 3392
rect 20628 3408 20680 3460
rect 22192 3408 22244 3460
rect 22376 3408 22428 3460
rect 26148 3476 26200 3528
rect 25872 3408 25924 3460
rect 26332 3476 26384 3528
rect 27436 3476 27488 3528
rect 27620 3476 27672 3528
rect 30288 3476 30340 3528
rect 30932 3519 30984 3528
rect 30932 3485 30941 3519
rect 30941 3485 30975 3519
rect 30975 3485 30984 3519
rect 30932 3476 30984 3485
rect 31208 3519 31260 3528
rect 31208 3485 31217 3519
rect 31217 3485 31251 3519
rect 31251 3485 31260 3519
rect 31208 3476 31260 3485
rect 31760 3476 31812 3528
rect 33324 3476 33376 3528
rect 34704 3476 34756 3528
rect 34980 3519 35032 3528
rect 34980 3485 34989 3519
rect 34989 3485 35023 3519
rect 35023 3485 35032 3519
rect 34980 3476 35032 3485
rect 29000 3451 29052 3460
rect 29000 3417 29009 3451
rect 29009 3417 29043 3451
rect 29043 3417 29052 3451
rect 29000 3408 29052 3417
rect 29276 3408 29328 3460
rect 22652 3340 22704 3392
rect 22744 3383 22796 3392
rect 22744 3349 22753 3383
rect 22753 3349 22787 3383
rect 22787 3349 22796 3383
rect 22744 3340 22796 3349
rect 23020 3340 23072 3392
rect 27344 3340 27396 3392
rect 28264 3383 28316 3392
rect 28264 3349 28273 3383
rect 28273 3349 28307 3383
rect 28307 3349 28316 3383
rect 28264 3340 28316 3349
rect 29184 3340 29236 3392
rect 33692 3408 33744 3460
rect 38844 3519 38896 3528
rect 38844 3485 38853 3519
rect 38853 3485 38887 3519
rect 38887 3485 38896 3519
rect 38844 3476 38896 3485
rect 36268 3408 36320 3460
rect 33416 3340 33468 3392
rect 33876 3340 33928 3392
rect 34152 3340 34204 3392
rect 34980 3340 35032 3392
rect 38384 3340 38436 3392
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 39010 3238 39062 3290
rect 39074 3238 39126 3290
rect 39138 3238 39190 3290
rect 39202 3238 39254 3290
rect 39266 3238 39318 3290
rect 3976 3136 4028 3188
rect 4344 3179 4396 3188
rect 4344 3145 4353 3179
rect 4353 3145 4387 3179
rect 4387 3145 4396 3179
rect 4344 3136 4396 3145
rect 1860 3068 1912 3120
rect 1216 3000 1268 3052
rect 2780 3000 2832 3052
rect 5356 3068 5408 3120
rect 6736 3136 6788 3188
rect 8392 3068 8444 3120
rect 388 2932 440 2984
rect 2688 2932 2740 2984
rect 3148 2975 3200 2984
rect 3148 2941 3157 2975
rect 3157 2941 3191 2975
rect 3191 2941 3200 2975
rect 3148 2932 3200 2941
rect 1124 2864 1176 2916
rect 3424 2907 3476 2916
rect 3424 2873 3433 2907
rect 3433 2873 3467 2907
rect 3467 2873 3476 2907
rect 3424 2864 3476 2873
rect 2504 2839 2556 2848
rect 2504 2805 2513 2839
rect 2513 2805 2547 2839
rect 2547 2805 2556 2839
rect 2504 2796 2556 2805
rect 2596 2796 2648 2848
rect 5080 3000 5132 3052
rect 6092 3000 6144 3052
rect 6276 3000 6328 3052
rect 11796 3136 11848 3188
rect 12624 3136 12676 3188
rect 17500 3136 17552 3188
rect 17776 3179 17828 3188
rect 17776 3145 17785 3179
rect 17785 3145 17819 3179
rect 17819 3145 17828 3179
rect 17776 3136 17828 3145
rect 18144 3179 18196 3188
rect 18144 3145 18153 3179
rect 18153 3145 18187 3179
rect 18187 3145 18196 3179
rect 18144 3136 18196 3145
rect 18236 3136 18288 3188
rect 20260 3136 20312 3188
rect 20352 3136 20404 3188
rect 23112 3179 23164 3188
rect 23112 3145 23121 3179
rect 23121 3145 23155 3179
rect 23155 3145 23164 3179
rect 23112 3136 23164 3145
rect 25596 3136 25648 3188
rect 26332 3179 26384 3188
rect 26332 3145 26341 3179
rect 26341 3145 26375 3179
rect 26375 3145 26384 3179
rect 26332 3136 26384 3145
rect 27712 3136 27764 3188
rect 11428 3068 11480 3120
rect 13268 3068 13320 3120
rect 21824 3068 21876 3120
rect 29276 3136 29328 3188
rect 30932 3136 30984 3188
rect 31300 3179 31352 3188
rect 31300 3145 31309 3179
rect 31309 3145 31343 3179
rect 31343 3145 31352 3179
rect 31300 3136 31352 3145
rect 33784 3136 33836 3188
rect 36544 3136 36596 3188
rect 39396 3179 39448 3188
rect 39396 3145 39405 3179
rect 39405 3145 39439 3179
rect 39439 3145 39448 3179
rect 39396 3136 39448 3145
rect 9864 3000 9916 3052
rect 10600 3000 10652 3052
rect 10692 3043 10744 3052
rect 10692 3009 10701 3043
rect 10701 3009 10735 3043
rect 10735 3009 10744 3043
rect 10692 3000 10744 3009
rect 12900 3000 12952 3052
rect 4804 2932 4856 2984
rect 4896 2975 4948 2984
rect 4896 2941 4905 2975
rect 4905 2941 4939 2975
rect 4939 2941 4948 2975
rect 4896 2932 4948 2941
rect 6368 2932 6420 2984
rect 9588 2932 9640 2984
rect 11796 2932 11848 2984
rect 13544 2932 13596 2984
rect 4160 2796 4212 2848
rect 4712 2796 4764 2848
rect 6552 2796 6604 2848
rect 7472 2796 7524 2848
rect 9772 2796 9824 2848
rect 10048 2796 10100 2848
rect 11336 2839 11388 2848
rect 11336 2805 11345 2839
rect 11345 2805 11379 2839
rect 11379 2805 11388 2839
rect 11336 2796 11388 2805
rect 14464 2864 14516 2916
rect 13728 2796 13780 2848
rect 15384 2932 15436 2984
rect 16028 3043 16080 3052
rect 16028 3009 16037 3043
rect 16037 3009 16071 3043
rect 16071 3009 16080 3043
rect 16028 3000 16080 3009
rect 16580 3000 16632 3052
rect 16948 3043 17000 3052
rect 16948 3009 16957 3043
rect 16957 3009 16991 3043
rect 16991 3009 17000 3043
rect 16948 3000 17000 3009
rect 16672 2975 16724 2984
rect 16672 2941 16681 2975
rect 16681 2941 16715 2975
rect 16715 2941 16724 2975
rect 16672 2932 16724 2941
rect 17500 2932 17552 2984
rect 14924 2796 14976 2848
rect 19432 3043 19484 3052
rect 19432 3009 19441 3043
rect 19441 3009 19475 3043
rect 19475 3009 19484 3043
rect 19432 3000 19484 3009
rect 22560 3043 22612 3052
rect 22560 3009 22569 3043
rect 22569 3009 22603 3043
rect 22603 3009 22612 3043
rect 22560 3000 22612 3009
rect 22836 3043 22888 3052
rect 22836 3009 22845 3043
rect 22845 3009 22879 3043
rect 22879 3009 22888 3043
rect 22836 3000 22888 3009
rect 19524 2932 19576 2984
rect 17592 2796 17644 2848
rect 19616 2839 19668 2848
rect 19616 2805 19625 2839
rect 19625 2805 19659 2839
rect 19659 2805 19668 2839
rect 19616 2796 19668 2805
rect 21824 2839 21876 2848
rect 21824 2805 21833 2839
rect 21833 2805 21867 2839
rect 21867 2805 21876 2839
rect 21824 2796 21876 2805
rect 23664 3000 23716 3052
rect 25044 3043 25096 3052
rect 25044 3009 25053 3043
rect 25053 3009 25087 3043
rect 25087 3009 25096 3043
rect 25872 3043 25924 3052
rect 25044 3000 25096 3009
rect 25872 3009 25881 3043
rect 25881 3009 25915 3043
rect 25915 3009 25924 3043
rect 25872 3000 25924 3009
rect 28264 3068 28316 3120
rect 24492 2932 24544 2984
rect 27436 3043 27488 3052
rect 27436 3009 27445 3043
rect 27445 3009 27479 3043
rect 27479 3009 27488 3043
rect 27436 3000 27488 3009
rect 29552 3000 29604 3052
rect 30840 3043 30892 3052
rect 30840 3009 30849 3043
rect 30849 3009 30883 3043
rect 30883 3009 30892 3043
rect 30840 3000 30892 3009
rect 26240 2932 26292 2984
rect 30748 2932 30800 2984
rect 31484 3043 31536 3052
rect 31484 3009 31493 3043
rect 31493 3009 31527 3043
rect 31527 3009 31536 3043
rect 31484 3000 31536 3009
rect 33784 3000 33836 3052
rect 34428 3000 34480 3052
rect 38384 3043 38436 3052
rect 38384 3009 38393 3043
rect 38393 3009 38427 3043
rect 38427 3009 38436 3043
rect 38384 3000 38436 3009
rect 38660 3000 38712 3052
rect 38936 3000 38988 3052
rect 30472 2839 30524 2848
rect 30472 2805 30481 2839
rect 30481 2805 30515 2839
rect 30515 2805 30524 2839
rect 30472 2796 30524 2805
rect 32956 2839 33008 2848
rect 32956 2805 32965 2839
rect 32965 2805 32999 2839
rect 32999 2805 33008 2839
rect 32956 2796 33008 2805
rect 38660 2839 38712 2848
rect 38660 2805 38669 2839
rect 38669 2805 38703 2839
rect 38703 2805 38712 2839
rect 38660 2796 38712 2805
rect 39028 2839 39080 2848
rect 39028 2805 39037 2839
rect 39037 2805 39071 2839
rect 39071 2805 39080 2839
rect 39028 2796 39080 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 37950 2694 38002 2746
rect 38014 2694 38066 2746
rect 38078 2694 38130 2746
rect 38142 2694 38194 2746
rect 38206 2694 38258 2746
rect 1216 2456 1268 2508
rect 4804 2592 4856 2644
rect 5908 2635 5960 2644
rect 5908 2601 5917 2635
rect 5917 2601 5951 2635
rect 5951 2601 5960 2635
rect 5908 2592 5960 2601
rect 10232 2592 10284 2644
rect 11888 2592 11940 2644
rect 12808 2592 12860 2644
rect 12992 2592 13044 2644
rect 16856 2592 16908 2644
rect 17408 2592 17460 2644
rect 4160 2524 4212 2576
rect 4712 2524 4764 2576
rect 5724 2524 5776 2576
rect 4252 2456 4304 2508
rect 4896 2499 4948 2508
rect 4896 2465 4905 2499
rect 4905 2465 4939 2499
rect 4939 2465 4948 2499
rect 4896 2456 4948 2465
rect 6184 2456 6236 2508
rect 1308 2388 1360 2440
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 3516 2388 3568 2440
rect 4712 2388 4764 2440
rect 5816 2320 5868 2372
rect 6368 2388 6420 2440
rect 9864 2524 9916 2576
rect 11060 2524 11112 2576
rect 9772 2456 9824 2508
rect 16120 2524 16172 2576
rect 16580 2524 16632 2576
rect 11336 2456 11388 2508
rect 6276 2320 6328 2372
rect 6644 2363 6696 2372
rect 6644 2329 6653 2363
rect 6653 2329 6687 2363
rect 6687 2329 6696 2363
rect 6644 2320 6696 2329
rect 7012 2363 7064 2372
rect 7012 2329 7021 2363
rect 7021 2329 7055 2363
rect 7055 2329 7064 2363
rect 7012 2320 7064 2329
rect 7288 2388 7340 2440
rect 7932 2388 7984 2440
rect 9404 2388 9456 2440
rect 10140 2388 10192 2440
rect 10876 2388 10928 2440
rect 11060 2388 11112 2440
rect 11704 2388 11756 2440
rect 12348 2388 12400 2440
rect 17500 2499 17552 2508
rect 17500 2465 17509 2499
rect 17509 2465 17543 2499
rect 17543 2465 17552 2499
rect 17500 2456 17552 2465
rect 21824 2592 21876 2644
rect 22284 2592 22336 2644
rect 22652 2592 22704 2644
rect 22928 2524 22980 2576
rect 23296 2567 23348 2576
rect 23296 2533 23305 2567
rect 23305 2533 23339 2567
rect 23339 2533 23348 2567
rect 23296 2524 23348 2533
rect 23388 2524 23440 2576
rect 7564 2320 7616 2372
rect 8668 2320 8720 2372
rect 9220 2363 9272 2372
rect 9220 2329 9229 2363
rect 9229 2329 9263 2363
rect 9263 2329 9272 2363
rect 9220 2320 9272 2329
rect 3700 2252 3752 2304
rect 6184 2295 6236 2304
rect 6184 2261 6193 2295
rect 6193 2261 6227 2295
rect 6227 2261 6236 2295
rect 6184 2252 6236 2261
rect 7656 2295 7708 2304
rect 7656 2261 7665 2295
rect 7665 2261 7699 2295
rect 7699 2261 7708 2295
rect 7656 2252 7708 2261
rect 8208 2295 8260 2304
rect 8208 2261 8217 2295
rect 8217 2261 8251 2295
rect 8251 2261 8260 2295
rect 8208 2252 8260 2261
rect 9680 2295 9732 2304
rect 9680 2261 9689 2295
rect 9689 2261 9723 2295
rect 9723 2261 9732 2295
rect 9680 2252 9732 2261
rect 10324 2252 10376 2304
rect 11612 2320 11664 2372
rect 11980 2363 12032 2372
rect 11980 2329 11989 2363
rect 11989 2329 12023 2363
rect 12023 2329 12032 2363
rect 11980 2320 12032 2329
rect 14924 2431 14976 2440
rect 14924 2397 14933 2431
rect 14933 2397 14967 2431
rect 14967 2397 14976 2431
rect 14924 2388 14976 2397
rect 15660 2431 15712 2440
rect 15660 2397 15669 2431
rect 15669 2397 15703 2431
rect 15703 2397 15712 2431
rect 15660 2388 15712 2397
rect 15752 2388 15804 2440
rect 16212 2388 16264 2440
rect 18144 2431 18196 2440
rect 18144 2397 18153 2431
rect 18153 2397 18187 2431
rect 18187 2397 18196 2431
rect 18144 2388 18196 2397
rect 17132 2320 17184 2372
rect 22744 2456 22796 2508
rect 18788 2388 18840 2440
rect 19432 2388 19484 2440
rect 20720 2388 20772 2440
rect 20904 2431 20956 2440
rect 20904 2397 20913 2431
rect 20913 2397 20947 2431
rect 20947 2397 20956 2431
rect 20904 2388 20956 2397
rect 21456 2388 21508 2440
rect 21824 2388 21876 2440
rect 22376 2388 22428 2440
rect 23480 2431 23532 2440
rect 23480 2397 23489 2431
rect 23489 2397 23523 2431
rect 23523 2397 23532 2431
rect 23480 2388 23532 2397
rect 29828 2524 29880 2576
rect 31484 2592 31536 2644
rect 33416 2592 33468 2644
rect 39396 2635 39448 2644
rect 39396 2601 39405 2635
rect 39405 2601 39439 2635
rect 39439 2601 39448 2635
rect 39396 2592 39448 2601
rect 24400 2431 24452 2440
rect 24400 2397 24409 2431
rect 24409 2397 24443 2431
rect 24443 2397 24452 2431
rect 24400 2388 24452 2397
rect 12992 2252 13044 2304
rect 13084 2252 13136 2304
rect 13820 2252 13872 2304
rect 14556 2252 14608 2304
rect 15384 2252 15436 2304
rect 16028 2252 16080 2304
rect 16764 2252 16816 2304
rect 17684 2252 17736 2304
rect 17776 2252 17828 2304
rect 18236 2252 18288 2304
rect 18972 2252 19024 2304
rect 19340 2295 19392 2304
rect 19340 2261 19349 2295
rect 19349 2261 19383 2295
rect 19383 2261 19392 2295
rect 19340 2252 19392 2261
rect 20444 2252 20496 2304
rect 20720 2252 20772 2304
rect 21364 2295 21416 2304
rect 21364 2261 21373 2295
rect 21373 2261 21407 2295
rect 21407 2261 21416 2295
rect 21364 2252 21416 2261
rect 22560 2320 22612 2372
rect 30472 2431 30524 2440
rect 30472 2397 30481 2431
rect 30481 2397 30515 2431
rect 30515 2397 30524 2431
rect 30472 2388 30524 2397
rect 32956 2456 33008 2508
rect 33600 2456 33652 2508
rect 39948 2524 40000 2576
rect 33416 2388 33468 2440
rect 38108 2431 38160 2440
rect 38108 2397 38117 2431
rect 38117 2397 38151 2431
rect 38151 2397 38160 2431
rect 38108 2388 38160 2397
rect 38476 2431 38528 2440
rect 38476 2397 38485 2431
rect 38485 2397 38519 2431
rect 38519 2397 38528 2431
rect 38476 2388 38528 2397
rect 38568 2388 38620 2440
rect 26332 2320 26384 2372
rect 24124 2252 24176 2304
rect 30288 2295 30340 2304
rect 30288 2261 30297 2295
rect 30297 2261 30331 2295
rect 30331 2261 30340 2295
rect 30288 2252 30340 2261
rect 30748 2252 30800 2304
rect 31300 2295 31352 2304
rect 31300 2261 31309 2295
rect 31309 2261 31343 2295
rect 31343 2261 31352 2295
rect 31300 2252 31352 2261
rect 37924 2295 37976 2304
rect 37924 2261 37933 2295
rect 37933 2261 37967 2295
rect 37967 2261 37976 2295
rect 37924 2252 37976 2261
rect 38292 2295 38344 2304
rect 38292 2261 38301 2295
rect 38301 2261 38335 2295
rect 38335 2261 38344 2295
rect 38292 2252 38344 2261
rect 38660 2295 38712 2304
rect 38660 2261 38669 2295
rect 38669 2261 38703 2295
rect 38703 2261 38712 2295
rect 38660 2252 38712 2261
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 39010 2150 39062 2202
rect 39074 2150 39126 2202
rect 39138 2150 39190 2202
rect 39202 2150 39254 2202
rect 39266 2150 39318 2202
rect 4804 2048 4856 2100
rect 7564 2048 7616 2100
rect 10968 2048 11020 2100
rect 20904 2048 20956 2100
rect 29828 2048 29880 2100
rect 32312 2048 32364 2100
rect 32956 2048 33008 2100
rect 38384 2048 38436 2100
rect 9680 1980 9732 2032
rect 25412 1980 25464 2032
rect 1676 1912 1728 1964
rect 19248 1912 19300 1964
rect 19616 1912 19668 1964
rect 38568 1912 38620 1964
rect 3700 1844 3752 1896
rect 11520 1844 11572 1896
rect 15660 1844 15712 1896
rect 24308 1844 24360 1896
rect 2872 1776 2924 1828
rect 21640 1776 21692 1828
rect 21916 1776 21968 1828
rect 23296 1776 23348 1828
rect 25596 1776 25648 1828
rect 27804 1776 27856 1828
rect 6184 1708 6236 1760
rect 12440 1708 12492 1760
rect 14832 1708 14884 1760
rect 24400 1708 24452 1760
rect 7656 1640 7708 1692
rect 14740 1640 14792 1692
rect 14924 1640 14976 1692
rect 29184 1640 29236 1692
rect 18144 1572 18196 1624
rect 29092 1572 29144 1624
rect 8208 1504 8260 1556
rect 16580 1504 16632 1556
rect 21732 1504 21784 1556
rect 38108 1504 38160 1556
rect 10784 1436 10836 1488
rect 19340 1436 19392 1488
rect 27068 1368 27120 1420
rect 29000 1368 29052 1420
rect 35716 1368 35768 1420
rect 38108 1368 38160 1420
rect 14464 1300 14516 1352
rect 32772 1300 32824 1352
rect 9956 1232 10008 1284
rect 39672 1232 39724 1284
rect 7564 1164 7616 1216
rect 21548 1164 21600 1216
rect 2504 1096 2556 1148
rect 29460 1096 29512 1148
rect 8576 1028 8628 1080
rect 35072 1028 35124 1080
rect 2688 960 2740 1012
rect 25044 960 25096 1012
rect 32220 960 32272 1012
rect 34244 960 34296 1012
rect 13360 892 13412 944
rect 37188 892 37240 944
rect 10508 824 10560 876
rect 26608 824 26660 876
rect 7012 756 7064 808
rect 38200 756 38252 808
rect 6644 688 6696 740
rect 33416 688 33468 740
rect 7840 620 7892 672
rect 23480 620 23532 672
rect 28632 8 28684 60
rect 39856 8 39908 60
<< metal2 >>
rect 3238 11194 3294 11250
rect 3514 11194 3570 11250
rect 3790 11194 3846 11250
rect 4066 11194 4122 11250
rect 4342 11194 4398 11250
rect 4618 11194 4674 11250
rect 4894 11194 4950 11250
rect 5170 11194 5226 11250
rect 5446 11194 5502 11250
rect 5722 11194 5778 11250
rect 5998 11194 6054 11250
rect 6274 11194 6330 11250
rect 6550 11194 6606 11250
rect 6826 11194 6882 11250
rect 7102 11194 7158 11250
rect 7378 11194 7434 11250
rect 7654 11194 7710 11250
rect 7930 11194 7986 11250
rect 8206 11194 8262 11250
rect 8482 11194 8538 11250
rect 8758 11194 8814 11250
rect 9034 11194 9090 11250
rect 9310 11194 9366 11250
rect 9586 11194 9642 11250
rect 9862 11194 9918 11250
rect 10138 11194 10194 11250
rect 10414 11194 10470 11250
rect 10690 11194 10746 11250
rect 10966 11194 11022 11250
rect 11242 11194 11298 11250
rect 11518 11194 11574 11250
rect 11794 11194 11850 11250
rect 12070 11194 12126 11250
rect 12346 11194 12402 11250
rect 12622 11194 12678 11250
rect 12898 11194 12954 11250
rect 13174 11194 13230 11250
rect 13450 11194 13506 11250
rect 13726 11194 13782 11250
rect 14002 11194 14058 11250
rect 14278 11194 14334 11250
rect 14554 11194 14610 11250
rect 14830 11194 14886 11250
rect 15106 11194 15162 11250
rect 15382 11194 15438 11250
rect 15658 11194 15714 11250
rect 15934 11194 15990 11250
rect 16210 11194 16266 11250
rect 16486 11194 16542 11250
rect 16762 11194 16818 11250
rect 17038 11194 17094 11250
rect 17314 11194 17370 11250
rect 17590 11194 17646 11250
rect 17866 11194 17922 11250
rect 18142 11194 18198 11250
rect 18418 11194 18474 11250
rect 18694 11194 18750 11250
rect 18970 11194 19026 11250
rect 19246 11194 19302 11250
rect 19522 11194 19578 11250
rect 19798 11194 19854 11250
rect 20074 11194 20130 11250
rect 20350 11194 20406 11250
rect 20626 11194 20682 11250
rect 20902 11194 20958 11250
rect 21178 11194 21234 11250
rect 21454 11194 21510 11250
rect 21730 11194 21786 11250
rect 22006 11194 22062 11250
rect 22282 11194 22338 11250
rect 22558 11194 22614 11250
rect 22834 11194 22890 11250
rect 23110 11194 23166 11250
rect 23386 11194 23442 11250
rect 23662 11194 23718 11250
rect 23938 11194 23994 11250
rect 24214 11194 24270 11250
rect 24490 11194 24546 11250
rect 24766 11194 24822 11250
rect 25042 11194 25098 11250
rect 25318 11194 25374 11250
rect 25594 11194 25650 11250
rect 25870 11194 25926 11250
rect 26146 11194 26202 11250
rect 26422 11194 26478 11250
rect 26698 11194 26754 11250
rect 26974 11194 27030 11250
rect 27250 11194 27306 11250
rect 27526 11194 27582 11250
rect 27802 11194 27858 11250
rect 28078 11194 28134 11250
rect 28354 11194 28410 11250
rect 28630 11194 28686 11250
rect 28906 11194 28962 11250
rect 29182 11194 29238 11250
rect 29458 11194 29514 11250
rect 29734 11194 29790 11250
rect 30010 11194 30066 11250
rect 30286 11194 30342 11250
rect 30562 11194 30618 11250
rect 30838 11194 30894 11250
rect 31114 11194 31170 11250
rect 31390 11194 31446 11250
rect 31666 11194 31722 11250
rect 31942 11194 31998 11250
rect 32218 11194 32274 11250
rect 32494 11194 32550 11250
rect 32770 11194 32826 11250
rect 33046 11194 33102 11250
rect 33322 11194 33378 11250
rect 33598 11194 33654 11250
rect 33874 11194 33930 11250
rect 34150 11194 34206 11250
rect 34426 11194 34482 11250
rect 34702 11194 34758 11250
rect 34978 11194 35034 11250
rect 35254 11194 35310 11250
rect 35530 11194 35586 11250
rect 35806 11194 35862 11250
rect 36082 11194 36138 11250
rect 36358 11194 36414 11250
rect 36634 11194 36690 11250
rect 36910 11194 36966 11250
rect 37186 11194 37242 11250
rect 37462 11194 37518 11250
rect 37738 11194 37794 11250
rect 2318 10160 2374 10169
rect 2318 10095 2374 10104
rect 478 9888 534 9897
rect 478 9823 534 9832
rect 492 8498 520 9823
rect 662 9616 718 9625
rect 662 9551 718 9560
rect 480 8492 532 8498
rect 480 8434 532 8440
rect 386 8256 442 8265
rect 386 8191 442 8200
rect 400 7818 428 8191
rect 676 7954 704 9551
rect 1214 9344 1270 9353
rect 1214 9279 1270 9288
rect 756 8424 808 8430
rect 756 8366 808 8372
rect 768 7993 796 8366
rect 754 7984 810 7993
rect 664 7948 716 7954
rect 754 7919 810 7928
rect 664 7890 716 7896
rect 388 7812 440 7818
rect 388 7754 440 7760
rect 1228 7750 1256 9279
rect 1676 9240 1728 9246
rect 1676 9182 1728 9188
rect 1308 8560 1360 8566
rect 1306 8528 1308 8537
rect 1360 8528 1362 8537
rect 1306 8463 1362 8472
rect 1688 8430 1716 9182
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 1216 7744 1268 7750
rect 754 7712 810 7721
rect 1216 7686 1268 7692
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 754 7647 810 7656
rect 768 7410 796 7647
rect 1964 7478 1992 7686
rect 940 7472 992 7478
rect 938 7440 940 7449
rect 1952 7472 2004 7478
rect 992 7440 994 7449
rect 756 7404 808 7410
rect 1952 7414 2004 7420
rect 938 7375 994 7384
rect 756 7346 808 7352
rect 1124 7336 1176 7342
rect 1124 7278 1176 7284
rect 1136 7177 1164 7278
rect 1122 7168 1178 7177
rect 1122 7103 1178 7112
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 204 6792 256 6798
rect 204 6734 256 6740
rect 216 6633 244 6734
rect 1584 6656 1636 6662
rect 202 6624 258 6633
rect 1584 6598 1636 6604
rect 202 6559 258 6568
rect 940 6384 992 6390
rect 938 6352 940 6361
rect 992 6352 994 6361
rect 756 6316 808 6322
rect 938 6287 994 6296
rect 756 6258 808 6264
rect 768 6089 796 6258
rect 754 6080 810 6089
rect 754 6015 810 6024
rect 1596 5914 1624 6598
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1676 6248 1728 6254
rect 1674 6216 1676 6225
rect 1728 6216 1730 6225
rect 1674 6151 1730 6160
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 754 5808 810 5817
rect 754 5743 810 5752
rect 1032 5772 1084 5778
rect 768 5710 796 5743
rect 1032 5714 1084 5720
rect 756 5704 808 5710
rect 756 5646 808 5652
rect 572 5636 624 5642
rect 572 5578 624 5584
rect 584 5545 612 5578
rect 570 5536 626 5545
rect 570 5471 626 5480
rect 940 5296 992 5302
rect 1044 5273 1072 5714
rect 940 5238 992 5244
rect 1030 5264 1086 5273
rect 388 5228 440 5234
rect 388 5170 440 5176
rect 400 5001 428 5170
rect 386 4992 442 5001
rect 386 4927 442 4936
rect 952 4729 980 5238
rect 1030 5199 1086 5208
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1596 4826 1624 4966
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1872 4758 1900 6258
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2332 5370 2360 10095
rect 2596 9988 2648 9994
rect 2596 9930 2648 9936
rect 2608 8022 2636 9930
rect 3252 9466 3280 11194
rect 3252 9438 3464 9466
rect 2688 9308 2740 9314
rect 2688 9250 2740 9256
rect 2596 8016 2648 8022
rect 2596 7958 2648 7964
rect 2700 6914 2728 9250
rect 2778 9072 2834 9081
rect 2778 9007 2834 9016
rect 2792 7886 2820 9007
rect 2870 8800 2926 8809
rect 2870 8735 2926 8744
rect 2884 7886 2912 8735
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 3436 8090 3464 9438
rect 3528 8090 3556 11194
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3620 8498 3648 9114
rect 3804 8634 3832 11194
rect 3974 10024 4030 10033
rect 3974 9959 4030 9968
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 3620 7449 3648 7822
rect 3606 7440 3662 7449
rect 2964 7404 3016 7410
rect 3606 7375 3662 7384
rect 2964 7346 3016 7352
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2884 7002 2912 7142
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 2608 6886 2728 6914
rect 2976 6905 3004 7346
rect 3608 7268 3660 7274
rect 3608 7210 3660 7216
rect 2962 6896 3018 6905
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2516 5166 2544 6394
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 1860 4752 1912 4758
rect 938 4720 994 4729
rect 1860 4694 1912 4700
rect 938 4655 994 4664
rect 572 4616 624 4622
rect 572 4558 624 4564
rect 584 3641 612 4558
rect 2516 4554 2544 5102
rect 756 4548 808 4554
rect 756 4490 808 4496
rect 2504 4548 2556 4554
rect 2504 4490 2556 4496
rect 768 4457 796 4490
rect 754 4448 810 4457
rect 754 4383 810 4392
rect 1952 4276 2004 4282
rect 1952 4218 2004 4224
rect 756 4208 808 4214
rect 754 4176 756 4185
rect 1964 4185 1992 4218
rect 808 4176 810 4185
rect 1950 4176 2006 4185
rect 754 4111 810 4120
rect 940 4140 992 4146
rect 1950 4111 2006 4120
rect 940 4082 992 4088
rect 952 3913 980 4082
rect 2504 4072 2556 4078
rect 2318 4040 2374 4049
rect 2504 4014 2556 4020
rect 2318 3975 2320 3984
rect 2372 3975 2374 3984
rect 2320 3946 2372 3952
rect 938 3904 994 3913
rect 938 3839 994 3848
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2516 3738 2544 4014
rect 2608 4010 2636 6886
rect 2962 6831 3018 6840
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 2792 5324 3188 5352
rect 2792 5250 2820 5324
rect 2700 5234 2820 5250
rect 2688 5228 2820 5234
rect 2740 5222 2820 5228
rect 2688 5170 2740 5176
rect 2792 4622 2820 5222
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2596 4004 2648 4010
rect 2596 3946 2648 3952
rect 2884 3942 2912 5170
rect 3160 5166 3188 5324
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3424 4752 3476 4758
rect 3424 4694 3476 4700
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 570 3632 626 3641
rect 570 3567 626 3576
rect 2502 3632 2558 3641
rect 3160 3602 3188 4014
rect 3436 3602 3464 4694
rect 3528 4078 3556 4966
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 2502 3567 2558 3576
rect 2872 3596 2924 3602
rect 204 3528 256 3534
rect 204 3470 256 3476
rect 2320 3528 2372 3534
rect 2320 3470 2372 3476
rect 216 3369 244 3470
rect 1308 3460 1360 3466
rect 1308 3402 1360 3408
rect 202 3360 258 3369
rect 202 3295 258 3304
rect 1320 3097 1348 3402
rect 1860 3120 1912 3126
rect 1306 3088 1362 3097
rect 1216 3052 1268 3058
rect 1860 3062 1912 3068
rect 1306 3023 1362 3032
rect 1216 2994 1268 3000
rect 388 2984 440 2990
rect 388 2926 440 2932
rect 400 2553 428 2926
rect 1124 2916 1176 2922
rect 1124 2858 1176 2864
rect 386 2544 442 2553
rect 386 2479 442 2488
rect 1136 2281 1164 2858
rect 1228 2825 1256 2994
rect 1214 2816 1270 2825
rect 1214 2751 1270 2760
rect 1216 2508 1268 2514
rect 1216 2450 1268 2456
rect 1122 2272 1178 2281
rect 1122 2207 1178 2216
rect 1228 1737 1256 2450
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1214 1728 1270 1737
rect 1214 1663 1270 1672
rect 1320 56 1348 2382
rect 1688 1970 1716 2382
rect 1872 2009 1900 3062
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 1858 2000 1914 2009
rect 1676 1964 1728 1970
rect 1858 1935 1914 1944
rect 1676 1906 1728 1912
rect 2056 56 2176 82
rect 1306 0 1362 56
rect 2042 54 2176 56
rect 2042 0 2098 54
rect 2148 42 2176 54
rect 2332 42 2360 3470
rect 2516 3398 2544 3567
rect 2872 3538 2924 3544
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2688 2984 2740 2990
rect 2688 2926 2740 2932
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 2516 1154 2544 2790
rect 2608 1465 2636 2790
rect 2594 1456 2650 1465
rect 2594 1391 2650 1400
rect 2504 1148 2556 1154
rect 2504 1090 2556 1096
rect 2700 1018 2728 2926
rect 2688 1012 2740 1018
rect 2688 954 2740 960
rect 2792 56 2820 2994
rect 2884 1834 2912 3538
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 3148 2984 3200 2990
rect 3146 2952 3148 2961
rect 3200 2952 3202 2961
rect 3146 2887 3202 2896
rect 3424 2916 3476 2922
rect 3424 2858 3476 2864
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 2872 1828 2924 1834
rect 2872 1770 2924 1776
rect 3436 921 3464 2858
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 3422 912 3478 921
rect 3422 847 3478 856
rect 3528 56 3556 2382
rect 3620 785 3648 7210
rect 3804 5166 3832 8298
rect 3988 7886 4016 9959
rect 4080 8090 4108 11194
rect 4252 10396 4304 10402
rect 4252 10338 4304 10344
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 4172 7478 4200 10202
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 3896 6458 3924 6734
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 4172 6390 4200 6734
rect 4160 6384 4212 6390
rect 4158 6352 4160 6361
rect 4212 6352 4214 6361
rect 4158 6287 4214 6296
rect 3884 6180 3936 6186
rect 3884 6122 3936 6128
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3700 2304 3752 2310
rect 3700 2246 3752 2252
rect 3712 1902 3740 2246
rect 3700 1896 3752 1902
rect 3700 1838 3752 1844
rect 3606 776 3662 785
rect 3606 711 3662 720
rect 3804 649 3832 3878
rect 3896 1329 3924 6122
rect 4172 5710 4200 6287
rect 4264 5930 4292 10338
rect 4356 8634 4384 11194
rect 4434 9752 4490 9761
rect 4434 9687 4490 9696
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4448 7970 4476 9687
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4540 8498 4568 9590
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4632 8090 4660 11194
rect 4908 8634 4936 11194
rect 5078 9208 5134 9217
rect 5078 9143 5134 9152
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5092 8498 5120 9143
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4448 7942 4568 7970
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4448 6390 4476 7686
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 4540 6322 4568 7942
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4264 5902 4476 5930
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4172 4146 4200 5510
rect 4342 5264 4398 5273
rect 4342 5199 4398 5208
rect 4356 4282 4384 5199
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4356 4146 4384 4218
rect 4448 4146 4476 5902
rect 4724 5370 4752 8434
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 4894 8392 4950 8401
rect 4816 7585 4844 8366
rect 4894 8327 4950 8336
rect 4908 7886 4936 8327
rect 5184 8090 5212 11194
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5080 8016 5132 8022
rect 5080 7958 5132 7964
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4802 7576 4858 7585
rect 4802 7511 4858 7520
rect 4896 7472 4948 7478
rect 4896 7414 4948 7420
rect 4908 7002 4936 7414
rect 5000 7002 5028 7822
rect 5092 7342 5120 7958
rect 5276 7698 5304 9522
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5184 7670 5304 7698
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 5080 6384 5132 6390
rect 5080 6326 5132 6332
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4908 5710 4936 6258
rect 5092 5846 5120 6326
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4896 5704 4948 5710
rect 4896 5646 4948 5652
rect 5078 5672 5134 5681
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4540 4729 4568 5170
rect 4526 4720 4582 4729
rect 4526 4655 4582 4664
rect 4540 4622 4568 4655
rect 4816 4622 4844 5646
rect 5078 5607 5134 5616
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3988 3194 4016 3878
rect 4448 3534 4476 4082
rect 4724 4078 4752 4422
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 4356 3194 4384 3334
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4816 3046 5028 3074
rect 5092 3058 5120 5607
rect 5184 3398 5212 7670
rect 5368 7546 5396 9046
rect 5460 8362 5488 11194
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5644 8498 5672 9318
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5736 8090 5764 11194
rect 5908 8900 5960 8906
rect 5908 8842 5960 8848
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5828 8498 5856 8774
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5540 7880 5592 7886
rect 5538 7848 5540 7857
rect 5592 7848 5594 7857
rect 5538 7783 5594 7792
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5276 4185 5304 7482
rect 5816 7336 5868 7342
rect 5816 7278 5868 7284
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5552 6798 5580 7142
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5460 6186 5488 6666
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5828 5409 5856 7278
rect 5920 6662 5948 8842
rect 6012 8566 6040 11194
rect 6182 9480 6238 9489
rect 6182 9415 6238 9424
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 6196 8498 6224 9415
rect 6288 8634 6316 11194
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6380 7886 6408 9386
rect 6564 8090 6592 11194
rect 6642 9888 6698 9897
rect 6642 9823 6698 9832
rect 6656 8634 6684 9823
rect 6734 9752 6790 9761
rect 6734 9687 6790 9696
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6642 8528 6698 8537
rect 6642 8463 6644 8472
rect 6696 8463 6698 8472
rect 6644 8434 6696 8440
rect 6748 8090 6776 9687
rect 6840 8430 6868 11194
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6826 7984 6882 7993
rect 6826 7919 6828 7928
rect 6880 7919 6882 7928
rect 6828 7890 6880 7896
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6012 7206 6040 7822
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6092 7472 6144 7478
rect 6092 7414 6144 7420
rect 6104 7342 6132 7414
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6460 7268 6512 7274
rect 6460 7210 6512 7216
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5814 5400 5870 5409
rect 5814 5335 5870 5344
rect 5262 4176 5318 4185
rect 5262 4111 5318 4120
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5368 3126 5396 3334
rect 5356 3120 5408 3126
rect 5460 3097 5488 4014
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5356 3062 5408 3068
rect 5446 3088 5502 3097
rect 4816 2990 4844 3046
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4172 2582 4200 2790
rect 4724 2689 4752 2790
rect 4710 2680 4766 2689
rect 4710 2615 4766 2624
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 4160 2576 4212 2582
rect 4160 2518 4212 2524
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4252 2508 4304 2514
rect 4252 2450 4304 2456
rect 3882 1320 3938 1329
rect 3882 1255 3938 1264
rect 3790 640 3846 649
rect 3790 575 3846 584
rect 4264 56 4292 2450
rect 4724 2446 4752 2518
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4816 2106 4844 2586
rect 4908 2514 4936 2926
rect 4896 2508 4948 2514
rect 4896 2450 4948 2456
rect 4804 2100 4856 2106
rect 4804 2042 4856 2048
rect 5000 56 5028 3046
rect 5080 3052 5132 3058
rect 5446 3023 5502 3032
rect 5080 2994 5132 3000
rect 5644 1057 5672 3674
rect 5724 3528 5776 3534
rect 5722 3496 5724 3505
rect 5776 3496 5778 3505
rect 5722 3431 5778 3440
rect 5724 2576 5776 2582
rect 5724 2518 5776 2524
rect 5630 1048 5686 1057
rect 5630 983 5686 992
rect 5736 56 5764 2518
rect 5828 2378 5856 5335
rect 5906 5128 5962 5137
rect 5906 5063 5962 5072
rect 5920 4690 5948 5063
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 6012 4554 6040 6802
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6104 5574 6132 5850
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6196 4622 6224 6054
rect 6288 5778 6316 6598
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6000 4548 6052 4554
rect 6000 4490 6052 4496
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 5920 2650 5948 3538
rect 6092 3052 6144 3058
rect 6196 3040 6224 4558
rect 6288 3210 6316 5714
rect 6380 5030 6408 6734
rect 6472 6458 6500 7210
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6460 6180 6512 6186
rect 6460 6122 6512 6128
rect 6472 5137 6500 6122
rect 6564 5710 6592 6190
rect 6656 5817 6684 7686
rect 6748 7478 6776 7686
rect 6736 7472 6788 7478
rect 6736 7414 6788 7420
rect 6642 5808 6698 5817
rect 6642 5743 6698 5752
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6458 5128 6514 5137
rect 6458 5063 6514 5072
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6564 4282 6592 5034
rect 6736 4548 6788 4554
rect 6736 4490 6788 4496
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6748 4146 6776 4490
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6564 3738 6592 4014
rect 6932 4010 6960 10066
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 7024 8498 7052 8910
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7116 7546 7144 11194
rect 7392 9761 7420 11194
rect 7378 9752 7434 9761
rect 7378 9687 7434 9696
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7300 8566 7328 9454
rect 7378 8936 7434 8945
rect 7378 8871 7434 8880
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 7392 8498 7420 8871
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 7012 7336 7064 7342
rect 7116 7313 7144 7346
rect 7012 7278 7064 7284
rect 7102 7304 7158 7313
rect 7024 6866 7052 7278
rect 7102 7239 7158 7248
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 7024 5642 7052 5850
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 7116 5545 7144 7142
rect 7208 6662 7236 8366
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7484 8090 7512 8230
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7668 8022 7696 11194
rect 7944 9518 7972 11194
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7380 7880 7432 7886
rect 7748 7880 7800 7886
rect 7380 7822 7432 7828
rect 7668 7840 7748 7868
rect 7300 6905 7328 7822
rect 7392 7313 7420 7822
rect 7564 7812 7616 7818
rect 7564 7754 7616 7760
rect 7576 7546 7604 7754
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7378 7304 7434 7313
rect 7378 7239 7434 7248
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7470 7168 7526 7177
rect 7286 6896 7342 6905
rect 7286 6831 7342 6840
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7286 6624 7342 6633
rect 7286 6559 7342 6568
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7208 5710 7236 6054
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7102 5536 7158 5545
rect 7102 5471 7158 5480
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7024 4826 7052 5170
rect 7300 5166 7328 6559
rect 7288 5160 7340 5166
rect 7286 5128 7288 5137
rect 7340 5128 7342 5137
rect 7286 5063 7342 5072
rect 7194 4992 7250 5001
rect 7194 4927 7250 4936
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 7208 4486 7236 4927
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 7024 4078 7052 4218
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6288 3182 6408 3210
rect 6748 3194 6776 3538
rect 6932 3534 6960 3946
rect 7208 3602 7236 4422
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7300 3942 7328 4218
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6144 3012 6224 3040
rect 6092 2994 6144 3000
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 6196 2514 6224 3012
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 6288 2378 6316 2994
rect 6380 2990 6408 3182
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6564 2689 6592 2790
rect 6550 2680 6606 2689
rect 6550 2615 6606 2624
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 6276 2372 6328 2378
rect 6276 2314 6328 2320
rect 6184 2304 6236 2310
rect 6184 2246 6236 2252
rect 6196 1766 6224 2246
rect 6184 1760 6236 1766
rect 6184 1702 6236 1708
rect 6380 1170 6408 2382
rect 6644 2372 6696 2378
rect 6644 2314 6696 2320
rect 7012 2372 7064 2378
rect 7012 2314 7064 2320
rect 6380 1142 6500 1170
rect 6472 56 6500 1142
rect 6656 746 6684 2314
rect 7024 814 7052 2314
rect 7300 1170 7328 2382
rect 7392 1193 7420 7142
rect 7470 7103 7526 7112
rect 7484 4826 7512 7103
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7576 6769 7604 6870
rect 7562 6760 7618 6769
rect 7562 6695 7618 6704
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7576 6186 7604 6598
rect 7668 6254 7696 7840
rect 7852 7868 7880 8434
rect 8220 8294 8248 11194
rect 8496 9897 8524 11194
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 8482 9888 8538 9897
rect 8482 9823 8538 9832
rect 8298 9616 8354 9625
rect 8298 9551 8354 9560
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 8024 7880 8076 7886
rect 7852 7840 8024 7868
rect 7748 7822 7800 7828
rect 8024 7822 8076 7828
rect 8036 7410 8064 7822
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 7748 7268 7800 7274
rect 7748 7210 7800 7216
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7668 5681 7696 6190
rect 7654 5672 7710 5681
rect 7654 5607 7710 5616
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7484 2854 7512 4422
rect 7576 4146 7604 5510
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7668 5137 7696 5170
rect 7654 5128 7710 5137
rect 7654 5063 7710 5072
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7668 4690 7696 4966
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7654 4584 7710 4593
rect 7654 4519 7656 4528
rect 7708 4519 7710 4528
rect 7656 4490 7708 4496
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7564 3528 7616 3534
rect 7668 3505 7696 3878
rect 7564 3470 7616 3476
rect 7654 3496 7710 3505
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7576 2378 7604 3470
rect 7654 3431 7710 3440
rect 7760 2553 7788 7210
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 8312 6882 8340 9551
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8496 8566 8524 9114
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8404 7177 8432 7754
rect 8496 7206 8524 8230
rect 8484 7200 8536 7206
rect 8390 7168 8446 7177
rect 8484 7142 8536 7148
rect 8390 7103 8446 7112
rect 8404 7018 8432 7103
rect 8404 6990 8524 7018
rect 8220 6854 8340 6882
rect 7932 6792 7984 6798
rect 7852 6740 7932 6746
rect 7852 6734 7984 6740
rect 7852 6718 7972 6734
rect 7852 6186 7880 6718
rect 7930 6488 7986 6497
rect 7930 6423 7932 6432
rect 7984 6423 7986 6432
rect 7932 6394 7984 6400
rect 8220 6202 8248 6854
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 7840 6180 7892 6186
rect 8220 6174 8340 6202
rect 7840 6122 7892 6128
rect 7852 4758 7880 6122
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 8206 5536 8262 5545
rect 7944 5302 7972 5510
rect 8206 5471 8262 5480
rect 7932 5296 7984 5302
rect 7932 5238 7984 5244
rect 8220 5137 8248 5471
rect 8206 5128 8262 5137
rect 8206 5063 8262 5072
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 8312 4758 8340 6174
rect 7840 4752 7892 4758
rect 7840 4694 7892 4700
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8312 4282 8340 4558
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8024 4004 8076 4010
rect 7852 3964 8024 3992
rect 7746 2544 7802 2553
rect 7746 2479 7802 2488
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 7564 2100 7616 2106
rect 7564 2042 7616 2048
rect 7576 1222 7604 2042
rect 7668 1698 7696 2246
rect 7656 1692 7708 1698
rect 7656 1634 7708 1640
rect 7564 1216 7616 1222
rect 7208 1142 7328 1170
rect 7378 1184 7434 1193
rect 7012 808 7064 814
rect 7012 750 7064 756
rect 6644 740 6696 746
rect 6644 682 6696 688
rect 7208 56 7236 1142
rect 7564 1158 7616 1164
rect 7378 1119 7434 1128
rect 7852 678 7880 3964
rect 8024 3946 8076 3952
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 8404 3126 8432 6734
rect 8496 6633 8524 6990
rect 8482 6624 8538 6633
rect 8482 6559 8538 6568
rect 8588 6338 8616 10406
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8680 7954 8708 9998
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8680 7750 8708 7890
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8680 7002 8708 7346
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8496 6310 8616 6338
rect 8680 6322 8708 6802
rect 8772 6662 8800 11194
rect 9048 8922 9076 11194
rect 9324 9674 9352 11194
rect 9324 9646 9444 9674
rect 8864 8894 9076 8922
rect 8864 8634 8892 8894
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9034 8392 9090 8401
rect 9034 8327 9090 8336
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 8956 8090 8984 8230
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8864 7392 8892 7890
rect 9048 7750 9076 8327
rect 9232 7886 9260 8434
rect 9220 7880 9272 7886
rect 9416 7868 9444 9646
rect 9494 9344 9550 9353
rect 9494 9279 9550 9288
rect 9508 8498 9536 9279
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9416 7840 9536 7868
rect 9220 7822 9272 7828
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 8944 7404 8996 7410
rect 8864 7364 8944 7392
rect 9508 7392 9536 7840
rect 8944 7346 8996 7352
rect 9416 7364 9536 7392
rect 9312 7200 9364 7206
rect 9140 7160 9312 7188
rect 9140 6866 9168 7160
rect 9312 7142 9364 7148
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9036 6792 9088 6798
rect 9312 6792 9364 6798
rect 9232 6752 9312 6780
rect 9232 6746 9260 6752
rect 9088 6740 9260 6746
rect 9036 6734 9260 6740
rect 9312 6734 9364 6740
rect 9048 6718 9260 6734
rect 9416 6662 9444 7364
rect 9496 7268 9548 7274
rect 9496 7210 9548 7216
rect 9508 7177 9536 7210
rect 9494 7168 9550 7177
rect 9494 7103 9550 7112
rect 9600 6798 9628 11194
rect 9680 9240 9732 9246
rect 9680 9182 9732 9188
rect 9692 9081 9720 9182
rect 9772 9104 9824 9110
rect 9678 9072 9734 9081
rect 9772 9046 9824 9052
rect 9678 9007 9734 9016
rect 9784 8786 9812 9046
rect 9876 8809 9904 11194
rect 9956 9852 10008 9858
rect 9956 9794 10008 9800
rect 9692 8758 9812 8786
rect 9862 8800 9918 8809
rect 9692 8634 9720 8758
rect 9862 8735 9918 8744
rect 9968 8634 9996 9794
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 10060 8634 10088 9658
rect 10152 9110 10180 11194
rect 10324 9308 10376 9314
rect 10324 9250 10376 9256
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 9692 8498 9996 8514
rect 10244 8498 10272 8978
rect 10336 8498 10364 9250
rect 9680 8492 9996 8498
rect 9732 8486 9996 8492
rect 9680 8434 9732 8440
rect 9968 8129 9996 8486
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 9770 8120 9826 8129
rect 9770 8055 9826 8064
rect 9954 8120 10010 8129
rect 10428 8090 10456 11194
rect 10600 10872 10652 10878
rect 10600 10814 10652 10820
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10520 8498 10548 8842
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 9954 8055 10010 8064
rect 10416 8084 10468 8090
rect 9784 7410 9812 8055
rect 10416 8026 10468 8032
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 9956 7812 10008 7818
rect 9956 7754 10008 7760
rect 9968 7721 9996 7754
rect 9954 7712 10010 7721
rect 9954 7647 10010 7656
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9968 7342 9996 7482
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 9692 6934 9720 7278
rect 10152 7041 10180 7346
rect 9954 7032 10010 7041
rect 9772 6996 9824 7002
rect 9954 6967 9956 6976
rect 9772 6938 9824 6944
rect 10008 6967 10010 6976
rect 10138 7032 10194 7041
rect 10138 6967 10194 6976
rect 9956 6938 10008 6944
rect 9680 6928 9732 6934
rect 9680 6870 9732 6876
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 8758 6488 8814 6497
rect 9010 6491 9318 6500
rect 8758 6423 8814 6432
rect 8772 6390 8800 6423
rect 8760 6384 8812 6390
rect 8760 6326 8812 6332
rect 9508 6322 9536 6666
rect 9784 6633 9812 6938
rect 10244 6916 10272 7890
rect 10416 7812 10468 7818
rect 10416 7754 10468 7760
rect 9954 6896 10010 6905
rect 9954 6831 10010 6840
rect 10152 6888 10272 6916
rect 9770 6624 9826 6633
rect 9770 6559 9826 6568
rect 9968 6361 9996 6831
rect 9954 6352 10010 6361
rect 8668 6316 8720 6322
rect 8496 5846 8524 6310
rect 8668 6258 8720 6264
rect 9496 6316 9548 6322
rect 9954 6287 10010 6296
rect 9496 6258 9548 6264
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8496 5302 8524 5646
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 7840 672 7892 678
rect 7840 614 7892 620
rect 7944 56 7972 2382
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 8220 1562 8248 2246
rect 8208 1556 8260 1562
rect 8208 1498 8260 1504
rect 8588 1086 8616 6054
rect 8680 4321 8708 6258
rect 10152 6254 10180 6888
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 9128 6248 9180 6254
rect 9772 6248 9824 6254
rect 9180 6196 9772 6202
rect 9128 6190 9824 6196
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 9140 6174 9812 6190
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9140 5710 9168 6054
rect 9128 5704 9180 5710
rect 9784 5681 9812 6174
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10152 5846 10180 6054
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 9128 5646 9180 5652
rect 9494 5672 9550 5681
rect 9494 5607 9550 5616
rect 9770 5672 9826 5681
rect 9770 5607 9826 5616
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8852 5568 8904 5574
rect 8852 5510 8904 5516
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 8772 5284 8800 5510
rect 8864 5409 8892 5510
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 8850 5400 8906 5409
rect 9010 5403 9318 5412
rect 8850 5335 8906 5344
rect 8852 5296 8904 5302
rect 8772 5256 8852 5284
rect 8852 5238 8904 5244
rect 9416 5137 9444 5510
rect 9508 5370 9536 5607
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 10046 5536 10102 5545
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9402 5128 9458 5137
rect 9402 5063 9458 5072
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 8760 4752 8812 4758
rect 8760 4694 8812 4700
rect 8666 4312 8722 4321
rect 8666 4247 8722 4256
rect 8772 4078 8800 4694
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 8772 3602 8800 4014
rect 8864 4010 8892 4966
rect 9784 4826 9812 5170
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 9312 4072 9364 4078
rect 9496 4072 9548 4078
rect 9312 4014 9364 4020
rect 9402 4040 9458 4049
rect 8852 4004 8904 4010
rect 8852 3946 8904 3952
rect 9324 3942 9352 4014
rect 9496 4014 9548 4020
rect 9680 4072 9732 4078
rect 9784 4049 9812 4490
rect 9862 4312 9918 4321
rect 9862 4247 9918 4256
rect 9680 4014 9732 4020
rect 9770 4040 9826 4049
rect 9402 3975 9458 3984
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9324 3641 9352 3878
rect 9310 3632 9366 3641
rect 8760 3596 8812 3602
rect 9310 3567 9366 3576
rect 8760 3538 8812 3544
rect 9416 3369 9444 3975
rect 9508 3738 9536 4014
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9402 3360 9458 3369
rect 9010 3292 9318 3301
rect 9402 3295 9458 3304
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 9508 2972 9536 3674
rect 9692 3398 9720 4014
rect 9770 3975 9826 3984
rect 9772 3936 9824 3942
rect 9770 3904 9772 3913
rect 9824 3904 9826 3913
rect 9770 3839 9826 3848
rect 9876 3720 9904 4247
rect 9784 3692 9904 3720
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9588 2984 9640 2990
rect 9508 2944 9588 2972
rect 9588 2926 9640 2932
rect 9784 2854 9812 3692
rect 9862 3632 9918 3641
rect 9862 3567 9864 3576
rect 9916 3567 9918 3576
rect 9864 3538 9916 3544
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9876 2582 9904 2994
rect 9864 2576 9916 2582
rect 9864 2518 9916 2524
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 9404 2440 9456 2446
rect 9218 2408 9274 2417
rect 8668 2372 8720 2378
rect 9404 2382 9456 2388
rect 9218 2343 9220 2352
rect 8668 2314 8720 2320
rect 9272 2343 9274 2352
rect 9220 2314 9272 2320
rect 8576 1080 8628 1086
rect 8576 1022 8628 1028
rect 8680 56 8708 2314
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 9416 56 9444 2382
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9692 2038 9720 2246
rect 9680 2032 9732 2038
rect 9680 1974 9732 1980
rect 9784 1465 9812 2450
rect 9770 1456 9826 1465
rect 9770 1391 9826 1400
rect 9968 1290 9996 5510
rect 10046 5471 10102 5480
rect 10060 5234 10088 5471
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 10060 4298 10088 4966
rect 10060 4270 10180 4298
rect 10152 3602 10180 4270
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10048 3528 10100 3534
rect 10244 3482 10272 6734
rect 10428 4865 10456 7754
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10520 5710 10548 6258
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10508 5296 10560 5302
rect 10508 5238 10560 5244
rect 10414 4856 10470 4865
rect 10414 4791 10470 4800
rect 10520 4486 10548 5238
rect 10612 4826 10640 10814
rect 10704 8294 10732 11194
rect 10784 10736 10836 10742
rect 10784 10678 10836 10684
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10704 6798 10732 7822
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10796 6662 10824 10678
rect 10876 9784 10928 9790
rect 10876 9726 10928 9732
rect 10888 8634 10916 9726
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10980 8378 11008 11194
rect 11256 9722 11284 11194
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11336 9308 11388 9314
rect 11336 9250 11388 9256
rect 11244 9104 11296 9110
rect 11058 9072 11114 9081
rect 11244 9046 11296 9052
rect 11058 9007 11114 9016
rect 11072 8548 11100 9007
rect 11256 8566 11284 9046
rect 11244 8560 11296 8566
rect 11072 8520 11192 8548
rect 10980 8350 11100 8378
rect 10966 8120 11022 8129
rect 10966 8055 11022 8064
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10704 4622 10732 5170
rect 10980 4826 11008 8055
rect 11072 7274 11100 8350
rect 11164 7886 11192 8520
rect 11244 8502 11296 8508
rect 11348 8498 11376 9250
rect 11428 9240 11480 9246
rect 11428 9182 11480 9188
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 11072 6361 11100 6666
rect 11058 6352 11114 6361
rect 11058 6287 11114 6296
rect 11164 5658 11192 7686
rect 11072 5630 11192 5658
rect 11072 5409 11100 5630
rect 11256 5574 11284 8366
rect 11336 8288 11388 8294
rect 11440 8265 11468 9182
rect 11532 8362 11560 11194
rect 11808 9790 11836 11194
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 11796 9784 11848 9790
rect 11796 9726 11848 9732
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11520 8356 11572 8362
rect 11520 8298 11572 8304
rect 11336 8230 11388 8236
rect 11426 8256 11482 8265
rect 11348 7546 11376 8230
rect 11426 8191 11482 8200
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11428 7744 11480 7750
rect 11428 7686 11480 7692
rect 11440 7546 11468 7686
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11532 7410 11560 7890
rect 11624 7562 11652 9318
rect 11716 8362 11744 9658
rect 11796 8900 11848 8906
rect 11796 8842 11848 8848
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 11624 7534 11744 7562
rect 11612 7472 11664 7478
rect 11612 7414 11664 7420
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11348 7002 11376 7346
rect 11624 7206 11652 7414
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11336 6996 11388 7002
rect 11336 6938 11388 6944
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11058 5400 11114 5409
rect 11164 5386 11192 5510
rect 11164 5358 11284 5386
rect 11348 5370 11376 6802
rect 11440 6798 11468 7142
rect 11532 6798 11560 7142
rect 11716 6882 11744 7534
rect 11624 6854 11744 6882
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11624 6644 11652 6854
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11532 6616 11652 6644
rect 11058 5335 11114 5344
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 10428 4146 10456 4422
rect 11164 4282 11192 4558
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11256 4146 11284 5358
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 11440 4282 11468 4966
rect 11428 4276 11480 4282
rect 11428 4218 11480 4224
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10414 3904 10470 3913
rect 10414 3839 10470 3848
rect 10428 3618 10456 3839
rect 10336 3602 10456 3618
rect 10324 3596 10456 3602
rect 10376 3590 10456 3596
rect 10324 3538 10376 3544
rect 10048 3470 10100 3476
rect 10060 2854 10088 3470
rect 10152 3454 10272 3482
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10152 2530 10180 3454
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 10244 2650 10272 3334
rect 10428 2774 10456 3590
rect 10336 2746 10456 2774
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10152 2502 10272 2530
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 9956 1284 10008 1290
rect 9956 1226 10008 1232
rect 10152 56 10180 2382
rect 10244 1737 10272 2502
rect 10336 2310 10364 2746
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 10230 1728 10286 1737
rect 10230 1663 10286 1672
rect 10520 882 10548 4014
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 10980 3738 11008 3946
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 11532 3670 11560 6616
rect 11716 6458 11744 6734
rect 11808 6662 11836 8842
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 11428 3392 11480 3398
rect 11428 3334 11480 3340
rect 10612 3058 10640 3334
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10704 2774 10732 2994
rect 10704 2746 10824 2774
rect 10796 1494 10824 2746
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 10784 1488 10836 1494
rect 10784 1430 10836 1436
rect 10508 876 10560 882
rect 10508 818 10560 824
rect 10888 56 10916 2382
rect 10980 2106 11008 3334
rect 11440 3126 11468 3334
rect 11428 3120 11480 3126
rect 11428 3062 11480 3068
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 11072 2446 11100 2518
rect 11348 2514 11376 2790
rect 11624 2774 11652 6190
rect 11794 5944 11850 5953
rect 11794 5879 11850 5888
rect 11808 5778 11836 5879
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 11900 5386 11928 10134
rect 12084 8634 12112 11194
rect 12164 9784 12216 9790
rect 12164 9726 12216 9732
rect 12176 8634 12204 9726
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12268 8498 12296 9522
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12360 8022 12388 11194
rect 12530 10432 12586 10441
rect 12530 10367 12586 10376
rect 12544 10033 12572 10367
rect 12530 10024 12586 10033
rect 12530 9959 12586 9968
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12452 8430 12480 9590
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12348 8016 12400 8022
rect 12348 7958 12400 7964
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 11992 7177 12020 7822
rect 12084 7721 12112 7822
rect 12070 7712 12126 7721
rect 12070 7647 12126 7656
rect 11978 7168 12034 7177
rect 11978 7103 12034 7112
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 11992 6458 12020 6802
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 12084 6254 12112 7647
rect 12162 7576 12218 7585
rect 12162 7511 12218 7520
rect 12176 7342 12204 7511
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12268 6730 12296 7822
rect 12636 7546 12664 11194
rect 12806 10024 12862 10033
rect 12806 9959 12862 9968
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12728 9042 12756 9318
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12820 8634 12848 9959
rect 12912 9722 12940 11194
rect 13188 10554 13216 11194
rect 13096 10526 13216 10554
rect 12990 10296 13046 10305
rect 12990 10231 13046 10240
rect 13004 9761 13032 10231
rect 13096 9790 13124 10526
rect 13084 9784 13136 9790
rect 12990 9752 13046 9761
rect 12900 9716 12952 9722
rect 13084 9726 13136 9732
rect 13174 9752 13230 9761
rect 12990 9687 13046 9696
rect 13174 9687 13230 9696
rect 12900 9658 12952 9664
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 13004 8838 13032 9590
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 13096 8566 13124 9522
rect 13188 8634 13216 9687
rect 13360 9240 13412 9246
rect 13360 9182 13412 9188
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 13280 8498 13308 8774
rect 13372 8498 13400 9182
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12820 7834 12848 8026
rect 12992 7880 13044 7886
rect 12912 7840 12992 7868
rect 12912 7834 12940 7840
rect 12728 7806 12940 7834
rect 12992 7822 13044 7828
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12544 7449 12572 7482
rect 12530 7440 12586 7449
rect 12440 7404 12492 7410
rect 12530 7375 12586 7384
rect 12624 7404 12676 7410
rect 12440 7346 12492 7352
rect 12624 7346 12676 7352
rect 12256 6724 12308 6730
rect 12176 6684 12256 6712
rect 12072 6248 12124 6254
rect 12072 6190 12124 6196
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11992 5778 12020 6054
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11808 5358 11928 5386
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11532 2746 11652 2774
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 10968 2100 11020 2106
rect 10968 2042 11020 2048
rect 11532 1902 11560 2746
rect 11716 2446 11744 3334
rect 11808 3194 11836 5358
rect 11888 5228 11940 5234
rect 11992 5216 12020 5510
rect 12176 5234 12204 6684
rect 12256 6666 12308 6672
rect 12452 6662 12480 7346
rect 12636 7002 12664 7346
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12636 6662 12664 6734
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 12360 6254 12388 6326
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12256 6180 12308 6186
rect 12256 6122 12308 6128
rect 12268 6066 12296 6122
rect 12268 6038 12388 6066
rect 12360 5914 12388 6038
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12268 5710 12296 5850
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12348 5636 12400 5642
rect 12348 5578 12400 5584
rect 11940 5188 12020 5216
rect 12164 5228 12216 5234
rect 11888 5170 11940 5176
rect 12164 5170 12216 5176
rect 12360 5166 12388 5578
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 12256 5092 12308 5098
rect 12256 5034 12308 5040
rect 12268 4826 12296 5034
rect 12452 4842 12480 6598
rect 12544 5370 12572 6598
rect 12728 5778 12756 7806
rect 13096 7478 13124 7822
rect 13084 7472 13136 7478
rect 13084 7414 13136 7420
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12360 4814 12480 4842
rect 12360 4298 12388 4814
rect 12360 4270 12480 4298
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11808 2990 11836 3130
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11900 2650 11928 3470
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 11980 2372 12032 2378
rect 11980 2314 12032 2320
rect 11520 1896 11572 1902
rect 11520 1838 11572 1844
rect 11624 56 11652 2314
rect 11992 1873 12020 2314
rect 11978 1864 12034 1873
rect 11978 1799 12034 1808
rect 12360 56 12388 2382
rect 12452 1766 12480 4270
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12636 3194 12664 3946
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12728 2774 12756 5714
rect 12820 3670 12848 7278
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 4622 12940 7142
rect 13188 6746 13216 8366
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13280 7478 13308 8026
rect 13372 7993 13400 8026
rect 13358 7984 13414 7993
rect 13358 7919 13414 7928
rect 13464 7546 13492 11194
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 13556 8566 13584 8842
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13544 8424 13596 8430
rect 13648 8401 13676 8434
rect 13544 8366 13596 8372
rect 13634 8392 13690 8401
rect 13556 8294 13584 8366
rect 13740 8362 13768 11194
rect 14016 10033 14044 11194
rect 14002 10024 14058 10033
rect 14002 9959 14058 9968
rect 14292 9761 14320 11194
rect 14464 9784 14516 9790
rect 14278 9752 14334 9761
rect 14464 9726 14516 9732
rect 14278 9687 14334 9696
rect 14096 9444 14148 9450
rect 14096 9386 14148 9392
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13634 8327 13690 8336
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13268 7472 13320 7478
rect 13268 7414 13320 7420
rect 13450 7440 13506 7449
rect 13450 7375 13506 7384
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13358 7304 13414 7313
rect 13280 6866 13308 7278
rect 13358 7239 13414 7248
rect 13372 7206 13400 7239
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13464 7154 13492 7375
rect 13464 7126 13584 7154
rect 13358 6896 13414 6905
rect 13268 6860 13320 6866
rect 13358 6831 13414 6840
rect 13268 6802 13320 6808
rect 13372 6798 13400 6831
rect 13096 6718 13216 6746
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13268 6724 13320 6730
rect 13096 6662 13124 6718
rect 13268 6666 13320 6672
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 12990 5944 13046 5953
rect 12990 5879 13046 5888
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 12808 3664 12860 3670
rect 12808 3606 12860 3612
rect 12912 3058 12940 4558
rect 13004 4010 13032 5879
rect 13188 5574 13216 6598
rect 13280 6390 13308 6666
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 13556 6322 13584 7126
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13176 5568 13228 5574
rect 13096 5528 13176 5556
rect 13096 5166 13124 5528
rect 13176 5510 13228 5516
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 13372 4570 13400 6258
rect 13464 4758 13492 6258
rect 13648 5642 13676 8230
rect 13726 7712 13782 7721
rect 13726 7647 13782 7656
rect 13740 7449 13768 7647
rect 13726 7440 13782 7449
rect 13832 7410 13860 8842
rect 14108 8362 14136 9386
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 13726 7375 13782 7384
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 14108 7342 14136 8026
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14096 7336 14148 7342
rect 13726 7304 13782 7313
rect 14200 7324 14228 7686
rect 14292 7546 14320 8434
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14384 8129 14412 8366
rect 14370 8120 14426 8129
rect 14370 8055 14426 8064
rect 14372 8016 14424 8022
rect 14372 7958 14424 7964
rect 14384 7750 14412 7958
rect 14372 7744 14424 7750
rect 14372 7686 14424 7692
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14476 7426 14504 9726
rect 14568 8634 14596 11194
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14648 9104 14700 9110
rect 14648 9046 14700 9052
rect 14660 8634 14688 9046
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14752 8362 14780 9862
rect 14740 8356 14792 8362
rect 14740 8298 14792 8304
rect 14844 7546 14872 11194
rect 15120 9926 15148 11194
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15396 9738 15424 11194
rect 14936 9710 15424 9738
rect 14936 8634 14964 9710
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 14924 8356 14976 8362
rect 14924 8298 14976 8304
rect 14936 7886 14964 8298
rect 15292 8288 15344 8294
rect 15290 8256 15292 8265
rect 15344 8256 15346 8265
rect 15290 8191 15346 8200
rect 15106 8120 15162 8129
rect 15106 8055 15162 8064
rect 15120 7954 15148 8055
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 15198 7848 15254 7857
rect 15198 7783 15254 7792
rect 15212 7750 15240 7783
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 14476 7398 14872 7426
rect 14556 7336 14608 7342
rect 14200 7296 14556 7324
rect 14096 7278 14148 7284
rect 14556 7278 14608 7284
rect 13726 7239 13782 7248
rect 13740 6934 13768 7239
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13818 7032 13874 7041
rect 13950 7035 14258 7044
rect 13818 6967 13874 6976
rect 14370 7032 14426 7041
rect 14370 6967 14426 6976
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 13832 6730 13860 6967
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 14200 6186 14228 6802
rect 14384 6390 14412 6967
rect 14462 6896 14518 6905
rect 14462 6831 14518 6840
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14384 6254 14412 6326
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 14476 6089 14504 6831
rect 14462 6080 14518 6089
rect 13950 6012 14258 6021
rect 14462 6015 14518 6024
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 14462 5944 14518 5953
rect 14462 5879 14518 5888
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13636 5636 13688 5642
rect 13636 5578 13688 5584
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13740 5370 13768 5510
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13726 4992 13782 5001
rect 13726 4927 13782 4936
rect 13542 4856 13598 4865
rect 13542 4791 13598 4800
rect 13452 4752 13504 4758
rect 13452 4694 13504 4700
rect 13372 4542 13492 4570
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 13096 4282 13124 4422
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 12992 4004 13044 4010
rect 12992 3946 13044 3952
rect 13188 3534 13216 4082
rect 13464 3942 13492 4542
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13280 3126 13308 3878
rect 13268 3120 13320 3126
rect 13268 3062 13320 3068
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 12728 2746 12848 2774
rect 12820 2650 12848 2746
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 13004 2310 13032 2586
rect 12992 2304 13044 2310
rect 12992 2246 13044 2252
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 12440 1760 12492 1766
rect 12440 1702 12492 1708
rect 13096 56 13124 2246
rect 13372 950 13400 3878
rect 13556 3738 13584 4791
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13648 4214 13676 4626
rect 13740 4622 13768 4927
rect 13832 4826 13860 5714
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 14280 5704 14332 5710
rect 14332 5652 14412 5658
rect 14280 5646 14412 5652
rect 13924 5234 13952 5646
rect 14292 5630 14412 5646
rect 14278 5536 14334 5545
rect 14278 5471 14334 5480
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 14292 4758 14320 5471
rect 14384 5370 14412 5630
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14384 5166 14412 5306
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 14280 4752 14332 4758
rect 14280 4694 14332 4700
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13820 4548 13872 4554
rect 13820 4490 13872 4496
rect 13832 4214 13860 4490
rect 13636 4208 13688 4214
rect 13636 4150 13688 4156
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 14200 4146 14228 4694
rect 14384 4690 14412 5102
rect 14372 4684 14424 4690
rect 14372 4626 14424 4632
rect 14476 4321 14504 5879
rect 14462 4312 14518 4321
rect 14462 4247 14518 4256
rect 14372 4208 14424 4214
rect 14372 4150 14424 4156
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13740 3602 13768 3946
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13556 2990 13584 3538
rect 14384 3369 14412 4150
rect 14568 3670 14596 7142
rect 14646 6896 14702 6905
rect 14646 6831 14702 6840
rect 14740 6860 14792 6866
rect 14660 6361 14688 6831
rect 14740 6802 14792 6808
rect 14646 6352 14702 6361
rect 14646 6287 14702 6296
rect 14752 5794 14780 6802
rect 14844 6730 14872 7398
rect 15396 7206 15424 8366
rect 15488 7546 15516 8910
rect 15476 7540 15528 7546
rect 15580 7528 15608 9590
rect 15672 8090 15700 11194
rect 15844 8560 15896 8566
rect 15844 8502 15896 8508
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15672 7721 15700 7890
rect 15658 7712 15714 7721
rect 15658 7647 15714 7656
rect 15580 7500 15700 7528
rect 15476 7482 15528 7488
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15384 7200 15436 7206
rect 14922 7168 14978 7177
rect 15384 7142 15436 7148
rect 14922 7103 14978 7112
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 14936 6338 14964 7103
rect 15488 7002 15516 7346
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15488 6633 15516 6734
rect 15474 6624 15530 6633
rect 15010 6556 15318 6565
rect 15474 6559 15530 6568
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 14936 6310 15056 6338
rect 14832 6180 14884 6186
rect 14832 6122 14884 6128
rect 14924 6180 14976 6186
rect 14924 6122 14976 6128
rect 14844 5846 14872 6122
rect 14936 5914 14964 6122
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 14660 5766 14780 5794
rect 14832 5840 14884 5846
rect 14832 5782 14884 5788
rect 14556 3664 14608 3670
rect 14556 3606 14608 3612
rect 14370 3360 14426 3369
rect 14370 3295 14426 3304
rect 14554 3224 14610 3233
rect 14554 3159 14610 3168
rect 13726 3088 13782 3097
rect 13726 3023 13782 3032
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 13740 2854 13768 3023
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 13820 2304 13872 2310
rect 13820 2246 13872 2252
rect 13360 944 13412 950
rect 13360 886 13412 892
rect 13832 56 13860 2246
rect 14476 1358 14504 2858
rect 14568 2825 14596 3159
rect 14554 2816 14610 2825
rect 14554 2751 14610 2760
rect 14660 2774 14688 5766
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14752 5234 14780 5646
rect 15028 5556 15056 6310
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15212 5710 15240 6190
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 14936 5528 15056 5556
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14752 4554 14780 5170
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 14740 4548 14792 4554
rect 14740 4490 14792 4496
rect 14660 2746 14780 2774
rect 14556 2304 14608 2310
rect 14556 2246 14608 2252
rect 14464 1352 14516 1358
rect 14464 1294 14516 1300
rect 14568 56 14596 2246
rect 14752 1698 14780 2746
rect 14844 1766 14872 4966
rect 14936 4593 14964 5528
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 15488 5273 15516 6258
rect 15290 5264 15346 5273
rect 15290 5199 15346 5208
rect 15474 5264 15530 5273
rect 15474 5199 15530 5208
rect 15016 5160 15068 5166
rect 15016 5102 15068 5108
rect 14922 4584 14978 4593
rect 14922 4519 14978 4528
rect 15028 4468 15056 5102
rect 15304 5098 15332 5199
rect 15292 5092 15344 5098
rect 15292 5034 15344 5040
rect 15476 4616 15528 4622
rect 15198 4584 15254 4593
rect 15476 4558 15528 4564
rect 15198 4519 15200 4528
rect 15252 4519 15254 4528
rect 15200 4490 15252 4496
rect 14936 4440 15056 4468
rect 14936 2854 14964 4440
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 15488 4146 15516 4558
rect 15580 4214 15608 7346
rect 15672 6662 15700 7500
rect 15764 7478 15792 8434
rect 15752 7472 15804 7478
rect 15752 7414 15804 7420
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15856 5953 15884 8502
rect 15948 7546 15976 11194
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 16040 7002 16068 8978
rect 16224 8634 16252 11194
rect 16394 9752 16450 9761
rect 16394 9687 16450 9696
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16132 7410 16160 8434
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16224 7750 16252 7822
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16210 7304 16266 7313
rect 16210 7239 16266 7248
rect 16224 7002 16252 7239
rect 16028 6996 16080 7002
rect 16028 6938 16080 6944
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 16316 6934 16344 8978
rect 16408 8634 16436 9687
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16500 8430 16528 11194
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16408 7313 16436 7686
rect 16488 7336 16540 7342
rect 16394 7304 16450 7313
rect 16488 7278 16540 7284
rect 16394 7239 16450 7248
rect 16304 6928 16356 6934
rect 16304 6870 16356 6876
rect 16316 6254 16344 6870
rect 16304 6248 16356 6254
rect 16304 6190 16356 6196
rect 15842 5944 15898 5953
rect 15842 5879 15898 5888
rect 16302 5672 16358 5681
rect 16302 5607 16358 5616
rect 16026 5400 16082 5409
rect 16026 5335 16082 5344
rect 16040 4865 16068 5335
rect 16316 4865 16344 5607
rect 16026 4856 16082 4865
rect 16026 4791 16082 4800
rect 16302 4856 16358 4865
rect 16302 4791 16358 4800
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 15856 4321 15884 4626
rect 16028 4616 16080 4622
rect 16316 4604 16344 4791
rect 16080 4576 16344 4604
rect 16028 4558 16080 4564
rect 15842 4312 15898 4321
rect 15842 4247 15898 4256
rect 15568 4208 15620 4214
rect 15568 4150 15620 4156
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 15010 3227 15318 3236
rect 15396 2990 15424 3470
rect 15764 3398 15792 4082
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16026 3632 16082 3641
rect 16026 3567 16082 3576
rect 15752 3392 15804 3398
rect 16040 3369 16068 3567
rect 16120 3392 16172 3398
rect 15752 3334 15804 3340
rect 16026 3360 16082 3369
rect 16120 3334 16172 3340
rect 16026 3295 16082 3304
rect 16028 3052 16080 3058
rect 16028 2994 16080 3000
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 14924 2848 14976 2854
rect 16040 2825 16068 2994
rect 14924 2790 14976 2796
rect 16026 2816 16082 2825
rect 16026 2751 16082 2760
rect 16132 2582 16160 3334
rect 16120 2576 16172 2582
rect 15750 2544 15806 2553
rect 16408 2553 16436 3878
rect 16500 3398 16528 7278
rect 16592 3942 16620 9522
rect 16776 8362 16804 11194
rect 17052 9761 17080 11194
rect 17224 10872 17276 10878
rect 17224 10814 17276 10820
rect 17236 10334 17264 10814
rect 17224 10328 17276 10334
rect 17224 10270 17276 10276
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17236 9926 17264 10066
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17038 9752 17094 9761
rect 17038 9687 17094 9696
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16684 5914 16712 6190
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16580 3528 16632 3534
rect 16632 3488 16712 3516
rect 16580 3470 16632 3476
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16592 2582 16620 2994
rect 16684 2990 16712 3488
rect 16776 3097 16804 7346
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16868 6866 16896 7278
rect 16960 6934 16988 9318
rect 16948 6928 17000 6934
rect 16948 6870 17000 6876
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 16960 6798 16988 6870
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16868 4434 16896 6258
rect 17052 5710 17080 9522
rect 17328 8634 17356 11194
rect 17408 10736 17460 10742
rect 17408 10678 17460 10684
rect 17420 10130 17448 10678
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17500 8560 17552 8566
rect 17500 8502 17552 8508
rect 17408 7812 17460 7818
rect 17408 7754 17460 7760
rect 17224 7744 17276 7750
rect 17224 7686 17276 7692
rect 17236 7410 17264 7686
rect 17420 7449 17448 7754
rect 17406 7440 17462 7449
rect 17224 7404 17276 7410
rect 17406 7375 17462 7384
rect 17224 7346 17276 7352
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17420 7002 17448 7142
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17420 6866 17448 6938
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17236 6322 17264 6734
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 17040 5704 17092 5710
rect 16946 5672 17002 5681
rect 17040 5646 17092 5652
rect 16946 5607 17002 5616
rect 17224 5636 17276 5642
rect 16960 5370 16988 5607
rect 17224 5578 17276 5584
rect 16948 5364 17000 5370
rect 16948 5306 17000 5312
rect 17236 5273 17264 5578
rect 17222 5264 17278 5273
rect 17222 5199 17278 5208
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 16960 4554 16988 5102
rect 16948 4548 17000 4554
rect 16948 4490 17000 4496
rect 17222 4448 17278 4457
rect 16868 4406 17172 4434
rect 16856 4208 16908 4214
rect 16856 4150 16908 4156
rect 16762 3088 16818 3097
rect 16762 3023 16818 3032
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 16868 2650 16896 4150
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 16960 3058 16988 3470
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 16580 2576 16632 2582
rect 16120 2518 16172 2524
rect 16394 2544 16450 2553
rect 15750 2479 15806 2488
rect 16580 2518 16632 2524
rect 16394 2479 16450 2488
rect 15764 2446 15792 2479
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 14832 1760 14884 1766
rect 14832 1702 14884 1708
rect 14936 1698 14964 2382
rect 15384 2304 15436 2310
rect 15384 2246 15436 2252
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 14740 1692 14792 1698
rect 14740 1634 14792 1640
rect 14924 1692 14976 1698
rect 14924 1634 14976 1640
rect 15396 1170 15424 2246
rect 15672 1902 15700 2382
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 15660 1896 15712 1902
rect 15660 1838 15712 1844
rect 15304 1142 15424 1170
rect 15304 56 15332 1142
rect 16040 56 16068 2246
rect 16224 649 16252 2382
rect 16592 1562 16620 2518
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 16580 1556 16632 1562
rect 16580 1498 16632 1504
rect 16210 640 16266 649
rect 16210 575 16266 584
rect 16776 56 16804 2246
rect 16960 785 16988 2994
rect 17144 2378 17172 4406
rect 17222 4383 17278 4392
rect 17236 4282 17264 4383
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17236 3602 17264 4014
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17420 2650 17448 3470
rect 17512 3194 17540 8502
rect 17604 8430 17632 11194
rect 17880 9110 17908 11194
rect 18052 9444 18104 9450
rect 18052 9386 18104 9392
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17590 7848 17646 7857
rect 17590 7783 17646 7792
rect 17604 7750 17632 7783
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 17604 7585 17632 7686
rect 17590 7576 17646 7585
rect 17590 7511 17646 7520
rect 17696 7041 17724 8570
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17682 7032 17738 7041
rect 17682 6967 17738 6976
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17696 4622 17724 5170
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 17604 3618 17632 4558
rect 17788 3738 17816 8434
rect 18064 7546 18092 9386
rect 18156 8498 18184 11194
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18432 7954 18460 11194
rect 18512 9104 18564 9110
rect 18512 9046 18564 9052
rect 18524 8106 18552 9046
rect 18708 8498 18736 11194
rect 18878 9752 18934 9761
rect 18878 9687 18934 9696
rect 18788 9104 18840 9110
rect 18788 9046 18840 9052
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18800 8294 18828 9046
rect 18788 8288 18840 8294
rect 18788 8230 18840 8236
rect 18524 8078 18644 8106
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18328 7812 18380 7818
rect 18328 7754 18380 7760
rect 18142 7576 18198 7585
rect 18052 7540 18104 7546
rect 18340 7546 18368 7754
rect 18142 7511 18198 7520
rect 18328 7540 18380 7546
rect 18052 7482 18104 7488
rect 17960 7472 18012 7478
rect 17960 7414 18012 7420
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 17880 7002 17908 7278
rect 17868 6996 17920 7002
rect 17868 6938 17920 6944
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17880 6458 17908 6802
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 17880 5817 17908 6054
rect 17866 5808 17922 5817
rect 17866 5743 17922 5752
rect 17972 4146 18000 7414
rect 18064 6780 18092 7482
rect 18156 7177 18184 7511
rect 18328 7482 18380 7488
rect 18236 7200 18288 7206
rect 18142 7168 18198 7177
rect 18236 7142 18288 7148
rect 18142 7103 18198 7112
rect 18144 6792 18196 6798
rect 18064 6752 18144 6780
rect 18144 6734 18196 6740
rect 18050 6216 18106 6225
rect 18050 6151 18106 6160
rect 18064 5817 18092 6151
rect 18050 5808 18106 5817
rect 18050 5743 18106 5752
rect 18248 5234 18276 7142
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 18432 5642 18460 6734
rect 18420 5636 18472 5642
rect 18420 5578 18472 5584
rect 18524 5574 18552 7822
rect 18616 7410 18644 8078
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18800 5914 18828 8230
rect 18892 7410 18920 9687
rect 18984 8022 19012 11194
rect 19154 10024 19210 10033
rect 19154 9959 19210 9968
rect 19062 8120 19118 8129
rect 19062 8055 19118 8064
rect 18972 8016 19024 8022
rect 18972 7958 19024 7964
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 18984 7478 19012 7822
rect 18972 7472 19024 7478
rect 18972 7414 19024 7420
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 19076 7342 19104 8055
rect 19168 7410 19196 9959
rect 19260 7886 19288 11194
rect 19536 9761 19564 11194
rect 19812 10033 19840 11194
rect 19798 10024 19854 10033
rect 19798 9959 19854 9968
rect 19522 9752 19578 9761
rect 19432 9716 19484 9722
rect 19522 9687 19578 9696
rect 20088 9674 20116 11194
rect 20364 9722 20392 11194
rect 20640 9738 20668 11194
rect 19432 9658 19484 9664
rect 19340 8832 19392 8838
rect 19444 8809 19472 9658
rect 19812 9646 20116 9674
rect 20352 9716 20404 9722
rect 20640 9710 20760 9738
rect 20352 9658 20404 9664
rect 19708 9580 19760 9586
rect 19708 9522 19760 9528
rect 19720 9246 19748 9522
rect 19616 9240 19668 9246
rect 19616 9182 19668 9188
rect 19708 9240 19760 9246
rect 19708 9182 19760 9188
rect 19628 9081 19656 9182
rect 19614 9072 19670 9081
rect 19614 9007 19670 9016
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19340 8774 19392 8780
rect 19430 8800 19486 8809
rect 19352 8129 19380 8774
rect 19430 8735 19486 8744
rect 19536 8242 19564 8910
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19720 8265 19748 8570
rect 19444 8214 19564 8242
rect 19706 8256 19762 8265
rect 19338 8120 19394 8129
rect 19444 8090 19472 8214
rect 19706 8191 19762 8200
rect 19706 8120 19762 8129
rect 19338 8055 19394 8064
rect 19432 8084 19484 8090
rect 19706 8055 19708 8064
rect 19432 8026 19484 8032
rect 19760 8055 19762 8064
rect 19708 8026 19760 8032
rect 19812 7886 19840 9646
rect 20074 8664 20130 8673
rect 20074 8599 20130 8608
rect 20088 8430 20116 8599
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20076 8424 20128 8430
rect 20076 8366 20128 8372
rect 20352 8288 20404 8294
rect 20352 8230 20404 8236
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 19950 8188 20258 8197
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 20364 8090 20392 8230
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 19904 7886 19932 8026
rect 19982 7984 20038 7993
rect 19982 7919 20038 7928
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 19260 6662 19288 7278
rect 18972 6656 19024 6662
rect 18892 6616 18972 6644
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18602 5536 18658 5545
rect 18892 5522 18920 6616
rect 18972 6598 19024 6604
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 18602 5471 18658 5480
rect 18800 5494 18920 5522
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 18064 4282 18092 5102
rect 18248 4622 18276 5170
rect 18616 5030 18644 5471
rect 18604 5024 18656 5030
rect 18604 4966 18656 4972
rect 18328 4752 18380 4758
rect 18328 4694 18380 4700
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 18340 4486 18368 4694
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18052 4276 18104 4282
rect 18052 4218 18104 4224
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 17776 3732 17828 3738
rect 17776 3674 17828 3680
rect 18144 3664 18196 3670
rect 17604 3590 17908 3618
rect 18144 3606 18196 3612
rect 17500 3188 17552 3194
rect 17500 3130 17552 3136
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 17512 2514 17540 2926
rect 17604 2854 17632 3590
rect 17880 3534 17908 3590
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17682 3224 17738 3233
rect 17788 3194 17816 3470
rect 18156 3369 18184 3606
rect 18616 3602 18644 3946
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 18142 3360 18198 3369
rect 18142 3295 18198 3304
rect 18156 3194 18184 3295
rect 18248 3194 18276 3538
rect 18326 3360 18382 3369
rect 18326 3295 18382 3304
rect 17682 3159 17738 3168
rect 17776 3188 17828 3194
rect 17592 2848 17644 2854
rect 17592 2790 17644 2796
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 17132 2372 17184 2378
rect 17132 2314 17184 2320
rect 17696 2310 17724 3159
rect 17776 3130 17828 3136
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18340 2825 18368 3295
rect 18326 2816 18382 2825
rect 18326 2751 18382 2760
rect 18800 2446 18828 5494
rect 18984 5234 19012 6258
rect 19246 5536 19302 5545
rect 19246 5471 19302 5480
rect 19260 5234 19288 5471
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 18984 4214 19012 5170
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 19352 4978 19380 7686
rect 19996 7562 20024 7919
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 19536 7546 20024 7562
rect 19524 7540 20024 7546
rect 19576 7534 20024 7540
rect 19524 7482 19576 7488
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 19812 6798 19840 7346
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 20364 6882 20392 7822
rect 20456 7546 20484 8230
rect 20548 8022 20576 8434
rect 20628 8356 20680 8362
rect 20628 8298 20680 8304
rect 20640 8022 20668 8298
rect 20536 8016 20588 8022
rect 20536 7958 20588 7964
rect 20628 8016 20680 8022
rect 20628 7958 20680 7964
rect 20534 7576 20590 7585
rect 20444 7540 20496 7546
rect 20534 7511 20536 7520
rect 20444 7482 20496 7488
rect 20588 7511 20590 7520
rect 20536 7482 20588 7488
rect 20732 7410 20760 9710
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20824 7410 20852 9658
rect 20916 8616 20944 11194
rect 21192 9874 21220 11194
rect 21192 9846 21404 9874
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 21180 8628 21232 8634
rect 20916 8588 21036 8616
rect 21008 8430 21036 8588
rect 21180 8570 21232 8576
rect 20996 8424 21048 8430
rect 20996 8366 21048 8372
rect 20994 8120 21050 8129
rect 20994 8055 21050 8064
rect 20904 7880 20956 7886
rect 21008 7857 21036 8055
rect 21192 7857 21220 8570
rect 21376 8498 21404 9846
rect 21364 8492 21416 8498
rect 21468 8480 21496 11194
rect 21548 9784 21600 9790
rect 21548 9726 21600 9732
rect 21560 8634 21588 9726
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21744 8566 21772 11194
rect 21916 9036 21968 9042
rect 21916 8978 21968 8984
rect 21928 8838 21956 8978
rect 21916 8832 21968 8838
rect 21916 8774 21968 8780
rect 22020 8634 22048 11194
rect 22192 9308 22244 9314
rect 22192 9250 22244 9256
rect 22100 9036 22152 9042
rect 22100 8978 22152 8984
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 21640 8560 21692 8566
rect 21640 8502 21692 8508
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 21548 8492 21600 8498
rect 21468 8452 21548 8480
rect 21364 8434 21416 8440
rect 21548 8434 21600 8440
rect 21652 8022 21680 8502
rect 22112 8362 22140 8978
rect 21916 8356 21968 8362
rect 21916 8298 21968 8304
rect 22100 8356 22152 8362
rect 22100 8298 22152 8304
rect 21640 8016 21692 8022
rect 21640 7958 21692 7964
rect 21548 7948 21600 7954
rect 21548 7890 21600 7896
rect 20904 7822 20956 7828
rect 20994 7848 21050 7857
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20916 7018 20944 7822
rect 20994 7783 21050 7792
rect 21178 7848 21234 7857
rect 21178 7783 21234 7792
rect 21560 7721 21588 7890
rect 21546 7712 21602 7721
rect 21010 7644 21318 7653
rect 21546 7647 21602 7656
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 20994 7032 21050 7041
rect 20720 6996 20772 7002
rect 20916 6990 20994 7018
rect 20994 6967 21050 6976
rect 20720 6938 20772 6944
rect 20628 6928 20680 6934
rect 20364 6876 20628 6882
rect 20364 6870 20680 6876
rect 20364 6854 20668 6870
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19800 6792 19852 6798
rect 19800 6734 19852 6740
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 19536 5545 19564 6734
rect 19706 6488 19762 6497
rect 19706 6423 19762 6432
rect 19720 6118 19748 6423
rect 19708 6112 19760 6118
rect 19708 6054 19760 6060
rect 19812 5778 19840 6734
rect 20180 6322 20208 6734
rect 20364 6458 20392 6854
rect 20444 6656 20496 6662
rect 20444 6598 20496 6604
rect 20626 6624 20682 6633
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20168 6316 20220 6322
rect 20168 6258 20220 6264
rect 20352 6180 20404 6186
rect 20352 6122 20404 6128
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 19522 5536 19578 5545
rect 19522 5471 19578 5480
rect 19430 5400 19486 5409
rect 19430 5335 19486 5344
rect 19444 5166 19472 5335
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19168 4758 19196 4966
rect 19352 4950 19472 4978
rect 19444 4826 19472 4950
rect 19536 4865 19564 5471
rect 19812 5188 20116 5216
rect 19812 5001 19840 5188
rect 19982 5128 20038 5137
rect 20088 5114 20116 5188
rect 20166 5128 20222 5137
rect 20088 5086 20166 5114
rect 19982 5063 19984 5072
rect 20036 5063 20038 5072
rect 20166 5063 20222 5072
rect 19984 5034 20036 5040
rect 19798 4992 19854 5001
rect 19798 4927 19854 4936
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19522 4856 19578 4865
rect 19950 4859 20258 4868
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19432 4820 19484 4826
rect 19522 4791 19578 4800
rect 19984 4820 20036 4826
rect 19432 4762 19484 4768
rect 19156 4752 19208 4758
rect 19156 4694 19208 4700
rect 19248 4752 19300 4758
rect 19248 4694 19300 4700
rect 19260 4622 19288 4694
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19248 4480 19300 4486
rect 19248 4422 19300 4428
rect 19062 4312 19118 4321
rect 19062 4247 19118 4256
rect 18972 4208 19024 4214
rect 18972 4150 19024 4156
rect 19076 3942 19104 4247
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 19168 3398 19196 4082
rect 19260 4078 19288 4422
rect 19352 4078 19380 4762
rect 19444 4622 19472 4762
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19430 4312 19486 4321
rect 19430 4247 19432 4256
rect 19484 4247 19486 4256
rect 19432 4218 19484 4224
rect 19430 4176 19486 4185
rect 19430 4111 19486 4120
rect 19248 4072 19300 4078
rect 19248 4014 19300 4020
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19294 3460 19346 3466
rect 19444 3448 19472 4111
rect 19346 3420 19472 3448
rect 19294 3402 19346 3408
rect 19156 3392 19208 3398
rect 19156 3334 19208 3340
rect 19168 2774 19196 3334
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19168 2746 19288 2774
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 16946 776 17002 785
rect 16946 711 17002 720
rect 17512 56 17632 82
rect 2148 14 2360 42
rect 2778 0 2834 56
rect 3514 0 3570 56
rect 4250 0 4306 56
rect 4986 0 5042 56
rect 5722 0 5778 56
rect 6458 0 6514 56
rect 7194 0 7250 56
rect 7930 0 7986 56
rect 8666 0 8722 56
rect 9402 0 9458 56
rect 10138 0 10194 56
rect 10874 0 10930 56
rect 11610 0 11666 56
rect 12346 0 12402 56
rect 13082 0 13138 56
rect 13818 0 13874 56
rect 14554 0 14610 56
rect 15290 0 15346 56
rect 16026 0 16082 56
rect 16762 0 16818 56
rect 17498 54 17632 56
rect 17498 0 17554 54
rect 17604 42 17632 54
rect 17788 42 17816 2246
rect 18156 1630 18184 2382
rect 18236 2304 18288 2310
rect 18236 2246 18288 2252
rect 18972 2304 19024 2310
rect 18972 2246 19024 2252
rect 18144 1624 18196 1630
rect 18144 1566 18196 1572
rect 18248 56 18276 2246
rect 18984 56 19012 2246
rect 19260 1970 19288 2746
rect 19444 2446 19472 2994
rect 19536 2990 19564 4791
rect 19984 4762 20036 4768
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19708 4276 19760 4282
rect 19708 4218 19760 4224
rect 19720 3534 19748 4218
rect 19904 4078 19932 4626
rect 19996 4214 20024 4762
rect 20076 4684 20128 4690
rect 20076 4626 20128 4632
rect 20088 4321 20116 4626
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 20074 4312 20130 4321
rect 20272 4282 20300 4558
rect 20074 4247 20130 4256
rect 20260 4276 20312 4282
rect 20260 4218 20312 4224
rect 19984 4208 20036 4214
rect 19984 4150 20036 4156
rect 19892 4072 19944 4078
rect 19892 4014 19944 4020
rect 19950 3836 20258 3845
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 19708 3528 19760 3534
rect 19708 3470 19760 3476
rect 20272 3194 20300 3674
rect 20364 3194 20392 6122
rect 20456 5302 20484 6598
rect 20626 6559 20682 6568
rect 20640 6225 20668 6559
rect 20732 6458 20760 6938
rect 20810 6896 20866 6905
rect 20810 6831 20866 6840
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20626 6216 20682 6225
rect 20824 6186 20852 6831
rect 21008 6662 21036 6967
rect 21652 6798 21680 7346
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 20904 6656 20956 6662
rect 20904 6598 20956 6604
rect 20996 6656 21048 6662
rect 20996 6598 21048 6604
rect 21456 6656 21508 6662
rect 21456 6598 21508 6604
rect 20916 6322 20944 6598
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 20904 6316 20956 6322
rect 20904 6258 20956 6264
rect 20626 6151 20682 6160
rect 20812 6180 20864 6186
rect 20812 6122 20864 6128
rect 21088 6112 21140 6118
rect 20640 6060 21088 6066
rect 20640 6054 21140 6060
rect 20640 6038 21128 6054
rect 20640 5846 20668 6038
rect 20902 5944 20958 5953
rect 20902 5879 20958 5888
rect 20628 5840 20680 5846
rect 20628 5782 20680 5788
rect 20812 5704 20864 5710
rect 20812 5646 20864 5652
rect 20824 5545 20852 5646
rect 20810 5536 20866 5545
rect 20810 5471 20866 5480
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20444 5296 20496 5302
rect 20444 5238 20496 5244
rect 20442 4856 20498 4865
rect 20442 4791 20498 4800
rect 20456 4457 20484 4791
rect 20640 4486 20668 5306
rect 20916 5030 20944 5879
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 21468 4826 21496 6598
rect 21548 5704 21600 5710
rect 21548 5646 21600 5652
rect 21560 5234 21588 5646
rect 21548 5228 21600 5234
rect 21548 5170 21600 5176
rect 21456 4820 21508 4826
rect 21456 4762 21508 4768
rect 21560 4622 21588 5170
rect 21548 4616 21600 4622
rect 21548 4558 21600 4564
rect 20628 4480 20680 4486
rect 20442 4448 20498 4457
rect 20628 4422 20680 4428
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 21456 4480 21508 4486
rect 21456 4422 21508 4428
rect 20442 4383 20498 4392
rect 20626 4312 20682 4321
rect 20626 4247 20682 4256
rect 20640 4010 20668 4247
rect 20628 4004 20680 4010
rect 20628 3946 20680 3952
rect 20442 3904 20498 3913
rect 20442 3839 20498 3848
rect 20456 3233 20484 3839
rect 20534 3768 20590 3777
rect 20534 3703 20590 3712
rect 20548 3505 20576 3703
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 20534 3496 20590 3505
rect 20640 3466 20668 3606
rect 20534 3431 20590 3440
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 20442 3224 20498 3233
rect 20260 3188 20312 3194
rect 20260 3130 20312 3136
rect 20352 3188 20404 3194
rect 20442 3159 20498 3168
rect 20352 3130 20404 3136
rect 19524 2984 19576 2990
rect 19524 2926 19576 2932
rect 19616 2848 19668 2854
rect 19616 2790 19668 2796
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 19248 1964 19300 1970
rect 19248 1906 19300 1912
rect 19352 1494 19380 2246
rect 19340 1488 19392 1494
rect 19340 1430 19392 1436
rect 19444 921 19472 2382
rect 19522 2000 19578 2009
rect 19628 1970 19656 2790
rect 19950 2748 20258 2757
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 20720 2440 20772 2446
rect 20824 2428 20852 4422
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 21468 2446 21496 4422
rect 20772 2400 20852 2428
rect 20904 2440 20956 2446
rect 20720 2382 20772 2388
rect 20904 2382 20956 2388
rect 21456 2440 21508 2446
rect 21456 2382 21508 2388
rect 20444 2304 20496 2310
rect 20444 2246 20496 2252
rect 20720 2304 20772 2310
rect 20720 2246 20772 2252
rect 19522 1935 19578 1944
rect 19616 1964 19668 1970
rect 19536 1737 19564 1935
rect 19616 1906 19668 1912
rect 19522 1728 19578 1737
rect 19522 1663 19578 1672
rect 19706 1728 19762 1737
rect 19706 1663 19762 1672
rect 19430 912 19486 921
rect 19430 847 19486 856
rect 19720 56 19748 1663
rect 20456 56 20484 2246
rect 20732 1737 20760 2246
rect 20916 2106 20944 2382
rect 21364 2304 21416 2310
rect 21364 2246 21416 2252
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 20904 2100 20956 2106
rect 20904 2042 20956 2048
rect 20718 1728 20774 1737
rect 20718 1663 20774 1672
rect 21192 56 21312 82
rect 17604 14 17816 42
rect 18234 0 18290 56
rect 18970 0 19026 56
rect 19706 0 19762 56
rect 20442 0 20498 56
rect 21178 54 21312 56
rect 21178 0 21234 54
rect 21284 42 21312 54
rect 21376 42 21404 2246
rect 21560 1222 21588 4558
rect 21652 1834 21680 6734
rect 21824 6724 21876 6730
rect 21824 6666 21876 6672
rect 21730 6624 21786 6633
rect 21730 6559 21786 6568
rect 21744 5642 21772 6559
rect 21732 5636 21784 5642
rect 21732 5578 21784 5584
rect 21732 5024 21784 5030
rect 21732 4966 21784 4972
rect 21640 1828 21692 1834
rect 21640 1770 21692 1776
rect 21744 1562 21772 4966
rect 21836 4282 21864 6666
rect 21824 4276 21876 4282
rect 21824 4218 21876 4224
rect 21928 3505 21956 8298
rect 22008 8288 22060 8294
rect 22008 8230 22060 8236
rect 22020 7886 22048 8230
rect 22204 8022 22232 9250
rect 22296 8548 22324 11194
rect 22572 8634 22600 11194
rect 22848 9625 22876 11194
rect 23124 10033 23152 11194
rect 23400 10305 23428 11194
rect 23386 10296 23442 10305
rect 23386 10231 23442 10240
rect 23110 10024 23166 10033
rect 23110 9959 23166 9968
rect 22834 9616 22890 9625
rect 22834 9551 22890 9560
rect 22652 9104 22704 9110
rect 22652 9046 22704 9052
rect 22664 8673 22692 9046
rect 23204 9036 23256 9042
rect 23204 8978 23256 8984
rect 22650 8664 22706 8673
rect 22560 8628 22612 8634
rect 22650 8599 22706 8608
rect 22560 8570 22612 8576
rect 22468 8560 22520 8566
rect 22296 8520 22468 8548
rect 22468 8502 22520 8508
rect 23112 8492 23164 8498
rect 23112 8434 23164 8440
rect 22376 8356 22428 8362
rect 22296 8316 22376 8344
rect 22192 8016 22244 8022
rect 22192 7958 22244 7964
rect 22008 7880 22060 7886
rect 22008 7822 22060 7828
rect 22100 7812 22152 7818
rect 22100 7754 22152 7760
rect 22008 7744 22060 7750
rect 22008 7686 22060 7692
rect 21914 3496 21970 3505
rect 21914 3431 21970 3440
rect 21822 3224 21878 3233
rect 21822 3159 21878 3168
rect 21836 3126 21864 3159
rect 21824 3120 21876 3126
rect 21824 3062 21876 3068
rect 21824 2848 21876 2854
rect 21824 2790 21876 2796
rect 21836 2650 21864 2790
rect 21824 2644 21876 2650
rect 21824 2586 21876 2592
rect 21824 2440 21876 2446
rect 22020 2428 22048 7686
rect 22112 7206 22140 7754
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 22204 7478 22232 7686
rect 22192 7472 22244 7478
rect 22192 7414 22244 7420
rect 22192 7336 22244 7342
rect 22192 7278 22244 7284
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 22204 4672 22232 7278
rect 22296 6118 22324 8316
rect 22376 8298 22428 8304
rect 22652 8356 22704 8362
rect 22652 8298 22704 8304
rect 22836 8356 22888 8362
rect 22836 8298 22888 8304
rect 22560 7948 22612 7954
rect 22560 7890 22612 7896
rect 22376 7812 22428 7818
rect 22376 7754 22428 7760
rect 22388 7478 22416 7754
rect 22376 7472 22428 7478
rect 22376 7414 22428 7420
rect 22572 6440 22600 7890
rect 22480 6412 22600 6440
rect 22284 6112 22336 6118
rect 22284 6054 22336 6060
rect 22376 5160 22428 5166
rect 22376 5102 22428 5108
rect 22284 4684 22336 4690
rect 22204 4644 22284 4672
rect 22284 4626 22336 4632
rect 22192 3936 22244 3942
rect 22296 3924 22324 4626
rect 22244 3896 22324 3924
rect 22192 3878 22244 3884
rect 22192 3664 22244 3670
rect 22192 3606 22244 3612
rect 22204 3466 22232 3606
rect 22192 3460 22244 3466
rect 22192 3402 22244 3408
rect 22296 2650 22324 3896
rect 22388 3466 22416 5102
rect 22480 4690 22508 6412
rect 22560 6316 22612 6322
rect 22560 6258 22612 6264
rect 22572 5234 22600 6258
rect 22664 5846 22692 8298
rect 22848 7750 22876 8298
rect 23124 8090 23152 8434
rect 23112 8084 23164 8090
rect 23112 8026 23164 8032
rect 22928 7948 22980 7954
rect 22928 7890 22980 7896
rect 23112 7948 23164 7954
rect 23216 7936 23244 8978
rect 23676 8430 23704 11194
rect 23952 9602 23980 11194
rect 23952 9574 24072 9602
rect 23296 8424 23348 8430
rect 23572 8424 23624 8430
rect 23296 8366 23348 8372
rect 23492 8384 23572 8412
rect 23308 8129 23336 8366
rect 23294 8120 23350 8129
rect 23294 8055 23350 8064
rect 23164 7908 23244 7936
rect 23112 7890 23164 7896
rect 22836 7744 22888 7750
rect 22836 7686 22888 7692
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22652 5840 22704 5846
rect 22652 5782 22704 5788
rect 22560 5228 22612 5234
rect 22560 5170 22612 5176
rect 22468 4684 22520 4690
rect 22468 4626 22520 4632
rect 22572 4146 22600 5170
rect 22560 4140 22612 4146
rect 22560 4082 22612 4088
rect 22572 4049 22600 4082
rect 22558 4040 22614 4049
rect 22558 3975 22614 3984
rect 22560 3528 22612 3534
rect 22756 3505 22784 7482
rect 22848 4758 22876 7686
rect 22836 4752 22888 4758
rect 22836 4694 22888 4700
rect 22836 4072 22888 4078
rect 22836 4014 22888 4020
rect 22848 3738 22876 4014
rect 22836 3732 22888 3738
rect 22836 3674 22888 3680
rect 22836 3596 22888 3602
rect 22836 3538 22888 3544
rect 22560 3470 22612 3476
rect 22742 3496 22798 3505
rect 22376 3460 22428 3466
rect 22376 3402 22428 3408
rect 22572 3058 22600 3470
rect 22742 3431 22798 3440
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 22744 3392 22796 3398
rect 22744 3334 22796 3340
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 22284 2644 22336 2650
rect 22284 2586 22336 2592
rect 22376 2440 22428 2446
rect 22020 2400 22376 2428
rect 21824 2382 21876 2388
rect 22376 2382 22428 2388
rect 21732 1556 21784 1562
rect 21732 1498 21784 1504
rect 21548 1216 21600 1222
rect 21548 1158 21600 1164
rect 21836 1057 21864 2382
rect 22572 2378 22600 2994
rect 22664 2774 22692 3334
rect 22756 3233 22784 3334
rect 22742 3224 22798 3233
rect 22742 3159 22798 3168
rect 22848 3058 22876 3538
rect 22836 3052 22888 3058
rect 22836 2994 22888 3000
rect 22664 2746 22784 2774
rect 22652 2644 22704 2650
rect 22652 2586 22704 2592
rect 22560 2372 22612 2378
rect 22560 2314 22612 2320
rect 21916 1828 21968 1834
rect 21916 1770 21968 1776
rect 21822 1048 21878 1057
rect 21822 983 21878 992
rect 21928 56 21956 1770
rect 22664 56 22692 2586
rect 22756 2514 22784 2746
rect 22940 2582 22968 7890
rect 23308 7410 23336 8055
rect 23296 7404 23348 7410
rect 23296 7346 23348 7352
rect 23492 6458 23520 8384
rect 23572 8366 23624 8372
rect 23664 8424 23716 8430
rect 23664 8366 23716 8372
rect 23848 8288 23900 8294
rect 23848 8230 23900 8236
rect 23572 7880 23624 7886
rect 23572 7822 23624 7828
rect 23584 7546 23612 7822
rect 23572 7540 23624 7546
rect 23572 7482 23624 7488
rect 23572 7336 23624 7342
rect 23572 7278 23624 7284
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23388 6248 23440 6254
rect 23388 6190 23440 6196
rect 23400 6100 23428 6190
rect 23400 6072 23520 6100
rect 23492 5778 23520 6072
rect 23584 5914 23612 7278
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 23572 5908 23624 5914
rect 23572 5850 23624 5856
rect 23676 5846 23704 6190
rect 23664 5840 23716 5846
rect 23664 5782 23716 5788
rect 23480 5772 23532 5778
rect 23480 5714 23532 5720
rect 23112 5636 23164 5642
rect 23112 5578 23164 5584
rect 23020 4684 23072 4690
rect 23020 4626 23072 4632
rect 23032 4282 23060 4626
rect 23020 4276 23072 4282
rect 23020 4218 23072 4224
rect 23020 3664 23072 3670
rect 23020 3606 23072 3612
rect 23032 3398 23060 3606
rect 23020 3392 23072 3398
rect 23020 3334 23072 3340
rect 23124 3194 23152 5578
rect 23572 5024 23624 5030
rect 23572 4966 23624 4972
rect 23584 4622 23612 4966
rect 23676 4865 23704 5782
rect 23768 5778 23796 6734
rect 23860 6390 23888 8230
rect 24044 8022 24072 9574
rect 24122 9072 24178 9081
rect 24122 9007 24178 9016
rect 24032 8016 24084 8022
rect 24032 7958 24084 7964
rect 23940 6452 23992 6458
rect 23940 6394 23992 6400
rect 23848 6384 23900 6390
rect 23848 6326 23900 6332
rect 23756 5772 23808 5778
rect 23756 5714 23808 5720
rect 23952 5642 23980 6394
rect 24032 6384 24084 6390
rect 24032 6326 24084 6332
rect 24044 5710 24072 6326
rect 24032 5704 24084 5710
rect 24032 5646 24084 5652
rect 23940 5636 23992 5642
rect 23940 5578 23992 5584
rect 24136 5030 24164 9007
rect 24228 7750 24256 11194
rect 24398 10432 24454 10441
rect 24398 10367 24454 10376
rect 24306 9208 24362 9217
rect 24306 9143 24362 9152
rect 24320 7750 24348 9143
rect 24412 8634 24440 10367
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 24504 8566 24532 11194
rect 24584 9988 24636 9994
rect 24584 9930 24636 9936
rect 24492 8560 24544 8566
rect 24492 8502 24544 8508
rect 24490 8256 24546 8265
rect 24490 8191 24546 8200
rect 24400 7880 24452 7886
rect 24400 7822 24452 7828
rect 24216 7744 24268 7750
rect 24216 7686 24268 7692
rect 24308 7744 24360 7750
rect 24308 7686 24360 7692
rect 24124 5024 24176 5030
rect 24124 4966 24176 4972
rect 23662 4856 23718 4865
rect 23662 4791 23718 4800
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 23676 4298 23704 4791
rect 23584 4270 23704 4298
rect 23584 3534 23612 4270
rect 23664 4140 23716 4146
rect 23664 4082 23716 4088
rect 23572 3528 23624 3534
rect 23572 3470 23624 3476
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 23676 3058 23704 4082
rect 23664 3052 23716 3058
rect 23664 2994 23716 3000
rect 22928 2576 22980 2582
rect 22928 2518 22980 2524
rect 23296 2576 23348 2582
rect 23296 2518 23348 2524
rect 23388 2576 23440 2582
rect 24412 2530 24440 7822
rect 24504 7342 24532 8191
rect 24596 7970 24624 9930
rect 24780 9897 24808 11194
rect 24950 10568 25006 10577
rect 24950 10503 25006 10512
rect 24766 9888 24822 9897
rect 24766 9823 24822 9832
rect 24674 9616 24730 9625
rect 24674 9551 24730 9560
rect 24688 8498 24716 9551
rect 24964 9500 24992 10503
rect 25056 9625 25084 11194
rect 25228 10260 25280 10266
rect 25228 10202 25280 10208
rect 25134 10024 25190 10033
rect 25134 9959 25190 9968
rect 25042 9616 25098 9625
rect 25042 9551 25098 9560
rect 24964 9472 25084 9500
rect 24860 9308 24912 9314
rect 24860 9250 24912 9256
rect 24872 8634 24900 9250
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 24676 8492 24728 8498
rect 24676 8434 24728 8440
rect 24768 8288 24820 8294
rect 24768 8230 24820 8236
rect 24596 7942 24716 7970
rect 24584 7880 24636 7886
rect 24584 7822 24636 7828
rect 24596 7546 24624 7822
rect 24688 7546 24716 7942
rect 24584 7540 24636 7546
rect 24584 7482 24636 7488
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 24492 7336 24544 7342
rect 24492 7278 24544 7284
rect 24504 6322 24532 7278
rect 24674 6896 24730 6905
rect 24674 6831 24730 6840
rect 24492 6316 24544 6322
rect 24492 6258 24544 6264
rect 24584 6248 24636 6254
rect 24584 6190 24636 6196
rect 24492 5772 24544 5778
rect 24492 5714 24544 5720
rect 24504 4622 24532 5714
rect 24596 5370 24624 6190
rect 24688 5817 24716 6831
rect 24674 5808 24730 5817
rect 24674 5743 24730 5752
rect 24584 5364 24636 5370
rect 24584 5306 24636 5312
rect 24780 5001 24808 8230
rect 24860 7948 24912 7954
rect 24860 7890 24912 7896
rect 24872 5953 24900 7890
rect 25056 7426 25084 9472
rect 25148 8498 25176 9959
rect 25240 9058 25268 10202
rect 25332 9217 25360 11194
rect 25410 10296 25466 10305
rect 25608 10266 25636 11194
rect 25410 10231 25466 10240
rect 25596 10260 25648 10266
rect 25318 9208 25374 9217
rect 25318 9143 25374 9152
rect 25240 9030 25360 9058
rect 25136 8492 25188 8498
rect 25136 8434 25188 8440
rect 25228 8288 25280 8294
rect 25228 8230 25280 8236
rect 24964 7398 25084 7426
rect 25136 7404 25188 7410
rect 24858 5944 24914 5953
rect 24858 5879 24914 5888
rect 24858 5808 24914 5817
rect 24858 5743 24914 5752
rect 24872 5098 24900 5743
rect 24964 5234 24992 7398
rect 25136 7346 25188 7352
rect 25148 7313 25176 7346
rect 25134 7304 25190 7313
rect 25056 7262 25134 7290
rect 25056 6322 25084 7262
rect 25134 7239 25190 7248
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 25044 6316 25096 6322
rect 25044 6258 25096 6264
rect 25148 6089 25176 6734
rect 25240 6662 25268 8230
rect 25228 6656 25280 6662
rect 25228 6598 25280 6604
rect 25134 6080 25190 6089
rect 25134 6015 25190 6024
rect 25228 5704 25280 5710
rect 25332 5692 25360 9030
rect 25424 8498 25452 10231
rect 25596 10202 25648 10208
rect 25884 9790 25912 11194
rect 25872 9784 25924 9790
rect 25872 9726 25924 9732
rect 25780 9172 25832 9178
rect 25780 9114 25832 9120
rect 25872 9172 25924 9178
rect 25872 9114 25924 9120
rect 25792 8634 25820 9114
rect 25780 8628 25832 8634
rect 25780 8570 25832 8576
rect 25412 8492 25464 8498
rect 25412 8434 25464 8440
rect 25780 8424 25832 8430
rect 25780 8366 25832 8372
rect 25504 8288 25556 8294
rect 25504 8230 25556 8236
rect 25412 7744 25464 7750
rect 25412 7686 25464 7692
rect 25424 6934 25452 7686
rect 25412 6928 25464 6934
rect 25412 6870 25464 6876
rect 25412 6792 25464 6798
rect 25412 6734 25464 6740
rect 25424 6497 25452 6734
rect 25410 6488 25466 6497
rect 25410 6423 25466 6432
rect 25280 5664 25360 5692
rect 25228 5646 25280 5652
rect 24952 5228 25004 5234
rect 24952 5170 25004 5176
rect 24860 5092 24912 5098
rect 24860 5034 24912 5040
rect 24766 4992 24822 5001
rect 24766 4927 24822 4936
rect 25332 4622 25360 5664
rect 24492 4616 24544 4622
rect 24492 4558 24544 4564
rect 25320 4616 25372 4622
rect 25320 4558 25372 4564
rect 24504 2990 24532 4558
rect 25332 4486 25360 4558
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 25320 4480 25372 4486
rect 25320 4422 25372 4428
rect 24780 4162 24808 4422
rect 25412 4276 25464 4282
rect 25412 4218 25464 4224
rect 25044 4208 25096 4214
rect 24964 4168 25044 4196
rect 24964 4162 24992 4168
rect 24780 4134 24992 4162
rect 25044 4150 25096 4156
rect 24858 4040 24914 4049
rect 24858 3975 24914 3984
rect 24676 3936 24728 3942
rect 24676 3878 24728 3884
rect 24492 2984 24544 2990
rect 24492 2926 24544 2932
rect 23388 2518 23440 2524
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 23308 1834 23336 2518
rect 23296 1828 23348 1834
rect 23296 1770 23348 1776
rect 23400 56 23428 2518
rect 24320 2502 24440 2530
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 23492 678 23520 2382
rect 24124 2304 24176 2310
rect 24124 2246 24176 2252
rect 23480 672 23532 678
rect 23480 614 23532 620
rect 24136 56 24164 2246
rect 24320 1902 24348 2502
rect 24400 2440 24452 2446
rect 24400 2382 24452 2388
rect 24308 1896 24360 1902
rect 24308 1838 24360 1844
rect 24412 1766 24440 2382
rect 24688 2009 24716 3878
rect 24674 2000 24730 2009
rect 24674 1935 24730 1944
rect 24400 1760 24452 1766
rect 24400 1702 24452 1708
rect 24872 56 24900 3975
rect 25044 3052 25096 3058
rect 25044 2994 25096 3000
rect 25056 1018 25084 2994
rect 25424 2038 25452 4218
rect 25516 4185 25544 8230
rect 25596 7880 25648 7886
rect 25596 7822 25648 7828
rect 25608 7410 25636 7822
rect 25596 7404 25648 7410
rect 25596 7346 25648 7352
rect 25792 7290 25820 8366
rect 25700 7262 25820 7290
rect 25596 5228 25648 5234
rect 25596 5170 25648 5176
rect 25608 4826 25636 5170
rect 25596 4820 25648 4826
rect 25596 4762 25648 4768
rect 25502 4176 25558 4185
rect 25502 4111 25558 4120
rect 25596 4072 25648 4078
rect 25596 4014 25648 4020
rect 25608 3194 25636 4014
rect 25700 3913 25728 7262
rect 25884 6882 25912 9114
rect 26160 8566 26188 11194
rect 26238 9888 26294 9897
rect 26238 9823 26294 9832
rect 26148 8560 26200 8566
rect 26148 8502 26200 8508
rect 26252 8498 26280 9823
rect 26330 9616 26386 9625
rect 26330 9551 26386 9560
rect 26344 8498 26372 9551
rect 26240 8492 26292 8498
rect 26240 8434 26292 8440
rect 26332 8492 26384 8498
rect 26332 8434 26384 8440
rect 26436 8362 26464 11194
rect 26516 10260 26568 10266
rect 26516 10202 26568 10208
rect 26528 8634 26556 10202
rect 26712 9625 26740 11194
rect 26698 9616 26754 9625
rect 26698 9551 26754 9560
rect 26700 9376 26752 9382
rect 26700 9318 26752 9324
rect 26608 8832 26660 8838
rect 26608 8774 26660 8780
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 26424 8356 26476 8362
rect 26424 8298 26476 8304
rect 26620 8294 26648 8774
rect 26712 8294 26740 9318
rect 26790 9208 26846 9217
rect 26790 9143 26846 9152
rect 26804 8498 26832 9143
rect 26988 8838 27016 11194
rect 27264 10690 27292 11194
rect 27264 10662 27384 10690
rect 26976 8832 27028 8838
rect 26976 8774 27028 8780
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 26882 8664 26938 8673
rect 27010 8667 27318 8676
rect 26882 8599 26938 8608
rect 27160 8628 27212 8634
rect 26792 8492 26844 8498
rect 26792 8434 26844 8440
rect 26516 8288 26568 8294
rect 26516 8230 26568 8236
rect 26608 8288 26660 8294
rect 26608 8230 26660 8236
rect 26700 8288 26752 8294
rect 26700 8230 26752 8236
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 26332 7744 26384 7750
rect 26330 7712 26332 7721
rect 26384 7712 26386 7721
rect 26330 7647 26386 7656
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 25884 6854 26004 6882
rect 25976 6610 26004 6854
rect 25792 6582 26004 6610
rect 25686 3904 25742 3913
rect 25686 3839 25742 3848
rect 25792 3777 25820 6582
rect 25962 6488 26018 6497
rect 26528 6458 26556 8230
rect 26896 7936 26924 8599
rect 27160 8570 27212 8576
rect 27172 8498 27200 8570
rect 27356 8566 27384 10662
rect 27436 9784 27488 9790
rect 27436 9726 27488 9732
rect 27344 8560 27396 8566
rect 27344 8502 27396 8508
rect 27448 8498 27476 9726
rect 27540 8634 27568 11194
rect 27618 9616 27674 9625
rect 27618 9551 27674 9560
rect 27528 8628 27580 8634
rect 27528 8570 27580 8576
rect 27068 8492 27120 8498
rect 27068 8434 27120 8440
rect 27160 8492 27212 8498
rect 27160 8434 27212 8440
rect 27436 8492 27488 8498
rect 27436 8434 27488 8440
rect 27080 8294 27108 8434
rect 27068 8288 27120 8294
rect 27068 8230 27120 8236
rect 27356 8078 27568 8106
rect 26896 7908 27108 7936
rect 26792 7880 26844 7886
rect 27080 7868 27108 7908
rect 27356 7886 27384 8078
rect 27436 8016 27488 8022
rect 27436 7958 27488 7964
rect 27160 7880 27212 7886
rect 27080 7840 27160 7868
rect 26792 7822 26844 7828
rect 27160 7822 27212 7828
rect 27344 7880 27396 7886
rect 27344 7822 27396 7828
rect 26608 7812 26660 7818
rect 26608 7754 26660 7760
rect 26620 6633 26648 7754
rect 26804 7546 26832 7822
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 26792 7540 26844 7546
rect 26792 7482 26844 7488
rect 26804 7410 26832 7482
rect 26792 7404 26844 7410
rect 26792 7346 26844 7352
rect 26606 6624 26662 6633
rect 26606 6559 26662 6568
rect 25962 6423 26018 6432
rect 26424 6452 26476 6458
rect 25872 6248 25924 6254
rect 25872 6190 25924 6196
rect 25884 4690 25912 6190
rect 25976 6118 26004 6423
rect 26424 6394 26476 6400
rect 26516 6452 26568 6458
rect 26516 6394 26568 6400
rect 26436 6338 26464 6394
rect 26436 6310 26648 6338
rect 26804 6322 26832 7346
rect 27160 7200 27212 7206
rect 27160 7142 27212 7148
rect 27172 6866 27200 7142
rect 27160 6860 27212 6866
rect 27160 6802 27212 6808
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 27356 6440 27384 7822
rect 27448 7002 27476 7958
rect 27540 7528 27568 8078
rect 27632 7886 27660 9551
rect 27816 8430 27844 11194
rect 28092 9654 28120 11194
rect 28080 9648 28132 9654
rect 28080 9590 28132 9596
rect 28080 9172 28132 9178
rect 28080 9114 28132 9120
rect 27804 8424 27856 8430
rect 27804 8366 27856 8372
rect 28092 8362 28120 9114
rect 28264 8832 28316 8838
rect 28264 8774 28316 8780
rect 28276 8498 28304 8774
rect 28264 8492 28316 8498
rect 28264 8434 28316 8440
rect 27712 8356 27764 8362
rect 27712 8298 27764 8304
rect 28080 8356 28132 8362
rect 28080 8298 28132 8304
rect 27724 8129 27752 8298
rect 27896 8288 27948 8294
rect 27896 8230 27948 8236
rect 27710 8120 27766 8129
rect 27710 8055 27766 8064
rect 27620 7880 27672 7886
rect 27620 7822 27672 7828
rect 27804 7812 27856 7818
rect 27804 7754 27856 7760
rect 27540 7500 27660 7528
rect 27526 7440 27582 7449
rect 27632 7410 27660 7500
rect 27526 7375 27582 7384
rect 27620 7404 27672 7410
rect 27436 6996 27488 7002
rect 27436 6938 27488 6944
rect 27540 6662 27568 7375
rect 27620 7346 27672 7352
rect 27528 6656 27580 6662
rect 27528 6598 27580 6604
rect 27528 6452 27580 6458
rect 27356 6412 27476 6440
rect 27066 6352 27122 6361
rect 26620 6118 26648 6310
rect 26792 6316 26844 6322
rect 27066 6287 27122 6296
rect 27342 6352 27398 6361
rect 27342 6287 27398 6296
rect 26792 6258 26844 6264
rect 26698 6216 26754 6225
rect 26698 6151 26754 6160
rect 25964 6112 26016 6118
rect 25964 6054 26016 6060
rect 26332 6112 26384 6118
rect 26332 6054 26384 6060
rect 26608 6112 26660 6118
rect 26608 6054 26660 6060
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 26344 5710 26372 6054
rect 26712 5710 26740 6151
rect 26792 5908 26844 5914
rect 26792 5850 26844 5856
rect 26332 5704 26384 5710
rect 26332 5646 26384 5652
rect 26700 5704 26752 5710
rect 26700 5646 26752 5652
rect 26056 5160 26108 5166
rect 26054 5128 26056 5137
rect 26108 5128 26110 5137
rect 26344 5098 26372 5646
rect 26424 5296 26476 5302
rect 26424 5238 26476 5244
rect 26054 5063 26110 5072
rect 26332 5092 26384 5098
rect 26332 5034 26384 5040
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 25872 4684 25924 4690
rect 25872 4626 25924 4632
rect 25884 4282 25912 4626
rect 26056 4480 26108 4486
rect 26056 4422 26108 4428
rect 26240 4480 26292 4486
rect 26240 4422 26292 4428
rect 26068 4282 26096 4422
rect 25872 4276 25924 4282
rect 25872 4218 25924 4224
rect 26056 4276 26108 4282
rect 26056 4218 26108 4224
rect 26252 4146 26280 4422
rect 26240 4140 26292 4146
rect 26240 4082 26292 4088
rect 26344 4010 26372 5034
rect 26436 4622 26464 5238
rect 26804 4690 26832 5850
rect 27080 5681 27108 6287
rect 27066 5672 27122 5681
rect 27066 5607 27122 5616
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 27160 5228 27212 5234
rect 27080 5188 27160 5216
rect 27080 4729 27108 5188
rect 27160 5170 27212 5176
rect 27066 4720 27122 4729
rect 26792 4684 26844 4690
rect 27066 4655 27122 4664
rect 26792 4626 26844 4632
rect 27080 4622 27108 4655
rect 26424 4616 26476 4622
rect 26424 4558 26476 4564
rect 27068 4616 27120 4622
rect 27068 4558 27120 4564
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 26332 4004 26384 4010
rect 26332 3946 26384 3952
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25778 3768 25834 3777
rect 25950 3771 26258 3780
rect 26344 3738 26372 3946
rect 26608 3936 26660 3942
rect 26608 3878 26660 3884
rect 25778 3703 25834 3712
rect 26332 3732 26384 3738
rect 26332 3674 26384 3680
rect 26148 3528 26200 3534
rect 26332 3528 26384 3534
rect 26200 3488 26280 3516
rect 26148 3470 26200 3476
rect 25872 3460 25924 3466
rect 25872 3402 25924 3408
rect 25596 3188 25648 3194
rect 25596 3130 25648 3136
rect 25884 3058 25912 3402
rect 25872 3052 25924 3058
rect 25872 2994 25924 3000
rect 26252 2990 26280 3488
rect 26332 3470 26384 3476
rect 26344 3194 26372 3470
rect 26332 3188 26384 3194
rect 26332 3130 26384 3136
rect 26240 2984 26292 2990
rect 26240 2926 26292 2932
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 26332 2372 26384 2378
rect 26332 2314 26384 2320
rect 25412 2032 25464 2038
rect 25412 1974 25464 1980
rect 25596 1828 25648 1834
rect 25596 1770 25648 1776
rect 25044 1012 25096 1018
rect 25044 954 25096 960
rect 25608 56 25636 1770
rect 26344 56 26372 2314
rect 26620 882 26648 3878
rect 27356 3398 27384 6287
rect 27448 5778 27476 6412
rect 27528 6394 27580 6400
rect 27540 6322 27568 6394
rect 27528 6316 27580 6322
rect 27528 6258 27580 6264
rect 27436 5772 27488 5778
rect 27436 5714 27488 5720
rect 27448 4622 27476 5714
rect 27540 5574 27568 6258
rect 27712 5704 27764 5710
rect 27632 5652 27712 5658
rect 27632 5646 27764 5652
rect 27632 5630 27752 5646
rect 27528 5568 27580 5574
rect 27528 5510 27580 5516
rect 27632 5386 27660 5630
rect 27540 5358 27660 5386
rect 27712 5364 27764 5370
rect 27540 4690 27568 5358
rect 27712 5306 27764 5312
rect 27724 5234 27752 5306
rect 27712 5228 27764 5234
rect 27712 5170 27764 5176
rect 27528 4684 27580 4690
rect 27528 4626 27580 4632
rect 27436 4616 27488 4622
rect 27436 4558 27488 4564
rect 27448 4486 27476 4558
rect 27712 4548 27764 4554
rect 27712 4490 27764 4496
rect 27436 4480 27488 4486
rect 27436 4422 27488 4428
rect 27528 4480 27580 4486
rect 27528 4422 27580 4428
rect 27436 4140 27488 4146
rect 27436 4082 27488 4088
rect 27448 3641 27476 4082
rect 27434 3632 27490 3641
rect 27434 3567 27490 3576
rect 27448 3534 27476 3567
rect 27436 3528 27488 3534
rect 27540 3516 27568 4422
rect 27620 3528 27672 3534
rect 27540 3488 27620 3516
rect 27436 3470 27488 3476
rect 27620 3470 27672 3476
rect 27344 3392 27396 3398
rect 27344 3334 27396 3340
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 27448 3058 27476 3470
rect 27724 3194 27752 4490
rect 27712 3188 27764 3194
rect 27712 3130 27764 3136
rect 27436 3052 27488 3058
rect 27436 2994 27488 3000
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 27816 1834 27844 7754
rect 27908 4214 27936 8230
rect 28368 7410 28396 11194
rect 28448 9512 28500 9518
rect 28448 9454 28500 9460
rect 28356 7404 28408 7410
rect 28356 7346 28408 7352
rect 28460 6458 28488 9454
rect 28644 8838 28672 11194
rect 28920 9874 28948 11194
rect 29000 10192 29052 10198
rect 29000 10134 29052 10140
rect 28828 9846 28948 9874
rect 28828 9625 28856 9846
rect 28908 9648 28960 9654
rect 28814 9616 28870 9625
rect 28724 9580 28776 9586
rect 28908 9590 28960 9596
rect 28814 9551 28870 9560
rect 28724 9522 28776 9528
rect 28632 8832 28684 8838
rect 28632 8774 28684 8780
rect 28736 8294 28764 9522
rect 28920 8566 28948 9590
rect 29012 8634 29040 10134
rect 29000 8628 29052 8634
rect 29000 8570 29052 8576
rect 28908 8560 28960 8566
rect 28908 8502 28960 8508
rect 29196 8430 29224 11194
rect 29472 8566 29500 11194
rect 29552 9852 29604 9858
rect 29552 9794 29604 9800
rect 29460 8560 29512 8566
rect 29460 8502 29512 8508
rect 29184 8424 29236 8430
rect 29184 8366 29236 8372
rect 28724 8288 28776 8294
rect 28724 8230 28776 8236
rect 28816 8288 28868 8294
rect 28816 8230 28868 8236
rect 28540 7812 28592 7818
rect 28540 7754 28592 7760
rect 28552 7206 28580 7754
rect 28540 7200 28592 7206
rect 28540 7142 28592 7148
rect 28724 6928 28776 6934
rect 28552 6888 28724 6916
rect 28448 6452 28500 6458
rect 28448 6394 28500 6400
rect 28552 5953 28580 6888
rect 28724 6870 28776 6876
rect 28724 6724 28776 6730
rect 28828 6712 28856 8230
rect 29092 7880 29144 7886
rect 29092 7822 29144 7828
rect 29368 7880 29420 7886
rect 29368 7822 29420 7828
rect 29460 7880 29512 7886
rect 29460 7822 29512 7828
rect 29000 7744 29052 7750
rect 29000 7686 29052 7692
rect 29012 7410 29040 7686
rect 29000 7404 29052 7410
rect 29000 7346 29052 7352
rect 29104 7392 29132 7822
rect 29184 7404 29236 7410
rect 29104 7364 29184 7392
rect 28908 7200 28960 7206
rect 28908 7142 28960 7148
rect 28776 6684 28856 6712
rect 28724 6666 28776 6672
rect 28632 6316 28684 6322
rect 28632 6258 28684 6264
rect 28538 5944 28594 5953
rect 28644 5914 28672 6258
rect 28724 6112 28776 6118
rect 28724 6054 28776 6060
rect 28736 5914 28764 6054
rect 28538 5879 28594 5888
rect 28632 5908 28684 5914
rect 28632 5850 28684 5856
rect 28724 5908 28776 5914
rect 28724 5850 28776 5856
rect 28264 5228 28316 5234
rect 28264 5170 28316 5176
rect 28080 5160 28132 5166
rect 27986 5128 28042 5137
rect 28080 5102 28132 5108
rect 27986 5063 28042 5072
rect 27896 4208 27948 4214
rect 27896 4150 27948 4156
rect 27804 1828 27856 1834
rect 27804 1770 27856 1776
rect 27068 1420 27120 1426
rect 27068 1362 27120 1368
rect 26608 876 26660 882
rect 26608 818 26660 824
rect 27080 56 27108 1362
rect 27816 56 27936 82
rect 21284 14 21404 42
rect 21914 0 21970 56
rect 22650 0 22706 56
rect 23386 0 23442 56
rect 24122 0 24178 56
rect 24858 0 24914 56
rect 25594 0 25650 56
rect 26330 0 26386 56
rect 27066 0 27122 56
rect 27802 54 27936 56
rect 27802 0 27858 54
rect 27908 42 27936 54
rect 28000 42 28028 5063
rect 28092 4622 28120 5102
rect 28080 4616 28132 4622
rect 28080 4558 28132 4564
rect 28172 4616 28224 4622
rect 28172 4558 28224 4564
rect 28092 4010 28120 4558
rect 28184 4146 28212 4558
rect 28172 4140 28224 4146
rect 28172 4082 28224 4088
rect 28080 4004 28132 4010
rect 28080 3946 28132 3952
rect 28276 3670 28304 5170
rect 28920 3942 28948 7142
rect 29104 7041 29132 7364
rect 29184 7346 29236 7352
rect 29380 7342 29408 7822
rect 29368 7336 29420 7342
rect 29368 7278 29420 7284
rect 29184 7268 29236 7274
rect 29184 7210 29236 7216
rect 29196 7154 29224 7210
rect 29368 7200 29420 7206
rect 29196 7148 29368 7154
rect 29196 7142 29420 7148
rect 29196 7126 29408 7142
rect 29090 7032 29146 7041
rect 29090 6967 29146 6976
rect 29090 6488 29146 6497
rect 29090 6423 29146 6432
rect 29104 6390 29132 6423
rect 29092 6384 29144 6390
rect 29092 6326 29144 6332
rect 29092 6112 29144 6118
rect 29092 6054 29144 6060
rect 29000 5772 29052 5778
rect 29000 5714 29052 5720
rect 29012 5273 29040 5714
rect 28998 5264 29054 5273
rect 28998 5199 29054 5208
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 29012 4282 29040 4558
rect 29000 4276 29052 4282
rect 29000 4218 29052 4224
rect 28908 3936 28960 3942
rect 28908 3878 28960 3884
rect 28264 3664 28316 3670
rect 28264 3606 28316 3612
rect 29000 3460 29052 3466
rect 29000 3402 29052 3408
rect 28264 3392 28316 3398
rect 28264 3334 28316 3340
rect 28276 3126 28304 3334
rect 28264 3120 28316 3126
rect 28264 3062 28316 3068
rect 29012 1426 29040 3402
rect 29104 1630 29132 6054
rect 29368 5772 29420 5778
rect 29368 5714 29420 5720
rect 29380 5642 29408 5714
rect 29368 5636 29420 5642
rect 29368 5578 29420 5584
rect 29182 5264 29238 5273
rect 29182 5199 29238 5208
rect 29196 4486 29224 5199
rect 29276 5160 29328 5166
rect 29276 5102 29328 5108
rect 29288 4622 29316 5102
rect 29472 5030 29500 7822
rect 29460 5024 29512 5030
rect 29460 4966 29512 4972
rect 29472 4690 29500 4966
rect 29460 4684 29512 4690
rect 29460 4626 29512 4632
rect 29564 4622 29592 9794
rect 29748 8634 29776 11194
rect 29828 10396 29880 10402
rect 29828 10338 29880 10344
rect 29736 8628 29788 8634
rect 29736 8570 29788 8576
rect 29840 8498 29868 10338
rect 30024 9654 30052 11194
rect 30300 9897 30328 11194
rect 30380 10124 30432 10130
rect 30380 10066 30432 10072
rect 30286 9888 30342 9897
rect 30286 9823 30342 9832
rect 30012 9648 30064 9654
rect 30012 9590 30064 9596
rect 30288 9104 30340 9110
rect 30288 9046 30340 9052
rect 29828 8492 29880 8498
rect 29828 8434 29880 8440
rect 29920 8356 29972 8362
rect 29920 8298 29972 8304
rect 29828 7880 29880 7886
rect 29828 7822 29880 7828
rect 29840 7585 29868 7822
rect 29826 7576 29882 7585
rect 29826 7511 29882 7520
rect 29840 7410 29868 7511
rect 29828 7404 29880 7410
rect 29828 7346 29880 7352
rect 29828 6996 29880 7002
rect 29828 6938 29880 6944
rect 29644 6316 29696 6322
rect 29644 6258 29696 6264
rect 29656 4826 29684 6258
rect 29644 4820 29696 4826
rect 29644 4762 29696 4768
rect 29276 4616 29328 4622
rect 29276 4558 29328 4564
rect 29552 4616 29604 4622
rect 29552 4558 29604 4564
rect 29184 4480 29236 4486
rect 29184 4422 29236 4428
rect 29458 3632 29514 3641
rect 29840 3602 29868 6938
rect 29932 6798 29960 8298
rect 30300 7721 30328 9046
rect 30392 8906 30420 10066
rect 30472 9036 30524 9042
rect 30472 8978 30524 8984
rect 30380 8900 30432 8906
rect 30380 8842 30432 8848
rect 30378 8800 30434 8809
rect 30378 8735 30434 8744
rect 30392 8265 30420 8735
rect 30484 8294 30512 8978
rect 30472 8288 30524 8294
rect 30378 8256 30434 8265
rect 30472 8230 30524 8236
rect 30378 8191 30434 8200
rect 30380 8084 30432 8090
rect 30380 8026 30432 8032
rect 30472 8084 30524 8090
rect 30472 8026 30524 8032
rect 30286 7712 30342 7721
rect 30286 7647 30342 7656
rect 30104 7268 30156 7274
rect 30104 7210 30156 7216
rect 30012 7200 30064 7206
rect 30012 7142 30064 7148
rect 30024 7002 30052 7142
rect 30012 6996 30064 7002
rect 30012 6938 30064 6944
rect 30116 6866 30144 7210
rect 30196 7200 30248 7206
rect 30196 7142 30248 7148
rect 30288 7200 30340 7206
rect 30288 7142 30340 7148
rect 30104 6860 30156 6866
rect 30104 6802 30156 6808
rect 30208 6798 30236 7142
rect 30300 6934 30328 7142
rect 30288 6928 30340 6934
rect 30288 6870 30340 6876
rect 30392 6866 30420 8026
rect 30484 7546 30512 8026
rect 30576 7546 30604 11194
rect 30748 10056 30800 10062
rect 30748 9998 30800 10004
rect 30656 8832 30708 8838
rect 30656 8774 30708 8780
rect 30668 8498 30696 8774
rect 30656 8492 30708 8498
rect 30656 8434 30708 8440
rect 30760 8294 30788 9998
rect 30748 8288 30800 8294
rect 30654 8256 30710 8265
rect 30748 8230 30800 8236
rect 30654 8191 30710 8200
rect 30472 7540 30524 7546
rect 30472 7482 30524 7488
rect 30564 7540 30616 7546
rect 30564 7482 30616 7488
rect 30564 7404 30616 7410
rect 30564 7346 30616 7352
rect 30472 7336 30524 7342
rect 30472 7278 30524 7284
rect 30380 6860 30432 6866
rect 30380 6802 30432 6808
rect 29920 6792 29972 6798
rect 29920 6734 29972 6740
rect 30196 6792 30248 6798
rect 30196 6734 30248 6740
rect 30378 6760 30434 6769
rect 29932 6322 29960 6734
rect 30378 6695 30434 6704
rect 30392 6662 30420 6695
rect 30288 6656 30340 6662
rect 30288 6598 30340 6604
rect 30380 6656 30432 6662
rect 30380 6598 30432 6604
rect 30300 6474 30328 6598
rect 30484 6474 30512 7278
rect 30576 6934 30604 7346
rect 30564 6928 30616 6934
rect 30564 6870 30616 6876
rect 30668 6662 30696 8191
rect 30748 7744 30800 7750
rect 30748 7686 30800 7692
rect 30760 7342 30788 7686
rect 30852 7546 30880 11194
rect 30930 9616 30986 9625
rect 30930 9551 30986 9560
rect 30944 8498 30972 9551
rect 31024 9240 31076 9246
rect 31024 9182 31076 9188
rect 30932 8492 30984 8498
rect 30932 8434 30984 8440
rect 30932 8288 30984 8294
rect 31036 8276 31064 9182
rect 30984 8248 31064 8276
rect 30932 8230 30984 8236
rect 31022 8120 31078 8129
rect 31022 8055 31078 8064
rect 30930 7712 30986 7721
rect 30930 7647 30986 7656
rect 30840 7540 30892 7546
rect 30840 7482 30892 7488
rect 30748 7336 30800 7342
rect 30748 7278 30800 7284
rect 30838 6896 30894 6905
rect 30838 6831 30894 6840
rect 30656 6656 30708 6662
rect 30656 6598 30708 6604
rect 30300 6446 30512 6474
rect 29920 6316 29972 6322
rect 29920 6258 29972 6264
rect 29918 6216 29974 6225
rect 29918 6151 29974 6160
rect 30196 6180 30248 6186
rect 29458 3567 29514 3576
rect 29828 3596 29880 3602
rect 29276 3460 29328 3466
rect 29276 3402 29328 3408
rect 29184 3392 29236 3398
rect 29184 3334 29236 3340
rect 29196 1698 29224 3334
rect 29288 3194 29316 3402
rect 29276 3188 29328 3194
rect 29276 3130 29328 3136
rect 29472 3074 29500 3567
rect 29828 3538 29880 3544
rect 29472 3058 29592 3074
rect 29472 3052 29604 3058
rect 29472 3046 29552 3052
rect 29184 1692 29236 1698
rect 29184 1634 29236 1640
rect 29092 1624 29144 1630
rect 29092 1566 29144 1572
rect 29000 1420 29052 1426
rect 29000 1362 29052 1368
rect 29472 1154 29500 3046
rect 29552 2994 29604 3000
rect 29828 2576 29880 2582
rect 29828 2518 29880 2524
rect 29840 2106 29868 2518
rect 29828 2100 29880 2106
rect 29828 2042 29880 2048
rect 29460 1148 29512 1154
rect 29460 1090 29512 1096
rect 28552 66 28672 82
rect 28552 60 28684 66
rect 28552 56 28632 60
rect 27908 14 28028 42
rect 28538 54 28632 56
rect 28538 0 28594 54
rect 29288 56 29408 82
rect 28632 2 28684 8
rect 29274 54 29408 56
rect 29274 0 29330 54
rect 29380 42 29408 54
rect 29932 42 29960 6151
rect 30196 6122 30248 6128
rect 30208 5846 30236 6122
rect 30196 5840 30248 5846
rect 30196 5782 30248 5788
rect 30288 5704 30340 5710
rect 30288 5646 30340 5652
rect 30392 5658 30420 6446
rect 30656 6248 30708 6254
rect 30656 6190 30708 6196
rect 30668 6089 30696 6190
rect 30654 6080 30710 6089
rect 30654 6015 30710 6024
rect 30668 5778 30696 6015
rect 30852 5914 30880 6831
rect 30944 6254 30972 7647
rect 30932 6248 30984 6254
rect 30932 6190 30984 6196
rect 30840 5908 30892 5914
rect 30840 5850 30892 5856
rect 30656 5772 30708 5778
rect 30656 5714 30708 5720
rect 30932 5772 30984 5778
rect 30932 5714 30984 5720
rect 30194 5536 30250 5545
rect 30194 5471 30250 5480
rect 30010 2952 30066 2961
rect 30010 2887 30066 2896
rect 30024 56 30052 2887
rect 30208 1873 30236 5471
rect 30300 4196 30328 5646
rect 30392 5630 30788 5658
rect 30484 5574 30512 5630
rect 30472 5568 30524 5574
rect 30472 5510 30524 5516
rect 30760 5250 30788 5630
rect 30944 5370 30972 5714
rect 31036 5370 31064 8055
rect 31128 7818 31156 11194
rect 31404 8430 31432 11194
rect 31484 9920 31536 9926
rect 31484 9862 31536 9868
rect 31300 8424 31352 8430
rect 31300 8366 31352 8372
rect 31392 8424 31444 8430
rect 31392 8366 31444 8372
rect 31496 8378 31524 9862
rect 31576 9648 31628 9654
rect 31576 9590 31628 9596
rect 31680 9602 31708 11194
rect 31758 9888 31814 9897
rect 31758 9823 31814 9832
rect 31772 9722 31800 9823
rect 31760 9716 31812 9722
rect 31760 9658 31812 9664
rect 31852 9648 31904 9654
rect 31680 9596 31852 9602
rect 31680 9590 31904 9596
rect 31588 8498 31616 9590
rect 31680 9574 31892 9590
rect 31760 9512 31812 9518
rect 31956 9500 31984 11194
rect 31760 9454 31812 9460
rect 31864 9472 31984 9500
rect 31668 8560 31720 8566
rect 31668 8502 31720 8508
rect 31576 8492 31628 8498
rect 31576 8434 31628 8440
rect 31680 8378 31708 8502
rect 31208 8356 31260 8362
rect 31208 8298 31260 8304
rect 31116 7812 31168 7818
rect 31116 7754 31168 7760
rect 31220 7546 31248 8298
rect 31116 7540 31168 7546
rect 31116 7482 31168 7488
rect 31208 7540 31260 7546
rect 31208 7482 31260 7488
rect 31128 7342 31156 7482
rect 31116 7336 31168 7342
rect 31116 7278 31168 7284
rect 31116 6792 31168 6798
rect 31116 6734 31168 6740
rect 31128 6458 31156 6734
rect 31116 6452 31168 6458
rect 31116 6394 31168 6400
rect 31312 6322 31340 8366
rect 31496 8350 31708 8378
rect 31668 8288 31720 8294
rect 31668 8230 31720 8236
rect 31680 8090 31708 8230
rect 31668 8084 31720 8090
rect 31668 8026 31720 8032
rect 31772 7886 31800 9454
rect 31864 7954 31892 9472
rect 31944 9376 31996 9382
rect 31944 9318 31996 9324
rect 31956 8634 31984 9318
rect 31944 8628 31996 8634
rect 31944 8570 31996 8576
rect 32232 8378 32260 11194
rect 32404 9172 32456 9178
rect 32404 9114 32456 9120
rect 32232 8350 32352 8378
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 32324 8090 32352 8350
rect 32312 8084 32364 8090
rect 32312 8026 32364 8032
rect 32416 8022 32444 9114
rect 32508 8634 32536 11194
rect 32680 9648 32732 9654
rect 32680 9590 32732 9596
rect 32586 9344 32642 9353
rect 32586 9279 32642 9288
rect 32496 8628 32548 8634
rect 32496 8570 32548 8576
rect 32404 8016 32456 8022
rect 32310 7984 32366 7993
rect 31852 7948 31904 7954
rect 32404 7958 32456 7964
rect 32310 7919 32366 7928
rect 31852 7890 31904 7896
rect 31392 7880 31444 7886
rect 31392 7822 31444 7828
rect 31760 7880 31812 7886
rect 31760 7822 31812 7828
rect 31404 7585 31432 7822
rect 31668 7744 31720 7750
rect 31668 7686 31720 7692
rect 31760 7744 31812 7750
rect 31760 7686 31812 7692
rect 31852 7744 31904 7750
rect 31852 7686 31904 7692
rect 32128 7744 32180 7750
rect 32128 7686 32180 7692
rect 31390 7576 31446 7585
rect 31390 7511 31446 7520
rect 31484 7540 31536 7546
rect 31484 7482 31536 7488
rect 31392 7268 31444 7274
rect 31392 7210 31444 7216
rect 31300 6316 31352 6322
rect 31300 6258 31352 6264
rect 31116 6248 31168 6254
rect 31116 6190 31168 6196
rect 31128 5574 31156 6190
rect 31208 6180 31260 6186
rect 31208 6122 31260 6128
rect 31220 5710 31248 6122
rect 31208 5704 31260 5710
rect 31208 5646 31260 5652
rect 31300 5704 31352 5710
rect 31300 5646 31352 5652
rect 31116 5568 31168 5574
rect 31220 5545 31248 5646
rect 31116 5510 31168 5516
rect 31206 5536 31262 5545
rect 31206 5471 31262 5480
rect 30932 5364 30984 5370
rect 30932 5306 30984 5312
rect 31024 5364 31076 5370
rect 31024 5306 31076 5312
rect 31312 5250 31340 5646
rect 31404 5302 31432 7210
rect 30564 5228 30616 5234
rect 30760 5222 31340 5250
rect 31392 5296 31444 5302
rect 31392 5238 31444 5244
rect 30564 5170 30616 5176
rect 30576 5001 30604 5170
rect 30562 4992 30618 5001
rect 30562 4927 30618 4936
rect 30472 4616 30524 4622
rect 30472 4558 30524 4564
rect 30380 4208 30432 4214
rect 30300 4168 30380 4196
rect 30380 4150 30432 4156
rect 30288 3528 30340 3534
rect 30288 3470 30340 3476
rect 30300 3369 30328 3470
rect 30286 3360 30342 3369
rect 30286 3295 30342 3304
rect 30392 2825 30420 4150
rect 30484 4078 30512 4558
rect 30564 4480 30616 4486
rect 30564 4422 30616 4428
rect 30576 4146 30604 4422
rect 30564 4140 30616 4146
rect 30564 4082 30616 4088
rect 30472 4072 30524 4078
rect 30472 4014 30524 4020
rect 30944 3890 30972 5222
rect 31496 5166 31524 7482
rect 31680 7426 31708 7686
rect 31772 7546 31800 7686
rect 31760 7540 31812 7546
rect 31760 7482 31812 7488
rect 31680 7398 31800 7426
rect 31772 6934 31800 7398
rect 31760 6928 31812 6934
rect 31760 6870 31812 6876
rect 31864 6610 31892 7686
rect 32140 7313 32168 7686
rect 32126 7304 32182 7313
rect 32126 7239 32182 7248
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 32220 6928 32272 6934
rect 32220 6870 32272 6876
rect 32036 6792 32088 6798
rect 32036 6734 32088 6740
rect 31680 6582 31892 6610
rect 31680 6361 31708 6582
rect 31850 6488 31906 6497
rect 31760 6452 31812 6458
rect 32048 6458 32076 6734
rect 31850 6423 31906 6432
rect 32036 6452 32088 6458
rect 31760 6394 31812 6400
rect 31666 6352 31722 6361
rect 31666 6287 31722 6296
rect 31772 6236 31800 6394
rect 31864 6254 31892 6423
rect 32036 6394 32088 6400
rect 31680 6208 31800 6236
rect 31852 6248 31904 6254
rect 31680 6089 31708 6208
rect 31852 6190 31904 6196
rect 32232 6118 32260 6870
rect 31852 6112 31904 6118
rect 31666 6080 31722 6089
rect 31852 6054 31904 6060
rect 32220 6112 32272 6118
rect 32220 6054 32272 6060
rect 31666 6015 31722 6024
rect 31576 5908 31628 5914
rect 31576 5850 31628 5856
rect 31484 5160 31536 5166
rect 31484 5102 31536 5108
rect 31484 4820 31536 4826
rect 31484 4762 31536 4768
rect 31390 4720 31446 4729
rect 31390 4655 31446 4664
rect 31022 4584 31078 4593
rect 31022 4519 31024 4528
rect 31076 4519 31078 4528
rect 31208 4548 31260 4554
rect 31024 4490 31076 4496
rect 31208 4490 31260 4496
rect 31220 4282 31248 4490
rect 31208 4276 31260 4282
rect 31208 4218 31260 4224
rect 31114 4176 31170 4185
rect 31114 4111 31170 4120
rect 30668 3862 30972 3890
rect 30470 3768 30526 3777
rect 30470 3703 30526 3712
rect 30484 3670 30512 3703
rect 30472 3664 30524 3670
rect 30472 3606 30524 3612
rect 30472 2848 30524 2854
rect 30378 2816 30434 2825
rect 30472 2790 30524 2796
rect 30378 2751 30434 2760
rect 30484 2446 30512 2790
rect 30472 2440 30524 2446
rect 30472 2382 30524 2388
rect 30288 2304 30340 2310
rect 30288 2246 30340 2252
rect 30194 1864 30250 1873
rect 30194 1799 30250 1808
rect 30300 1601 30328 2246
rect 30286 1592 30342 1601
rect 30286 1527 30342 1536
rect 30668 1465 30696 3862
rect 30748 3596 30800 3602
rect 30800 3556 30880 3584
rect 30748 3538 30800 3544
rect 30852 3058 30880 3556
rect 30932 3528 30984 3534
rect 30932 3470 30984 3476
rect 30944 3194 30972 3470
rect 30932 3188 30984 3194
rect 30932 3130 30984 3136
rect 30840 3052 30892 3058
rect 30840 2994 30892 3000
rect 30748 2984 30800 2990
rect 30748 2926 30800 2932
rect 30760 2825 30788 2926
rect 30746 2816 30802 2825
rect 30746 2751 30802 2760
rect 30760 2310 30788 2751
rect 30748 2304 30800 2310
rect 30748 2246 30800 2252
rect 30654 1456 30710 1465
rect 30654 1391 30710 1400
rect 30760 56 30880 82
rect 29380 14 29960 42
rect 30010 0 30066 56
rect 30746 54 30880 56
rect 30746 0 30802 54
rect 30852 42 30880 54
rect 31128 42 31156 4111
rect 31208 3936 31260 3942
rect 31208 3878 31260 3884
rect 31220 3534 31248 3878
rect 31208 3528 31260 3534
rect 31208 3470 31260 3476
rect 31220 2394 31248 3470
rect 31300 3188 31352 3194
rect 31300 3130 31352 3136
rect 31312 3097 31340 3130
rect 31298 3088 31354 3097
rect 31298 3023 31354 3032
rect 31404 2417 31432 4655
rect 31496 4593 31524 4762
rect 31482 4584 31538 4593
rect 31482 4519 31538 4528
rect 31484 3052 31536 3058
rect 31484 2994 31536 3000
rect 31496 2650 31524 2994
rect 31484 2644 31536 2650
rect 31484 2586 31536 2592
rect 31588 2530 31616 5850
rect 31680 4536 31708 6015
rect 31864 5778 31892 6054
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 32324 5794 32352 7919
rect 32404 7880 32456 7886
rect 32404 7822 32456 7828
rect 32416 7546 32444 7822
rect 32404 7540 32456 7546
rect 32404 7482 32456 7488
rect 32600 7426 32628 9279
rect 32692 7886 32720 9590
rect 32784 8362 32812 11194
rect 32864 9308 32916 9314
rect 32864 9250 32916 9256
rect 32772 8356 32824 8362
rect 32772 8298 32824 8304
rect 32680 7880 32732 7886
rect 32680 7822 32732 7828
rect 32680 7744 32732 7750
rect 32680 7686 32732 7692
rect 32692 7546 32720 7686
rect 32680 7540 32732 7546
rect 32680 7482 32732 7488
rect 32416 7398 32628 7426
rect 32416 6458 32444 7398
rect 32496 7336 32548 7342
rect 32692 7290 32720 7482
rect 32496 7278 32548 7284
rect 32404 6452 32456 6458
rect 32404 6394 32456 6400
rect 32508 6186 32536 7278
rect 32600 7262 32720 7290
rect 32600 6866 32628 7262
rect 32680 7200 32732 7206
rect 32680 7142 32732 7148
rect 32692 7041 32720 7142
rect 32678 7032 32734 7041
rect 32678 6967 32734 6976
rect 32876 6882 32904 9250
rect 33060 8838 33088 11194
rect 33336 9092 33364 11194
rect 33336 9064 33456 9092
rect 33048 8832 33100 8838
rect 33048 8774 33100 8780
rect 33010 8732 33318 8741
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 33010 8667 33318 8676
rect 33428 8430 33456 9064
rect 33416 8424 33468 8430
rect 33416 8366 33468 8372
rect 33612 8090 33640 11194
rect 33888 8838 33916 11194
rect 33784 8832 33836 8838
rect 33784 8774 33836 8780
rect 33876 8832 33928 8838
rect 33876 8774 33928 8780
rect 33796 8634 33824 8774
rect 34164 8634 34192 11194
rect 34336 8832 34388 8838
rect 34336 8774 34388 8780
rect 33784 8628 33836 8634
rect 33784 8570 33836 8576
rect 34152 8628 34204 8634
rect 34152 8570 34204 8576
rect 33784 8492 33836 8498
rect 33784 8434 33836 8440
rect 33600 8084 33652 8090
rect 33600 8026 33652 8032
rect 32954 7848 33010 7857
rect 32954 7783 33010 7792
rect 32968 7750 32996 7783
rect 32956 7744 33008 7750
rect 32956 7686 33008 7692
rect 33010 7644 33318 7653
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 32588 6860 32640 6866
rect 32588 6802 32640 6808
rect 32692 6854 32904 6882
rect 32588 6316 32640 6322
rect 32588 6258 32640 6264
rect 32496 6180 32548 6186
rect 32496 6122 32548 6128
rect 31852 5772 31904 5778
rect 32324 5766 32444 5794
rect 31852 5714 31904 5720
rect 32312 5704 32364 5710
rect 32312 5646 32364 5652
rect 31852 5364 31904 5370
rect 31772 5324 31852 5352
rect 31772 4690 31800 5324
rect 31852 5306 31904 5312
rect 32324 5234 32352 5646
rect 32312 5228 32364 5234
rect 32312 5170 32364 5176
rect 31852 5024 31904 5030
rect 31852 4966 31904 4972
rect 32312 5024 32364 5030
rect 32312 4966 32364 4972
rect 31864 4690 31892 4966
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 32324 4758 32352 4966
rect 32312 4752 32364 4758
rect 31942 4720 31998 4729
rect 31760 4684 31812 4690
rect 31760 4626 31812 4632
rect 31852 4684 31904 4690
rect 32312 4694 32364 4700
rect 31942 4655 31998 4664
rect 31852 4626 31904 4632
rect 31852 4548 31904 4554
rect 31680 4508 31852 4536
rect 31852 4490 31904 4496
rect 31760 4208 31812 4214
rect 31760 4150 31812 4156
rect 31666 3768 31722 3777
rect 31666 3703 31668 3712
rect 31720 3703 31722 3712
rect 31668 3674 31720 3680
rect 31772 3534 31800 4150
rect 31864 3602 31892 4490
rect 31956 4486 31984 4655
rect 31944 4480 31996 4486
rect 31944 4422 31996 4428
rect 32416 4298 32444 5766
rect 32508 5710 32536 6122
rect 32496 5704 32548 5710
rect 32496 5646 32548 5652
rect 32232 4270 32444 4298
rect 32232 4214 32260 4270
rect 32220 4208 32272 4214
rect 32600 4162 32628 6258
rect 32692 5574 32720 6854
rect 32772 6792 32824 6798
rect 32772 6734 32824 6740
rect 32864 6792 32916 6798
rect 32864 6734 32916 6740
rect 32784 6390 32812 6734
rect 32876 6458 32904 6734
rect 33508 6656 33560 6662
rect 33508 6598 33560 6604
rect 33010 6556 33318 6565
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 32864 6452 32916 6458
rect 32864 6394 32916 6400
rect 32772 6384 32824 6390
rect 32772 6326 32824 6332
rect 33520 6322 33548 6598
rect 33508 6316 33560 6322
rect 33508 6258 33560 6264
rect 32772 6248 32824 6254
rect 32772 6190 32824 6196
rect 32784 5914 32812 6190
rect 32772 5908 32824 5914
rect 32772 5850 32824 5856
rect 33416 5704 33468 5710
rect 33416 5646 33468 5652
rect 32680 5568 32732 5574
rect 32680 5510 32732 5516
rect 32692 5370 32720 5510
rect 33010 5468 33318 5477
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 33010 5403 33318 5412
rect 32680 5364 32732 5370
rect 32680 5306 32732 5312
rect 32772 5296 32824 5302
rect 32772 5238 32824 5244
rect 32680 5160 32732 5166
rect 32680 5102 32732 5108
rect 32692 4826 32720 5102
rect 32680 4820 32732 4826
rect 32680 4762 32732 4768
rect 32692 4690 32720 4762
rect 32784 4690 32812 5238
rect 32680 4684 32732 4690
rect 32680 4626 32732 4632
rect 32772 4684 32824 4690
rect 32772 4626 32824 4632
rect 32956 4616 33008 4622
rect 32876 4576 32956 4604
rect 32876 4282 32904 4576
rect 32956 4558 33008 4564
rect 33010 4380 33318 4389
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 32864 4276 32916 4282
rect 32864 4218 32916 4224
rect 33428 4162 33456 5646
rect 33692 4616 33744 4622
rect 33692 4558 33744 4564
rect 33600 4480 33652 4486
rect 33600 4422 33652 4428
rect 32220 4150 32272 4156
rect 32324 4134 32628 4162
rect 33336 4134 33456 4162
rect 33508 4140 33560 4146
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 32036 3664 32088 3670
rect 32036 3606 32088 3612
rect 31852 3596 31904 3602
rect 31852 3538 31904 3544
rect 31760 3528 31812 3534
rect 31760 3470 31812 3476
rect 32048 3369 32076 3606
rect 32034 3360 32090 3369
rect 32034 3295 32090 3304
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 31496 2502 31616 2530
rect 31390 2408 31446 2417
rect 31220 2366 31340 2394
rect 31312 2310 31340 2366
rect 31390 2343 31446 2352
rect 31300 2304 31352 2310
rect 31300 2246 31352 2252
rect 31496 56 31524 2502
rect 32324 2106 32352 4134
rect 33336 3942 33364 4134
rect 33508 4082 33560 4088
rect 33416 4072 33468 4078
rect 33416 4014 33468 4020
rect 32772 3936 32824 3942
rect 32772 3878 32824 3884
rect 33324 3936 33376 3942
rect 33324 3878 33376 3884
rect 32312 2100 32364 2106
rect 32312 2042 32364 2048
rect 32784 1358 32812 3878
rect 33428 3738 33456 4014
rect 33324 3732 33376 3738
rect 33324 3674 33376 3680
rect 33416 3732 33468 3738
rect 33416 3674 33468 3680
rect 33336 3534 33364 3674
rect 33324 3528 33376 3534
rect 33324 3470 33376 3476
rect 33428 3398 33456 3674
rect 33520 3641 33548 4082
rect 33506 3632 33562 3641
rect 33506 3567 33562 3576
rect 33416 3392 33468 3398
rect 33416 3334 33468 3340
rect 33010 3292 33318 3301
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 32956 2848 33008 2854
rect 32956 2790 33008 2796
rect 32968 2514 32996 2790
rect 33428 2650 33456 3334
rect 33416 2644 33468 2650
rect 33416 2586 33468 2592
rect 33612 2514 33640 4422
rect 33704 4282 33732 4558
rect 33692 4276 33744 4282
rect 33692 4218 33744 4224
rect 33692 3936 33744 3942
rect 33692 3878 33744 3884
rect 33704 3602 33732 3878
rect 33692 3596 33744 3602
rect 33692 3538 33744 3544
rect 33692 3460 33744 3466
rect 33692 3402 33744 3408
rect 32956 2508 33008 2514
rect 32956 2450 33008 2456
rect 33600 2508 33652 2514
rect 33600 2450 33652 2456
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 33010 2204 33318 2213
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 32956 2100 33008 2106
rect 32956 2042 33008 2048
rect 32772 1352 32824 1358
rect 32772 1294 32824 1300
rect 32220 1012 32272 1018
rect 32220 954 32272 960
rect 32232 56 32260 954
rect 32968 56 32996 2042
rect 33428 746 33456 2382
rect 33416 740 33468 746
rect 33416 682 33468 688
rect 33704 56 33732 3402
rect 33796 3194 33824 8434
rect 34348 8362 34376 8774
rect 34336 8356 34388 8362
rect 34336 8298 34388 8304
rect 34440 8090 34468 11194
rect 34520 8832 34572 8838
rect 34520 8774 34572 8780
rect 34532 8566 34560 8774
rect 34716 8634 34744 11194
rect 34704 8628 34756 8634
rect 34704 8570 34756 8576
rect 34520 8560 34572 8566
rect 34520 8502 34572 8508
rect 34520 8424 34572 8430
rect 34520 8366 34572 8372
rect 34794 8392 34850 8401
rect 34428 8084 34480 8090
rect 34428 8026 34480 8032
rect 33876 7880 33928 7886
rect 33876 7822 33928 7828
rect 34152 7880 34204 7886
rect 34152 7822 34204 7828
rect 34334 7848 34390 7857
rect 33888 3942 33916 7822
rect 34164 7478 34192 7822
rect 34334 7783 34390 7792
rect 34348 7750 34376 7783
rect 34336 7744 34388 7750
rect 34336 7686 34388 7692
rect 34152 7472 34204 7478
rect 34152 7414 34204 7420
rect 34244 7404 34296 7410
rect 34244 7346 34296 7352
rect 33968 6316 34020 6322
rect 33968 6258 34020 6264
rect 33980 5681 34008 6258
rect 33966 5672 34022 5681
rect 34022 5630 34192 5658
rect 33966 5607 34022 5616
rect 33968 5092 34020 5098
rect 33968 5034 34020 5040
rect 33980 4758 34008 5034
rect 33968 4752 34020 4758
rect 33968 4694 34020 4700
rect 34060 4276 34112 4282
rect 34060 4218 34112 4224
rect 34072 4146 34100 4218
rect 34060 4140 34112 4146
rect 34060 4082 34112 4088
rect 33876 3936 33928 3942
rect 33876 3878 33928 3884
rect 34164 3398 34192 5630
rect 33876 3392 33928 3398
rect 33876 3334 33928 3340
rect 34152 3392 34204 3398
rect 34152 3334 34204 3340
rect 33784 3188 33836 3194
rect 33784 3130 33836 3136
rect 33784 3052 33836 3058
rect 33888 3040 33916 3334
rect 33836 3012 33916 3040
rect 33784 2994 33836 3000
rect 34256 1018 34284 7346
rect 34336 4208 34388 4214
rect 34336 4150 34388 4156
rect 34348 2774 34376 4150
rect 34428 4072 34480 4078
rect 34428 4014 34480 4020
rect 34440 3738 34468 4014
rect 34532 3738 34560 8366
rect 34992 8362 35020 11194
rect 35070 9208 35126 9217
rect 35070 9143 35126 9152
rect 34794 8327 34850 8336
rect 34980 8356 35032 8362
rect 34704 6316 34756 6322
rect 34704 6258 34756 6264
rect 34428 3732 34480 3738
rect 34428 3674 34480 3680
rect 34520 3732 34572 3738
rect 34520 3674 34572 3680
rect 34440 3058 34468 3674
rect 34716 3534 34744 6258
rect 34808 4758 34836 8327
rect 34980 8298 35032 8304
rect 34888 8288 34940 8294
rect 34888 8230 34940 8236
rect 34900 7342 34928 8230
rect 34888 7336 34940 7342
rect 34888 7278 34940 7284
rect 35084 5030 35112 9143
rect 35268 8362 35296 11194
rect 35348 8968 35400 8974
rect 35348 8910 35400 8916
rect 35360 8498 35388 8910
rect 35438 8528 35494 8537
rect 35348 8492 35400 8498
rect 35438 8463 35494 8472
rect 35348 8434 35400 8440
rect 35256 8356 35308 8362
rect 35256 8298 35308 8304
rect 35348 8016 35400 8022
rect 35348 7958 35400 7964
rect 35164 7880 35216 7886
rect 35164 7822 35216 7828
rect 35072 5024 35124 5030
rect 35072 4966 35124 4972
rect 34796 4752 34848 4758
rect 34796 4694 34848 4700
rect 34980 4752 35032 4758
rect 34980 4694 35032 4700
rect 34992 4622 35020 4694
rect 34980 4616 35032 4622
rect 34980 4558 35032 4564
rect 35176 4185 35204 7822
rect 35256 5296 35308 5302
rect 35256 5238 35308 5244
rect 35268 4554 35296 5238
rect 35256 4548 35308 4554
rect 35256 4490 35308 4496
rect 35162 4176 35218 4185
rect 35162 4111 35218 4120
rect 35256 4140 35308 4146
rect 35256 4082 35308 4088
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 34980 3528 35032 3534
rect 35268 3482 35296 4082
rect 34980 3470 35032 3476
rect 34992 3398 35020 3470
rect 35084 3454 35296 3482
rect 34980 3392 35032 3398
rect 34980 3334 35032 3340
rect 34428 3052 34480 3058
rect 34428 2994 34480 3000
rect 34348 2746 34468 2774
rect 34244 1012 34296 1018
rect 34244 954 34296 960
rect 34440 56 34468 2746
rect 35084 1086 35112 3454
rect 35360 2774 35388 7958
rect 35452 6458 35480 8463
rect 35544 8090 35572 11194
rect 35820 8634 35848 11194
rect 35808 8628 35860 8634
rect 35808 8570 35860 8576
rect 35716 8492 35768 8498
rect 35716 8434 35768 8440
rect 35808 8492 35860 8498
rect 35808 8434 35860 8440
rect 35624 8424 35676 8430
rect 35624 8366 35676 8372
rect 35532 8084 35584 8090
rect 35532 8026 35584 8032
rect 35532 7880 35584 7886
rect 35532 7822 35584 7828
rect 35544 6848 35572 7822
rect 35636 7750 35664 8366
rect 35624 7744 35676 7750
rect 35624 7686 35676 7692
rect 35544 6820 35664 6848
rect 35532 6724 35584 6730
rect 35532 6666 35584 6672
rect 35440 6452 35492 6458
rect 35440 6394 35492 6400
rect 35544 6390 35572 6666
rect 35532 6384 35584 6390
rect 35532 6326 35584 6332
rect 35440 6112 35492 6118
rect 35440 6054 35492 6060
rect 35452 5778 35480 6054
rect 35440 5772 35492 5778
rect 35440 5714 35492 5720
rect 35532 5568 35584 5574
rect 35532 5510 35584 5516
rect 35544 4486 35572 5510
rect 35636 4808 35664 6820
rect 35728 5574 35756 8434
rect 35820 7546 35848 8434
rect 36096 8090 36124 11194
rect 36372 8362 36400 11194
rect 36452 10464 36504 10470
rect 36452 10406 36504 10412
rect 36360 8356 36412 8362
rect 36360 8298 36412 8304
rect 36084 8084 36136 8090
rect 36084 8026 36136 8032
rect 36084 7948 36136 7954
rect 36084 7890 36136 7896
rect 36176 7948 36228 7954
rect 36176 7890 36228 7896
rect 35900 7880 35952 7886
rect 35900 7822 35952 7828
rect 35808 7540 35860 7546
rect 35808 7482 35860 7488
rect 35912 5658 35940 7822
rect 36096 6458 36124 7890
rect 36084 6452 36136 6458
rect 36084 6394 36136 6400
rect 35992 6316 36044 6322
rect 35992 6258 36044 6264
rect 36004 5914 36032 6258
rect 35992 5908 36044 5914
rect 35992 5850 36044 5856
rect 35912 5630 36032 5658
rect 35716 5568 35768 5574
rect 35716 5510 35768 5516
rect 35900 5228 35952 5234
rect 35900 5170 35952 5176
rect 35912 4826 35940 5170
rect 35900 4820 35952 4826
rect 35636 4780 35756 4808
rect 35624 4684 35676 4690
rect 35624 4626 35676 4632
rect 35532 4480 35584 4486
rect 35532 4422 35584 4428
rect 35636 4282 35664 4626
rect 35624 4276 35676 4282
rect 35624 4218 35676 4224
rect 35176 2746 35388 2774
rect 35072 1080 35124 1086
rect 35072 1022 35124 1028
rect 35176 56 35204 2746
rect 35728 1426 35756 4780
rect 35900 4762 35952 4768
rect 36004 3738 36032 5630
rect 35992 3732 36044 3738
rect 35992 3674 36044 3680
rect 35716 1420 35768 1426
rect 35716 1362 35768 1368
rect 35912 56 36032 82
rect 30852 14 31156 42
rect 31482 0 31538 56
rect 32218 0 32274 56
rect 32954 0 33010 56
rect 33690 0 33746 56
rect 34426 0 34482 56
rect 35162 0 35218 56
rect 35898 54 36032 56
rect 35898 0 35954 54
rect 36004 42 36032 54
rect 36188 42 36216 7890
rect 36360 7880 36412 7886
rect 36360 7822 36412 7828
rect 36372 7750 36400 7822
rect 36360 7744 36412 7750
rect 36360 7686 36412 7692
rect 36464 5914 36492 10406
rect 36544 8968 36596 8974
rect 36544 8910 36596 8916
rect 36452 5908 36504 5914
rect 36452 5850 36504 5856
rect 36452 4684 36504 4690
rect 36452 4626 36504 4632
rect 36266 4584 36322 4593
rect 36266 4519 36322 4528
rect 36280 3466 36308 4519
rect 36464 4282 36492 4626
rect 36452 4276 36504 4282
rect 36452 4218 36504 4224
rect 36268 3460 36320 3466
rect 36268 3402 36320 3408
rect 36556 3194 36584 8910
rect 36648 8090 36676 11194
rect 36924 8634 36952 11194
rect 37004 8832 37056 8838
rect 37004 8774 37056 8780
rect 36912 8628 36964 8634
rect 36912 8570 36964 8576
rect 36728 8492 36780 8498
rect 36728 8434 36780 8440
rect 36820 8492 36872 8498
rect 36820 8434 36872 8440
rect 36636 8084 36688 8090
rect 36636 8026 36688 8032
rect 36636 7880 36688 7886
rect 36634 7848 36636 7857
rect 36688 7848 36690 7857
rect 36634 7783 36690 7792
rect 36636 7472 36688 7478
rect 36636 7414 36688 7420
rect 36544 3188 36596 3194
rect 36544 3130 36596 3136
rect 36648 56 36676 7414
rect 36740 4758 36768 8434
rect 36832 4826 36860 8434
rect 36912 7336 36964 7342
rect 36912 7278 36964 7284
rect 36924 5273 36952 7278
rect 37016 6730 37044 8774
rect 37096 8560 37148 8566
rect 37096 8502 37148 8508
rect 37108 7546 37136 8502
rect 37200 8362 37228 11194
rect 37476 8566 37504 11194
rect 37648 10260 37700 10266
rect 37648 10202 37700 10208
rect 37554 9752 37610 9761
rect 37554 9687 37610 9696
rect 37464 8560 37516 8566
rect 37464 8502 37516 8508
rect 37280 8492 37332 8498
rect 37280 8434 37332 8440
rect 37188 8356 37240 8362
rect 37188 8298 37240 8304
rect 37292 8090 37320 8434
rect 37280 8084 37332 8090
rect 37280 8026 37332 8032
rect 37372 7948 37424 7954
rect 37372 7890 37424 7896
rect 37096 7540 37148 7546
rect 37096 7482 37148 7488
rect 37004 6724 37056 6730
rect 37004 6666 37056 6672
rect 36910 5264 36966 5273
rect 36910 5199 36966 5208
rect 36820 4820 36872 4826
rect 36820 4762 36872 4768
rect 36728 4752 36780 4758
rect 36728 4694 36780 4700
rect 37188 4684 37240 4690
rect 37188 4626 37240 4632
rect 37200 950 37228 4626
rect 37280 4548 37332 4554
rect 37280 4490 37332 4496
rect 37292 1329 37320 4490
rect 37278 1320 37334 1329
rect 37278 1255 37334 1264
rect 37188 944 37240 950
rect 37188 886 37240 892
rect 37384 56 37412 7890
rect 37464 7812 37516 7818
rect 37464 7754 37516 7760
rect 37476 7274 37504 7754
rect 37568 7750 37596 9687
rect 37660 7834 37688 10202
rect 37752 8022 37780 11194
rect 38474 10160 38530 10169
rect 38474 10095 38530 10104
rect 38290 9888 38346 9897
rect 38290 9823 38346 9832
rect 37832 8492 37884 8498
rect 37832 8434 37884 8440
rect 37844 8090 37872 8434
rect 37950 8188 38258 8197
rect 37950 8186 37956 8188
rect 38012 8186 38036 8188
rect 38092 8186 38116 8188
rect 38172 8186 38196 8188
rect 38252 8186 38258 8188
rect 38012 8134 38014 8186
rect 38194 8134 38196 8186
rect 37950 8132 37956 8134
rect 38012 8132 38036 8134
rect 38092 8132 38116 8134
rect 38172 8132 38196 8134
rect 38252 8132 38258 8134
rect 37950 8123 38258 8132
rect 37832 8084 37884 8090
rect 37832 8026 37884 8032
rect 37740 8016 37792 8022
rect 37740 7958 37792 7964
rect 37832 7880 37884 7886
rect 37660 7806 37780 7834
rect 37832 7822 37884 7828
rect 37556 7744 37608 7750
rect 37556 7686 37608 7692
rect 37648 7404 37700 7410
rect 37648 7346 37700 7352
rect 37464 7268 37516 7274
rect 37464 7210 37516 7216
rect 37660 6225 37688 7346
rect 37752 7274 37780 7806
rect 37740 7268 37792 7274
rect 37740 7210 37792 7216
rect 37844 7002 37872 7822
rect 38200 7744 38252 7750
rect 38200 7686 38252 7692
rect 38212 7342 38240 7686
rect 38304 7546 38332 9823
rect 38488 7886 38516 10095
rect 39670 9616 39726 9625
rect 39670 9551 39726 9560
rect 38750 9344 38806 9353
rect 38750 9279 38806 9288
rect 38658 8528 38714 8537
rect 38568 8492 38620 8498
rect 38658 8463 38714 8472
rect 38568 8434 38620 8440
rect 38476 7880 38528 7886
rect 38476 7822 38528 7828
rect 38292 7540 38344 7546
rect 38292 7482 38344 7488
rect 38384 7404 38436 7410
rect 38384 7346 38436 7352
rect 38200 7336 38252 7342
rect 38200 7278 38252 7284
rect 37950 7100 38258 7109
rect 37950 7098 37956 7100
rect 38012 7098 38036 7100
rect 38092 7098 38116 7100
rect 38172 7098 38196 7100
rect 38252 7098 38258 7100
rect 38012 7046 38014 7098
rect 38194 7046 38196 7098
rect 37950 7044 37956 7046
rect 38012 7044 38036 7046
rect 38092 7044 38116 7046
rect 38172 7044 38196 7046
rect 38252 7044 38258 7046
rect 37950 7035 38258 7044
rect 37832 6996 37884 7002
rect 37832 6938 37884 6944
rect 38016 6792 38068 6798
rect 38016 6734 38068 6740
rect 37832 6656 37884 6662
rect 37832 6598 37884 6604
rect 37646 6216 37702 6225
rect 37646 6151 37702 6160
rect 37844 5137 37872 6598
rect 38028 6186 38056 6734
rect 38292 6724 38344 6730
rect 38292 6666 38344 6672
rect 38016 6180 38068 6186
rect 38016 6122 38068 6128
rect 37950 6012 38258 6021
rect 37950 6010 37956 6012
rect 38012 6010 38036 6012
rect 38092 6010 38116 6012
rect 38172 6010 38196 6012
rect 38252 6010 38258 6012
rect 38012 5958 38014 6010
rect 38194 5958 38196 6010
rect 37950 5956 37956 5958
rect 38012 5956 38036 5958
rect 38092 5956 38116 5958
rect 38172 5956 38196 5958
rect 38252 5956 38258 5958
rect 37950 5947 38258 5956
rect 37830 5128 37886 5137
rect 37830 5063 37886 5072
rect 37950 4924 38258 4933
rect 37950 4922 37956 4924
rect 38012 4922 38036 4924
rect 38092 4922 38116 4924
rect 38172 4922 38196 4924
rect 38252 4922 38258 4924
rect 38012 4870 38014 4922
rect 38194 4870 38196 4922
rect 37950 4868 37956 4870
rect 38012 4868 38036 4870
rect 38092 4868 38116 4870
rect 38172 4868 38196 4870
rect 38252 4868 38258 4870
rect 37950 4859 38258 4868
rect 37556 4140 37608 4146
rect 37556 4082 37608 4088
rect 37568 4049 37596 4082
rect 37554 4040 37610 4049
rect 37554 3975 37610 3984
rect 37950 3836 38258 3845
rect 37950 3834 37956 3836
rect 38012 3834 38036 3836
rect 38092 3834 38116 3836
rect 38172 3834 38196 3836
rect 38252 3834 38258 3836
rect 38012 3782 38014 3834
rect 38194 3782 38196 3834
rect 37950 3780 37956 3782
rect 38012 3780 38036 3782
rect 38092 3780 38116 3782
rect 38172 3780 38196 3782
rect 38252 3780 38258 3782
rect 37950 3771 38258 3780
rect 37950 2748 38258 2757
rect 37950 2746 37956 2748
rect 38012 2746 38036 2748
rect 38092 2746 38116 2748
rect 38172 2746 38196 2748
rect 38252 2746 38258 2748
rect 38012 2694 38014 2746
rect 38194 2694 38196 2746
rect 37950 2692 37956 2694
rect 38012 2692 38036 2694
rect 38092 2692 38116 2694
rect 38172 2692 38196 2694
rect 38252 2692 38258 2694
rect 37950 2683 38258 2692
rect 38108 2440 38160 2446
rect 38304 2394 38332 6666
rect 38396 3398 38424 7346
rect 38476 6656 38528 6662
rect 38476 6598 38528 6604
rect 38488 5642 38516 6598
rect 38476 5636 38528 5642
rect 38476 5578 38528 5584
rect 38580 5370 38608 8434
rect 38672 8090 38700 8463
rect 38660 8084 38712 8090
rect 38660 8026 38712 8032
rect 38764 7546 38792 9279
rect 38936 8900 38988 8906
rect 38936 8842 38988 8848
rect 38948 8634 38976 8842
rect 39578 8800 39634 8809
rect 39010 8732 39318 8741
rect 39578 8735 39634 8744
rect 39010 8730 39016 8732
rect 39072 8730 39096 8732
rect 39152 8730 39176 8732
rect 39232 8730 39256 8732
rect 39312 8730 39318 8732
rect 39072 8678 39074 8730
rect 39254 8678 39256 8730
rect 39010 8676 39016 8678
rect 39072 8676 39096 8678
rect 39152 8676 39176 8678
rect 39232 8676 39256 8678
rect 39312 8676 39318 8678
rect 39010 8667 39318 8676
rect 38936 8628 38988 8634
rect 38936 8570 38988 8576
rect 39396 8356 39448 8362
rect 39396 8298 39448 8304
rect 39408 7993 39436 8298
rect 39486 8256 39542 8265
rect 39486 8191 39542 8200
rect 39394 7984 39450 7993
rect 39394 7919 39450 7928
rect 38844 7880 38896 7886
rect 38844 7822 38896 7828
rect 38752 7540 38804 7546
rect 38752 7482 38804 7488
rect 38856 7206 38884 7822
rect 38936 7744 38988 7750
rect 39396 7744 39448 7750
rect 38936 7686 38988 7692
rect 39394 7712 39396 7721
rect 39448 7712 39450 7721
rect 38948 7449 38976 7686
rect 39010 7644 39318 7653
rect 39394 7647 39450 7656
rect 39010 7642 39016 7644
rect 39072 7642 39096 7644
rect 39152 7642 39176 7644
rect 39232 7642 39256 7644
rect 39312 7642 39318 7644
rect 39072 7590 39074 7642
rect 39254 7590 39256 7642
rect 39010 7588 39016 7590
rect 39072 7588 39096 7590
rect 39152 7588 39176 7590
rect 39232 7588 39256 7590
rect 39312 7588 39318 7590
rect 39010 7579 39318 7588
rect 39500 7478 39528 8191
rect 39592 7546 39620 8735
rect 39580 7540 39632 7546
rect 39580 7482 39632 7488
rect 39488 7472 39540 7478
rect 38934 7440 38990 7449
rect 39488 7414 39540 7420
rect 38934 7375 38990 7384
rect 38844 7200 38896 7206
rect 38844 7142 38896 7148
rect 39394 7168 39450 7177
rect 39394 7103 39450 7112
rect 38936 6860 38988 6866
rect 38936 6802 38988 6808
rect 38752 6724 38804 6730
rect 38752 6666 38804 6672
rect 38660 6656 38712 6662
rect 38660 6598 38712 6604
rect 38672 6361 38700 6598
rect 38658 6352 38714 6361
rect 38658 6287 38714 6296
rect 38764 5386 38792 6666
rect 38948 6322 38976 6802
rect 39408 6662 39436 7103
rect 39684 6730 39712 9551
rect 39854 9072 39910 9081
rect 39854 9007 39910 9016
rect 39672 6724 39724 6730
rect 39672 6666 39724 6672
rect 39396 6656 39448 6662
rect 39396 6598 39448 6604
rect 39670 6624 39726 6633
rect 39010 6556 39318 6565
rect 39670 6559 39726 6568
rect 39010 6554 39016 6556
rect 39072 6554 39096 6556
rect 39152 6554 39176 6556
rect 39232 6554 39256 6556
rect 39312 6554 39318 6556
rect 39072 6502 39074 6554
rect 39254 6502 39256 6554
rect 39010 6500 39016 6502
rect 39072 6500 39096 6502
rect 39152 6500 39176 6502
rect 39232 6500 39256 6502
rect 39312 6500 39318 6502
rect 39010 6491 39318 6500
rect 38936 6316 38988 6322
rect 38936 6258 38988 6264
rect 39580 6180 39632 6186
rect 39580 6122 39632 6128
rect 39028 6112 39080 6118
rect 39026 6080 39028 6089
rect 39080 6080 39082 6089
rect 39026 6015 39082 6024
rect 38842 5808 38898 5817
rect 38842 5743 38898 5752
rect 39394 5808 39450 5817
rect 39394 5743 39450 5752
rect 38856 5710 38884 5743
rect 38844 5704 38896 5710
rect 38844 5646 38896 5652
rect 39010 5468 39318 5477
rect 39010 5466 39016 5468
rect 39072 5466 39096 5468
rect 39152 5466 39176 5468
rect 39232 5466 39256 5468
rect 39312 5466 39318 5468
rect 39072 5414 39074 5466
rect 39254 5414 39256 5466
rect 39010 5412 39016 5414
rect 39072 5412 39096 5414
rect 39152 5412 39176 5414
rect 39232 5412 39256 5414
rect 39312 5412 39318 5414
rect 39010 5403 39318 5412
rect 38568 5364 38620 5370
rect 38568 5306 38620 5312
rect 38672 5358 38792 5386
rect 39408 5370 39436 5743
rect 39396 5364 39448 5370
rect 38672 5098 38700 5358
rect 39396 5306 39448 5312
rect 39394 5264 39450 5273
rect 38752 5228 38804 5234
rect 39394 5199 39450 5208
rect 38752 5170 38804 5176
rect 38660 5092 38712 5098
rect 38660 5034 38712 5040
rect 38476 4616 38528 4622
rect 38476 4558 38528 4564
rect 38568 4616 38620 4622
rect 38568 4558 38620 4564
rect 38488 4214 38516 4558
rect 38476 4208 38528 4214
rect 38476 4150 38528 4156
rect 38384 3392 38436 3398
rect 38384 3334 38436 3340
rect 38384 3052 38436 3058
rect 38384 2994 38436 3000
rect 38396 2961 38424 2994
rect 38382 2952 38438 2961
rect 38382 2887 38438 2896
rect 38580 2632 38608 4558
rect 38660 3596 38712 3602
rect 38660 3538 38712 3544
rect 38672 3058 38700 3538
rect 38660 3052 38712 3058
rect 38660 2994 38712 3000
rect 38660 2848 38712 2854
rect 38660 2790 38712 2796
rect 38108 2382 38160 2388
rect 37924 2304 37976 2310
rect 37924 2246 37976 2252
rect 37936 2009 37964 2246
rect 37922 2000 37978 2009
rect 37922 1935 37978 1944
rect 38120 1562 38148 2382
rect 38212 2366 38332 2394
rect 38396 2604 38608 2632
rect 38108 1556 38160 1562
rect 38108 1498 38160 1504
rect 38108 1420 38160 1426
rect 38108 1362 38160 1368
rect 38120 56 38148 1362
rect 38212 814 38240 2366
rect 38292 2304 38344 2310
rect 38292 2246 38344 2252
rect 38304 1737 38332 2246
rect 38396 2106 38424 2604
rect 38672 2553 38700 2790
rect 38764 2774 38792 5170
rect 39028 5024 39080 5030
rect 39026 4992 39028 5001
rect 39080 4992 39082 5001
rect 39026 4927 39082 4936
rect 39408 4826 39436 5199
rect 39396 4820 39448 4826
rect 39396 4762 39448 4768
rect 39486 4720 39542 4729
rect 39486 4655 39542 4664
rect 39010 4380 39318 4389
rect 39010 4378 39016 4380
rect 39072 4378 39096 4380
rect 39152 4378 39176 4380
rect 39232 4378 39256 4380
rect 39312 4378 39318 4380
rect 39072 4326 39074 4378
rect 39254 4326 39256 4378
rect 39010 4324 39016 4326
rect 39072 4324 39096 4326
rect 39152 4324 39176 4326
rect 39232 4324 39256 4326
rect 39312 4324 39318 4326
rect 39010 4315 39318 4324
rect 39394 4176 39450 4185
rect 38936 4140 38988 4146
rect 39394 4111 39450 4120
rect 38936 4082 38988 4088
rect 38948 3670 38976 4082
rect 39028 3936 39080 3942
rect 39026 3904 39028 3913
rect 39080 3904 39082 3913
rect 39026 3839 39082 3848
rect 39408 3738 39436 4111
rect 39500 4010 39528 4655
rect 39488 4004 39540 4010
rect 39488 3946 39540 3952
rect 39396 3732 39448 3738
rect 39396 3674 39448 3680
rect 38936 3664 38988 3670
rect 38936 3606 38988 3612
rect 39394 3632 39450 3641
rect 39394 3567 39450 3576
rect 38844 3528 38896 3534
rect 38842 3496 38844 3505
rect 38896 3496 38898 3505
rect 38842 3431 38898 3440
rect 39010 3292 39318 3301
rect 39010 3290 39016 3292
rect 39072 3290 39096 3292
rect 39152 3290 39176 3292
rect 39232 3290 39256 3292
rect 39312 3290 39318 3292
rect 39072 3238 39074 3290
rect 39254 3238 39256 3290
rect 39010 3236 39016 3238
rect 39072 3236 39096 3238
rect 39152 3236 39176 3238
rect 39232 3236 39256 3238
rect 39312 3236 39318 3238
rect 39010 3227 39318 3236
rect 39408 3194 39436 3567
rect 39396 3188 39448 3194
rect 39396 3130 39448 3136
rect 39394 3088 39450 3097
rect 38936 3052 38988 3058
rect 39394 3023 39450 3032
rect 38936 2994 38988 3000
rect 38764 2746 38884 2774
rect 38474 2544 38530 2553
rect 38474 2479 38530 2488
rect 38658 2544 38714 2553
rect 38658 2479 38714 2488
rect 38488 2446 38516 2479
rect 38476 2440 38528 2446
rect 38476 2382 38528 2388
rect 38568 2440 38620 2446
rect 38568 2382 38620 2388
rect 38384 2100 38436 2106
rect 38384 2042 38436 2048
rect 38580 1970 38608 2382
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 38568 1964 38620 1970
rect 38568 1906 38620 1912
rect 38290 1728 38346 1737
rect 38290 1663 38346 1672
rect 38672 1465 38700 2246
rect 38658 1456 38714 1465
rect 38658 1391 38714 1400
rect 38200 808 38252 814
rect 38200 750 38252 756
rect 38856 56 38884 2746
rect 38948 1193 38976 2994
rect 39028 2848 39080 2854
rect 39026 2816 39028 2825
rect 39080 2816 39082 2825
rect 39026 2751 39082 2760
rect 39408 2650 39436 3023
rect 39396 2644 39448 2650
rect 39396 2586 39448 2592
rect 39010 2204 39318 2213
rect 39010 2202 39016 2204
rect 39072 2202 39096 2204
rect 39152 2202 39176 2204
rect 39232 2202 39256 2204
rect 39312 2202 39318 2204
rect 39072 2150 39074 2202
rect 39254 2150 39256 2202
rect 39010 2148 39016 2150
rect 39072 2148 39096 2150
rect 39152 2148 39176 2150
rect 39232 2148 39256 2150
rect 39312 2148 39318 2150
rect 39010 2139 39318 2148
rect 38934 1184 38990 1193
rect 38934 1119 38990 1128
rect 39592 56 39620 6122
rect 39684 5914 39712 6559
rect 39868 6458 39896 9007
rect 40040 7268 40092 7274
rect 40040 7210 40092 7216
rect 40052 6905 40080 7210
rect 40038 6896 40094 6905
rect 40038 6831 40094 6840
rect 39856 6452 39908 6458
rect 39856 6394 39908 6400
rect 39856 6248 39908 6254
rect 39856 6190 39908 6196
rect 39672 5908 39724 5914
rect 39672 5850 39724 5856
rect 39672 5228 39724 5234
rect 39672 5170 39724 5176
rect 39684 1290 39712 5170
rect 39672 1284 39724 1290
rect 39672 1226 39724 1232
rect 39868 66 39896 6190
rect 39948 5840 40000 5846
rect 39948 5782 40000 5788
rect 39960 5545 39988 5782
rect 39946 5536 40002 5545
rect 39946 5471 40002 5480
rect 39948 4752 40000 4758
rect 39948 4694 40000 4700
rect 39960 4457 39988 4694
rect 39946 4448 40002 4457
rect 39946 4383 40002 4392
rect 39948 3664 40000 3670
rect 39948 3606 40000 3612
rect 39960 3369 39988 3606
rect 39946 3360 40002 3369
rect 39946 3295 40002 3304
rect 39948 2576 40000 2582
rect 39948 2518 40000 2524
rect 39960 2281 39988 2518
rect 39946 2272 40002 2281
rect 39946 2207 40002 2216
rect 39856 60 39908 66
rect 36004 14 36216 42
rect 36634 0 36690 56
rect 37370 0 37426 56
rect 38106 0 38162 56
rect 38842 0 38898 56
rect 39578 0 39634 56
rect 39856 2 39908 8
<< via2 >>
rect 2318 10104 2374 10160
rect 478 9832 534 9888
rect 662 9560 718 9616
rect 386 8200 442 8256
rect 1214 9288 1270 9344
rect 754 7928 810 7984
rect 1306 8508 1308 8528
rect 1308 8508 1360 8528
rect 1360 8508 1362 8528
rect 1306 8472 1362 8508
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 754 7656 810 7712
rect 938 7420 940 7440
rect 940 7420 992 7440
rect 992 7420 994 7440
rect 938 7384 994 7420
rect 1122 7112 1178 7168
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 202 6568 258 6624
rect 938 6332 940 6352
rect 940 6332 992 6352
rect 992 6332 994 6352
rect 938 6296 994 6332
rect 754 6024 810 6080
rect 1674 6196 1676 6216
rect 1676 6196 1728 6216
rect 1728 6196 1730 6216
rect 1674 6160 1730 6196
rect 754 5752 810 5808
rect 570 5480 626 5536
rect 386 4936 442 4992
rect 1030 5208 1086 5264
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 2778 9016 2834 9072
rect 2870 8744 2926 8800
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 3974 9968 4030 10024
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 3606 7384 3662 7440
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 938 4664 994 4720
rect 754 4392 810 4448
rect 754 4156 756 4176
rect 756 4156 808 4176
rect 808 4156 810 4176
rect 754 4120 810 4156
rect 1950 4120 2006 4176
rect 2318 4004 2374 4040
rect 2318 3984 2320 4004
rect 2320 3984 2372 4004
rect 2372 3984 2374 4004
rect 938 3848 994 3904
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 2962 6840 3018 6896
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 570 3576 626 3632
rect 2502 3576 2558 3632
rect 202 3304 258 3360
rect 1306 3032 1362 3088
rect 386 2488 442 2544
rect 1214 2760 1270 2816
rect 1122 2216 1178 2272
rect 1214 1672 1270 1728
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 1858 1944 1914 2000
rect 2594 1400 2650 1456
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 3146 2932 3148 2952
rect 3148 2932 3200 2952
rect 3200 2932 3202 2952
rect 3146 2896 3202 2932
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 3422 856 3478 912
rect 4158 6332 4160 6352
rect 4160 6332 4212 6352
rect 4212 6332 4214 6352
rect 4158 6296 4214 6332
rect 3606 720 3662 776
rect 4434 9696 4490 9752
rect 5078 9152 5134 9208
rect 4342 5208 4398 5264
rect 4894 8336 4950 8392
rect 4802 7520 4858 7576
rect 4526 4664 4582 4720
rect 5078 5616 5134 5672
rect 5538 7828 5540 7848
rect 5540 7828 5592 7848
rect 5592 7828 5594 7848
rect 5538 7792 5594 7828
rect 6182 9424 6238 9480
rect 6642 9832 6698 9888
rect 6734 9696 6790 9752
rect 6642 8492 6698 8528
rect 6642 8472 6644 8492
rect 6644 8472 6696 8492
rect 6696 8472 6698 8492
rect 6826 7948 6882 7984
rect 6826 7928 6828 7948
rect 6828 7928 6880 7948
rect 6880 7928 6882 7948
rect 5814 5344 5870 5400
rect 5262 4120 5318 4176
rect 4710 2624 4766 2680
rect 3882 1264 3938 1320
rect 3790 584 3846 640
rect 5446 3032 5502 3088
rect 5722 3476 5724 3496
rect 5724 3476 5776 3496
rect 5776 3476 5778 3496
rect 5722 3440 5778 3476
rect 5630 992 5686 1048
rect 5906 5072 5962 5128
rect 6642 5752 6698 5808
rect 6458 5072 6514 5128
rect 7378 9696 7434 9752
rect 7378 8880 7434 8936
rect 7102 7248 7158 7304
rect 7378 7248 7434 7304
rect 7286 6840 7342 6896
rect 7286 6568 7342 6624
rect 7102 5480 7158 5536
rect 7286 5108 7288 5128
rect 7288 5108 7340 5128
rect 7340 5108 7342 5128
rect 7286 5072 7342 5108
rect 7194 4936 7250 4992
rect 6550 2624 6606 2680
rect 7470 7112 7526 7168
rect 7562 6704 7618 6760
rect 8482 9832 8538 9888
rect 8298 9560 8354 9616
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 7654 5616 7710 5672
rect 7654 5072 7710 5128
rect 7654 4548 7710 4584
rect 7654 4528 7656 4548
rect 7656 4528 7708 4548
rect 7708 4528 7710 4548
rect 7654 3440 7710 3496
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 8390 7112 8446 7168
rect 7930 6452 7986 6488
rect 7930 6432 7932 6452
rect 7932 6432 7984 6452
rect 7984 6432 7986 6452
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 8206 5480 8262 5536
rect 8206 5072 8262 5128
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 7746 2488 7802 2544
rect 7378 1128 7434 1184
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 8482 6568 8538 6624
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 9034 8336 9090 8392
rect 9494 9288 9550 9344
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 9494 7112 9550 7168
rect 9678 9016 9734 9072
rect 9862 8744 9918 8800
rect 9770 8064 9826 8120
rect 9954 8064 10010 8120
rect 9954 7656 10010 7712
rect 9954 6996 10010 7032
rect 9954 6976 9956 6996
rect 9956 6976 10008 6996
rect 10008 6976 10010 6996
rect 10138 6976 10194 7032
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 8758 6432 8814 6488
rect 9954 6840 10010 6896
rect 9770 6568 9826 6624
rect 9954 6296 10010 6352
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 9494 5616 9550 5672
rect 9770 5616 9826 5672
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 8850 5344 8906 5400
rect 9402 5072 9458 5128
rect 8666 4256 8722 4312
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 9402 3984 9458 4040
rect 9862 4256 9918 4312
rect 9310 3576 9366 3632
rect 9402 3304 9458 3360
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 9770 3984 9826 4040
rect 9770 3884 9772 3904
rect 9772 3884 9824 3904
rect 9824 3884 9826 3904
rect 9770 3848 9826 3884
rect 9862 3596 9918 3632
rect 9862 3576 9864 3596
rect 9864 3576 9916 3596
rect 9916 3576 9918 3596
rect 9218 2372 9274 2408
rect 9218 2352 9220 2372
rect 9220 2352 9272 2372
rect 9272 2352 9274 2372
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 9770 1400 9826 1456
rect 10046 5480 10102 5536
rect 10414 4800 10470 4856
rect 11058 9016 11114 9072
rect 10966 8064 11022 8120
rect 11058 6296 11114 6352
rect 11426 8200 11482 8256
rect 11058 5344 11114 5400
rect 10414 3848 10470 3904
rect 10230 1672 10286 1728
rect 11794 5888 11850 5944
rect 12530 10376 12586 10432
rect 12530 9968 12586 10024
rect 12070 7656 12126 7712
rect 11978 7112 12034 7168
rect 12162 7520 12218 7576
rect 12806 9968 12862 10024
rect 12990 10240 13046 10296
rect 12990 9696 13046 9752
rect 13174 9696 13230 9752
rect 12530 7384 12586 7440
rect 11978 1808 12034 1864
rect 13358 7928 13414 7984
rect 13634 8336 13690 8392
rect 14002 9968 14058 10024
rect 14278 9696 14334 9752
rect 13450 7384 13506 7440
rect 13358 7248 13414 7304
rect 13358 6840 13414 6896
rect 12990 5888 13046 5944
rect 13726 7656 13782 7712
rect 13726 7384 13782 7440
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 13726 7248 13782 7304
rect 14370 8064 14426 8120
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 15290 8236 15292 8256
rect 15292 8236 15344 8256
rect 15344 8236 15346 8256
rect 15290 8200 15346 8236
rect 15106 8064 15162 8120
rect 15198 7792 15254 7848
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 13818 6976 13874 7032
rect 14370 6976 14426 7032
rect 14462 6840 14518 6896
rect 14462 6024 14518 6080
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 14462 5888 14518 5944
rect 13726 4936 13782 4992
rect 13542 4800 13598 4856
rect 14278 5480 14334 5536
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 14462 4256 14518 4312
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 14646 6840 14702 6896
rect 14646 6296 14702 6352
rect 15658 7656 15714 7712
rect 14922 7112 14978 7168
rect 15474 6568 15530 6624
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 14370 3304 14426 3360
rect 14554 3168 14610 3224
rect 13726 3032 13782 3088
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 14554 2760 14610 2816
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 15290 5208 15346 5264
rect 15474 5208 15530 5264
rect 14922 4528 14978 4584
rect 15198 4548 15254 4584
rect 15198 4528 15200 4548
rect 15200 4528 15252 4548
rect 15252 4528 15254 4548
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 16394 9696 16450 9752
rect 16210 7248 16266 7304
rect 16394 7248 16450 7304
rect 15842 5888 15898 5944
rect 16302 5616 16358 5672
rect 16026 5344 16082 5400
rect 16026 4800 16082 4856
rect 16302 4800 16358 4856
rect 15842 4256 15898 4312
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 16026 3576 16082 3632
rect 16026 3304 16082 3360
rect 16026 2760 16082 2816
rect 15750 2488 15806 2544
rect 17038 9696 17094 9752
rect 17406 7384 17462 7440
rect 16946 5616 17002 5672
rect 17222 5208 17278 5264
rect 16762 3032 16818 3088
rect 16394 2488 16450 2544
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 16210 584 16266 640
rect 17222 4392 17278 4448
rect 17590 7792 17646 7848
rect 17590 7520 17646 7576
rect 17682 6976 17738 7032
rect 18878 9696 18934 9752
rect 18142 7520 18198 7576
rect 17866 5752 17922 5808
rect 18142 7112 18198 7168
rect 18050 6160 18106 6216
rect 18050 5752 18106 5808
rect 19154 9968 19210 10024
rect 19062 8064 19118 8120
rect 19798 9968 19854 10024
rect 19522 9696 19578 9752
rect 19614 9016 19670 9072
rect 19430 8744 19486 8800
rect 19338 8064 19394 8120
rect 19706 8200 19762 8256
rect 19706 8084 19762 8120
rect 19706 8064 19708 8084
rect 19708 8064 19760 8084
rect 19760 8064 19762 8084
rect 20074 8608 20130 8664
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 19982 7928 20038 7984
rect 18602 5480 18658 5536
rect 17682 3168 17738 3224
rect 18142 3304 18198 3360
rect 18326 3304 18382 3360
rect 18326 2760 18382 2816
rect 19246 5480 19302 5536
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 20534 7540 20590 7576
rect 20534 7520 20536 7540
rect 20536 7520 20588 7540
rect 20588 7520 20590 7540
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 20994 8064 21050 8120
rect 20994 7792 21050 7848
rect 21178 7792 21234 7848
rect 21546 7656 21602 7712
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 20994 6976 21050 7032
rect 19706 6432 19762 6488
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 19522 5480 19578 5536
rect 19430 5344 19486 5400
rect 19982 5092 20038 5128
rect 19982 5072 19984 5092
rect 19984 5072 20036 5092
rect 20036 5072 20038 5092
rect 20166 5072 20222 5128
rect 19798 4936 19854 4992
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 19522 4800 19578 4856
rect 19062 4256 19118 4312
rect 19430 4276 19486 4312
rect 19430 4256 19432 4276
rect 19432 4256 19484 4276
rect 19484 4256 19486 4276
rect 19430 4120 19486 4176
rect 16946 720 17002 776
rect 20074 4256 20130 4312
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 20626 6568 20682 6624
rect 20810 6840 20866 6896
rect 20626 6160 20682 6216
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 20902 5888 20958 5944
rect 20810 5480 20866 5536
rect 20442 4800 20498 4856
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 20442 4392 20498 4448
rect 20626 4256 20682 4312
rect 20442 3848 20498 3904
rect 20534 3712 20590 3768
rect 20534 3440 20590 3496
rect 20442 3168 20498 3224
rect 19522 1944 19578 2000
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 19522 1672 19578 1728
rect 19706 1672 19762 1728
rect 19430 856 19486 912
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 20718 1672 20774 1728
rect 21730 6568 21786 6624
rect 23386 10240 23442 10296
rect 23110 9968 23166 10024
rect 22834 9560 22890 9616
rect 22650 8608 22706 8664
rect 21914 3440 21970 3496
rect 21822 3168 21878 3224
rect 23294 8064 23350 8120
rect 22558 3984 22614 4040
rect 22742 3440 22798 3496
rect 22742 3168 22798 3224
rect 21822 992 21878 1048
rect 24122 9016 24178 9072
rect 24398 10376 24454 10432
rect 24306 9152 24362 9208
rect 24490 8200 24546 8256
rect 23662 4800 23718 4856
rect 24950 10512 25006 10568
rect 24766 9832 24822 9888
rect 24674 9560 24730 9616
rect 25134 9968 25190 10024
rect 25042 9560 25098 9616
rect 24674 6840 24730 6896
rect 24674 5752 24730 5808
rect 25410 10240 25466 10296
rect 25318 9152 25374 9208
rect 24858 5888 24914 5944
rect 24858 5752 24914 5808
rect 25134 7248 25190 7304
rect 25134 6024 25190 6080
rect 25410 6432 25466 6488
rect 24766 4936 24822 4992
rect 24858 3984 24914 4040
rect 24674 1944 24730 2000
rect 25502 4120 25558 4176
rect 26238 9832 26294 9888
rect 26330 9560 26386 9616
rect 26698 9560 26754 9616
rect 26790 9152 26846 9208
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 26882 8608 26938 8664
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 26330 7692 26332 7712
rect 26332 7692 26384 7712
rect 26384 7692 26386 7712
rect 26330 7656 26386 7692
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 25686 3848 25742 3904
rect 25962 6432 26018 6488
rect 27618 9560 27674 9616
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 26606 6568 26662 6624
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 27710 8064 27766 8120
rect 27526 7384 27582 7440
rect 27066 6296 27122 6352
rect 27342 6296 27398 6352
rect 26698 6160 26754 6216
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 26054 5108 26056 5128
rect 26056 5108 26108 5128
rect 26108 5108 26110 5128
rect 26054 5072 26110 5108
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 27066 5616 27122 5672
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27066 4664 27122 4720
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 25778 3712 25834 3768
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 27434 3576 27490 3632
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 28814 9560 28870 9616
rect 28538 5888 28594 5944
rect 27986 5072 28042 5128
rect 29090 6976 29146 7032
rect 29090 6432 29146 6488
rect 28998 5208 29054 5264
rect 29182 5208 29238 5264
rect 30286 9832 30342 9888
rect 29826 7520 29882 7576
rect 29458 3576 29514 3632
rect 30378 8744 30434 8800
rect 30378 8200 30434 8256
rect 30286 7656 30342 7712
rect 30654 8200 30710 8256
rect 30378 6704 30434 6760
rect 30930 9560 30986 9616
rect 31022 8064 31078 8120
rect 30930 7656 30986 7712
rect 30838 6840 30894 6896
rect 29918 6160 29974 6216
rect 30654 6024 30710 6080
rect 30194 5480 30250 5536
rect 30010 2896 30066 2952
rect 31758 9832 31814 9888
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 32586 9288 32642 9344
rect 32310 7928 32366 7984
rect 31390 7520 31446 7576
rect 31206 5480 31262 5536
rect 30562 4936 30618 4992
rect 30286 3304 30342 3360
rect 32126 7248 32182 7304
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 31850 6432 31906 6488
rect 31666 6296 31722 6352
rect 31666 6024 31722 6080
rect 31390 4664 31446 4720
rect 31022 4548 31078 4584
rect 31022 4528 31024 4548
rect 31024 4528 31076 4548
rect 31076 4528 31078 4548
rect 31114 4120 31170 4176
rect 30470 3712 30526 3768
rect 30378 2760 30434 2816
rect 30194 1808 30250 1864
rect 30286 1536 30342 1592
rect 30746 2760 30802 2816
rect 30654 1400 30710 1456
rect 31298 3032 31354 3088
rect 31482 4528 31538 4584
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 32678 6976 32734 7032
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 32954 7792 33010 7848
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 31942 4664 31998 4720
rect 31666 3732 31722 3768
rect 31666 3712 31668 3732
rect 31668 3712 31720 3732
rect 31720 3712 31722 3732
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 32034 3304 32090 3360
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 31390 2352 31446 2408
rect 33506 3576 33562 3632
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
rect 34334 7792 34390 7848
rect 33966 5616 34022 5672
rect 34794 8336 34850 8392
rect 35070 9152 35126 9208
rect 35438 8472 35494 8528
rect 35162 4120 35218 4176
rect 36266 4528 36322 4584
rect 36634 7828 36636 7848
rect 36636 7828 36688 7848
rect 36688 7828 36690 7848
rect 36634 7792 36690 7828
rect 37554 9696 37610 9752
rect 36910 5208 36966 5264
rect 37278 1264 37334 1320
rect 38474 10104 38530 10160
rect 38290 9832 38346 9888
rect 37956 8186 38012 8188
rect 38036 8186 38092 8188
rect 38116 8186 38172 8188
rect 38196 8186 38252 8188
rect 37956 8134 38002 8186
rect 38002 8134 38012 8186
rect 38036 8134 38066 8186
rect 38066 8134 38078 8186
rect 38078 8134 38092 8186
rect 38116 8134 38130 8186
rect 38130 8134 38142 8186
rect 38142 8134 38172 8186
rect 38196 8134 38206 8186
rect 38206 8134 38252 8186
rect 37956 8132 38012 8134
rect 38036 8132 38092 8134
rect 38116 8132 38172 8134
rect 38196 8132 38252 8134
rect 39670 9560 39726 9616
rect 38750 9288 38806 9344
rect 38658 8472 38714 8528
rect 37956 7098 38012 7100
rect 38036 7098 38092 7100
rect 38116 7098 38172 7100
rect 38196 7098 38252 7100
rect 37956 7046 38002 7098
rect 38002 7046 38012 7098
rect 38036 7046 38066 7098
rect 38066 7046 38078 7098
rect 38078 7046 38092 7098
rect 38116 7046 38130 7098
rect 38130 7046 38142 7098
rect 38142 7046 38172 7098
rect 38196 7046 38206 7098
rect 38206 7046 38252 7098
rect 37956 7044 38012 7046
rect 38036 7044 38092 7046
rect 38116 7044 38172 7046
rect 38196 7044 38252 7046
rect 37646 6160 37702 6216
rect 37956 6010 38012 6012
rect 38036 6010 38092 6012
rect 38116 6010 38172 6012
rect 38196 6010 38252 6012
rect 37956 5958 38002 6010
rect 38002 5958 38012 6010
rect 38036 5958 38066 6010
rect 38066 5958 38078 6010
rect 38078 5958 38092 6010
rect 38116 5958 38130 6010
rect 38130 5958 38142 6010
rect 38142 5958 38172 6010
rect 38196 5958 38206 6010
rect 38206 5958 38252 6010
rect 37956 5956 38012 5958
rect 38036 5956 38092 5958
rect 38116 5956 38172 5958
rect 38196 5956 38252 5958
rect 37830 5072 37886 5128
rect 37956 4922 38012 4924
rect 38036 4922 38092 4924
rect 38116 4922 38172 4924
rect 38196 4922 38252 4924
rect 37956 4870 38002 4922
rect 38002 4870 38012 4922
rect 38036 4870 38066 4922
rect 38066 4870 38078 4922
rect 38078 4870 38092 4922
rect 38116 4870 38130 4922
rect 38130 4870 38142 4922
rect 38142 4870 38172 4922
rect 38196 4870 38206 4922
rect 38206 4870 38252 4922
rect 37956 4868 38012 4870
rect 38036 4868 38092 4870
rect 38116 4868 38172 4870
rect 38196 4868 38252 4870
rect 37554 3984 37610 4040
rect 37956 3834 38012 3836
rect 38036 3834 38092 3836
rect 38116 3834 38172 3836
rect 38196 3834 38252 3836
rect 37956 3782 38002 3834
rect 38002 3782 38012 3834
rect 38036 3782 38066 3834
rect 38066 3782 38078 3834
rect 38078 3782 38092 3834
rect 38116 3782 38130 3834
rect 38130 3782 38142 3834
rect 38142 3782 38172 3834
rect 38196 3782 38206 3834
rect 38206 3782 38252 3834
rect 37956 3780 38012 3782
rect 38036 3780 38092 3782
rect 38116 3780 38172 3782
rect 38196 3780 38252 3782
rect 37956 2746 38012 2748
rect 38036 2746 38092 2748
rect 38116 2746 38172 2748
rect 38196 2746 38252 2748
rect 37956 2694 38002 2746
rect 38002 2694 38012 2746
rect 38036 2694 38066 2746
rect 38066 2694 38078 2746
rect 38078 2694 38092 2746
rect 38116 2694 38130 2746
rect 38130 2694 38142 2746
rect 38142 2694 38172 2746
rect 38196 2694 38206 2746
rect 38206 2694 38252 2746
rect 37956 2692 38012 2694
rect 38036 2692 38092 2694
rect 38116 2692 38172 2694
rect 38196 2692 38252 2694
rect 39578 8744 39634 8800
rect 39016 8730 39072 8732
rect 39096 8730 39152 8732
rect 39176 8730 39232 8732
rect 39256 8730 39312 8732
rect 39016 8678 39062 8730
rect 39062 8678 39072 8730
rect 39096 8678 39126 8730
rect 39126 8678 39138 8730
rect 39138 8678 39152 8730
rect 39176 8678 39190 8730
rect 39190 8678 39202 8730
rect 39202 8678 39232 8730
rect 39256 8678 39266 8730
rect 39266 8678 39312 8730
rect 39016 8676 39072 8678
rect 39096 8676 39152 8678
rect 39176 8676 39232 8678
rect 39256 8676 39312 8678
rect 39486 8200 39542 8256
rect 39394 7928 39450 7984
rect 39394 7692 39396 7712
rect 39396 7692 39448 7712
rect 39448 7692 39450 7712
rect 39394 7656 39450 7692
rect 39016 7642 39072 7644
rect 39096 7642 39152 7644
rect 39176 7642 39232 7644
rect 39256 7642 39312 7644
rect 39016 7590 39062 7642
rect 39062 7590 39072 7642
rect 39096 7590 39126 7642
rect 39126 7590 39138 7642
rect 39138 7590 39152 7642
rect 39176 7590 39190 7642
rect 39190 7590 39202 7642
rect 39202 7590 39232 7642
rect 39256 7590 39266 7642
rect 39266 7590 39312 7642
rect 39016 7588 39072 7590
rect 39096 7588 39152 7590
rect 39176 7588 39232 7590
rect 39256 7588 39312 7590
rect 38934 7384 38990 7440
rect 39394 7112 39450 7168
rect 38658 6296 38714 6352
rect 39854 9016 39910 9072
rect 39670 6568 39726 6624
rect 39016 6554 39072 6556
rect 39096 6554 39152 6556
rect 39176 6554 39232 6556
rect 39256 6554 39312 6556
rect 39016 6502 39062 6554
rect 39062 6502 39072 6554
rect 39096 6502 39126 6554
rect 39126 6502 39138 6554
rect 39138 6502 39152 6554
rect 39176 6502 39190 6554
rect 39190 6502 39202 6554
rect 39202 6502 39232 6554
rect 39256 6502 39266 6554
rect 39266 6502 39312 6554
rect 39016 6500 39072 6502
rect 39096 6500 39152 6502
rect 39176 6500 39232 6502
rect 39256 6500 39312 6502
rect 39026 6060 39028 6080
rect 39028 6060 39080 6080
rect 39080 6060 39082 6080
rect 39026 6024 39082 6060
rect 38842 5752 38898 5808
rect 39394 5752 39450 5808
rect 39016 5466 39072 5468
rect 39096 5466 39152 5468
rect 39176 5466 39232 5468
rect 39256 5466 39312 5468
rect 39016 5414 39062 5466
rect 39062 5414 39072 5466
rect 39096 5414 39126 5466
rect 39126 5414 39138 5466
rect 39138 5414 39152 5466
rect 39176 5414 39190 5466
rect 39190 5414 39202 5466
rect 39202 5414 39232 5466
rect 39256 5414 39266 5466
rect 39266 5414 39312 5466
rect 39016 5412 39072 5414
rect 39096 5412 39152 5414
rect 39176 5412 39232 5414
rect 39256 5412 39312 5414
rect 39394 5208 39450 5264
rect 38382 2896 38438 2952
rect 37922 1944 37978 2000
rect 39026 4972 39028 4992
rect 39028 4972 39080 4992
rect 39080 4972 39082 4992
rect 39026 4936 39082 4972
rect 39486 4664 39542 4720
rect 39016 4378 39072 4380
rect 39096 4378 39152 4380
rect 39176 4378 39232 4380
rect 39256 4378 39312 4380
rect 39016 4326 39062 4378
rect 39062 4326 39072 4378
rect 39096 4326 39126 4378
rect 39126 4326 39138 4378
rect 39138 4326 39152 4378
rect 39176 4326 39190 4378
rect 39190 4326 39202 4378
rect 39202 4326 39232 4378
rect 39256 4326 39266 4378
rect 39266 4326 39312 4378
rect 39016 4324 39072 4326
rect 39096 4324 39152 4326
rect 39176 4324 39232 4326
rect 39256 4324 39312 4326
rect 39394 4120 39450 4176
rect 39026 3884 39028 3904
rect 39028 3884 39080 3904
rect 39080 3884 39082 3904
rect 39026 3848 39082 3884
rect 39394 3576 39450 3632
rect 38842 3476 38844 3496
rect 38844 3476 38896 3496
rect 38896 3476 38898 3496
rect 38842 3440 38898 3476
rect 39016 3290 39072 3292
rect 39096 3290 39152 3292
rect 39176 3290 39232 3292
rect 39256 3290 39312 3292
rect 39016 3238 39062 3290
rect 39062 3238 39072 3290
rect 39096 3238 39126 3290
rect 39126 3238 39138 3290
rect 39138 3238 39152 3290
rect 39176 3238 39190 3290
rect 39190 3238 39202 3290
rect 39202 3238 39232 3290
rect 39256 3238 39266 3290
rect 39266 3238 39312 3290
rect 39016 3236 39072 3238
rect 39096 3236 39152 3238
rect 39176 3236 39232 3238
rect 39256 3236 39312 3238
rect 39394 3032 39450 3088
rect 38474 2488 38530 2544
rect 38658 2488 38714 2544
rect 38290 1672 38346 1728
rect 38658 1400 38714 1456
rect 39026 2796 39028 2816
rect 39028 2796 39080 2816
rect 39080 2796 39082 2816
rect 39026 2760 39082 2796
rect 39016 2202 39072 2204
rect 39096 2202 39152 2204
rect 39176 2202 39232 2204
rect 39256 2202 39312 2204
rect 39016 2150 39062 2202
rect 39062 2150 39072 2202
rect 39096 2150 39126 2202
rect 39126 2150 39138 2202
rect 39138 2150 39152 2202
rect 39176 2150 39190 2202
rect 39190 2150 39202 2202
rect 39202 2150 39232 2202
rect 39256 2150 39266 2202
rect 39266 2150 39312 2202
rect 39016 2148 39072 2150
rect 39096 2148 39152 2150
rect 39176 2148 39232 2150
rect 39256 2148 39312 2150
rect 38934 1128 38990 1184
rect 40038 6840 40094 6896
rect 39946 5480 40002 5536
rect 39946 4392 40002 4448
rect 39946 3304 40002 3360
rect 39946 2216 40002 2272
<< metal3 >>
rect 24945 10570 25011 10573
rect 22050 10568 25011 10570
rect 22050 10512 24950 10568
rect 25006 10512 25011 10568
rect 22050 10510 25011 10512
rect 12525 10434 12591 10437
rect 22050 10434 22110 10510
rect 24945 10507 25011 10510
rect 24393 10434 24459 10437
rect 12525 10432 22110 10434
rect 12525 10376 12530 10432
rect 12586 10376 22110 10432
rect 12525 10374 22110 10376
rect 23246 10432 24459 10434
rect 23246 10376 24398 10432
rect 24454 10376 24459 10432
rect 23246 10374 24459 10376
rect 12525 10371 12591 10374
rect 12985 10298 13051 10301
rect 23246 10298 23306 10374
rect 24393 10371 24459 10374
rect 12985 10296 23306 10298
rect 12985 10240 12990 10296
rect 13046 10240 23306 10296
rect 12985 10238 23306 10240
rect 23381 10298 23447 10301
rect 25405 10298 25471 10301
rect 23381 10296 25471 10298
rect 23381 10240 23386 10296
rect 23442 10240 25410 10296
rect 25466 10240 25471 10296
rect 23381 10238 25471 10240
rect 12985 10235 13051 10238
rect 23381 10235 23447 10238
rect 25405 10235 25471 10238
rect 2313 10162 2379 10165
rect 38469 10162 38535 10165
rect 2313 10160 38535 10162
rect 2313 10104 2318 10160
rect 2374 10104 38474 10160
rect 38530 10104 38535 10160
rect 2313 10102 38535 10104
rect 2313 10099 2379 10102
rect 38469 10099 38535 10102
rect 3969 10026 4035 10029
rect 12525 10026 12591 10029
rect 3969 10024 12591 10026
rect 3969 9968 3974 10024
rect 4030 9968 12530 10024
rect 12586 9968 12591 10024
rect 3969 9966 12591 9968
rect 3969 9963 4035 9966
rect 12525 9963 12591 9966
rect 12801 10026 12867 10029
rect 13997 10026 14063 10029
rect 12801 10024 14063 10026
rect 12801 9968 12806 10024
rect 12862 9968 14002 10024
rect 14058 9968 14063 10024
rect 12801 9966 14063 9968
rect 12801 9963 12867 9966
rect 13997 9963 14063 9966
rect 19149 10026 19215 10029
rect 19793 10026 19859 10029
rect 19149 10024 19859 10026
rect 19149 9968 19154 10024
rect 19210 9968 19798 10024
rect 19854 9968 19859 10024
rect 19149 9966 19859 9968
rect 19149 9963 19215 9966
rect 19793 9963 19859 9966
rect 23105 10026 23171 10029
rect 25129 10026 25195 10029
rect 23105 10024 25195 10026
rect 23105 9968 23110 10024
rect 23166 9968 25134 10024
rect 25190 9968 25195 10024
rect 23105 9966 25195 9968
rect 23105 9963 23171 9966
rect 25129 9963 25195 9966
rect 0 9890 120 9920
rect 473 9890 539 9893
rect 0 9888 539 9890
rect 0 9832 478 9888
rect 534 9832 539 9888
rect 0 9830 539 9832
rect 0 9800 120 9830
rect 473 9827 539 9830
rect 6637 9890 6703 9893
rect 8477 9890 8543 9893
rect 24761 9890 24827 9893
rect 26233 9890 26299 9893
rect 6637 9888 8543 9890
rect 6637 9832 6642 9888
rect 6698 9832 8482 9888
rect 8538 9832 8543 9888
rect 6637 9830 8543 9832
rect 6637 9827 6703 9830
rect 8477 9827 8543 9830
rect 8710 9830 22110 9890
rect 4429 9754 4495 9757
rect 6729 9754 6795 9757
rect 7373 9754 7439 9757
rect 8710 9754 8770 9830
rect 12985 9754 13051 9757
rect 4429 9752 6608 9754
rect 4429 9696 4434 9752
rect 4490 9696 6608 9752
rect 4429 9694 6608 9696
rect 4429 9691 4495 9694
rect 0 9618 120 9648
rect 657 9618 723 9621
rect 0 9616 723 9618
rect 0 9560 662 9616
rect 718 9560 723 9616
rect 0 9558 723 9560
rect 6548 9618 6608 9694
rect 6729 9752 7439 9754
rect 6729 9696 6734 9752
rect 6790 9696 7378 9752
rect 7434 9696 7439 9752
rect 6729 9694 7439 9696
rect 6729 9691 6795 9694
rect 7373 9691 7439 9694
rect 7606 9694 8770 9754
rect 8894 9752 13051 9754
rect 8894 9696 12990 9752
rect 13046 9696 13051 9752
rect 8894 9694 13051 9696
rect 7606 9618 7666 9694
rect 6548 9558 7666 9618
rect 8293 9618 8359 9621
rect 8894 9618 8954 9694
rect 12985 9691 13051 9694
rect 13169 9754 13235 9757
rect 14273 9754 14339 9757
rect 13169 9752 14339 9754
rect 13169 9696 13174 9752
rect 13230 9696 14278 9752
rect 14334 9696 14339 9752
rect 13169 9694 14339 9696
rect 13169 9691 13235 9694
rect 14273 9691 14339 9694
rect 16389 9754 16455 9757
rect 17033 9754 17099 9757
rect 16389 9752 17099 9754
rect 16389 9696 16394 9752
rect 16450 9696 17038 9752
rect 17094 9696 17099 9752
rect 16389 9694 17099 9696
rect 16389 9691 16455 9694
rect 17033 9691 17099 9694
rect 18873 9754 18939 9757
rect 19517 9754 19583 9757
rect 18873 9752 19583 9754
rect 18873 9696 18878 9752
rect 18934 9696 19522 9752
rect 19578 9696 19583 9752
rect 18873 9694 19583 9696
rect 22050 9754 22110 9830
rect 24761 9888 26299 9890
rect 24761 9832 24766 9888
rect 24822 9832 26238 9888
rect 26294 9832 26299 9888
rect 24761 9830 26299 9832
rect 24761 9827 24827 9830
rect 26233 9827 26299 9830
rect 30281 9890 30347 9893
rect 31753 9890 31819 9893
rect 30281 9888 31819 9890
rect 30281 9832 30286 9888
rect 30342 9832 31758 9888
rect 31814 9832 31819 9888
rect 30281 9830 31819 9832
rect 30281 9827 30347 9830
rect 31753 9827 31819 9830
rect 38285 9890 38351 9893
rect 40880 9890 41000 9920
rect 38285 9888 41000 9890
rect 38285 9832 38290 9888
rect 38346 9832 41000 9888
rect 38285 9830 41000 9832
rect 38285 9827 38351 9830
rect 40880 9800 41000 9830
rect 37549 9754 37615 9757
rect 22050 9752 37615 9754
rect 22050 9696 37554 9752
rect 37610 9696 37615 9752
rect 22050 9694 37615 9696
rect 18873 9691 18939 9694
rect 19517 9691 19583 9694
rect 37549 9691 37615 9694
rect 8293 9616 8954 9618
rect 8293 9560 8298 9616
rect 8354 9560 8954 9616
rect 8293 9558 8954 9560
rect 22829 9618 22895 9621
rect 24669 9618 24735 9621
rect 22829 9616 24735 9618
rect 22829 9560 22834 9616
rect 22890 9560 24674 9616
rect 24730 9560 24735 9616
rect 22829 9558 24735 9560
rect 0 9528 120 9558
rect 657 9555 723 9558
rect 8293 9555 8359 9558
rect 22829 9555 22895 9558
rect 24669 9555 24735 9558
rect 25037 9618 25103 9621
rect 26325 9618 26391 9621
rect 25037 9616 26391 9618
rect 25037 9560 25042 9616
rect 25098 9560 26330 9616
rect 26386 9560 26391 9616
rect 25037 9558 26391 9560
rect 25037 9555 25103 9558
rect 26325 9555 26391 9558
rect 26693 9618 26759 9621
rect 27613 9618 27679 9621
rect 26693 9616 27679 9618
rect 26693 9560 26698 9616
rect 26754 9560 27618 9616
rect 27674 9560 27679 9616
rect 26693 9558 27679 9560
rect 26693 9555 26759 9558
rect 27613 9555 27679 9558
rect 28809 9618 28875 9621
rect 30925 9618 30991 9621
rect 28809 9616 30991 9618
rect 28809 9560 28814 9616
rect 28870 9560 30930 9616
rect 30986 9560 30991 9616
rect 28809 9558 30991 9560
rect 28809 9555 28875 9558
rect 30925 9555 30991 9558
rect 39665 9618 39731 9621
rect 40880 9618 41000 9648
rect 39665 9616 41000 9618
rect 39665 9560 39670 9616
rect 39726 9560 41000 9616
rect 39665 9558 41000 9560
rect 39665 9555 39731 9558
rect 40880 9528 41000 9558
rect 6177 9482 6243 9485
rect 6177 9480 31770 9482
rect 6177 9424 6182 9480
rect 6238 9424 31770 9480
rect 6177 9422 31770 9424
rect 6177 9419 6243 9422
rect 0 9346 120 9376
rect 1209 9346 1275 9349
rect 0 9344 1275 9346
rect 0 9288 1214 9344
rect 1270 9288 1275 9344
rect 0 9286 1275 9288
rect 0 9256 120 9286
rect 1209 9283 1275 9286
rect 9489 9346 9555 9349
rect 31710 9346 31770 9422
rect 32581 9346 32647 9349
rect 9489 9344 26986 9346
rect 9489 9288 9494 9344
rect 9550 9288 26986 9344
rect 9489 9286 26986 9288
rect 31710 9344 32647 9346
rect 31710 9288 32586 9344
rect 32642 9288 32647 9344
rect 31710 9286 32647 9288
rect 9489 9283 9555 9286
rect 5073 9210 5139 9213
rect 24301 9210 24367 9213
rect 5073 9208 24367 9210
rect 5073 9152 5078 9208
rect 5134 9152 24306 9208
rect 24362 9152 24367 9208
rect 5073 9150 24367 9152
rect 5073 9147 5139 9150
rect 24301 9147 24367 9150
rect 25313 9210 25379 9213
rect 26785 9210 26851 9213
rect 25313 9208 26851 9210
rect 25313 9152 25318 9208
rect 25374 9152 26790 9208
rect 26846 9152 26851 9208
rect 25313 9150 26851 9152
rect 26926 9210 26986 9286
rect 32581 9283 32647 9286
rect 38745 9346 38811 9349
rect 40880 9346 41000 9376
rect 38745 9344 41000 9346
rect 38745 9288 38750 9344
rect 38806 9288 41000 9344
rect 38745 9286 41000 9288
rect 38745 9283 38811 9286
rect 40880 9256 41000 9286
rect 35065 9210 35131 9213
rect 26926 9208 35131 9210
rect 26926 9152 35070 9208
rect 35126 9152 35131 9208
rect 26926 9150 35131 9152
rect 25313 9147 25379 9150
rect 26785 9147 26851 9150
rect 35065 9147 35131 9150
rect 0 9074 120 9104
rect 2773 9074 2839 9077
rect 0 9072 2839 9074
rect 0 9016 2778 9072
rect 2834 9016 2839 9072
rect 0 9014 2839 9016
rect 0 8984 120 9014
rect 2773 9011 2839 9014
rect 9673 9074 9739 9077
rect 11053 9074 11119 9077
rect 9673 9072 11119 9074
rect 9673 9016 9678 9072
rect 9734 9016 11058 9072
rect 11114 9016 11119 9072
rect 9673 9014 11119 9016
rect 9673 9011 9739 9014
rect 11053 9011 11119 9014
rect 19609 9074 19675 9077
rect 24117 9074 24183 9077
rect 19609 9072 24183 9074
rect 19609 9016 19614 9072
rect 19670 9016 24122 9072
rect 24178 9016 24183 9072
rect 19609 9014 24183 9016
rect 19609 9011 19675 9014
rect 24117 9011 24183 9014
rect 39849 9074 39915 9077
rect 40880 9074 41000 9104
rect 39849 9072 41000 9074
rect 39849 9016 39854 9072
rect 39910 9016 41000 9072
rect 39849 9014 41000 9016
rect 39849 9011 39915 9014
rect 40880 8984 41000 9014
rect 7373 8938 7439 8941
rect 7373 8936 30298 8938
rect 7373 8880 7378 8936
rect 7434 8880 30298 8936
rect 7373 8878 30298 8880
rect 7373 8875 7439 8878
rect 0 8802 120 8832
rect 2865 8802 2931 8805
rect 0 8800 2931 8802
rect 0 8744 2870 8800
rect 2926 8744 2931 8800
rect 0 8742 2931 8744
rect 0 8712 120 8742
rect 2865 8739 2931 8742
rect 9857 8802 9923 8805
rect 9990 8802 9996 8804
rect 9857 8800 9996 8802
rect 9857 8744 9862 8800
rect 9918 8744 9996 8800
rect 9857 8742 9996 8744
rect 9857 8739 9923 8742
rect 9990 8740 9996 8742
rect 10060 8740 10066 8804
rect 19425 8802 19491 8805
rect 20662 8802 20668 8804
rect 19425 8800 20668 8802
rect 19425 8744 19430 8800
rect 19486 8744 20668 8800
rect 19425 8742 20668 8744
rect 19425 8739 19491 8742
rect 20662 8740 20668 8742
rect 20732 8740 20738 8804
rect 30238 8802 30298 8878
rect 30373 8802 30439 8805
rect 30238 8800 30439 8802
rect 30238 8744 30378 8800
rect 30434 8744 30439 8800
rect 30238 8742 30439 8744
rect 30373 8739 30439 8742
rect 39573 8802 39639 8805
rect 40880 8802 41000 8832
rect 39573 8800 41000 8802
rect 39573 8744 39578 8800
rect 39634 8744 41000 8800
rect 39573 8742 41000 8744
rect 39573 8739 39639 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 33006 8671 33322 8672
rect 39006 8736 39322 8737
rect 39006 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39322 8736
rect 40880 8712 41000 8742
rect 39006 8671 39322 8672
rect 19742 8604 19748 8668
rect 19812 8666 19818 8668
rect 20069 8666 20135 8669
rect 19812 8664 20135 8666
rect 19812 8608 20074 8664
rect 20130 8608 20135 8664
rect 19812 8606 20135 8608
rect 19812 8604 19818 8606
rect 20069 8603 20135 8606
rect 22645 8666 22711 8669
rect 26877 8666 26943 8669
rect 22645 8664 26943 8666
rect 22645 8608 22650 8664
rect 22706 8608 26882 8664
rect 26938 8608 26943 8664
rect 22645 8606 26943 8608
rect 22645 8603 22711 8606
rect 26877 8603 26943 8606
rect 0 8530 120 8560
rect 1301 8530 1367 8533
rect 0 8528 1367 8530
rect 0 8472 1306 8528
rect 1362 8472 1367 8528
rect 0 8470 1367 8472
rect 0 8440 120 8470
rect 1301 8467 1367 8470
rect 6637 8530 6703 8533
rect 35433 8530 35499 8533
rect 6637 8528 35499 8530
rect 6637 8472 6642 8528
rect 6698 8472 35438 8528
rect 35494 8472 35499 8528
rect 6637 8470 35499 8472
rect 6637 8467 6703 8470
rect 35433 8467 35499 8470
rect 38653 8530 38719 8533
rect 40880 8530 41000 8560
rect 38653 8528 41000 8530
rect 38653 8472 38658 8528
rect 38714 8472 41000 8528
rect 38653 8470 41000 8472
rect 38653 8467 38719 8470
rect 40880 8440 41000 8470
rect 4889 8394 4955 8397
rect 9029 8394 9095 8397
rect 4889 8392 9095 8394
rect 4889 8336 4894 8392
rect 4950 8336 9034 8392
rect 9090 8336 9095 8392
rect 4889 8334 9095 8336
rect 4889 8331 4955 8334
rect 9029 8331 9095 8334
rect 13629 8394 13695 8397
rect 34789 8394 34855 8397
rect 13629 8392 34855 8394
rect 13629 8336 13634 8392
rect 13690 8336 34794 8392
rect 34850 8336 34855 8392
rect 13629 8334 34855 8336
rect 13629 8331 13695 8334
rect 34789 8331 34855 8334
rect 0 8258 120 8288
rect 381 8258 447 8261
rect 11421 8258 11487 8261
rect 0 8256 447 8258
rect 0 8200 386 8256
rect 442 8200 447 8256
rect 0 8198 447 8200
rect 0 8168 120 8198
rect 381 8195 447 8198
rect 9768 8256 11487 8258
rect 9768 8200 11426 8256
rect 11482 8200 11487 8256
rect 9768 8198 11487 8200
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 9768 8125 9828 8198
rect 11421 8195 11487 8198
rect 15285 8258 15351 8261
rect 19701 8258 19767 8261
rect 15285 8256 19767 8258
rect 15285 8200 15290 8256
rect 15346 8200 19706 8256
rect 19762 8200 19767 8256
rect 15285 8198 19767 8200
rect 15285 8195 15351 8198
rect 19701 8195 19767 8198
rect 20478 8196 20484 8260
rect 20548 8258 20554 8260
rect 24485 8258 24551 8261
rect 20548 8256 24551 8258
rect 20548 8200 24490 8256
rect 24546 8200 24551 8256
rect 20548 8198 24551 8200
rect 20548 8196 20554 8198
rect 24485 8195 24551 8198
rect 30373 8258 30439 8261
rect 30649 8258 30715 8261
rect 30373 8256 30715 8258
rect 30373 8200 30378 8256
rect 30434 8200 30654 8256
rect 30710 8200 30715 8256
rect 30373 8198 30715 8200
rect 30373 8195 30439 8198
rect 30649 8195 30715 8198
rect 39481 8258 39547 8261
rect 40880 8258 41000 8288
rect 39481 8256 41000 8258
rect 39481 8200 39486 8256
rect 39542 8200 41000 8256
rect 39481 8198 41000 8200
rect 39481 8195 39547 8198
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 37946 8192 38262 8193
rect 37946 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38262 8192
rect 40880 8168 41000 8198
rect 37946 8127 38262 8128
rect 9765 8120 9831 8125
rect 9765 8064 9770 8120
rect 9826 8064 9831 8120
rect 9765 8059 9831 8064
rect 9949 8122 10015 8125
rect 10961 8122 11027 8125
rect 9949 8120 11027 8122
rect 9949 8064 9954 8120
rect 10010 8064 10966 8120
rect 11022 8064 11027 8120
rect 9949 8062 11027 8064
rect 9949 8059 10015 8062
rect 10961 8059 11027 8062
rect 14365 8122 14431 8125
rect 15101 8122 15167 8125
rect 19057 8122 19123 8125
rect 14365 8120 19123 8122
rect 14365 8064 14370 8120
rect 14426 8064 15106 8120
rect 15162 8064 19062 8120
rect 19118 8064 19123 8120
rect 14365 8062 19123 8064
rect 14365 8059 14431 8062
rect 15101 8059 15167 8062
rect 19057 8059 19123 8062
rect 19333 8122 19399 8125
rect 19558 8122 19564 8124
rect 19333 8120 19564 8122
rect 19333 8064 19338 8120
rect 19394 8064 19564 8120
rect 19333 8062 19564 8064
rect 19333 8059 19399 8062
rect 19558 8060 19564 8062
rect 19628 8060 19634 8124
rect 19701 8120 19767 8125
rect 19701 8064 19706 8120
rect 19762 8064 19767 8120
rect 19701 8059 19767 8064
rect 20989 8122 21055 8125
rect 23289 8122 23355 8125
rect 20989 8120 23355 8122
rect 20989 8064 20994 8120
rect 21050 8064 23294 8120
rect 23350 8064 23355 8120
rect 20989 8062 23355 8064
rect 20989 8059 21055 8062
rect 23289 8059 23355 8062
rect 27705 8122 27771 8125
rect 31017 8122 31083 8125
rect 27705 8120 31083 8122
rect 27705 8064 27710 8120
rect 27766 8064 31022 8120
rect 31078 8064 31083 8120
rect 27705 8062 31083 8064
rect 27705 8059 27771 8062
rect 31017 8059 31083 8062
rect 0 7986 120 8016
rect 749 7986 815 7989
rect 0 7984 815 7986
rect 0 7928 754 7984
rect 810 7928 815 7984
rect 0 7926 815 7928
rect 0 7896 120 7926
rect 749 7923 815 7926
rect 6821 7986 6887 7989
rect 13353 7986 13419 7989
rect 19704 7986 19764 8059
rect 6821 7984 13419 7986
rect 6821 7928 6826 7984
rect 6882 7928 13358 7984
rect 13414 7928 13419 7984
rect 6821 7926 13419 7928
rect 6821 7923 6887 7926
rect 13353 7923 13419 7926
rect 13678 7926 19764 7986
rect 19977 7986 20043 7989
rect 32305 7986 32371 7989
rect 19977 7984 32371 7986
rect 19977 7928 19982 7984
rect 20038 7928 32310 7984
rect 32366 7928 32371 7984
rect 19977 7926 32371 7928
rect 5533 7850 5599 7853
rect 13678 7850 13738 7926
rect 19977 7923 20043 7926
rect 32305 7923 32371 7926
rect 39389 7986 39455 7989
rect 40880 7986 41000 8016
rect 39389 7984 41000 7986
rect 39389 7928 39394 7984
rect 39450 7928 41000 7984
rect 39389 7926 41000 7928
rect 39389 7923 39455 7926
rect 40880 7896 41000 7926
rect 15193 7850 15259 7853
rect 5533 7848 13738 7850
rect 5533 7792 5538 7848
rect 5594 7792 13738 7848
rect 5533 7790 13738 7792
rect 13862 7848 15259 7850
rect 13862 7792 15198 7848
rect 15254 7792 15259 7848
rect 13862 7790 15259 7792
rect 5533 7787 5599 7790
rect 0 7714 120 7744
rect 749 7714 815 7717
rect 0 7712 815 7714
rect 0 7656 754 7712
rect 810 7656 815 7712
rect 0 7654 815 7656
rect 0 7624 120 7654
rect 749 7651 815 7654
rect 9949 7712 10015 7717
rect 9949 7656 9954 7712
rect 10010 7656 10015 7712
rect 9949 7651 10015 7656
rect 12065 7714 12131 7717
rect 13721 7714 13787 7717
rect 12065 7712 13787 7714
rect 12065 7656 12070 7712
rect 12126 7656 13726 7712
rect 13782 7656 13787 7712
rect 12065 7654 13787 7656
rect 12065 7651 12131 7654
rect 13721 7651 13787 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 4797 7578 4863 7581
rect 8702 7578 8708 7580
rect 4797 7576 8708 7578
rect 4797 7520 4802 7576
rect 4858 7520 8708 7576
rect 4797 7518 8708 7520
rect 4797 7515 4863 7518
rect 8702 7516 8708 7518
rect 8772 7516 8778 7580
rect 9952 7578 10012 7651
rect 12157 7578 12223 7581
rect 13862 7578 13922 7790
rect 15193 7787 15259 7790
rect 17585 7850 17651 7853
rect 20989 7850 21055 7853
rect 17585 7848 21055 7850
rect 17585 7792 17590 7848
rect 17646 7792 20994 7848
rect 21050 7792 21055 7848
rect 17585 7790 21055 7792
rect 17585 7787 17651 7790
rect 20989 7787 21055 7790
rect 21173 7850 21239 7853
rect 32949 7850 33015 7853
rect 21173 7848 33015 7850
rect 21173 7792 21178 7848
rect 21234 7792 32954 7848
rect 33010 7792 33015 7848
rect 21173 7790 33015 7792
rect 21173 7787 21239 7790
rect 32949 7787 33015 7790
rect 34329 7850 34395 7853
rect 36629 7850 36695 7853
rect 34329 7848 36695 7850
rect 34329 7792 34334 7848
rect 34390 7792 36634 7848
rect 36690 7792 36695 7848
rect 34329 7790 36695 7792
rect 34329 7787 34395 7790
rect 36629 7787 36695 7790
rect 15653 7714 15719 7717
rect 20478 7714 20484 7716
rect 15653 7712 20484 7714
rect 15653 7656 15658 7712
rect 15714 7656 20484 7712
rect 15653 7654 20484 7656
rect 15653 7651 15719 7654
rect 20478 7652 20484 7654
rect 20548 7652 20554 7716
rect 21541 7714 21607 7717
rect 26325 7714 26391 7717
rect 21541 7712 26391 7714
rect 21541 7656 21546 7712
rect 21602 7656 26330 7712
rect 26386 7656 26391 7712
rect 21541 7654 26391 7656
rect 21541 7651 21607 7654
rect 26325 7651 26391 7654
rect 30281 7714 30347 7717
rect 30925 7714 30991 7717
rect 30281 7712 30991 7714
rect 30281 7656 30286 7712
rect 30342 7656 30930 7712
rect 30986 7656 30991 7712
rect 30281 7654 30991 7656
rect 30281 7651 30347 7654
rect 30925 7651 30991 7654
rect 39389 7714 39455 7717
rect 40880 7714 41000 7744
rect 39389 7712 41000 7714
rect 39389 7656 39394 7712
rect 39450 7656 41000 7712
rect 39389 7654 41000 7656
rect 39389 7651 39455 7654
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 33006 7583 33322 7584
rect 39006 7648 39322 7649
rect 39006 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39322 7648
rect 40880 7624 41000 7654
rect 39006 7583 39322 7584
rect 17585 7578 17651 7581
rect 9952 7576 12223 7578
rect 9952 7520 12162 7576
rect 12218 7520 12223 7576
rect 9952 7518 12223 7520
rect 12157 7515 12223 7518
rect 12390 7518 13922 7578
rect 16254 7576 17651 7578
rect 16254 7520 17590 7576
rect 17646 7520 17651 7576
rect 16254 7518 17651 7520
rect 0 7442 120 7472
rect 933 7442 999 7445
rect 0 7440 999 7442
rect 0 7384 938 7440
rect 994 7384 999 7440
rect 0 7382 999 7384
rect 0 7352 120 7382
rect 933 7379 999 7382
rect 3601 7442 3667 7445
rect 12390 7442 12450 7518
rect 3601 7440 12450 7442
rect 3601 7384 3606 7440
rect 3662 7384 12450 7440
rect 3601 7382 12450 7384
rect 12525 7442 12591 7445
rect 13445 7442 13511 7445
rect 12525 7440 13511 7442
rect 12525 7384 12530 7440
rect 12586 7384 13450 7440
rect 13506 7384 13511 7440
rect 12525 7382 13511 7384
rect 3601 7379 3667 7382
rect 12525 7379 12591 7382
rect 13445 7379 13511 7382
rect 13721 7442 13787 7445
rect 16254 7442 16314 7518
rect 17585 7515 17651 7518
rect 18137 7578 18203 7581
rect 20529 7578 20595 7581
rect 18137 7576 20595 7578
rect 18137 7520 18142 7576
rect 18198 7520 20534 7576
rect 20590 7520 20595 7576
rect 18137 7518 20595 7520
rect 18137 7515 18203 7518
rect 20529 7515 20595 7518
rect 29821 7578 29887 7581
rect 31385 7578 31451 7581
rect 29821 7576 31451 7578
rect 29821 7520 29826 7576
rect 29882 7520 31390 7576
rect 31446 7520 31451 7576
rect 29821 7518 31451 7520
rect 29821 7515 29887 7518
rect 31385 7515 31451 7518
rect 13721 7440 16314 7442
rect 13721 7384 13726 7440
rect 13782 7384 16314 7440
rect 13721 7382 16314 7384
rect 17401 7442 17467 7445
rect 27521 7442 27587 7445
rect 17401 7440 27587 7442
rect 17401 7384 17406 7440
rect 17462 7384 27526 7440
rect 27582 7384 27587 7440
rect 17401 7382 27587 7384
rect 13721 7379 13787 7382
rect 17401 7379 17467 7382
rect 27521 7379 27587 7382
rect 38929 7442 38995 7445
rect 40880 7442 41000 7472
rect 38929 7440 41000 7442
rect 38929 7384 38934 7440
rect 38990 7384 41000 7440
rect 38929 7382 41000 7384
rect 38929 7379 38995 7382
rect 40880 7352 41000 7382
rect 7097 7304 7163 7309
rect 7097 7248 7102 7304
rect 7158 7248 7163 7304
rect 7097 7243 7163 7248
rect 7373 7306 7439 7309
rect 13353 7306 13419 7309
rect 7373 7304 13419 7306
rect 7373 7248 7378 7304
rect 7434 7248 13358 7304
rect 13414 7248 13419 7304
rect 7373 7246 13419 7248
rect 7373 7243 7439 7246
rect 13353 7243 13419 7246
rect 13721 7306 13787 7309
rect 16205 7306 16271 7309
rect 13721 7304 16271 7306
rect 13721 7248 13726 7304
rect 13782 7248 16210 7304
rect 16266 7248 16271 7304
rect 13721 7246 16271 7248
rect 13721 7243 13787 7246
rect 16205 7243 16271 7246
rect 16389 7306 16455 7309
rect 25129 7306 25195 7309
rect 32121 7306 32187 7309
rect 16389 7304 25195 7306
rect 16389 7248 16394 7304
rect 16450 7248 25134 7304
rect 25190 7248 25195 7304
rect 16389 7246 25195 7248
rect 16389 7243 16455 7246
rect 25129 7243 25195 7246
rect 25822 7304 32187 7306
rect 25822 7248 32126 7304
rect 32182 7248 32187 7304
rect 25822 7246 32187 7248
rect 0 7170 120 7200
rect 1117 7170 1183 7173
rect 0 7168 1183 7170
rect 0 7112 1122 7168
rect 1178 7112 1183 7168
rect 0 7110 1183 7112
rect 7100 7170 7160 7243
rect 7465 7170 7531 7173
rect 7100 7168 7531 7170
rect 7100 7112 7470 7168
rect 7526 7112 7531 7168
rect 7100 7110 7531 7112
rect 0 7080 120 7110
rect 1117 7107 1183 7110
rect 7465 7107 7531 7110
rect 8385 7170 8451 7173
rect 9489 7170 9555 7173
rect 8385 7168 9555 7170
rect 8385 7112 8390 7168
rect 8446 7112 9494 7168
rect 9550 7112 9555 7168
rect 8385 7110 9555 7112
rect 8385 7107 8451 7110
rect 9489 7107 9555 7110
rect 11973 7170 12039 7173
rect 12382 7170 12388 7172
rect 11973 7168 12388 7170
rect 11973 7112 11978 7168
rect 12034 7112 12388 7168
rect 11973 7110 12388 7112
rect 11973 7107 12039 7110
rect 12382 7108 12388 7110
rect 12452 7108 12458 7172
rect 14917 7170 14983 7173
rect 18137 7170 18203 7173
rect 14917 7168 18203 7170
rect 14917 7112 14922 7168
rect 14978 7112 18142 7168
rect 18198 7112 18203 7168
rect 14917 7110 18203 7112
rect 14917 7107 14983 7110
rect 18137 7107 18203 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 9949 7036 10015 7037
rect 9949 7034 9996 7036
rect 9904 7032 9996 7034
rect 9904 6976 9954 7032
rect 9904 6974 9996 6976
rect 9949 6972 9996 6974
rect 10060 6972 10066 7036
rect 10133 7034 10199 7037
rect 13813 7034 13879 7037
rect 10133 7032 13879 7034
rect 10133 6976 10138 7032
rect 10194 6976 13818 7032
rect 13874 6976 13879 7032
rect 10133 6974 13879 6976
rect 9949 6971 10015 6972
rect 10133 6971 10199 6974
rect 13813 6971 13879 6974
rect 14365 7034 14431 7037
rect 17677 7034 17743 7037
rect 14365 7032 17743 7034
rect 14365 6976 14370 7032
rect 14426 6976 17682 7032
rect 17738 6976 17743 7032
rect 14365 6974 17743 6976
rect 14365 6971 14431 6974
rect 17677 6971 17743 6974
rect 20989 7034 21055 7037
rect 25822 7034 25882 7246
rect 32121 7243 32187 7246
rect 39389 7170 39455 7173
rect 40880 7170 41000 7200
rect 39389 7168 41000 7170
rect 39389 7112 39394 7168
rect 39450 7112 41000 7168
rect 39389 7110 41000 7112
rect 39389 7107 39455 7110
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 37946 7104 38262 7105
rect 37946 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38262 7104
rect 40880 7080 41000 7110
rect 37946 7039 38262 7040
rect 29085 7034 29151 7037
rect 32673 7034 32739 7037
rect 20989 7032 25882 7034
rect 20989 6976 20994 7032
rect 21050 6976 25882 7032
rect 20989 6974 25882 6976
rect 26374 7032 29151 7034
rect 26374 6976 29090 7032
rect 29146 6976 29151 7032
rect 26374 6974 29151 6976
rect 20989 6971 21055 6974
rect 0 6898 120 6928
rect 2957 6898 3023 6901
rect 0 6896 3023 6898
rect 0 6840 2962 6896
rect 3018 6840 3023 6896
rect 0 6838 3023 6840
rect 0 6808 120 6838
rect 2957 6835 3023 6838
rect 7281 6898 7347 6901
rect 9949 6898 10015 6901
rect 13353 6898 13419 6901
rect 14457 6898 14523 6901
rect 7281 6896 9874 6898
rect 7281 6840 7286 6896
rect 7342 6840 9874 6896
rect 7281 6838 9874 6840
rect 7281 6835 7347 6838
rect 7557 6762 7623 6765
rect 9814 6762 9874 6838
rect 9949 6896 13419 6898
rect 9949 6840 9954 6896
rect 10010 6840 13358 6896
rect 13414 6840 13419 6896
rect 9949 6838 13419 6840
rect 9949 6835 10015 6838
rect 13353 6835 13419 6838
rect 13494 6896 14523 6898
rect 13494 6840 14462 6896
rect 14518 6840 14523 6896
rect 13494 6838 14523 6840
rect 13494 6762 13554 6838
rect 14457 6835 14523 6838
rect 14641 6898 14707 6901
rect 20805 6898 20871 6901
rect 14641 6896 20871 6898
rect 14641 6840 14646 6896
rect 14702 6840 20810 6896
rect 20866 6840 20871 6896
rect 14641 6838 20871 6840
rect 14641 6835 14707 6838
rect 20805 6835 20871 6838
rect 24669 6898 24735 6901
rect 26374 6898 26434 6974
rect 29085 6971 29151 6974
rect 32446 7032 32739 7034
rect 32446 6976 32678 7032
rect 32734 6976 32739 7032
rect 32446 6974 32739 6976
rect 24669 6896 26434 6898
rect 24669 6840 24674 6896
rect 24730 6840 26434 6896
rect 24669 6838 26434 6840
rect 30833 6898 30899 6901
rect 32446 6898 32506 6974
rect 32673 6971 32739 6974
rect 30833 6896 32506 6898
rect 30833 6840 30838 6896
rect 30894 6840 32506 6896
rect 30833 6838 32506 6840
rect 40033 6898 40099 6901
rect 40880 6898 41000 6928
rect 40033 6896 41000 6898
rect 40033 6840 40038 6896
rect 40094 6840 41000 6896
rect 40033 6838 41000 6840
rect 24669 6835 24735 6838
rect 30833 6835 30899 6838
rect 40033 6835 40099 6838
rect 40880 6808 41000 6838
rect 30373 6762 30439 6765
rect 7557 6760 9506 6762
rect 7557 6704 7562 6760
rect 7618 6704 9506 6760
rect 7557 6702 9506 6704
rect 9814 6702 13554 6762
rect 13678 6760 30439 6762
rect 13678 6704 30378 6760
rect 30434 6704 30439 6760
rect 13678 6702 30439 6704
rect 7557 6699 7623 6702
rect 0 6626 120 6656
rect 197 6626 263 6629
rect 0 6624 263 6626
rect 0 6568 202 6624
rect 258 6568 263 6624
rect 0 6566 263 6568
rect 0 6536 120 6566
rect 197 6563 263 6566
rect 7281 6626 7347 6629
rect 8477 6626 8543 6629
rect 7281 6624 8543 6626
rect 7281 6568 7286 6624
rect 7342 6568 8482 6624
rect 8538 6568 8543 6624
rect 7281 6566 8543 6568
rect 7281 6563 7347 6566
rect 8477 6563 8543 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 7925 6490 7991 6493
rect 8753 6490 8819 6493
rect 7925 6488 8819 6490
rect 7925 6432 7930 6488
rect 7986 6432 8758 6488
rect 8814 6432 8819 6488
rect 7925 6430 8819 6432
rect 9446 6490 9506 6702
rect 9765 6626 9831 6629
rect 13678 6626 13738 6702
rect 30373 6699 30439 6702
rect 9765 6624 13738 6626
rect 9765 6568 9770 6624
rect 9826 6568 13738 6624
rect 9765 6566 13738 6568
rect 15469 6626 15535 6629
rect 20621 6626 20687 6629
rect 15469 6624 20687 6626
rect 15469 6568 15474 6624
rect 15530 6568 20626 6624
rect 20682 6568 20687 6624
rect 15469 6566 20687 6568
rect 9765 6563 9831 6566
rect 15469 6563 15535 6566
rect 20621 6563 20687 6566
rect 21725 6626 21791 6629
rect 26601 6626 26667 6629
rect 21725 6624 26667 6626
rect 21725 6568 21730 6624
rect 21786 6568 26606 6624
rect 26662 6568 26667 6624
rect 21725 6566 26667 6568
rect 21725 6563 21791 6566
rect 26601 6563 26667 6566
rect 39665 6626 39731 6629
rect 40880 6626 41000 6656
rect 39665 6624 41000 6626
rect 39665 6568 39670 6624
rect 39726 6568 41000 6624
rect 39665 6566 41000 6568
rect 39665 6563 39731 6566
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 33006 6495 33322 6496
rect 39006 6560 39322 6561
rect 39006 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39322 6560
rect 40880 6536 41000 6566
rect 39006 6495 39322 6496
rect 9446 6430 14842 6490
rect 7925 6427 7991 6430
rect 8753 6427 8819 6430
rect 0 6354 120 6384
rect 933 6354 999 6357
rect 0 6352 999 6354
rect 0 6296 938 6352
rect 994 6296 999 6352
rect 0 6294 999 6296
rect 0 6264 120 6294
rect 933 6291 999 6294
rect 4153 6354 4219 6357
rect 9949 6354 10015 6357
rect 4153 6352 10015 6354
rect 4153 6296 4158 6352
rect 4214 6296 9954 6352
rect 10010 6296 10015 6352
rect 4153 6294 10015 6296
rect 4153 6291 4219 6294
rect 9949 6291 10015 6294
rect 11053 6354 11119 6357
rect 14641 6354 14707 6357
rect 11053 6352 14707 6354
rect 11053 6296 11058 6352
rect 11114 6296 14646 6352
rect 14702 6296 14707 6352
rect 11053 6294 14707 6296
rect 14782 6354 14842 6430
rect 19558 6428 19564 6492
rect 19628 6490 19634 6492
rect 19701 6490 19767 6493
rect 19628 6488 19767 6490
rect 19628 6432 19706 6488
rect 19762 6432 19767 6488
rect 19628 6430 19767 6432
rect 19628 6428 19634 6430
rect 19701 6427 19767 6430
rect 25405 6490 25471 6493
rect 25957 6490 26023 6493
rect 25405 6488 26023 6490
rect 25405 6432 25410 6488
rect 25466 6432 25962 6488
rect 26018 6432 26023 6488
rect 25405 6430 26023 6432
rect 25405 6427 25471 6430
rect 25957 6427 26023 6430
rect 29085 6490 29151 6493
rect 31845 6490 31911 6493
rect 29085 6488 31911 6490
rect 29085 6432 29090 6488
rect 29146 6432 31850 6488
rect 31906 6432 31911 6488
rect 29085 6430 31911 6432
rect 29085 6427 29151 6430
rect 31845 6427 31911 6430
rect 27061 6354 27127 6357
rect 14782 6352 27127 6354
rect 14782 6296 27066 6352
rect 27122 6296 27127 6352
rect 14782 6294 27127 6296
rect 11053 6291 11119 6294
rect 14641 6291 14707 6294
rect 27061 6291 27127 6294
rect 27337 6354 27403 6357
rect 31661 6354 31727 6357
rect 27337 6352 31727 6354
rect 27337 6296 27342 6352
rect 27398 6296 31666 6352
rect 31722 6296 31727 6352
rect 27337 6294 31727 6296
rect 27337 6291 27403 6294
rect 31661 6291 31727 6294
rect 38653 6354 38719 6357
rect 40880 6354 41000 6384
rect 38653 6352 41000 6354
rect 38653 6296 38658 6352
rect 38714 6296 41000 6352
rect 38653 6294 41000 6296
rect 38653 6291 38719 6294
rect 40880 6264 41000 6294
rect 1669 6218 1735 6221
rect 18045 6218 18111 6221
rect 20621 6218 20687 6221
rect 26693 6218 26759 6221
rect 1669 6216 18111 6218
rect 1669 6160 1674 6216
rect 1730 6160 18050 6216
rect 18106 6160 18111 6216
rect 1669 6158 18111 6160
rect 1669 6155 1735 6158
rect 18045 6155 18111 6158
rect 18278 6158 20546 6218
rect 0 6082 120 6112
rect 749 6082 815 6085
rect 0 6080 815 6082
rect 0 6024 754 6080
rect 810 6024 815 6080
rect 0 6022 815 6024
rect 0 5992 120 6022
rect 749 6019 815 6022
rect 14457 6082 14523 6085
rect 18278 6082 18338 6158
rect 14457 6080 18338 6082
rect 14457 6024 14462 6080
rect 14518 6024 18338 6080
rect 14457 6022 18338 6024
rect 20486 6082 20546 6158
rect 20621 6216 26759 6218
rect 20621 6160 20626 6216
rect 20682 6160 26698 6216
rect 26754 6160 26759 6216
rect 20621 6158 26759 6160
rect 20621 6155 20687 6158
rect 26693 6155 26759 6158
rect 29913 6218 29979 6221
rect 37641 6218 37707 6221
rect 29913 6216 37707 6218
rect 29913 6160 29918 6216
rect 29974 6160 37646 6216
rect 37702 6160 37707 6216
rect 29913 6158 37707 6160
rect 29913 6155 29979 6158
rect 37641 6155 37707 6158
rect 25129 6082 25195 6085
rect 20486 6080 25195 6082
rect 20486 6024 25134 6080
rect 25190 6024 25195 6080
rect 20486 6022 25195 6024
rect 14457 6019 14523 6022
rect 25129 6019 25195 6022
rect 30649 6082 30715 6085
rect 31661 6082 31727 6085
rect 30649 6080 31727 6082
rect 30649 6024 30654 6080
rect 30710 6024 31666 6080
rect 31722 6024 31727 6080
rect 30649 6022 31727 6024
rect 30649 6019 30715 6022
rect 31661 6019 31727 6022
rect 39021 6082 39087 6085
rect 40880 6082 41000 6112
rect 39021 6080 41000 6082
rect 39021 6024 39026 6080
rect 39082 6024 41000 6080
rect 39021 6022 41000 6024
rect 39021 6019 39087 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 37946 6016 38262 6017
rect 37946 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38262 6016
rect 40880 5992 41000 6022
rect 37946 5951 38262 5952
rect 11789 5946 11855 5949
rect 12985 5946 13051 5949
rect 11789 5944 13051 5946
rect 11789 5888 11794 5944
rect 11850 5888 12990 5944
rect 13046 5888 13051 5944
rect 11789 5886 13051 5888
rect 11789 5883 11855 5886
rect 12985 5883 13051 5886
rect 14457 5946 14523 5949
rect 15837 5946 15903 5949
rect 14457 5944 15903 5946
rect 14457 5888 14462 5944
rect 14518 5888 15842 5944
rect 15898 5888 15903 5944
rect 14457 5886 15903 5888
rect 14457 5883 14523 5886
rect 15837 5883 15903 5886
rect 20897 5946 20963 5949
rect 24853 5946 24919 5949
rect 28533 5946 28599 5949
rect 20897 5944 24919 5946
rect 20897 5888 20902 5944
rect 20958 5888 24858 5944
rect 24914 5888 24919 5944
rect 20897 5886 24919 5888
rect 20897 5883 20963 5886
rect 24853 5883 24919 5886
rect 26328 5944 28599 5946
rect 26328 5888 28538 5944
rect 28594 5888 28599 5944
rect 26328 5886 28599 5888
rect 0 5810 120 5840
rect 749 5810 815 5813
rect 0 5808 815 5810
rect 0 5752 754 5808
rect 810 5752 815 5808
rect 0 5750 815 5752
rect 0 5720 120 5750
rect 749 5747 815 5750
rect 6637 5810 6703 5813
rect 17861 5810 17927 5813
rect 6637 5808 17927 5810
rect 6637 5752 6642 5808
rect 6698 5752 17866 5808
rect 17922 5752 17927 5808
rect 6637 5750 17927 5752
rect 6637 5747 6703 5750
rect 17861 5747 17927 5750
rect 18045 5810 18111 5813
rect 24669 5810 24735 5813
rect 18045 5808 24735 5810
rect 18045 5752 18050 5808
rect 18106 5752 24674 5808
rect 24730 5752 24735 5808
rect 18045 5750 24735 5752
rect 18045 5747 18111 5750
rect 24669 5747 24735 5750
rect 24853 5810 24919 5813
rect 26328 5810 26388 5886
rect 28533 5883 28599 5886
rect 38837 5810 38903 5813
rect 24853 5808 26388 5810
rect 24853 5752 24858 5808
rect 24914 5752 26388 5808
rect 24853 5750 26388 5752
rect 26926 5808 38903 5810
rect 26926 5752 38842 5808
rect 38898 5752 38903 5808
rect 26926 5750 38903 5752
rect 24853 5747 24919 5750
rect 5073 5674 5139 5677
rect 7649 5674 7715 5677
rect 5073 5672 7715 5674
rect 5073 5616 5078 5672
rect 5134 5616 7654 5672
rect 7710 5616 7715 5672
rect 5073 5614 7715 5616
rect 5073 5611 5139 5614
rect 7649 5611 7715 5614
rect 8702 5612 8708 5676
rect 8772 5674 8778 5676
rect 9489 5674 9555 5677
rect 8772 5672 9555 5674
rect 8772 5616 9494 5672
rect 9550 5616 9555 5672
rect 8772 5614 9555 5616
rect 8772 5612 8778 5614
rect 9489 5611 9555 5614
rect 9765 5674 9831 5677
rect 16297 5674 16363 5677
rect 9765 5672 16363 5674
rect 9765 5616 9770 5672
rect 9826 5616 16302 5672
rect 16358 5616 16363 5672
rect 9765 5614 16363 5616
rect 9765 5611 9831 5614
rect 16297 5611 16363 5614
rect 16941 5674 17007 5677
rect 26926 5674 26986 5750
rect 38837 5747 38903 5750
rect 39389 5810 39455 5813
rect 40880 5810 41000 5840
rect 39389 5808 41000 5810
rect 39389 5752 39394 5808
rect 39450 5752 41000 5808
rect 39389 5750 41000 5752
rect 39389 5747 39455 5750
rect 40880 5720 41000 5750
rect 16941 5672 26986 5674
rect 16941 5616 16946 5672
rect 17002 5616 26986 5672
rect 16941 5614 26986 5616
rect 27061 5674 27127 5677
rect 33961 5674 34027 5677
rect 27061 5672 34027 5674
rect 27061 5616 27066 5672
rect 27122 5616 33966 5672
rect 34022 5616 34027 5672
rect 27061 5614 34027 5616
rect 16941 5611 17007 5614
rect 27061 5611 27127 5614
rect 33961 5611 34027 5614
rect 0 5538 120 5568
rect 565 5538 631 5541
rect 0 5536 631 5538
rect 0 5480 570 5536
rect 626 5480 631 5536
rect 0 5478 631 5480
rect 0 5448 120 5478
rect 565 5475 631 5478
rect 7097 5538 7163 5541
rect 8201 5538 8267 5541
rect 7097 5536 8267 5538
rect 7097 5480 7102 5536
rect 7158 5480 8206 5536
rect 8262 5480 8267 5536
rect 7097 5478 8267 5480
rect 7097 5475 7163 5478
rect 8201 5475 8267 5478
rect 10041 5538 10107 5541
rect 14273 5538 14339 5541
rect 10041 5536 14339 5538
rect 10041 5480 10046 5536
rect 10102 5480 14278 5536
rect 14334 5480 14339 5536
rect 10041 5478 14339 5480
rect 10041 5475 10107 5478
rect 14273 5475 14339 5478
rect 18597 5538 18663 5541
rect 19241 5538 19307 5541
rect 18597 5536 19307 5538
rect 18597 5480 18602 5536
rect 18658 5480 19246 5536
rect 19302 5480 19307 5536
rect 18597 5478 19307 5480
rect 18597 5475 18663 5478
rect 19241 5475 19307 5478
rect 19517 5538 19583 5541
rect 20805 5538 20871 5541
rect 19517 5536 20871 5538
rect 19517 5480 19522 5536
rect 19578 5480 20810 5536
rect 20866 5480 20871 5536
rect 19517 5478 20871 5480
rect 19517 5475 19583 5478
rect 20805 5475 20871 5478
rect 30189 5538 30255 5541
rect 31201 5538 31267 5541
rect 30189 5536 31267 5538
rect 30189 5480 30194 5536
rect 30250 5480 31206 5536
rect 31262 5480 31267 5536
rect 30189 5478 31267 5480
rect 30189 5475 30255 5478
rect 31201 5475 31267 5478
rect 39941 5538 40007 5541
rect 40880 5538 41000 5568
rect 39941 5536 41000 5538
rect 39941 5480 39946 5536
rect 40002 5480 41000 5536
rect 39941 5478 41000 5480
rect 39941 5475 40007 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 33006 5407 33322 5408
rect 39006 5472 39322 5473
rect 39006 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39322 5472
rect 40880 5448 41000 5478
rect 39006 5407 39322 5408
rect 5809 5402 5875 5405
rect 8845 5402 8911 5405
rect 5809 5400 8911 5402
rect 5809 5344 5814 5400
rect 5870 5344 8850 5400
rect 8906 5344 8911 5400
rect 5809 5342 8911 5344
rect 5809 5339 5875 5342
rect 8845 5339 8911 5342
rect 11053 5402 11119 5405
rect 16021 5402 16087 5405
rect 19425 5402 19491 5405
rect 19742 5402 19748 5404
rect 11053 5400 14842 5402
rect 11053 5344 11058 5400
rect 11114 5344 14842 5400
rect 11053 5342 14842 5344
rect 11053 5339 11119 5342
rect 0 5266 120 5296
rect 1025 5266 1091 5269
rect 0 5264 1091 5266
rect 0 5208 1030 5264
rect 1086 5208 1091 5264
rect 0 5206 1091 5208
rect 0 5176 120 5206
rect 1025 5203 1091 5206
rect 4337 5266 4403 5269
rect 4337 5264 14658 5266
rect 4337 5208 4342 5264
rect 4398 5208 14658 5264
rect 4337 5206 14658 5208
rect 4337 5203 4403 5206
rect 5901 5130 5967 5133
rect 6453 5130 6519 5133
rect 7281 5130 7347 5133
rect 5901 5128 7347 5130
rect 5901 5072 5906 5128
rect 5962 5072 6458 5128
rect 6514 5072 7286 5128
rect 7342 5072 7347 5128
rect 5901 5070 7347 5072
rect 5901 5067 5967 5070
rect 6453 5067 6519 5070
rect 7281 5067 7347 5070
rect 7649 5128 7715 5133
rect 7649 5072 7654 5128
rect 7710 5072 7715 5128
rect 7649 5067 7715 5072
rect 8201 5130 8267 5133
rect 9397 5130 9463 5133
rect 8201 5128 9276 5130
rect 8201 5072 8206 5128
rect 8262 5072 9276 5128
rect 8201 5070 9276 5072
rect 8201 5067 8267 5070
rect 0 4994 120 5024
rect 381 4994 447 4997
rect 0 4992 447 4994
rect 0 4936 386 4992
rect 442 4936 447 4992
rect 0 4934 447 4936
rect 0 4904 120 4934
rect 381 4931 447 4934
rect 7189 4994 7255 4997
rect 7652 4994 7712 5067
rect 7189 4992 7712 4994
rect 7189 4936 7194 4992
rect 7250 4936 7712 4992
rect 7189 4934 7712 4936
rect 9216 4994 9276 5070
rect 9397 5128 14520 5130
rect 9397 5072 9402 5128
rect 9458 5072 14520 5128
rect 9397 5070 14520 5072
rect 9397 5067 9463 5070
rect 13721 4994 13787 4997
rect 9216 4992 13787 4994
rect 9216 4936 13726 4992
rect 13782 4936 13787 4992
rect 9216 4934 13787 4936
rect 7189 4931 7255 4934
rect 13721 4931 13787 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 10409 4858 10475 4861
rect 13537 4858 13603 4861
rect 10409 4856 13603 4858
rect 10409 4800 10414 4856
rect 10470 4800 13542 4856
rect 13598 4800 13603 4856
rect 10409 4798 13603 4800
rect 14460 4858 14520 5070
rect 14598 4994 14658 5206
rect 14782 5130 14842 5342
rect 16021 5400 19748 5402
rect 16021 5344 16026 5400
rect 16082 5344 19430 5400
rect 19486 5344 19748 5400
rect 16021 5342 19748 5344
rect 16021 5339 16087 5342
rect 19425 5339 19491 5342
rect 19742 5340 19748 5342
rect 19812 5340 19818 5404
rect 15285 5266 15351 5269
rect 15469 5266 15535 5269
rect 15285 5264 15535 5266
rect 15285 5208 15290 5264
rect 15346 5208 15474 5264
rect 15530 5208 15535 5264
rect 15285 5206 15535 5208
rect 15285 5203 15351 5206
rect 15469 5203 15535 5206
rect 17217 5266 17283 5269
rect 28993 5266 29059 5269
rect 17217 5264 29059 5266
rect 17217 5208 17222 5264
rect 17278 5208 28998 5264
rect 29054 5208 29059 5264
rect 17217 5206 29059 5208
rect 17217 5203 17283 5206
rect 28993 5203 29059 5206
rect 29177 5266 29243 5269
rect 36905 5266 36971 5269
rect 29177 5264 36971 5266
rect 29177 5208 29182 5264
rect 29238 5208 36910 5264
rect 36966 5208 36971 5264
rect 29177 5206 36971 5208
rect 29177 5203 29243 5206
rect 36905 5203 36971 5206
rect 39389 5266 39455 5269
rect 40880 5266 41000 5296
rect 39389 5264 41000 5266
rect 39389 5208 39394 5264
rect 39450 5208 41000 5264
rect 39389 5206 41000 5208
rect 39389 5203 39455 5206
rect 40880 5176 41000 5206
rect 19977 5130 20043 5133
rect 14782 5128 20043 5130
rect 14782 5072 19982 5128
rect 20038 5072 20043 5128
rect 14782 5070 20043 5072
rect 19977 5067 20043 5070
rect 20161 5130 20227 5133
rect 26049 5130 26115 5133
rect 27981 5130 28047 5133
rect 37825 5130 37891 5133
rect 20161 5128 20546 5130
rect 20161 5072 20166 5128
rect 20222 5072 20546 5128
rect 20161 5070 20546 5072
rect 20161 5067 20227 5070
rect 19793 4994 19859 4997
rect 14598 4992 19859 4994
rect 14598 4936 19798 4992
rect 19854 4936 19859 4992
rect 14598 4934 19859 4936
rect 20486 4994 20546 5070
rect 26049 5128 26802 5130
rect 26049 5072 26054 5128
rect 26110 5072 26802 5128
rect 26049 5070 26802 5072
rect 26049 5067 26115 5070
rect 24761 4994 24827 4997
rect 20486 4992 24827 4994
rect 20486 4936 24766 4992
rect 24822 4936 24827 4992
rect 20486 4934 24827 4936
rect 26742 4994 26802 5070
rect 27981 5128 37891 5130
rect 27981 5072 27986 5128
rect 28042 5072 37830 5128
rect 37886 5072 37891 5128
rect 27981 5070 37891 5072
rect 27981 5067 28047 5070
rect 37825 5067 37891 5070
rect 30557 4994 30623 4997
rect 26742 4992 30623 4994
rect 26742 4936 30562 4992
rect 30618 4936 30623 4992
rect 26742 4934 30623 4936
rect 19793 4931 19859 4934
rect 24761 4931 24827 4934
rect 30557 4931 30623 4934
rect 39021 4994 39087 4997
rect 40880 4994 41000 5024
rect 39021 4992 41000 4994
rect 39021 4936 39026 4992
rect 39082 4936 41000 4992
rect 39021 4934 41000 4936
rect 39021 4931 39087 4934
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 37946 4928 38262 4929
rect 37946 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38262 4928
rect 40880 4904 41000 4934
rect 37946 4863 38262 4864
rect 16021 4858 16087 4861
rect 14460 4856 16087 4858
rect 14460 4800 16026 4856
rect 16082 4800 16087 4856
rect 14460 4798 16087 4800
rect 10409 4795 10475 4798
rect 13537 4795 13603 4798
rect 16021 4795 16087 4798
rect 16297 4858 16363 4861
rect 19517 4858 19583 4861
rect 16297 4856 19583 4858
rect 16297 4800 16302 4856
rect 16358 4800 19522 4856
rect 19578 4800 19583 4856
rect 16297 4798 19583 4800
rect 16297 4795 16363 4798
rect 19517 4795 19583 4798
rect 20437 4858 20503 4861
rect 23657 4858 23723 4861
rect 20437 4856 23723 4858
rect 20437 4800 20442 4856
rect 20498 4800 23662 4856
rect 23718 4800 23723 4856
rect 20437 4798 23723 4800
rect 20437 4795 20503 4798
rect 23657 4795 23723 4798
rect 0 4722 120 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 120 4662
rect 933 4659 999 4662
rect 4521 4722 4587 4725
rect 27061 4722 27127 4725
rect 4521 4720 27127 4722
rect 4521 4664 4526 4720
rect 4582 4664 27066 4720
rect 27122 4664 27127 4720
rect 4521 4662 27127 4664
rect 4521 4659 4587 4662
rect 27061 4659 27127 4662
rect 31385 4722 31451 4725
rect 31937 4722 32003 4725
rect 31385 4720 32003 4722
rect 31385 4664 31390 4720
rect 31446 4664 31942 4720
rect 31998 4664 32003 4720
rect 31385 4662 32003 4664
rect 31385 4659 31451 4662
rect 31937 4659 32003 4662
rect 39481 4722 39547 4725
rect 40880 4722 41000 4752
rect 39481 4720 41000 4722
rect 39481 4664 39486 4720
rect 39542 4664 41000 4720
rect 39481 4662 41000 4664
rect 39481 4659 39547 4662
rect 40880 4632 41000 4662
rect 7649 4586 7715 4589
rect 14917 4586 14983 4589
rect 7649 4584 12450 4586
rect 7649 4528 7654 4584
rect 7710 4528 12450 4584
rect 7649 4526 12450 4528
rect 7649 4523 7715 4526
rect 0 4450 120 4480
rect 749 4450 815 4453
rect 0 4448 815 4450
rect 0 4392 754 4448
rect 810 4392 815 4448
rect 0 4390 815 4392
rect 12390 4450 12450 4526
rect 14414 4584 14983 4586
rect 14414 4528 14922 4584
rect 14978 4528 14983 4584
rect 14414 4526 14983 4528
rect 14414 4450 14474 4526
rect 14917 4523 14983 4526
rect 15193 4586 15259 4589
rect 31017 4586 31083 4589
rect 15193 4584 31083 4586
rect 15193 4528 15198 4584
rect 15254 4528 31022 4584
rect 31078 4528 31083 4584
rect 15193 4526 31083 4528
rect 15193 4523 15259 4526
rect 31017 4523 31083 4526
rect 31477 4586 31543 4589
rect 36261 4586 36327 4589
rect 31477 4584 36327 4586
rect 31477 4528 31482 4584
rect 31538 4528 36266 4584
rect 36322 4528 36327 4584
rect 31477 4526 36327 4528
rect 31477 4523 31543 4526
rect 36261 4523 36327 4526
rect 12390 4390 14474 4450
rect 17217 4450 17283 4453
rect 20437 4450 20503 4453
rect 17217 4448 20503 4450
rect 17217 4392 17222 4448
rect 17278 4392 20442 4448
rect 20498 4392 20503 4448
rect 17217 4390 20503 4392
rect 0 4360 120 4390
rect 749 4387 815 4390
rect 17217 4387 17283 4390
rect 20437 4387 20503 4390
rect 39941 4450 40007 4453
rect 40880 4450 41000 4480
rect 39941 4448 41000 4450
rect 39941 4392 39946 4448
rect 40002 4392 41000 4448
rect 39941 4390 41000 4392
rect 39941 4387 40007 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 33006 4319 33322 4320
rect 39006 4384 39322 4385
rect 39006 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39322 4384
rect 40880 4360 41000 4390
rect 39006 4319 39322 4320
rect 8661 4314 8727 4317
rect 5076 4312 8727 4314
rect 5076 4256 8666 4312
rect 8722 4256 8727 4312
rect 5076 4254 8727 4256
rect 0 4178 120 4208
rect 749 4178 815 4181
rect 0 4176 815 4178
rect 0 4120 754 4176
rect 810 4120 815 4176
rect 0 4118 815 4120
rect 0 4088 120 4118
rect 749 4115 815 4118
rect 1945 4178 2011 4181
rect 5076 4178 5136 4254
rect 8661 4251 8727 4254
rect 9857 4314 9923 4317
rect 14457 4314 14523 4317
rect 9857 4312 14523 4314
rect 9857 4256 9862 4312
rect 9918 4256 14462 4312
rect 14518 4256 14523 4312
rect 9857 4254 14523 4256
rect 9857 4251 9923 4254
rect 14457 4251 14523 4254
rect 15837 4314 15903 4317
rect 19057 4314 19123 4317
rect 15837 4312 19123 4314
rect 15837 4256 15842 4312
rect 15898 4256 19062 4312
rect 19118 4256 19123 4312
rect 15837 4254 19123 4256
rect 15837 4251 15903 4254
rect 19057 4251 19123 4254
rect 19425 4314 19491 4317
rect 20069 4314 20135 4317
rect 20621 4316 20687 4317
rect 20621 4314 20668 4316
rect 19425 4312 20135 4314
rect 19425 4256 19430 4312
rect 19486 4256 20074 4312
rect 20130 4256 20135 4312
rect 19425 4254 20135 4256
rect 20576 4312 20668 4314
rect 20576 4256 20626 4312
rect 20576 4254 20668 4256
rect 19425 4251 19491 4254
rect 20069 4251 20135 4254
rect 20621 4252 20668 4254
rect 20732 4252 20738 4316
rect 20621 4251 20687 4252
rect 1945 4176 5136 4178
rect 1945 4120 1950 4176
rect 2006 4120 5136 4176
rect 1945 4118 5136 4120
rect 5257 4178 5323 4181
rect 19425 4178 19491 4181
rect 25497 4178 25563 4181
rect 5257 4176 16498 4178
rect 5257 4120 5262 4176
rect 5318 4120 16498 4176
rect 5257 4118 16498 4120
rect 1945 4115 2011 4118
rect 5257 4115 5323 4118
rect 2313 4042 2379 4045
rect 9397 4042 9463 4045
rect 2313 4040 9463 4042
rect 2313 3984 2318 4040
rect 2374 3984 9402 4040
rect 9458 3984 9463 4040
rect 2313 3982 9463 3984
rect 2313 3979 2379 3982
rect 9397 3979 9463 3982
rect 9765 4042 9831 4045
rect 16438 4042 16498 4118
rect 19425 4176 25563 4178
rect 19425 4120 19430 4176
rect 19486 4120 25502 4176
rect 25558 4120 25563 4176
rect 19425 4118 25563 4120
rect 19425 4115 19491 4118
rect 25497 4115 25563 4118
rect 31109 4178 31175 4181
rect 35157 4178 35223 4181
rect 31109 4176 35223 4178
rect 31109 4120 31114 4176
rect 31170 4120 35162 4176
rect 35218 4120 35223 4176
rect 31109 4118 35223 4120
rect 31109 4115 31175 4118
rect 35157 4115 35223 4118
rect 39389 4178 39455 4181
rect 40880 4178 41000 4208
rect 39389 4176 41000 4178
rect 39389 4120 39394 4176
rect 39450 4120 41000 4176
rect 39389 4118 41000 4120
rect 39389 4115 39455 4118
rect 40880 4088 41000 4118
rect 22553 4042 22619 4045
rect 9765 4040 16314 4042
rect 9765 3984 9770 4040
rect 9826 3984 16314 4040
rect 9765 3982 16314 3984
rect 16438 4040 22619 4042
rect 16438 3984 22558 4040
rect 22614 3984 22619 4040
rect 16438 3982 22619 3984
rect 9765 3979 9831 3982
rect 0 3906 120 3936
rect 933 3906 999 3909
rect 0 3904 999 3906
rect 0 3848 938 3904
rect 994 3848 999 3904
rect 0 3846 999 3848
rect 0 3816 120 3846
rect 933 3843 999 3846
rect 9765 3906 9831 3909
rect 10409 3906 10475 3909
rect 9765 3904 10475 3906
rect 9765 3848 9770 3904
rect 9826 3848 10414 3904
rect 10470 3848 10475 3904
rect 9765 3846 10475 3848
rect 9765 3843 9831 3846
rect 10409 3843 10475 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 0 3634 120 3664
rect 565 3634 631 3637
rect 0 3632 631 3634
rect 0 3576 570 3632
rect 626 3576 631 3632
rect 0 3574 631 3576
rect 0 3544 120 3574
rect 565 3571 631 3574
rect 2497 3634 2563 3637
rect 9305 3634 9371 3637
rect 2497 3632 9371 3634
rect 2497 3576 2502 3632
rect 2558 3576 9310 3632
rect 9366 3576 9371 3632
rect 2497 3574 9371 3576
rect 2497 3571 2563 3574
rect 9305 3571 9371 3574
rect 9857 3634 9923 3637
rect 16021 3634 16087 3637
rect 9857 3632 16087 3634
rect 9857 3576 9862 3632
rect 9918 3576 16026 3632
rect 16082 3576 16087 3632
rect 9857 3574 16087 3576
rect 16254 3634 16314 3982
rect 22553 3979 22619 3982
rect 24853 4042 24919 4045
rect 37549 4042 37615 4045
rect 24853 4040 37615 4042
rect 24853 3984 24858 4040
rect 24914 3984 37554 4040
rect 37610 3984 37615 4040
rect 24853 3982 37615 3984
rect 24853 3979 24919 3982
rect 37549 3979 37615 3982
rect 20437 3906 20503 3909
rect 25681 3906 25747 3909
rect 20437 3904 25747 3906
rect 20437 3848 20442 3904
rect 20498 3848 25686 3904
rect 25742 3848 25747 3904
rect 20437 3846 25747 3848
rect 20437 3843 20503 3846
rect 25681 3843 25747 3846
rect 39021 3906 39087 3909
rect 40880 3906 41000 3936
rect 39021 3904 41000 3906
rect 39021 3848 39026 3904
rect 39082 3848 41000 3904
rect 39021 3846 41000 3848
rect 39021 3843 39087 3846
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 37946 3840 38262 3841
rect 37946 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38262 3840
rect 40880 3816 41000 3846
rect 37946 3775 38262 3776
rect 20529 3770 20595 3773
rect 25773 3770 25839 3773
rect 20529 3768 25839 3770
rect 20529 3712 20534 3768
rect 20590 3712 25778 3768
rect 25834 3712 25839 3768
rect 20529 3710 25839 3712
rect 20529 3707 20595 3710
rect 25773 3707 25839 3710
rect 30465 3770 30531 3773
rect 31661 3770 31727 3773
rect 30465 3768 31727 3770
rect 30465 3712 30470 3768
rect 30526 3712 31666 3768
rect 31722 3712 31727 3768
rect 30465 3710 31727 3712
rect 30465 3707 30531 3710
rect 31661 3707 31727 3710
rect 27429 3634 27495 3637
rect 16254 3632 27495 3634
rect 16254 3576 27434 3632
rect 27490 3576 27495 3632
rect 16254 3574 27495 3576
rect 9857 3571 9923 3574
rect 16021 3571 16087 3574
rect 27429 3571 27495 3574
rect 29453 3634 29519 3637
rect 33501 3634 33567 3637
rect 29453 3632 33567 3634
rect 29453 3576 29458 3632
rect 29514 3576 33506 3632
rect 33562 3576 33567 3632
rect 29453 3574 33567 3576
rect 29453 3571 29519 3574
rect 33501 3571 33567 3574
rect 39389 3634 39455 3637
rect 40880 3634 41000 3664
rect 39389 3632 41000 3634
rect 39389 3576 39394 3632
rect 39450 3576 41000 3632
rect 39389 3574 41000 3576
rect 39389 3571 39455 3574
rect 40880 3544 41000 3574
rect 5717 3498 5783 3501
rect 7649 3498 7715 3501
rect 20529 3498 20595 3501
rect 21909 3498 21975 3501
rect 5717 3496 20595 3498
rect 5717 3440 5722 3496
rect 5778 3440 7654 3496
rect 7710 3440 20534 3496
rect 20590 3440 20595 3496
rect 5717 3438 20595 3440
rect 5717 3435 5783 3438
rect 7649 3435 7715 3438
rect 20529 3435 20595 3438
rect 20670 3496 21975 3498
rect 20670 3440 21914 3496
rect 21970 3440 21975 3496
rect 20670 3438 21975 3440
rect 0 3362 120 3392
rect 197 3362 263 3365
rect 0 3360 263 3362
rect 0 3304 202 3360
rect 258 3304 263 3360
rect 0 3302 263 3304
rect 0 3272 120 3302
rect 197 3299 263 3302
rect 9397 3362 9463 3365
rect 14365 3362 14431 3365
rect 9397 3360 14431 3362
rect 9397 3304 9402 3360
rect 9458 3304 14370 3360
rect 14426 3304 14431 3360
rect 9397 3302 14431 3304
rect 9397 3299 9463 3302
rect 14365 3299 14431 3302
rect 16021 3362 16087 3365
rect 18137 3362 18203 3365
rect 16021 3360 18203 3362
rect 16021 3304 16026 3360
rect 16082 3304 18142 3360
rect 18198 3304 18203 3360
rect 16021 3302 18203 3304
rect 16021 3299 16087 3302
rect 18137 3299 18203 3302
rect 18321 3362 18387 3365
rect 20670 3362 20730 3438
rect 21909 3435 21975 3438
rect 22737 3498 22803 3501
rect 38837 3498 38903 3501
rect 22737 3496 38903 3498
rect 22737 3440 22742 3496
rect 22798 3440 38842 3496
rect 38898 3440 38903 3496
rect 22737 3438 38903 3440
rect 22737 3435 22803 3438
rect 38837 3435 38903 3438
rect 18321 3360 20730 3362
rect 18321 3304 18326 3360
rect 18382 3304 20730 3360
rect 18321 3302 20730 3304
rect 30281 3362 30347 3365
rect 32029 3362 32095 3365
rect 30281 3360 32095 3362
rect 30281 3304 30286 3360
rect 30342 3304 32034 3360
rect 32090 3304 32095 3360
rect 30281 3302 32095 3304
rect 18321 3299 18387 3302
rect 30281 3299 30347 3302
rect 32029 3299 32095 3302
rect 39941 3362 40007 3365
rect 40880 3362 41000 3392
rect 39941 3360 41000 3362
rect 39941 3304 39946 3360
rect 40002 3304 41000 3360
rect 39941 3302 41000 3304
rect 39941 3299 40007 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 33006 3231 33322 3232
rect 39006 3296 39322 3297
rect 39006 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39322 3296
rect 40880 3272 41000 3302
rect 39006 3231 39322 3232
rect 14549 3226 14615 3229
rect 17677 3226 17743 3229
rect 20437 3226 20503 3229
rect 12390 3224 14615 3226
rect 12390 3168 14554 3224
rect 14610 3168 14615 3224
rect 12390 3166 14615 3168
rect 0 3090 120 3120
rect 1301 3090 1367 3093
rect 0 3088 1367 3090
rect 0 3032 1306 3088
rect 1362 3032 1367 3088
rect 0 3030 1367 3032
rect 0 3000 120 3030
rect 1301 3027 1367 3030
rect 5441 3090 5507 3093
rect 12390 3090 12450 3166
rect 14549 3163 14615 3166
rect 15518 3224 20503 3226
rect 15518 3168 17682 3224
rect 17738 3168 20442 3224
rect 20498 3168 20503 3224
rect 15518 3166 20503 3168
rect 5441 3088 12450 3090
rect 5441 3032 5446 3088
rect 5502 3032 12450 3088
rect 5441 3030 12450 3032
rect 13721 3090 13787 3093
rect 15518 3090 15578 3166
rect 17677 3163 17743 3166
rect 20437 3163 20503 3166
rect 21817 3226 21883 3229
rect 22737 3226 22803 3229
rect 21817 3224 22803 3226
rect 21817 3168 21822 3224
rect 21878 3168 22742 3224
rect 22798 3168 22803 3224
rect 21817 3166 22803 3168
rect 21817 3163 21883 3166
rect 22737 3163 22803 3166
rect 13721 3088 15578 3090
rect 13721 3032 13726 3088
rect 13782 3032 15578 3088
rect 13721 3030 15578 3032
rect 16757 3090 16823 3093
rect 31293 3090 31359 3093
rect 16757 3088 31359 3090
rect 16757 3032 16762 3088
rect 16818 3032 31298 3088
rect 31354 3032 31359 3088
rect 16757 3030 31359 3032
rect 5441 3027 5507 3030
rect 13721 3027 13787 3030
rect 16757 3027 16823 3030
rect 31293 3027 31359 3030
rect 39389 3090 39455 3093
rect 40880 3090 41000 3120
rect 39389 3088 41000 3090
rect 39389 3032 39394 3088
rect 39450 3032 41000 3088
rect 39389 3030 41000 3032
rect 39389 3027 39455 3030
rect 40880 3000 41000 3030
rect 3141 2954 3207 2957
rect 30005 2954 30071 2957
rect 38377 2954 38443 2957
rect 3141 2952 29930 2954
rect 3141 2896 3146 2952
rect 3202 2896 29930 2952
rect 3141 2894 29930 2896
rect 3141 2891 3207 2894
rect 0 2818 120 2848
rect 1209 2818 1275 2821
rect 0 2816 1275 2818
rect 0 2760 1214 2816
rect 1270 2760 1275 2816
rect 0 2758 1275 2760
rect 0 2728 120 2758
rect 1209 2755 1275 2758
rect 14549 2818 14615 2821
rect 16021 2818 16087 2821
rect 18321 2818 18387 2821
rect 14549 2816 18387 2818
rect 14549 2760 14554 2816
rect 14610 2760 16026 2816
rect 16082 2760 18326 2816
rect 18382 2760 18387 2816
rect 14549 2758 18387 2760
rect 29870 2818 29930 2894
rect 30005 2952 38443 2954
rect 30005 2896 30010 2952
rect 30066 2896 38382 2952
rect 38438 2896 38443 2952
rect 30005 2894 38443 2896
rect 30005 2891 30071 2894
rect 38377 2891 38443 2894
rect 30373 2818 30439 2821
rect 30741 2818 30807 2821
rect 29870 2816 30807 2818
rect 29870 2760 30378 2816
rect 30434 2760 30746 2816
rect 30802 2760 30807 2816
rect 29870 2758 30807 2760
rect 14549 2755 14615 2758
rect 16021 2755 16087 2758
rect 18321 2755 18387 2758
rect 30373 2755 30439 2758
rect 30741 2755 30807 2758
rect 39021 2818 39087 2821
rect 40880 2818 41000 2848
rect 39021 2816 41000 2818
rect 39021 2760 39026 2816
rect 39082 2760 41000 2816
rect 39021 2758 41000 2760
rect 39021 2755 39087 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 37946 2752 38262 2753
rect 37946 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38262 2752
rect 40880 2728 41000 2758
rect 37946 2687 38262 2688
rect 4705 2682 4771 2685
rect 6545 2682 6611 2685
rect 4705 2680 6611 2682
rect 4705 2624 4710 2680
rect 4766 2624 6550 2680
rect 6606 2624 6611 2680
rect 4705 2622 6611 2624
rect 4705 2619 4771 2622
rect 6545 2619 6611 2622
rect 0 2546 120 2576
rect 381 2546 447 2549
rect 0 2544 447 2546
rect 0 2488 386 2544
rect 442 2488 447 2544
rect 0 2486 447 2488
rect 0 2456 120 2486
rect 381 2483 447 2486
rect 7741 2546 7807 2549
rect 15745 2546 15811 2549
rect 7741 2544 15811 2546
rect 7741 2488 7746 2544
rect 7802 2488 15750 2544
rect 15806 2488 15811 2544
rect 7741 2486 15811 2488
rect 7741 2483 7807 2486
rect 15745 2483 15811 2486
rect 16389 2546 16455 2549
rect 38469 2546 38535 2549
rect 16389 2544 38535 2546
rect 16389 2488 16394 2544
rect 16450 2488 38474 2544
rect 38530 2488 38535 2544
rect 16389 2486 38535 2488
rect 16389 2483 16455 2486
rect 38469 2483 38535 2486
rect 38653 2546 38719 2549
rect 40880 2546 41000 2576
rect 38653 2544 41000 2546
rect 38653 2488 38658 2544
rect 38714 2488 41000 2544
rect 38653 2486 41000 2488
rect 38653 2483 38719 2486
rect 40880 2456 41000 2486
rect 9213 2410 9279 2413
rect 31385 2410 31451 2413
rect 9213 2408 31451 2410
rect 9213 2352 9218 2408
rect 9274 2352 31390 2408
rect 31446 2352 31451 2408
rect 9213 2350 31451 2352
rect 9213 2347 9279 2350
rect 31385 2347 31451 2350
rect 0 2274 120 2304
rect 1117 2274 1183 2277
rect 0 2272 1183 2274
rect 0 2216 1122 2272
rect 1178 2216 1183 2272
rect 0 2214 1183 2216
rect 0 2184 120 2214
rect 1117 2211 1183 2214
rect 39941 2274 40007 2277
rect 40880 2274 41000 2304
rect 39941 2272 41000 2274
rect 39941 2216 39946 2272
rect 40002 2216 41000 2272
rect 39941 2214 41000 2216
rect 39941 2211 40007 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 33006 2143 33322 2144
rect 39006 2208 39322 2209
rect 39006 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39322 2208
rect 40880 2184 41000 2214
rect 39006 2143 39322 2144
rect 0 2002 120 2032
rect 1853 2002 1919 2005
rect 0 2000 1919 2002
rect 0 1944 1858 2000
rect 1914 1944 1919 2000
rect 0 1942 1919 1944
rect 0 1912 120 1942
rect 1853 1939 1919 1942
rect 19517 2002 19583 2005
rect 24669 2002 24735 2005
rect 19517 2000 24735 2002
rect 19517 1944 19522 2000
rect 19578 1944 24674 2000
rect 24730 1944 24735 2000
rect 19517 1942 24735 1944
rect 19517 1939 19583 1942
rect 24669 1939 24735 1942
rect 37917 2002 37983 2005
rect 40880 2002 41000 2032
rect 37917 2000 41000 2002
rect 37917 1944 37922 2000
rect 37978 1944 41000 2000
rect 37917 1942 41000 1944
rect 37917 1939 37983 1942
rect 40880 1912 41000 1942
rect 11973 1866 12039 1869
rect 30189 1866 30255 1869
rect 11973 1864 30255 1866
rect 11973 1808 11978 1864
rect 12034 1808 30194 1864
rect 30250 1808 30255 1864
rect 11973 1806 30255 1808
rect 11973 1803 12039 1806
rect 30189 1803 30255 1806
rect 0 1730 120 1760
rect 1209 1730 1275 1733
rect 0 1728 1275 1730
rect 0 1672 1214 1728
rect 1270 1672 1275 1728
rect 0 1670 1275 1672
rect 0 1640 120 1670
rect 1209 1667 1275 1670
rect 10225 1730 10291 1733
rect 19517 1730 19583 1733
rect 10225 1728 19583 1730
rect 10225 1672 10230 1728
rect 10286 1672 19522 1728
rect 19578 1672 19583 1728
rect 10225 1670 19583 1672
rect 10225 1667 10291 1670
rect 19517 1667 19583 1670
rect 19701 1730 19767 1733
rect 20713 1730 20779 1733
rect 19701 1728 20779 1730
rect 19701 1672 19706 1728
rect 19762 1672 20718 1728
rect 20774 1672 20779 1728
rect 19701 1670 20779 1672
rect 19701 1667 19767 1670
rect 20713 1667 20779 1670
rect 38285 1730 38351 1733
rect 40880 1730 41000 1760
rect 38285 1728 41000 1730
rect 38285 1672 38290 1728
rect 38346 1672 41000 1728
rect 38285 1670 41000 1672
rect 38285 1667 38351 1670
rect 40880 1640 41000 1670
rect 12198 1532 12204 1596
rect 12268 1594 12274 1596
rect 30281 1594 30347 1597
rect 12268 1592 30347 1594
rect 12268 1536 30286 1592
rect 30342 1536 30347 1592
rect 12268 1534 30347 1536
rect 12268 1532 12274 1534
rect 30281 1531 30347 1534
rect 0 1458 120 1488
rect 2589 1458 2655 1461
rect 0 1456 2655 1458
rect 0 1400 2594 1456
rect 2650 1400 2655 1456
rect 0 1398 2655 1400
rect 0 1368 120 1398
rect 2589 1395 2655 1398
rect 9765 1458 9831 1461
rect 30649 1458 30715 1461
rect 9765 1456 30715 1458
rect 9765 1400 9770 1456
rect 9826 1400 30654 1456
rect 30710 1400 30715 1456
rect 9765 1398 30715 1400
rect 9765 1395 9831 1398
rect 30649 1395 30715 1398
rect 38653 1458 38719 1461
rect 40880 1458 41000 1488
rect 38653 1456 41000 1458
rect 38653 1400 38658 1456
rect 38714 1400 41000 1456
rect 38653 1398 41000 1400
rect 38653 1395 38719 1398
rect 40880 1368 41000 1398
rect 3877 1322 3943 1325
rect 37273 1322 37339 1325
rect 3877 1320 37339 1322
rect 3877 1264 3882 1320
rect 3938 1264 37278 1320
rect 37334 1264 37339 1320
rect 3877 1262 37339 1264
rect 3877 1259 3943 1262
rect 37273 1259 37339 1262
rect 7373 1186 7439 1189
rect 38929 1186 38995 1189
rect 7373 1184 38995 1186
rect 7373 1128 7378 1184
rect 7434 1128 38934 1184
rect 38990 1128 38995 1184
rect 7373 1126 38995 1128
rect 7373 1123 7439 1126
rect 38929 1123 38995 1126
rect 5625 1050 5691 1053
rect 21817 1050 21883 1053
rect 5625 1048 21883 1050
rect 5625 992 5630 1048
rect 5686 992 21822 1048
rect 21878 992 21883 1048
rect 5625 990 21883 992
rect 5625 987 5691 990
rect 21817 987 21883 990
rect 3417 914 3483 917
rect 19425 914 19491 917
rect 3417 912 19491 914
rect 3417 856 3422 912
rect 3478 856 19430 912
rect 19486 856 19491 912
rect 3417 854 19491 856
rect 3417 851 3483 854
rect 19425 851 19491 854
rect 3601 778 3667 781
rect 16941 778 17007 781
rect 3601 776 17007 778
rect 3601 720 3606 776
rect 3662 720 16946 776
rect 17002 720 17007 776
rect 3601 718 17007 720
rect 3601 715 3667 718
rect 16941 715 17007 718
rect 3785 642 3851 645
rect 16205 642 16271 645
rect 3785 640 16271 642
rect 3785 584 3790 640
rect 3846 584 16210 640
rect 16266 584 16271 640
rect 3785 582 16271 584
rect 3785 579 3851 582
rect 16205 579 16271 582
<< via3 >>
rect 9996 8740 10060 8804
rect 20668 8740 20732 8804
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 39012 8732 39076 8736
rect 39012 8676 39016 8732
rect 39016 8676 39072 8732
rect 39072 8676 39076 8732
rect 39012 8672 39076 8676
rect 39092 8732 39156 8736
rect 39092 8676 39096 8732
rect 39096 8676 39152 8732
rect 39152 8676 39156 8732
rect 39092 8672 39156 8676
rect 39172 8732 39236 8736
rect 39172 8676 39176 8732
rect 39176 8676 39232 8732
rect 39232 8676 39236 8732
rect 39172 8672 39236 8676
rect 39252 8732 39316 8736
rect 39252 8676 39256 8732
rect 39256 8676 39312 8732
rect 39312 8676 39316 8732
rect 39252 8672 39316 8676
rect 19748 8604 19812 8668
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 20484 8196 20548 8260
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 37952 8188 38016 8192
rect 37952 8132 37956 8188
rect 37956 8132 38012 8188
rect 38012 8132 38016 8188
rect 37952 8128 38016 8132
rect 38032 8188 38096 8192
rect 38032 8132 38036 8188
rect 38036 8132 38092 8188
rect 38092 8132 38096 8188
rect 38032 8128 38096 8132
rect 38112 8188 38176 8192
rect 38112 8132 38116 8188
rect 38116 8132 38172 8188
rect 38172 8132 38176 8188
rect 38112 8128 38176 8132
rect 38192 8188 38256 8192
rect 38192 8132 38196 8188
rect 38196 8132 38252 8188
rect 38252 8132 38256 8188
rect 38192 8128 38256 8132
rect 19564 8060 19628 8124
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 8708 7516 8772 7580
rect 20484 7652 20548 7716
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 39012 7644 39076 7648
rect 39012 7588 39016 7644
rect 39016 7588 39072 7644
rect 39072 7588 39076 7644
rect 39012 7584 39076 7588
rect 39092 7644 39156 7648
rect 39092 7588 39096 7644
rect 39096 7588 39152 7644
rect 39152 7588 39156 7644
rect 39092 7584 39156 7588
rect 39172 7644 39236 7648
rect 39172 7588 39176 7644
rect 39176 7588 39232 7644
rect 39232 7588 39236 7644
rect 39172 7584 39236 7588
rect 39252 7644 39316 7648
rect 39252 7588 39256 7644
rect 39256 7588 39312 7644
rect 39312 7588 39316 7644
rect 39252 7584 39316 7588
rect 12388 7108 12452 7172
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 9996 7032 10060 7036
rect 9996 6976 10010 7032
rect 10010 6976 10060 7032
rect 9996 6972 10060 6976
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 37952 7100 38016 7104
rect 37952 7044 37956 7100
rect 37956 7044 38012 7100
rect 38012 7044 38016 7100
rect 37952 7040 38016 7044
rect 38032 7100 38096 7104
rect 38032 7044 38036 7100
rect 38036 7044 38092 7100
rect 38092 7044 38096 7100
rect 38032 7040 38096 7044
rect 38112 7100 38176 7104
rect 38112 7044 38116 7100
rect 38116 7044 38172 7100
rect 38172 7044 38176 7100
rect 38112 7040 38176 7044
rect 38192 7100 38256 7104
rect 38192 7044 38196 7100
rect 38196 7044 38252 7100
rect 38252 7044 38256 7100
rect 38192 7040 38256 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 39012 6556 39076 6560
rect 39012 6500 39016 6556
rect 39016 6500 39072 6556
rect 39072 6500 39076 6556
rect 39012 6496 39076 6500
rect 39092 6556 39156 6560
rect 39092 6500 39096 6556
rect 39096 6500 39152 6556
rect 39152 6500 39156 6556
rect 39092 6496 39156 6500
rect 39172 6556 39236 6560
rect 39172 6500 39176 6556
rect 39176 6500 39232 6556
rect 39232 6500 39236 6556
rect 39172 6496 39236 6500
rect 39252 6556 39316 6560
rect 39252 6500 39256 6556
rect 39256 6500 39312 6556
rect 39312 6500 39316 6556
rect 39252 6496 39316 6500
rect 19564 6428 19628 6492
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 37952 6012 38016 6016
rect 37952 5956 37956 6012
rect 37956 5956 38012 6012
rect 38012 5956 38016 6012
rect 37952 5952 38016 5956
rect 38032 6012 38096 6016
rect 38032 5956 38036 6012
rect 38036 5956 38092 6012
rect 38092 5956 38096 6012
rect 38032 5952 38096 5956
rect 38112 6012 38176 6016
rect 38112 5956 38116 6012
rect 38116 5956 38172 6012
rect 38172 5956 38176 6012
rect 38112 5952 38176 5956
rect 38192 6012 38256 6016
rect 38192 5956 38196 6012
rect 38196 5956 38252 6012
rect 38252 5956 38256 6012
rect 38192 5952 38256 5956
rect 8708 5612 8772 5676
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 39012 5468 39076 5472
rect 39012 5412 39016 5468
rect 39016 5412 39072 5468
rect 39072 5412 39076 5468
rect 39012 5408 39076 5412
rect 39092 5468 39156 5472
rect 39092 5412 39096 5468
rect 39096 5412 39152 5468
rect 39152 5412 39156 5468
rect 39092 5408 39156 5412
rect 39172 5468 39236 5472
rect 39172 5412 39176 5468
rect 39176 5412 39232 5468
rect 39232 5412 39236 5468
rect 39172 5408 39236 5412
rect 39252 5468 39316 5472
rect 39252 5412 39256 5468
rect 39256 5412 39312 5468
rect 39312 5412 39316 5468
rect 39252 5408 39316 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19748 5340 19812 5404
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 37952 4924 38016 4928
rect 37952 4868 37956 4924
rect 37956 4868 38012 4924
rect 38012 4868 38016 4924
rect 37952 4864 38016 4868
rect 38032 4924 38096 4928
rect 38032 4868 38036 4924
rect 38036 4868 38092 4924
rect 38092 4868 38096 4924
rect 38032 4864 38096 4868
rect 38112 4924 38176 4928
rect 38112 4868 38116 4924
rect 38116 4868 38172 4924
rect 38172 4868 38176 4924
rect 38112 4864 38176 4868
rect 38192 4924 38256 4928
rect 38192 4868 38196 4924
rect 38196 4868 38252 4924
rect 38252 4868 38256 4924
rect 38192 4864 38256 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 39012 4380 39076 4384
rect 39012 4324 39016 4380
rect 39016 4324 39072 4380
rect 39072 4324 39076 4380
rect 39012 4320 39076 4324
rect 39092 4380 39156 4384
rect 39092 4324 39096 4380
rect 39096 4324 39152 4380
rect 39152 4324 39156 4380
rect 39092 4320 39156 4324
rect 39172 4380 39236 4384
rect 39172 4324 39176 4380
rect 39176 4324 39232 4380
rect 39232 4324 39236 4380
rect 39172 4320 39236 4324
rect 39252 4380 39316 4384
rect 39252 4324 39256 4380
rect 39256 4324 39312 4380
rect 39312 4324 39316 4380
rect 39252 4320 39316 4324
rect 20668 4312 20732 4316
rect 20668 4256 20682 4312
rect 20682 4256 20732 4312
rect 20668 4252 20732 4256
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 37952 3836 38016 3840
rect 37952 3780 37956 3836
rect 37956 3780 38012 3836
rect 38012 3780 38016 3836
rect 37952 3776 38016 3780
rect 38032 3836 38096 3840
rect 38032 3780 38036 3836
rect 38036 3780 38092 3836
rect 38092 3780 38096 3836
rect 38032 3776 38096 3780
rect 38112 3836 38176 3840
rect 38112 3780 38116 3836
rect 38116 3780 38172 3836
rect 38172 3780 38176 3836
rect 38112 3776 38176 3780
rect 38192 3836 38256 3840
rect 38192 3780 38196 3836
rect 38196 3780 38252 3836
rect 38252 3780 38256 3836
rect 38192 3776 38256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 39012 3292 39076 3296
rect 39012 3236 39016 3292
rect 39016 3236 39072 3292
rect 39072 3236 39076 3292
rect 39012 3232 39076 3236
rect 39092 3292 39156 3296
rect 39092 3236 39096 3292
rect 39096 3236 39152 3292
rect 39152 3236 39156 3292
rect 39092 3232 39156 3236
rect 39172 3292 39236 3296
rect 39172 3236 39176 3292
rect 39176 3236 39232 3292
rect 39232 3236 39236 3292
rect 39172 3232 39236 3236
rect 39252 3292 39316 3296
rect 39252 3236 39256 3292
rect 39256 3236 39312 3292
rect 39312 3236 39316 3292
rect 39252 3232 39316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 37952 2748 38016 2752
rect 37952 2692 37956 2748
rect 37956 2692 38012 2748
rect 38012 2692 38016 2748
rect 37952 2688 38016 2692
rect 38032 2748 38096 2752
rect 38032 2692 38036 2748
rect 38036 2692 38092 2748
rect 38092 2692 38096 2748
rect 38032 2688 38096 2692
rect 38112 2748 38176 2752
rect 38112 2692 38116 2748
rect 38116 2692 38172 2748
rect 38172 2692 38176 2748
rect 38112 2688 38176 2692
rect 38192 2748 38256 2752
rect 38192 2692 38196 2748
rect 38196 2692 38252 2748
rect 38252 2692 38256 2748
rect 38192 2688 38256 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
rect 39012 2204 39076 2208
rect 39012 2148 39016 2204
rect 39016 2148 39072 2204
rect 39072 2148 39076 2204
rect 39012 2144 39076 2148
rect 39092 2204 39156 2208
rect 39092 2148 39096 2204
rect 39096 2148 39152 2204
rect 39152 2148 39156 2204
rect 39092 2144 39156 2148
rect 39172 2204 39236 2208
rect 39172 2148 39176 2204
rect 39176 2148 39232 2204
rect 39232 2148 39236 2204
rect 39172 2144 39236 2148
rect 39252 2204 39316 2208
rect 39252 2148 39256 2204
rect 39256 2148 39312 2204
rect 39312 2148 39316 2204
rect 39252 2144 39316 2148
rect 12204 1532 12268 1596
<< metal4 >>
rect 1944 8192 2264 11250
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 8736 3324 11250
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11250
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 9004 8736 9324 11250
rect 9995 8804 10061 8805
rect 9995 8740 9996 8804
rect 10060 8740 10061 8804
rect 9995 8739 10061 8740
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 8707 7580 8773 7581
rect 8707 7516 8708 7580
rect 8772 7516 8773 7580
rect 8707 7515 8773 7516
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 8710 5677 8770 7515
rect 9004 6560 9324 7584
rect 9998 7037 10058 8739
rect 13944 8192 14264 11250
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 12387 7172 12453 7173
rect 12387 7108 12388 7172
rect 12452 7170 12453 7172
rect 12452 7110 12634 7170
rect 12452 7108 12453 7110
rect 12387 7107 12453 7108
rect 9995 7036 10061 7037
rect 9995 6972 9996 7036
rect 10060 6972 10061 7036
rect 9995 6971 10061 6972
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 8707 5676 8773 5677
rect 8707 5612 8708 5676
rect 8772 5612 8773 5676
rect 8707 5611 8773 5612
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 12574 2790 12634 7110
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 12206 2730 12634 2790
rect 13944 7104 14264 8128
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 12206 1597 12266 2730
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 12203 1596 12269 1597
rect 12203 1532 12204 1596
rect 12268 1532 12269 1596
rect 12203 1531 12269 1532
rect 13944 0 14264 2688
rect 15004 8736 15324 11250
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 19747 8668 19813 8669
rect 19747 8604 19748 8668
rect 19812 8604 19813 8668
rect 19747 8603 19813 8604
rect 19563 8124 19629 8125
rect 19563 8060 19564 8124
rect 19628 8060 19629 8124
rect 19563 8059 19629 8060
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 19566 6493 19626 8059
rect 19563 6492 19629 6493
rect 19563 6428 19564 6492
rect 19628 6428 19629 6492
rect 19563 6427 19629 6428
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 19750 5405 19810 8603
rect 19944 8192 20264 11250
rect 20667 8804 20733 8805
rect 20667 8740 20668 8804
rect 20732 8740 20733 8804
rect 20667 8739 20733 8740
rect 20483 8260 20549 8261
rect 20483 8196 20484 8260
rect 20548 8196 20549 8260
rect 20483 8195 20549 8196
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 20486 7717 20546 8195
rect 20483 7716 20549 7717
rect 20483 7652 20484 7716
rect 20548 7652 20549 7716
rect 20483 7651 20549 7652
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 19747 5404 19813 5405
rect 19747 5340 19748 5404
rect 19812 5340 19813 5404
rect 19747 5339 19813 5340
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 20670 4317 20730 8739
rect 21004 8736 21324 11250
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 21004 6560 21324 7584
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 20667 4316 20733 4317
rect 20667 4252 20668 4316
rect 20732 4252 20733 4316
rect 20667 4251 20733 4252
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19944 0 20264 2688
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25944 8192 26264 11250
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25944 0 26264 2688
rect 27004 8736 27324 11250
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 31944 8192 32264 11250
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 0 32264 2688
rect 33004 8736 33324 11250
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
rect 37944 8192 38264 11250
rect 37944 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38264 8192
rect 37944 7104 38264 8128
rect 37944 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38264 7104
rect 37944 6016 38264 7040
rect 37944 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38264 6016
rect 37944 4928 38264 5952
rect 37944 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38264 4928
rect 37944 3840 38264 4864
rect 37944 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38264 3840
rect 37944 2752 38264 3776
rect 37944 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38264 2752
rect 37944 0 38264 2688
rect 39004 8736 39324 11250
rect 39004 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39324 8736
rect 39004 7648 39324 8672
rect 39004 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39324 7648
rect 39004 6560 39324 7584
rect 39004 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39324 6560
rect 39004 5472 39324 6496
rect 39004 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39324 5472
rect 39004 4384 39324 5408
rect 39004 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39324 4384
rect 39004 3296 39324 4320
rect 39004 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39324 3296
rect 39004 2208 39324 3232
rect 39004 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39324 2208
rect 39004 0 39324 2144
use sky130_fd_sc_hd__mux4_1  _000_
timestamp -3599
transform 1 0 11960 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _001_
timestamp -3599
transform 1 0 31648 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _002_
timestamp -3599
transform 1 0 6348 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _003_
timestamp -3599
transform 1 0 19964 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _004_
timestamp -3599
transform 1 0 22356 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _005_
timestamp -3599
transform 1 0 31740 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _006_
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _007_
timestamp -3599
transform 1 0 17204 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _008_
timestamp -3599
transform 1 0 14260 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _009_
timestamp -3599
transform -1 0 30912 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _010_
timestamp -3599
transform -1 0 5428 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _011_
timestamp -3599
transform -1 0 9936 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _012_
timestamp -3599
transform 1 0 22356 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _013_
timestamp -3599
transform -1 0 32200 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _014_
timestamp -3599
transform 1 0 9476 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _015_
timestamp -3599
transform 1 0 19320 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _016_
timestamp -3599
transform -1 0 20148 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _017_
timestamp -3599
transform 1 0 11500 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _018_
timestamp -3599
transform -1 0 31740 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _019_
timestamp -3599
transform 1 0 17112 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _020_
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _021_
timestamp -3599
transform 1 0 2852 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _022_
timestamp -3599
transform 1 0 29532 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _023_
timestamp -3599
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _024_
timestamp -3599
transform 1 0 17296 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _025_
timestamp -3599
transform 1 0 17756 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _026_
timestamp -3599
transform 1 0 35052 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _027_
timestamp -3599
transform 1 0 25576 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _028_
timestamp -3599
transform 1 0 20608 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _029_
timestamp -3599
transform 1 0 6164 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _030_
timestamp -3599
transform 1 0 32108 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _031_
timestamp -3599
transform 1 0 11408 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _032_
timestamp -3599
transform 1 0 18676 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _033_
timestamp -3599
transform -1 0 11684 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _034_
timestamp -3599
transform 1 0 30452 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _035_
timestamp -3599
transform 1 0 23000 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _036_
timestamp -3599
transform 1 0 5428 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _037_
timestamp -3599
transform 1 0 2668 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _038_
timestamp -3599
transform 1 0 28612 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _039_
timestamp -3599
transform 1 0 12328 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _040_
timestamp -3599
transform 1 0 16376 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _041_
timestamp -3599
transform 1 0 17020 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _042_
timestamp -3599
transform 1 0 35880 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _043_
timestamp -3599
transform 1 0 24932 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _044_
timestamp -3599
transform -1 0 20700 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _045_
timestamp -3599
transform 1 0 5336 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _046_
timestamp -3599
transform 1 0 31096 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _047_
timestamp -3599
transform 1 0 12236 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _048_
timestamp -3599
transform -1 0 15272 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _049_
timestamp -3599
transform 1 0 15640 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _050_
timestamp -3599
transform -1 0 36064 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _051_
timestamp -3599
transform 1 0 25852 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _052_
timestamp -3599
transform 1 0 18124 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _053_
timestamp -3599
transform 1 0 8464 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _054_
timestamp -3599
transform 1 0 32200 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _055_
timestamp -3599
transform 1 0 13984 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _056_
timestamp -3599
transform -1 0 20608 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _057_
timestamp -3599
transform -1 0 11408 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _058_
timestamp -3599
transform -1 0 30912 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _059_
timestamp -3599
transform -1 0 24196 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _060_
timestamp -3599
transform 1 0 20332 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _061_
timestamp -3599
transform 1 0 6992 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _062_
timestamp -3599
transform 1 0 30176 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _063_
timestamp -3599
transform -1 0 12972 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _064_
timestamp -3599
transform 1 0 18032 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _065_
timestamp -3599
transform 1 0 9292 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _066_
timestamp -3599
transform 1 0 30268 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _067_
timestamp -3599
transform 1 0 12052 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dlxtp_1  _068_
timestamp -3599
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _069_
timestamp -3599
transform 1 0 9936 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _070_
timestamp -3599
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _071_
timestamp -3599
transform 1 0 26404 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _072_
timestamp -3599
transform -1 0 23828 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _073_
timestamp -3599
transform -1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _074_
timestamp -3599
transform 1 0 15456 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _075_
timestamp -3599
transform 1 0 16928 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _076_
timestamp -3599
transform -1 0 13064 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _077_
timestamp -3599
transform 1 0 29624 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _078_
timestamp -3599
transform 1 0 5888 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _079_
timestamp -3599
transform 1 0 19412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _080_
timestamp -3599
transform -1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _081_
timestamp -3599
transform 1 0 29900 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _082_
timestamp -3599
transform -1 0 17204 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _083_
timestamp -3599
transform -1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _084_
timestamp -3599
transform -1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _085_
timestamp -3599
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _086_
timestamp -3599
transform 1 0 7268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _087_
timestamp -3599
transform 1 0 6716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _088_
timestamp -3599
transform 1 0 24748 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _089_
timestamp -3599
transform 1 0 34500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _090_
timestamp -3599
transform 1 0 14536 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _091_
timestamp -3599
transform 1 0 13156 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _092_
timestamp -3599
transform -1 0 15824 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _093_
timestamp -3599
transform 1 0 20792 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _094_
timestamp -3599
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _095_
timestamp -3599
transform 1 0 19688 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _096_
timestamp -3599
transform 1 0 24748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _097_
timestamp -3599
transform 1 0 34868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _098_
timestamp -3599
transform -1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _099_
timestamp -3599
transform -1 0 23368 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _100_
timestamp -3599
transform 1 0 7728 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _101_
timestamp -3599
transform 1 0 9108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _102_
timestamp -3599
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _103_
timestamp -3599
transform 1 0 3864 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _104_
timestamp -3599
transform -1 0 24564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _105_
timestamp -3599
transform 1 0 27232 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _106_
timestamp -3599
transform -1 0 13616 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _107_
timestamp -3599
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _108_
timestamp -3599
transform 1 0 10212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _109_
timestamp -3599
transform 1 0 30728 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _110_
timestamp -3599
transform 1 0 4876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _111_
timestamp -3599
transform 1 0 19504 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _112_
timestamp -3599
transform 1 0 24472 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _113_
timestamp -3599
transform 1 0 33764 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _114_
timestamp -3599
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _115_
timestamp -3599
transform -1 0 23460 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _116_
timestamp -3599
transform 1 0 10396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _117_
timestamp -3599
transform 1 0 27232 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _118_
timestamp -3599
transform 1 0 2024 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _119_
timestamp -3599
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _120_
timestamp -3599
transform 1 0 15824 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _121_
timestamp -3599
transform -1 0 34040 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _122_
timestamp -3599
transform -1 0 13524 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _123_
timestamp -3599
transform 1 0 13892 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _124_
timestamp -3599
transform 1 0 15824 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _125_
timestamp -3599
transform -1 0 22356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _126_
timestamp -3599
transform 1 0 6624 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _127_
timestamp -3599
transform -1 0 20424 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _128_
timestamp -3599
transform 1 0 25944 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _129_
timestamp -3599
transform 1 0 29348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _130_
timestamp -3599
transform 1 0 21988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _131_
timestamp -3599
transform 1 0 22172 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _132_
timestamp -3599
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _133_
timestamp -3599
transform 1 0 7728 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _134_
timestamp -3599
transform -1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _135_
timestamp -3599
transform -1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _136_
timestamp -3599
transform 1 0 27508 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _137_
timestamp -3599
transform 1 0 27876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _138_
timestamp -3599
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _139_
timestamp -3599
transform 1 0 14352 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _140_
timestamp -3599
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _141_
timestamp -3599
transform -1 0 29440 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _142_
timestamp -3599
transform 1 0 7176 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _143_
timestamp -3599
transform 1 0 8372 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _144_
timestamp -3599
transform 1 0 28520 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _145_
timestamp -3599
transform 1 0 30912 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _146_
timestamp -3599
transform -1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _147_
timestamp -3599
transform 1 0 22356 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _148_
timestamp -3599
transform 1 0 19228 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _149_
timestamp -3599
transform -1 0 27416 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _150_
timestamp -3599
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _151_
timestamp -3599
transform 1 0 6256 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _152_
timestamp -3599
transform 1 0 25208 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _153_
timestamp -3599
transform -1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _154_
timestamp -3599
transform -1 0 13248 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _155_
timestamp -3599
transform 1 0 10304 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _157_
timestamp -3599
transform 1 0 15640 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _158_
timestamp -3599
transform 1 0 21068 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _160_
timestamp -3599
transform 1 0 19412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _161_
timestamp -3599
transform 1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp -3599
transform -1 0 33764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _163_
timestamp -3599
transform 1 0 22080 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _164_
timestamp -3599
transform 1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _165_
timestamp -3599
transform 1 0 7636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp -3599
transform 1 0 8280 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _167_
timestamp -3599
transform 1 0 27048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _168_
timestamp -3599
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _169_
timestamp -3599
transform 1 0 27324 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _170_
timestamp -3599
transform 1 0 27416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _171_
timestamp -3599
transform 1 0 13156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp -3599
transform -1 0 16928 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _173_
timestamp -3599
transform 1 0 10396 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _174_
timestamp -3599
transform -1 0 30084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _175_
timestamp -3599
transform 1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _176_
timestamp -3599
transform 1 0 9016 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _177_
timestamp -3599
transform 1 0 28980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp -3599
transform -1 0 33948 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _179_
timestamp -3599
transform 1 0 22908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _180_
timestamp -3599
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _181_
timestamp -3599
transform 1 0 10672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _182_
timestamp -3599
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _183_
timestamp -3599
transform 1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp -3599
transform 1 0 4324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _185_
timestamp -3599
transform 1 0 25116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _186_
timestamp -3599
transform -1 0 35236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _187_
timestamp -3599
transform 1 0 13524 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp -3599
transform 1 0 10580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _189_
timestamp -3599
transform -1 0 31280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp -3599
transform 1 0 34040 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _191_
timestamp -3599
transform 1 0 34684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp -3599
transform 1 0 38180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp -3599
transform 1 0 38548 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp -3599
transform 1 0 37444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp -3599
transform 1 0 38180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp -3599
transform 1 0 35052 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp -3599
transform 1 0 37996 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp -3599
transform -1 0 35604 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp -3599
transform 1 0 38548 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp -3599
transform 1 0 35972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp -3599
transform 1 0 38272 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp -3599
transform 1 0 37352 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _203_
timestamp -3599
transform -1 0 37352 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp -3599
transform -1 0 34408 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp -3599
transform 1 0 38180 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _206_
timestamp -3599
transform -1 0 35604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _207_
timestamp -3599
transform 1 0 38548 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _208_
timestamp -3599
transform -1 0 37904 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _209_
timestamp -3599
transform 1 0 15180 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _210_
timestamp -3599
transform -1 0 32476 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _211_
timestamp -3599
transform 1 0 10948 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _212_
timestamp -3599
transform -1 0 20240 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp -3599
transform 1 0 12972 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _214_
timestamp -3599
transform -1 0 30636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _215_
timestamp -3599
transform 1 0 6440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _216_
timestamp -3599
transform -1 0 19964 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _217_
timestamp -3599
transform -1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _218_
timestamp -3599
transform -1 0 31372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp -3599
transform 1 0 11684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _220_
timestamp -3599
transform -1 0 20884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp -3599
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _222_
timestamp -3599
transform -1 0 32384 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp -3599
transform 1 0 8096 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _224_
timestamp -3599
transform -1 0 18124 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _225_
timestamp -3599
transform -1 0 25392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _226_
timestamp -3599
transform -1 0 35972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _227_
timestamp -3599
transform -1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _228_
timestamp -3599
transform 1 0 15272 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _229_
timestamp -3599
transform 1 0 11592 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _230_
timestamp -3599
transform -1 0 31464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _231_
timestamp -3599
transform -1 0 4876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _232_
timestamp -3599
transform -1 0 21252 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _233_
timestamp -3599
transform -1 0 24932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _234_
timestamp -3599
transform -1 0 35788 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _235_
timestamp -3599
transform -1 0 17480 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _236_
timestamp -3599
transform 1 0 16100 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _237_
timestamp -3599
transform 1 0 11224 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _238_
timestamp -3599
transform -1 0 28980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _239_
timestamp -3599
transform 1 0 2392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp -3599
transform -1 0 5796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _241_
timestamp -3599
transform 1 0 22080 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _242_
timestamp -3599
transform -1 0 30544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _243_
timestamp -3599
transform -1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _244_
timestamp -3599
transform 1 0 18400 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _245_
timestamp -3599
transform -1 0 11408 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _246_
timestamp -3599
transform -1 0 32660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _247_
timestamp -3599
transform 1 0 4968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _248_
timestamp -3599
transform 1 0 20700 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _249_
timestamp -3599
transform -1 0 25208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _250_
timestamp -3599
transform -1 0 35052 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _251_
timestamp -3599
transform 1 0 17572 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp -3599
transform 1 0 16744 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _253_
timestamp -3599
transform -1 0 11776 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _254_
timestamp -3599
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _255_
timestamp -3599
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp -3599
transform -1 0 5428 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _257_
timestamp -3599
transform 1 0 17020 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _258_
timestamp -3599
transform -1 0 31556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _259_
timestamp -3599
transform 1 0 9200 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp -3599
transform 1 0 20148 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _261_
timestamp -3599
transform 1 0 37536 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform 1 0 39008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform -1 0 38180 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform -1 0 13616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform -1 0 6624 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  fanout35
timestamp -3599
transform 1 0 26036 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp -3599
transform 1 0 28152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout37
timestamp -3599
transform 1 0 28888 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout38
timestamp -3599
transform 1 0 7820 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout39
timestamp -3599
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp -3599
transform 1 0 26128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout41
timestamp -3599
transform 1 0 33120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout42
timestamp -3599
transform 1 0 9936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout43
timestamp -3599
transform 1 0 6440 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp -3599
transform 1 0 29072 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout45
timestamp -3599
transform 1 0 27876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23
timestamp -3599
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72
timestamp -3599
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp -3599
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp -3599
transform 1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94
timestamp -3599
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp -3599
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119
timestamp -3599
transform 1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_126
timestamp -3599
transform 1 0 12696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_130
timestamp -3599
transform 1 0 13064 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135
timestamp -3599
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp -3599
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp -3599
transform 1 0 14444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp -3599
transform 1 0 14996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_159
timestamp -3599
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp -3599
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_186
timestamp -3599
transform 1 0 18216 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_191
timestamp -3599
transform 1 0 18676 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_197
timestamp -3599
transform 1 0 19228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_210
timestamp -3599
transform 1 0 20424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp -3599
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp -3599
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp -3599
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_257
timestamp 1636964856
transform 1 0 24748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_269
timestamp -3599
transform 1 0 25852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -3599
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636964856
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636964856
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -3599
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_309
timestamp -3599
transform 1 0 29532 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_320
timestamp -3599
transform 1 0 30544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp -3599
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_337
timestamp -3599
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_345
timestamp -3599
transform 1 0 32844 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_352
timestamp 1636964856
transform 1 0 33488 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1636964856
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1636964856
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp -3599
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_393
timestamp -3599
transform 1 0 37260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_397
timestamp -3599
transform 1 0 37628 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_17
timestamp -3599
transform 1 0 2668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_32
timestamp -3599
transform 1 0 4048 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp -3599
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_72
timestamp 1636964856
transform 1 0 7728 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_84
timestamp -3599
transform 1 0 8832 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_122
timestamp -3599
transform 1 0 12328 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_139
timestamp -3599
transform 1 0 13892 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_145
timestamp -3599
transform 1 0 14444 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -3599
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_190
timestamp -3599
transform 1 0 18584 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_198
timestamp -3599
transform 1 0 19320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_214
timestamp -3599
transform 1 0 20792 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp -3599
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_240
timestamp 1636964856
transform 1 0 23184 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_252
timestamp -3599
transform 1 0 24288 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_256
timestamp -3599
transform 1 0 24656 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp -3599
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp -3599
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_285
timestamp -3599
transform 1 0 27324 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_289
timestamp 1636964856
transform 1 0 27692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_301
timestamp -3599
transform 1 0 28796 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp -3599
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp -3599
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_337
timestamp -3599
transform 1 0 32108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_345
timestamp -3599
transform 1 0 32844 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636964856
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636964856
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp -3599
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp -3599
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp -3599
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_401
timestamp -3599
transform 1 0 37996 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636964856
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_41
timestamp -3599
transform 1 0 4876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_45
timestamp -3599
transform 1 0 5244 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_64
timestamp -3599
transform 1 0 6992 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp -3599
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_121
timestamp -3599
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp -3599
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636964856
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_156
timestamp -3599
transform 1 0 15456 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_162
timestamp -3599
transform 1 0 16008 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_178
timestamp -3599
transform 1 0 17480 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_182
timestamp 1636964856
transform 1 0 17848 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp -3599
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_197
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_210
timestamp 1636964856
transform 1 0 20424 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_222
timestamp -3599
transform 1 0 21528 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_231
timestamp -3599
transform 1 0 22356 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp -3599
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp -3599
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636964856
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_265
timestamp -3599
transform 1 0 25484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_269
timestamp -3599
transform 1 0 25852 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_282
timestamp -3599
transform 1 0 27048 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_296
timestamp -3599
transform 1 0 28336 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp -3599
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_309
timestamp -3599
transform 1 0 29532 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_338
timestamp 1636964856
transform 1 0 32200 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_350
timestamp 1636964856
transform 1 0 33304 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp -3599
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_371
timestamp -3599
transform 1 0 35236 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_382
timestamp 1636964856
transform 1 0 36248 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_394
timestamp 1636964856
transform 1 0 37352 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_406
timestamp -3599
transform 1 0 38456 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_10
timestamp -3599
transform 1 0 2024 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp -3599
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -3599
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_78
timestamp -3599
transform 1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp -3599
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636964856
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_125
timestamp -3599
transform 1 0 12604 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_134
timestamp -3599
transform 1 0 13432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_138
timestamp -3599
transform 1 0 13800 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_151
timestamp -3599
transform 1 0 14996 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_157
timestamp -3599
transform 1 0 15548 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp -3599
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -3599
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636964856
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_181
timestamp -3599
transform 1 0 17756 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_187
timestamp -3599
transform 1 0 18308 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_200
timestamp -3599
transform 1 0 19504 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_215
timestamp -3599
transform 1 0 20884 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp -3599
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_249
timestamp -3599
transform 1 0 24012 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_255
timestamp -3599
transform 1 0 24564 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_268
timestamp 1636964856
transform 1 0 25760 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636964856
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_305
timestamp -3599
transform 1 0 29164 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_313
timestamp -3599
transform 1 0 29900 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636964856
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_349
timestamp -3599
transform 1 0 33212 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_379
timestamp 1636964856
transform 1 0 35972 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp -3599
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_393
timestamp -3599
transform 1 0 37260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_400
timestamp -3599
transform 1 0 37904 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_408
timestamp -3599
transform 1 0 38640 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_22
timestamp -3599
transform 1 0 3128 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_41
timestamp -3599
transform 1 0 4876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_49
timestamp -3599
transform 1 0 5612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_73
timestamp -3599
transform 1 0 7820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_79
timestamp -3599
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -3599
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636964856
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_97
timestamp -3599
transform 1 0 10028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_110
timestamp -3599
transform 1 0 11224 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_118
timestamp -3599
transform 1 0 11960 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_132
timestamp -3599
transform 1 0 13248 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_141
timestamp -3599
transform 1 0 14076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_147
timestamp -3599
transform 1 0 14628 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_172
timestamp -3599
transform 1 0 16928 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_176
timestamp -3599
transform 1 0 17296 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp -3599
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp -3599
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_197
timestamp -3599
transform 1 0 19228 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_253
timestamp -3599
transform 1 0 24380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_275
timestamp -3599
transform 1 0 26404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_281
timestamp -3599
transform 1 0 26956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_288
timestamp -3599
transform 1 0 27600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp -3599
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_309
timestamp -3599
transform 1 0 29532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_329
timestamp -3599
transform 1 0 31372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp -3599
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp -3599
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_365
timestamp -3599
transform 1 0 34684 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_387
timestamp 1636964856
transform 1 0 36708 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_399
timestamp -3599
transform 1 0 37812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_403
timestamp -3599
transform 1 0 38180 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636964856
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_39
timestamp -3599
transform 1 0 4692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_43
timestamp -3599
transform 1 0 5060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp -3599
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_61
timestamp -3599
transform 1 0 6716 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_91
timestamp -3599
transform 1 0 9476 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_95
timestamp -3599
transform 1 0 9844 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp -3599
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_117
timestamp -3599
transform 1 0 11868 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_139
timestamp -3599
transform 1 0 13892 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_143
timestamp -3599
transform 1 0 14260 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_208
timestamp -3599
transform 1 0 20240 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_216
timestamp -3599
transform 1 0 20976 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp -3599
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp -3599
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_243
timestamp 1636964856
transform 1 0 23460 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_255
timestamp -3599
transform 1 0 24564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_262
timestamp -3599
transform 1 0 25208 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_270
timestamp -3599
transform 1 0 25944 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_275
timestamp -3599
transform 1 0 26404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp -3599
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_293
timestamp -3599
transform 1 0 28060 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_310
timestamp 1636964856
transform 1 0 29624 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_322
timestamp 1636964856
transform 1 0 30728 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp -3599
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_341
timestamp 1636964856
transform 1 0 32476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_353
timestamp 1636964856
transform 1 0 33580 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_365
timestamp -3599
transform 1 0 34684 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_373
timestamp -3599
transform 1 0 35420 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_377
timestamp 1636964856
transform 1 0 35788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_389
timestamp -3599
transform 1 0 36892 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636964856
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp -3599
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_12
timestamp 1636964856
transform 1 0 2208 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp -3599
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_45
timestamp -3599
transform 1 0 5244 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_53
timestamp -3599
transform 1 0 5980 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_68
timestamp 1636964856
transform 1 0 7360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp -3599
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp -3599
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_90
timestamp -3599
transform 1 0 9384 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_98
timestamp -3599
transform 1 0 10120 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_105
timestamp -3599
transform 1 0 10764 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_130
timestamp -3599
transform 1 0 13064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp -3599
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636964856
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636964856
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636964856
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp -3599
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp -3599
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636964856
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_209
timestamp -3599
transform 1 0 20332 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp -3599
transform 1 0 20700 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_226
timestamp 1636964856
transform 1 0 21896 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_238
timestamp 1636964856
transform 1 0 23000 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp -3599
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_265
timestamp -3599
transform 1 0 25484 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_273
timestamp -3599
transform 1 0 26220 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_309
timestamp -3599
transform 1 0 29532 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_347
timestamp 1636964856
transform 1 0 33028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_359
timestamp -3599
transform 1 0 34132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp -3599
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_365
timestamp -3599
transform 1 0 34684 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_380
timestamp 1636964856
transform 1 0 36064 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_392
timestamp -3599
transform 1 0 37168 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_400
timestamp -3599
transform 1 0 37904 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_404
timestamp -3599
transform 1 0 38272 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_10
timestamp 1636964856
transform 1 0 2024 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_22
timestamp -3599
transform 1 0 3128 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_26
timestamp -3599
transform 1 0 3496 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_31
timestamp -3599
transform 1 0 3956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp -3599
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -3599
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_77
timestamp -3599
transform 1 0 8188 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_82
timestamp -3599
transform 1 0 8648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_86
timestamp -3599
transform 1 0 9016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp -3599
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp -3599
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_117
timestamp -3599
transform 1 0 11868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_130
timestamp -3599
transform 1 0 13064 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp -3599
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_181
timestamp -3599
transform 1 0 17756 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_194
timestamp -3599
transform 1 0 18952 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_202
timestamp -3599
transform 1 0 19688 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp -3599
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp -3599
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_225
timestamp -3599
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_255
timestamp -3599
transform 1 0 24564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp -3599
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp -3599
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_299
timestamp -3599
transform 1 0 28612 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_324
timestamp -3599
transform 1 0 30912 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp -3599
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_340
timestamp -3599
transform 1 0 32384 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_348
timestamp -3599
transform 1 0 33120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_361
timestamp -3599
transform 1 0 34316 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_379
timestamp 1636964856
transform 1 0 35972 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp -3599
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1636964856
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp -3599
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_13
timestamp 1636964856
transform 1 0 2300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp -3599
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_42
timestamp -3599
transform 1 0 4968 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_51
timestamp -3599
transform 1 0 5796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_57
timestamp -3599
transform 1 0 6348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_62
timestamp -3599
transform 1 0 6808 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_70
timestamp -3599
transform 1 0 7544 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_89
timestamp -3599
transform 1 0 9292 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_94
timestamp -3599
transform 1 0 9752 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_107
timestamp -3599
transform 1 0 10948 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_116
timestamp -3599
transform 1 0 11776 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_132
timestamp -3599
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp -3599
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_154
timestamp -3599
transform 1 0 15272 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_162
timestamp -3599
transform 1 0 16008 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp -3599
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_221
timestamp -3599
transform 1 0 21436 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_229
timestamp -3599
transform 1 0 22172 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_242
timestamp -3599
transform 1 0 23368 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp -3599
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_253
timestamp -3599
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_264
timestamp 1636964856
transform 1 0 25392 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_276
timestamp 1636964856
transform 1 0 26496 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_288
timestamp -3599
transform 1 0 27600 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_296
timestamp -3599
transform 1 0 28336 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_302
timestamp -3599
transform 1 0 28888 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_321
timestamp -3599
transform 1 0 30636 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_330
timestamp -3599
transform 1 0 31464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_353
timestamp -3599
transform 1 0 33580 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_361
timestamp -3599
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1636964856
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1636964856
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_389
timestamp -3599
transform 1 0 36892 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_400
timestamp -3599
transform 1 0 37904 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_23
timestamp 1636964856
transform 1 0 3220 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_35
timestamp -3599
transform 1 0 4324 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_43
timestamp -3599
transform 1 0 5060 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_70
timestamp -3599
transform 1 0 7544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_139
timestamp -3599
transform 1 0 13892 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_149
timestamp -3599
transform 1 0 14812 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_157
timestamp -3599
transform 1 0 15548 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_161
timestamp -3599
transform 1 0 15916 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp -3599
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_169
timestamp -3599
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp -3599
transform 1 0 18400 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_211
timestamp -3599
transform 1 0 20516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_219
timestamp -3599
transform 1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp -3599
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_225
timestamp -3599
transform 1 0 21804 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_241
timestamp -3599
transform 1 0 23276 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_251
timestamp -3599
transform 1 0 24196 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_259
timestamp -3599
transform 1 0 24932 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_264
timestamp 1636964856
transform 1 0 25392 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp -3599
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_296
timestamp -3599
transform 1 0 28336 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_300
timestamp -3599
transform 1 0 28704 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_308
timestamp -3599
transform 1 0 29440 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_315
timestamp -3599
transform 1 0 30084 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp -3599
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_346
timestamp 1636964856
transform 1 0 32936 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_358
timestamp 1636964856
transform 1 0 34040 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_370
timestamp -3599
transform 1 0 35144 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_375
timestamp 1636964856
transform 1 0 35604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_387
timestamp -3599
transform 1 0 36708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp -3599
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp -3599
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_37
timestamp -3599
transform 1 0 4508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_43
timestamp -3599
transform 1 0 5060 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_49
timestamp -3599
transform 1 0 5612 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_113
timestamp -3599
transform 1 0 11500 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_172
timestamp -3599
transform 1 0 16928 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp -3599
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_226
timestamp -3599
transform 1 0 21896 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_289
timestamp -3599
transform 1 0 27692 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_295
timestamp -3599
transform 1 0 28244 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_309
timestamp -3599
transform 1 0 29532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_352
timestamp -3599
transform 1 0 33488 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_358
timestamp -3599
transform 1 0 34040 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp -3599
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_379
timestamp -3599
transform 1 0 35972 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_385
timestamp -3599
transform 1 0 36524 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_397
timestamp -3599
transform 1 0 37628 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_23
timestamp -3599
transform 1 0 3220 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_81
timestamp -3599
transform 1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp -3599
transform 1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_218
timestamp -3599
transform 1 0 21160 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp -3599
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_237
timestamp -3599
transform 1 0 22908 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_250
timestamp -3599
transform 1 0 24104 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp -3599
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_363
timestamp -3599
transform 1 0 34500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp -3599
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_409
timestamp -3599
transform 1 0 38732 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp -3599
transform 1 0 3496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp -3599
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input6
timestamp -3599
transform 1 0 1932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp -3599
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp -3599
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp -3599
transform -1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp -3599
transform 1 0 2300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp -3599
transform 1 0 2852 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp -3599
transform 1 0 2116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp -3599
transform 1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp -3599
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp -3599
transform 1 0 2300 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input19
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp -3599
transform 1 0 3036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp -3599
transform 1 0 2668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp -3599
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input23
timestamp -3599
transform 1 0 3772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp -3599
transform 1 0 2300 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input26
timestamp -3599
transform 1 0 3220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp -3599
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input29
timestamp -3599
transform 1 0 2576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input31
timestamp -3599
transform 1 0 1748 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp -3599
transform 1 0 1748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp -3599
transform -1 0 2576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp -3599
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input36
timestamp -3599
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp -3599
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp -3599
transform -1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp -3599
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input40
timestamp -3599
transform 1 0 12420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp -3599
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp -3599
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp -3599
transform -1 0 4876 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input44
timestamp -3599
transform -1 0 4600 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp -3599
transform 1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input46
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp -3599
transform -1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp -3599
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp -3599
transform 1 0 18124 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp -3599
transform -1 0 18216 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp -3599
transform 1 0 18216 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp -3599
transform -1 0 19136 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input53
timestamp -3599
transform -1 0 21528 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp -3599
transform -1 0 22080 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input55
timestamp -3599
transform 1 0 22080 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input56
timestamp -3599
transform 1 0 22356 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp -3599
transform 1 0 23828 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp -3599
transform -1 0 24656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input59
timestamp -3599
transform 1 0 24656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp -3599
transform -1 0 25208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp -3599
transform -1 0 18216 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input62
timestamp -3599
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input63
timestamp -3599
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp -3599
transform -1 0 19412 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp -3599
transform -1 0 19688 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp -3599
transform -1 0 21252 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp -3599
transform 1 0 20700 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp -3599
transform -1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp -3599
transform 1 0 25208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input70
timestamp -3599
transform 1 0 27508 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp -3599
transform 1 0 27784 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp -3599
transform -1 0 27692 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp -3599
transform -1 0 28336 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp -3599
transform -1 0 28612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input75
timestamp -3599
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input76
timestamp -3599
transform -1 0 25760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input77
timestamp -3599
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp -3599
transform 1 0 24932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input79
timestamp -3599
transform -1 0 26036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input80
timestamp -3599
transform -1 0 26312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp -3599
transform -1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input82
timestamp -3599
transform -1 0 26864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input83
timestamp -3599
transform -1 0 27232 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input84
timestamp -3599
transform -1 0 27508 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input85
timestamp -3599
transform -1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp -3599
transform -1 0 31556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input87
timestamp -3599
transform -1 0 31832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input88
timestamp -3599
transform -1 0 32384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input89
timestamp -3599
transform 1 0 32108 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp -3599
transform 1 0 32660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input91
timestamp -3599
transform -1 0 33212 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input92
timestamp -3599
transform -1 0 29440 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp -3599
transform -1 0 28704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input94
timestamp -3599
transform -1 0 30728 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input95
timestamp -3599
transform -1 0 31004 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input96
timestamp -3599
transform 1 0 29532 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp -3599
transform 1 0 31004 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input98
timestamp -3599
transform -1 0 31556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input99
timestamp -3599
transform -1 0 31832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input100
timestamp -3599
transform -1 0 32108 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform 1 0 38456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform 1 0 39192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform 1 0 38824 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform 1 0 39192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp -3599
transform 1 0 38824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp -3599
transform 1 0 39192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp -3599
transform 1 0 38824 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp -3599
transform 1 0 39192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp -3599
transform 1 0 38824 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp -3599
transform 1 0 38456 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp -3599
transform 1 0 39192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp -3599
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp -3599
transform 1 0 37720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp -3599
transform 1 0 39192 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp -3599
transform 1 0 38824 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp -3599
transform 1 0 39192 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp -3599
transform 1 0 39192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp -3599
transform 1 0 38824 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp -3599
transform 1 0 38456 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp -3599
transform 1 0 39192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp -3599
transform 1 0 39192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp -3599
transform 1 0 38456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp -3599
transform 1 0 37720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp -3599
transform 1 0 38824 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp -3599
transform 1 0 38088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp -3599
transform 1 0 38824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp -3599
transform 1 0 38456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp -3599
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp -3599
transform 1 0 39192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp -3599
transform 1 0 38824 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp -3599
transform 1 0 39192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp -3599
transform 1 0 38824 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp -3599
transform 1 0 33028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp -3599
transform -1 0 36524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp -3599
transform -1 0 35972 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp -3599
transform -1 0 36892 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp -3599
transform -1 0 36524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp -3599
transform 1 0 37260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp -3599
transform 1 0 36708 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp -3599
transform -1 0 37996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp -3599
transform 1 0 37996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp -3599
transform -1 0 38732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp -3599
transform 1 0 37812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp -3599
transform -1 0 33764 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp -3599
transform -1 0 34132 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp -3599
transform -1 0 34500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp -3599
transform -1 0 34040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp -3599
transform -1 0 35052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp -3599
transform -1 0 35420 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp -3599
transform -1 0 35052 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp -3599
transform -1 0 35788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp -3599
transform 1 0 35788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp -3599
transform -1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp -3599
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp -3599
transform -1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp -3599
transform -1 0 21620 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp -3599
transform 1 0 23092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp -3599
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp -3599
transform -1 0 24196 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp -3599
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp -3599
transform -1 0 14996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp -3599
transform -1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp -3599
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp -3599
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp -3599
transform -1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp -3599
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp -3599
transform -1 0 19136 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp -3599
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp -3599
transform -1 0 3680 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp -3599
transform -1 0 4140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp -3599
transform -1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp -3599
transform -1 0 4508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp -3599
transform -1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp -3599
transform -1 0 5060 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp -3599
transform -1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp -3599
transform -1 0 5612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp -3599
transform -1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp -3599
transform -1 0 6072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp -3599
transform -1 0 5520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp -3599
transform -1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp -3599
transform -1 0 6440 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp -3599
transform -1 0 6256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp -3599
transform -1 0 7544 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp -3599
transform 1 0 6624 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp -3599
transform -1 0 7360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp -3599
transform -1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp -3599
transform -1 0 7728 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp -3599
transform -1 0 7084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp -3599
transform -1 0 9292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp -3599
transform 1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp -3599
transform 1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp -3599
transform -1 0 11408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp -3599
transform -1 0 12052 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp -3599
transform 1 0 13156 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp -3599
transform -1 0 11960 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp -3599
transform -1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp -3599
transform 1 0 9384 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp -3599
transform -1 0 10672 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp -3599
transform -1 0 10304 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp -3599
transform -1 0 9568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp -3599
transform -1 0 10396 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp -3599
transform -1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp -3599
transform -1 0 11408 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp -3599
transform -1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp -3599
transform 1 0 11960 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp -3599
transform 1 0 16008 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp -3599
transform 1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp -3599
transform -1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp -3599
transform -1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp -3599
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp -3599
transform -1 0 17296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp -3599
transform -1 0 13892 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp -3599
transform 1 0 12328 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp -3599
transform -1 0 13064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp -3599
transform -1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp -3599
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp -3599
transform -1 0 15272 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp -3599
transform -1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp -3599
transform 1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp -3599
transform -1 0 15824 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output221
timestamp -3599
transform -1 0 33488 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 39836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 39836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 39836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 39836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 39836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 39836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 39836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 39836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 39836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 39836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  S_CPU_IF_222
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_38
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -3599
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_45
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_48
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_49
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_50
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -3599
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_52
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_53
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_54
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_55
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_56
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_57
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_58
timestamp -3599
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_59
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_60
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_61
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_62
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_63
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_65
timestamp -3599
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_66
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_67
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_68
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_69
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_70
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_71
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp -3599
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_73
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_74
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_75
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_76
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp -3599
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_83
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_84
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_85
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp -3599
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_87
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_88
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_92
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_93
timestamp -3599
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_95
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_96
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_97
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_98
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_99
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_100
timestamp -3599
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_101
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_102
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_103
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_104
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_105
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp -3599
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_108
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_109
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_110
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_111
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_112
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_113
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_114
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_115
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_116
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_117
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_118
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_119
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp -3599
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_121
timestamp -3599
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 17590 11194 17646 11250 0 FreeSans 224 0 0 0 Co
port 0 nsew signal output
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[0]
port 1 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[10]
port 2 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[11]
port 3 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[12]
port 4 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[13]
port 5 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[14]
port 6 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[15]
port 7 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[16]
port 8 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[17]
port 9 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[18]
port 10 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[19]
port 11 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[1]
port 12 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[20]
port 13 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[21]
port 14 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[22]
port 15 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[23]
port 16 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[24]
port 17 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[25]
port 18 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[26]
port 19 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[27]
port 20 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[28]
port 21 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[29]
port 22 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[2]
port 23 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[30]
port 24 nsew signal input
flabel metal3 s 0 9800 120 9920 0 FreeSans 480 0 0 0 FrameData[31]
port 25 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[3]
port 26 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[4]
port 27 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[5]
port 28 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[6]
port 29 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[7]
port 30 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[8]
port 31 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[9]
port 32 nsew signal input
flabel metal3 s 40880 1368 41000 1488 0 FreeSans 480 0 0 0 FrameData_O[0]
port 33 nsew signal output
flabel metal3 s 40880 4088 41000 4208 0 FreeSans 480 0 0 0 FrameData_O[10]
port 34 nsew signal output
flabel metal3 s 40880 4360 41000 4480 0 FreeSans 480 0 0 0 FrameData_O[11]
port 35 nsew signal output
flabel metal3 s 40880 4632 41000 4752 0 FreeSans 480 0 0 0 FrameData_O[12]
port 36 nsew signal output
flabel metal3 s 40880 4904 41000 5024 0 FreeSans 480 0 0 0 FrameData_O[13]
port 37 nsew signal output
flabel metal3 s 40880 5176 41000 5296 0 FreeSans 480 0 0 0 FrameData_O[14]
port 38 nsew signal output
flabel metal3 s 40880 5448 41000 5568 0 FreeSans 480 0 0 0 FrameData_O[15]
port 39 nsew signal output
flabel metal3 s 40880 5720 41000 5840 0 FreeSans 480 0 0 0 FrameData_O[16]
port 40 nsew signal output
flabel metal3 s 40880 5992 41000 6112 0 FreeSans 480 0 0 0 FrameData_O[17]
port 41 nsew signal output
flabel metal3 s 40880 6264 41000 6384 0 FreeSans 480 0 0 0 FrameData_O[18]
port 42 nsew signal output
flabel metal3 s 40880 6536 41000 6656 0 FreeSans 480 0 0 0 FrameData_O[19]
port 43 nsew signal output
flabel metal3 s 40880 1640 41000 1760 0 FreeSans 480 0 0 0 FrameData_O[1]
port 44 nsew signal output
flabel metal3 s 40880 6808 41000 6928 0 FreeSans 480 0 0 0 FrameData_O[20]
port 45 nsew signal output
flabel metal3 s 40880 7080 41000 7200 0 FreeSans 480 0 0 0 FrameData_O[21]
port 46 nsew signal output
flabel metal3 s 40880 7352 41000 7472 0 FreeSans 480 0 0 0 FrameData_O[22]
port 47 nsew signal output
flabel metal3 s 40880 7624 41000 7744 0 FreeSans 480 0 0 0 FrameData_O[23]
port 48 nsew signal output
flabel metal3 s 40880 7896 41000 8016 0 FreeSans 480 0 0 0 FrameData_O[24]
port 49 nsew signal output
flabel metal3 s 40880 8168 41000 8288 0 FreeSans 480 0 0 0 FrameData_O[25]
port 50 nsew signal output
flabel metal3 s 40880 8440 41000 8560 0 FreeSans 480 0 0 0 FrameData_O[26]
port 51 nsew signal output
flabel metal3 s 40880 8712 41000 8832 0 FreeSans 480 0 0 0 FrameData_O[27]
port 52 nsew signal output
flabel metal3 s 40880 8984 41000 9104 0 FreeSans 480 0 0 0 FrameData_O[28]
port 53 nsew signal output
flabel metal3 s 40880 9256 41000 9376 0 FreeSans 480 0 0 0 FrameData_O[29]
port 54 nsew signal output
flabel metal3 s 40880 1912 41000 2032 0 FreeSans 480 0 0 0 FrameData_O[2]
port 55 nsew signal output
flabel metal3 s 40880 9528 41000 9648 0 FreeSans 480 0 0 0 FrameData_O[30]
port 56 nsew signal output
flabel metal3 s 40880 9800 41000 9920 0 FreeSans 480 0 0 0 FrameData_O[31]
port 57 nsew signal output
flabel metal3 s 40880 2184 41000 2304 0 FreeSans 480 0 0 0 FrameData_O[3]
port 58 nsew signal output
flabel metal3 s 40880 2456 41000 2576 0 FreeSans 480 0 0 0 FrameData_O[4]
port 59 nsew signal output
flabel metal3 s 40880 2728 41000 2848 0 FreeSans 480 0 0 0 FrameData_O[5]
port 60 nsew signal output
flabel metal3 s 40880 3000 41000 3120 0 FreeSans 480 0 0 0 FrameData_O[6]
port 61 nsew signal output
flabel metal3 s 40880 3272 41000 3392 0 FreeSans 480 0 0 0 FrameData_O[7]
port 62 nsew signal output
flabel metal3 s 40880 3544 41000 3664 0 FreeSans 480 0 0 0 FrameData_O[8]
port 63 nsew signal output
flabel metal3 s 40880 3816 41000 3936 0 FreeSans 480 0 0 0 FrameData_O[9]
port 64 nsew signal output
flabel metal2 s 25594 0 25650 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 65 nsew signal input
flabel metal2 s 32954 0 33010 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 66 nsew signal input
flabel metal2 s 33690 0 33746 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 67 nsew signal input
flabel metal2 s 34426 0 34482 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 68 nsew signal input
flabel metal2 s 35162 0 35218 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 69 nsew signal input
flabel metal2 s 35898 0 35954 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 70 nsew signal input
flabel metal2 s 36634 0 36690 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 71 nsew signal input
flabel metal2 s 37370 0 37426 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 72 nsew signal input
flabel metal2 s 38106 0 38162 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 73 nsew signal input
flabel metal2 s 38842 0 38898 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 74 nsew signal input
flabel metal2 s 39578 0 39634 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 75 nsew signal input
flabel metal2 s 26330 0 26386 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 76 nsew signal input
flabel metal2 s 27066 0 27122 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 77 nsew signal input
flabel metal2 s 27802 0 27858 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 78 nsew signal input
flabel metal2 s 28538 0 28594 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 79 nsew signal input
flabel metal2 s 29274 0 29330 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 80 nsew signal input
flabel metal2 s 30010 0 30066 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 81 nsew signal input
flabel metal2 s 30746 0 30802 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 82 nsew signal input
flabel metal2 s 31482 0 31538 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 83 nsew signal input
flabel metal2 s 32218 0 32274 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 84 nsew signal input
flabel metal2 s 32494 11194 32550 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 85 nsew signal output
flabel metal2 s 35254 11194 35310 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 86 nsew signal output
flabel metal2 s 35530 11194 35586 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 87 nsew signal output
flabel metal2 s 35806 11194 35862 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 88 nsew signal output
flabel metal2 s 36082 11194 36138 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 89 nsew signal output
flabel metal2 s 36358 11194 36414 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 90 nsew signal output
flabel metal2 s 36634 11194 36690 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 91 nsew signal output
flabel metal2 s 36910 11194 36966 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 92 nsew signal output
flabel metal2 s 37186 11194 37242 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 93 nsew signal output
flabel metal2 s 37462 11194 37518 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 94 nsew signal output
flabel metal2 s 37738 11194 37794 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 95 nsew signal output
flabel metal2 s 32770 11194 32826 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 96 nsew signal output
flabel metal2 s 33046 11194 33102 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 97 nsew signal output
flabel metal2 s 33322 11194 33378 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 98 nsew signal output
flabel metal2 s 33598 11194 33654 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 99 nsew signal output
flabel metal2 s 33874 11194 33930 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 100 nsew signal output
flabel metal2 s 34150 11194 34206 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 101 nsew signal output
flabel metal2 s 34426 11194 34482 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 102 nsew signal output
flabel metal2 s 34702 11194 34758 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 103 nsew signal output
flabel metal2 s 34978 11194 35034 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 104 nsew signal output
flabel metal2 s 13082 0 13138 56 0 FreeSans 224 0 0 0 I_top0
port 105 nsew signal output
flabel metal2 s 13818 0 13874 56 0 FreeSans 224 0 0 0 I_top1
port 106 nsew signal output
flabel metal2 s 20442 0 20498 56 0 FreeSans 224 0 0 0 I_top10
port 107 nsew signal output
flabel metal2 s 21178 0 21234 56 0 FreeSans 224 0 0 0 I_top11
port 108 nsew signal output
flabel metal2 s 21914 0 21970 56 0 FreeSans 224 0 0 0 I_top12
port 109 nsew signal output
flabel metal2 s 22650 0 22706 56 0 FreeSans 224 0 0 0 I_top13
port 110 nsew signal output
flabel metal2 s 23386 0 23442 56 0 FreeSans 224 0 0 0 I_top14
port 111 nsew signal output
flabel metal2 s 24122 0 24178 56 0 FreeSans 224 0 0 0 I_top15
port 112 nsew signal output
flabel metal2 s 14554 0 14610 56 0 FreeSans 224 0 0 0 I_top2
port 113 nsew signal output
flabel metal2 s 15290 0 15346 56 0 FreeSans 224 0 0 0 I_top3
port 114 nsew signal output
flabel metal2 s 16026 0 16082 56 0 FreeSans 224 0 0 0 I_top4
port 115 nsew signal output
flabel metal2 s 16762 0 16818 56 0 FreeSans 224 0 0 0 I_top5
port 116 nsew signal output
flabel metal2 s 17498 0 17554 56 0 FreeSans 224 0 0 0 I_top6
port 117 nsew signal output
flabel metal2 s 18234 0 18290 56 0 FreeSans 224 0 0 0 I_top7
port 118 nsew signal output
flabel metal2 s 18970 0 19026 56 0 FreeSans 224 0 0 0 I_top8
port 119 nsew signal output
flabel metal2 s 19706 0 19762 56 0 FreeSans 224 0 0 0 I_top9
port 120 nsew signal output
flabel metal2 s 3238 11194 3294 11250 0 FreeSans 224 0 0 0 N1BEG[0]
port 121 nsew signal output
flabel metal2 s 3514 11194 3570 11250 0 FreeSans 224 0 0 0 N1BEG[1]
port 122 nsew signal output
flabel metal2 s 3790 11194 3846 11250 0 FreeSans 224 0 0 0 N1BEG[2]
port 123 nsew signal output
flabel metal2 s 4066 11194 4122 11250 0 FreeSans 224 0 0 0 N1BEG[3]
port 124 nsew signal output
flabel metal2 s 4342 11194 4398 11250 0 FreeSans 224 0 0 0 N2BEG[0]
port 125 nsew signal output
flabel metal2 s 4618 11194 4674 11250 0 FreeSans 224 0 0 0 N2BEG[1]
port 126 nsew signal output
flabel metal2 s 4894 11194 4950 11250 0 FreeSans 224 0 0 0 N2BEG[2]
port 127 nsew signal output
flabel metal2 s 5170 11194 5226 11250 0 FreeSans 224 0 0 0 N2BEG[3]
port 128 nsew signal output
flabel metal2 s 5446 11194 5502 11250 0 FreeSans 224 0 0 0 N2BEG[4]
port 129 nsew signal output
flabel metal2 s 5722 11194 5778 11250 0 FreeSans 224 0 0 0 N2BEG[5]
port 130 nsew signal output
flabel metal2 s 5998 11194 6054 11250 0 FreeSans 224 0 0 0 N2BEG[6]
port 131 nsew signal output
flabel metal2 s 6274 11194 6330 11250 0 FreeSans 224 0 0 0 N2BEG[7]
port 132 nsew signal output
flabel metal2 s 6550 11194 6606 11250 0 FreeSans 224 0 0 0 N2BEGb[0]
port 133 nsew signal output
flabel metal2 s 6826 11194 6882 11250 0 FreeSans 224 0 0 0 N2BEGb[1]
port 134 nsew signal output
flabel metal2 s 7102 11194 7158 11250 0 FreeSans 224 0 0 0 N2BEGb[2]
port 135 nsew signal output
flabel metal2 s 7378 11194 7434 11250 0 FreeSans 224 0 0 0 N2BEGb[3]
port 136 nsew signal output
flabel metal2 s 7654 11194 7710 11250 0 FreeSans 224 0 0 0 N2BEGb[4]
port 137 nsew signal output
flabel metal2 s 7930 11194 7986 11250 0 FreeSans 224 0 0 0 N2BEGb[5]
port 138 nsew signal output
flabel metal2 s 8206 11194 8262 11250 0 FreeSans 224 0 0 0 N2BEGb[6]
port 139 nsew signal output
flabel metal2 s 8482 11194 8538 11250 0 FreeSans 224 0 0 0 N2BEGb[7]
port 140 nsew signal output
flabel metal2 s 8758 11194 8814 11250 0 FreeSans 224 0 0 0 N4BEG[0]
port 141 nsew signal output
flabel metal2 s 11518 11194 11574 11250 0 FreeSans 224 0 0 0 N4BEG[10]
port 142 nsew signal output
flabel metal2 s 11794 11194 11850 11250 0 FreeSans 224 0 0 0 N4BEG[11]
port 143 nsew signal output
flabel metal2 s 12070 11194 12126 11250 0 FreeSans 224 0 0 0 N4BEG[12]
port 144 nsew signal output
flabel metal2 s 12346 11194 12402 11250 0 FreeSans 224 0 0 0 N4BEG[13]
port 145 nsew signal output
flabel metal2 s 12622 11194 12678 11250 0 FreeSans 224 0 0 0 N4BEG[14]
port 146 nsew signal output
flabel metal2 s 12898 11194 12954 11250 0 FreeSans 224 0 0 0 N4BEG[15]
port 147 nsew signal output
flabel metal2 s 9034 11194 9090 11250 0 FreeSans 224 0 0 0 N4BEG[1]
port 148 nsew signal output
flabel metal2 s 9310 11194 9366 11250 0 FreeSans 224 0 0 0 N4BEG[2]
port 149 nsew signal output
flabel metal2 s 9586 11194 9642 11250 0 FreeSans 224 0 0 0 N4BEG[3]
port 150 nsew signal output
flabel metal2 s 9862 11194 9918 11250 0 FreeSans 224 0 0 0 N4BEG[4]
port 151 nsew signal output
flabel metal2 s 10138 11194 10194 11250 0 FreeSans 224 0 0 0 N4BEG[5]
port 152 nsew signal output
flabel metal2 s 10414 11194 10470 11250 0 FreeSans 224 0 0 0 N4BEG[6]
port 153 nsew signal output
flabel metal2 s 10690 11194 10746 11250 0 FreeSans 224 0 0 0 N4BEG[7]
port 154 nsew signal output
flabel metal2 s 10966 11194 11022 11250 0 FreeSans 224 0 0 0 N4BEG[8]
port 155 nsew signal output
flabel metal2 s 11242 11194 11298 11250 0 FreeSans 224 0 0 0 N4BEG[9]
port 156 nsew signal output
flabel metal2 s 13174 11194 13230 11250 0 FreeSans 224 0 0 0 NN4BEG[0]
port 157 nsew signal output
flabel metal2 s 15934 11194 15990 11250 0 FreeSans 224 0 0 0 NN4BEG[10]
port 158 nsew signal output
flabel metal2 s 16210 11194 16266 11250 0 FreeSans 224 0 0 0 NN4BEG[11]
port 159 nsew signal output
flabel metal2 s 16486 11194 16542 11250 0 FreeSans 224 0 0 0 NN4BEG[12]
port 160 nsew signal output
flabel metal2 s 16762 11194 16818 11250 0 FreeSans 224 0 0 0 NN4BEG[13]
port 161 nsew signal output
flabel metal2 s 17038 11194 17094 11250 0 FreeSans 224 0 0 0 NN4BEG[14]
port 162 nsew signal output
flabel metal2 s 17314 11194 17370 11250 0 FreeSans 224 0 0 0 NN4BEG[15]
port 163 nsew signal output
flabel metal2 s 13450 11194 13506 11250 0 FreeSans 224 0 0 0 NN4BEG[1]
port 164 nsew signal output
flabel metal2 s 13726 11194 13782 11250 0 FreeSans 224 0 0 0 NN4BEG[2]
port 165 nsew signal output
flabel metal2 s 14002 11194 14058 11250 0 FreeSans 224 0 0 0 NN4BEG[3]
port 166 nsew signal output
flabel metal2 s 14278 11194 14334 11250 0 FreeSans 224 0 0 0 NN4BEG[4]
port 167 nsew signal output
flabel metal2 s 14554 11194 14610 11250 0 FreeSans 224 0 0 0 NN4BEG[5]
port 168 nsew signal output
flabel metal2 s 14830 11194 14886 11250 0 FreeSans 224 0 0 0 NN4BEG[6]
port 169 nsew signal output
flabel metal2 s 15106 11194 15162 11250 0 FreeSans 224 0 0 0 NN4BEG[7]
port 170 nsew signal output
flabel metal2 s 15382 11194 15438 11250 0 FreeSans 224 0 0 0 NN4BEG[8]
port 171 nsew signal output
flabel metal2 s 15658 11194 15714 11250 0 FreeSans 224 0 0 0 NN4BEG[9]
port 172 nsew signal output
flabel metal2 s 1306 0 1362 56 0 FreeSans 224 0 0 0 O_top0
port 173 nsew signal input
flabel metal2 s 2042 0 2098 56 0 FreeSans 224 0 0 0 O_top1
port 174 nsew signal input
flabel metal2 s 8666 0 8722 56 0 FreeSans 224 0 0 0 O_top10
port 175 nsew signal input
flabel metal2 s 9402 0 9458 56 0 FreeSans 224 0 0 0 O_top11
port 176 nsew signal input
flabel metal2 s 10138 0 10194 56 0 FreeSans 224 0 0 0 O_top12
port 177 nsew signal input
flabel metal2 s 10874 0 10930 56 0 FreeSans 224 0 0 0 O_top13
port 178 nsew signal input
flabel metal2 s 11610 0 11666 56 0 FreeSans 224 0 0 0 O_top14
port 179 nsew signal input
flabel metal2 s 12346 0 12402 56 0 FreeSans 224 0 0 0 O_top15
port 180 nsew signal input
flabel metal2 s 2778 0 2834 56 0 FreeSans 224 0 0 0 O_top2
port 181 nsew signal input
flabel metal2 s 3514 0 3570 56 0 FreeSans 224 0 0 0 O_top3
port 182 nsew signal input
flabel metal2 s 4250 0 4306 56 0 FreeSans 224 0 0 0 O_top4
port 183 nsew signal input
flabel metal2 s 4986 0 5042 56 0 FreeSans 224 0 0 0 O_top5
port 184 nsew signal input
flabel metal2 s 5722 0 5778 56 0 FreeSans 224 0 0 0 O_top6
port 185 nsew signal input
flabel metal2 s 6458 0 6514 56 0 FreeSans 224 0 0 0 O_top7
port 186 nsew signal input
flabel metal2 s 7194 0 7250 56 0 FreeSans 224 0 0 0 O_top8
port 187 nsew signal input
flabel metal2 s 7930 0 7986 56 0 FreeSans 224 0 0 0 O_top9
port 188 nsew signal input
flabel metal2 s 17866 11194 17922 11250 0 FreeSans 224 0 0 0 S1END[0]
port 189 nsew signal input
flabel metal2 s 18142 11194 18198 11250 0 FreeSans 224 0 0 0 S1END[1]
port 190 nsew signal input
flabel metal2 s 18418 11194 18474 11250 0 FreeSans 224 0 0 0 S1END[2]
port 191 nsew signal input
flabel metal2 s 18694 11194 18750 11250 0 FreeSans 224 0 0 0 S1END[3]
port 192 nsew signal input
flabel metal2 s 21178 11194 21234 11250 0 FreeSans 224 0 0 0 S2END[0]
port 193 nsew signal input
flabel metal2 s 21454 11194 21510 11250 0 FreeSans 224 0 0 0 S2END[1]
port 194 nsew signal input
flabel metal2 s 21730 11194 21786 11250 0 FreeSans 224 0 0 0 S2END[2]
port 195 nsew signal input
flabel metal2 s 22006 11194 22062 11250 0 FreeSans 224 0 0 0 S2END[3]
port 196 nsew signal input
flabel metal2 s 22282 11194 22338 11250 0 FreeSans 224 0 0 0 S2END[4]
port 197 nsew signal input
flabel metal2 s 22558 11194 22614 11250 0 FreeSans 224 0 0 0 S2END[5]
port 198 nsew signal input
flabel metal2 s 22834 11194 22890 11250 0 FreeSans 224 0 0 0 S2END[6]
port 199 nsew signal input
flabel metal2 s 23110 11194 23166 11250 0 FreeSans 224 0 0 0 S2END[7]
port 200 nsew signal input
flabel metal2 s 18970 11194 19026 11250 0 FreeSans 224 0 0 0 S2MID[0]
port 201 nsew signal input
flabel metal2 s 19246 11194 19302 11250 0 FreeSans 224 0 0 0 S2MID[1]
port 202 nsew signal input
flabel metal2 s 19522 11194 19578 11250 0 FreeSans 224 0 0 0 S2MID[2]
port 203 nsew signal input
flabel metal2 s 19798 11194 19854 11250 0 FreeSans 224 0 0 0 S2MID[3]
port 204 nsew signal input
flabel metal2 s 20074 11194 20130 11250 0 FreeSans 224 0 0 0 S2MID[4]
port 205 nsew signal input
flabel metal2 s 20350 11194 20406 11250 0 FreeSans 224 0 0 0 S2MID[5]
port 206 nsew signal input
flabel metal2 s 20626 11194 20682 11250 0 FreeSans 224 0 0 0 S2MID[6]
port 207 nsew signal input
flabel metal2 s 20902 11194 20958 11250 0 FreeSans 224 0 0 0 S2MID[7]
port 208 nsew signal input
flabel metal2 s 23386 11194 23442 11250 0 FreeSans 224 0 0 0 S4END[0]
port 209 nsew signal input
flabel metal2 s 26146 11194 26202 11250 0 FreeSans 224 0 0 0 S4END[10]
port 210 nsew signal input
flabel metal2 s 26422 11194 26478 11250 0 FreeSans 224 0 0 0 S4END[11]
port 211 nsew signal input
flabel metal2 s 26698 11194 26754 11250 0 FreeSans 224 0 0 0 S4END[12]
port 212 nsew signal input
flabel metal2 s 26974 11194 27030 11250 0 FreeSans 224 0 0 0 S4END[13]
port 213 nsew signal input
flabel metal2 s 27250 11194 27306 11250 0 FreeSans 224 0 0 0 S4END[14]
port 214 nsew signal input
flabel metal2 s 27526 11194 27582 11250 0 FreeSans 224 0 0 0 S4END[15]
port 215 nsew signal input
flabel metal2 s 23662 11194 23718 11250 0 FreeSans 224 0 0 0 S4END[1]
port 216 nsew signal input
flabel metal2 s 23938 11194 23994 11250 0 FreeSans 224 0 0 0 S4END[2]
port 217 nsew signal input
flabel metal2 s 24214 11194 24270 11250 0 FreeSans 224 0 0 0 S4END[3]
port 218 nsew signal input
flabel metal2 s 24490 11194 24546 11250 0 FreeSans 224 0 0 0 S4END[4]
port 219 nsew signal input
flabel metal2 s 24766 11194 24822 11250 0 FreeSans 224 0 0 0 S4END[5]
port 220 nsew signal input
flabel metal2 s 25042 11194 25098 11250 0 FreeSans 224 0 0 0 S4END[6]
port 221 nsew signal input
flabel metal2 s 25318 11194 25374 11250 0 FreeSans 224 0 0 0 S4END[7]
port 222 nsew signal input
flabel metal2 s 25594 11194 25650 11250 0 FreeSans 224 0 0 0 S4END[8]
port 223 nsew signal input
flabel metal2 s 25870 11194 25926 11250 0 FreeSans 224 0 0 0 S4END[9]
port 224 nsew signal input
flabel metal2 s 27802 11194 27858 11250 0 FreeSans 224 0 0 0 SS4END[0]
port 225 nsew signal input
flabel metal2 s 30562 11194 30618 11250 0 FreeSans 224 0 0 0 SS4END[10]
port 226 nsew signal input
flabel metal2 s 30838 11194 30894 11250 0 FreeSans 224 0 0 0 SS4END[11]
port 227 nsew signal input
flabel metal2 s 31114 11194 31170 11250 0 FreeSans 224 0 0 0 SS4END[12]
port 228 nsew signal input
flabel metal2 s 31390 11194 31446 11250 0 FreeSans 224 0 0 0 SS4END[13]
port 229 nsew signal input
flabel metal2 s 31666 11194 31722 11250 0 FreeSans 224 0 0 0 SS4END[14]
port 230 nsew signal input
flabel metal2 s 31942 11194 31998 11250 0 FreeSans 224 0 0 0 SS4END[15]
port 231 nsew signal input
flabel metal2 s 28078 11194 28134 11250 0 FreeSans 224 0 0 0 SS4END[1]
port 232 nsew signal input
flabel metal2 s 28354 11194 28410 11250 0 FreeSans 224 0 0 0 SS4END[2]
port 233 nsew signal input
flabel metal2 s 28630 11194 28686 11250 0 FreeSans 224 0 0 0 SS4END[3]
port 234 nsew signal input
flabel metal2 s 28906 11194 28962 11250 0 FreeSans 224 0 0 0 SS4END[4]
port 235 nsew signal input
flabel metal2 s 29182 11194 29238 11250 0 FreeSans 224 0 0 0 SS4END[5]
port 236 nsew signal input
flabel metal2 s 29458 11194 29514 11250 0 FreeSans 224 0 0 0 SS4END[6]
port 237 nsew signal input
flabel metal2 s 29734 11194 29790 11250 0 FreeSans 224 0 0 0 SS4END[7]
port 238 nsew signal input
flabel metal2 s 30010 11194 30066 11250 0 FreeSans 224 0 0 0 SS4END[8]
port 239 nsew signal input
flabel metal2 s 30286 11194 30342 11250 0 FreeSans 224 0 0 0 SS4END[9]
port 240 nsew signal input
flabel metal2 s 24858 0 24914 56 0 FreeSans 224 0 0 0 UserCLK
port 241 nsew signal input
flabel metal2 s 32218 11194 32274 11250 0 FreeSans 224 0 0 0 UserCLKo
port 242 nsew signal output
flabel metal4 s 3004 0 3324 11250 0 FreeSans 1920 90 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 3004 11190 3324 11250 0 FreeSans 480 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11250 0 FreeSans 1920 90 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 9004 11190 9324 11250 0 FreeSans 480 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11250 0 FreeSans 1920 90 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 15004 11190 15324 11250 0 FreeSans 480 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11250 0 FreeSans 1920 90 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 21004 11190 21324 11250 0 FreeSans 480 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11250 0 FreeSans 1920 90 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 27004 11190 27324 11250 0 FreeSans 480 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11250 0 FreeSans 1920 90 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 33004 11190 33324 11250 0 FreeSans 480 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 39004 0 39324 11250 0 FreeSans 1920 90 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 39004 0 39324 60 0 FreeSans 480 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 39004 11190 39324 11250 0 FreeSans 480 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11250 0 FreeSans 1920 90 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 1944 11190 2264 11250 0 FreeSans 480 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 7944 0 8264 11250 0 FreeSans 1920 90 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 7944 11190 8264 11250 0 FreeSans 480 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 13944 0 14264 11250 0 FreeSans 1920 90 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 13944 11190 14264 11250 0 FreeSans 480 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 19944 0 20264 11250 0 FreeSans 1920 90 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 19944 11190 20264 11250 0 FreeSans 480 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 25944 0 26264 11250 0 FreeSans 1920 90 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 25944 11190 26264 11250 0 FreeSans 480 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 31944 0 32264 11250 0 FreeSans 1920 90 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 31944 11190 32264 11250 0 FreeSans 480 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 37944 0 38264 11250 0 FreeSans 1920 90 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 37944 0 38264 60 0 FreeSans 480 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal4 s 37944 11190 38264 11250 0 FreeSans 480 0 0 0 VPWR
port 244 nsew power bidirectional
rlabel metal1 20470 8704 20470 8704 0 VGND
rlabel metal1 20470 8160 20470 8160 0 VPWR
rlabel metal3 1356 1428 1356 1428 0 FrameData[0]
rlabel metal3 436 4148 436 4148 0 FrameData[10]
rlabel metal3 436 4420 436 4420 0 FrameData[11]
rlabel metal3 528 4692 528 4692 0 FrameData[12]
rlabel metal3 252 4964 252 4964 0 FrameData[13]
rlabel metal3 574 5236 574 5236 0 FrameData[14]
rlabel metal3 344 5508 344 5508 0 FrameData[15]
rlabel metal3 436 5780 436 5780 0 FrameData[16]
rlabel metal3 436 6052 436 6052 0 FrameData[17]
rlabel metal3 528 6324 528 6324 0 FrameData[18]
rlabel metal3 160 6596 160 6596 0 FrameData[19]
rlabel metal3 666 1700 666 1700 0 FrameData[1]
rlabel metal2 2990 7123 2990 7123 0 FrameData[20]
rlabel metal3 620 7140 620 7140 0 FrameData[21]
rlabel metal3 528 7412 528 7412 0 FrameData[22]
rlabel metal3 436 7684 436 7684 0 FrameData[23]
rlabel metal3 436 7956 436 7956 0 FrameData[24]
rlabel metal3 252 8228 252 8228 0 FrameData[25]
rlabel metal3 712 8500 712 8500 0 FrameData[26]
rlabel metal2 2898 8313 2898 8313 0 FrameData[27]
rlabel metal2 2806 8449 2806 8449 0 FrameData[28]
rlabel metal3 666 9316 666 9316 0 FrameData[29]
rlabel metal3 988 1972 988 1972 0 FrameData[2]
rlabel metal3 390 9588 390 9588 0 FrameData[30]
rlabel metal3 298 9860 298 9860 0 FrameData[31]
rlabel metal3 620 2244 620 2244 0 FrameData[3]
rlabel metal3 252 2516 252 2516 0 FrameData[4]
rlabel metal3 666 2788 666 2788 0 FrameData[5]
rlabel metal3 712 3060 712 3060 0 FrameData[6]
rlabel metal3 160 3332 160 3332 0 FrameData[7]
rlabel metal3 344 3604 344 3604 0 FrameData[8]
rlabel metal3 528 3876 528 3876 0 FrameData[9]
rlabel metal3 39798 1428 39798 1428 0 FrameData_O[0]
rlabel metal2 39422 3927 39422 3927 0 FrameData_O[10]
rlabel metal3 40442 4420 40442 4420 0 FrameData_O[11]
rlabel metal1 39468 3978 39468 3978 0 FrameData_O[12]
rlabel metal3 39982 4964 39982 4964 0 FrameData_O[13]
rlabel metal2 39422 5015 39422 5015 0 FrameData_O[14]
rlabel metal3 40442 5508 40442 5508 0 FrameData_O[15]
rlabel metal2 39422 5559 39422 5559 0 FrameData_O[16]
rlabel metal3 39982 6052 39982 6052 0 FrameData_O[17]
rlabel metal3 39798 6324 39798 6324 0 FrameData_O[18]
rlabel metal1 39560 5882 39560 5882 0 FrameData_O[19]
rlabel metal3 39614 1700 39614 1700 0 FrameData_O[1]
rlabel metal3 40488 6868 40488 6868 0 FrameData_O[20]
rlabel metal2 39422 6885 39422 6885 0 FrameData_O[21]
rlabel metal3 39936 7412 39936 7412 0 FrameData_O[22]
rlabel metal3 40166 7684 40166 7684 0 FrameData_O[23]
rlabel metal3 40166 7956 40166 7956 0 FrameData_O[24]
rlabel metal1 39054 7480 39054 7480 0 FrameData_O[25]
rlabel metal2 38686 8279 38686 8279 0 FrameData_O[26]
rlabel metal1 39514 7514 39514 7514 0 FrameData_O[27]
rlabel metal1 39652 6426 39652 6426 0 FrameData_O[28]
rlabel metal1 38732 7514 38732 7514 0 FrameData_O[29]
rlabel metal3 39430 1972 39430 1972 0 FrameData_O[2]
rlabel metal1 39054 6664 39054 6664 0 FrameData_O[30]
rlabel metal2 38318 8687 38318 8687 0 FrameData_O[31]
rlabel metal3 40442 2244 40442 2244 0 FrameData_O[3]
rlabel metal3 39798 2516 39798 2516 0 FrameData_O[4]
rlabel metal3 39982 2788 39982 2788 0 FrameData_O[5]
rlabel metal3 40166 3060 40166 3060 0 FrameData_O[6]
rlabel metal3 40442 3332 40442 3332 0 FrameData_O[7]
rlabel metal2 39422 3383 39422 3383 0 FrameData_O[8]
rlabel metal3 39982 3876 39982 3876 0 FrameData_O[9]
rlabel metal2 25622 922 25622 922 0 FrameStrobe[0]
rlabel metal2 32982 1058 32982 1058 0 FrameStrobe[10]
rlabel metal1 34960 3434 34960 3434 0 FrameStrobe[11]
rlabel metal2 34454 1401 34454 1401 0 FrameStrobe[12]
rlabel metal2 35190 1401 35190 1401 0 FrameStrobe[13]
rlabel metal2 35926 55 35926 55 0 FrameStrobe[14]
rlabel metal1 35420 7446 35420 7446 0 FrameStrobe[15]
rlabel metal1 37904 7922 37904 7922 0 FrameStrobe[16]
rlabel metal2 38134 718 38134 718 0 FrameStrobe[17]
rlabel metal2 38870 1401 38870 1401 0 FrameStrobe[18]
rlabel metal1 38824 6154 38824 6154 0 FrameStrobe[19]
rlabel metal2 26358 1194 26358 1194 0 FrameStrobe[1]
rlabel metal2 27094 718 27094 718 0 FrameStrobe[2]
rlabel metal2 27830 55 27830 55 0 FrameStrobe[3]
rlabel metal2 28566 55 28566 55 0 FrameStrobe[4]
rlabel metal2 29302 55 29302 55 0 FrameStrobe[5]
rlabel metal2 38410 2975 38410 2975 0 FrameStrobe[6]
rlabel metal2 30774 55 30774 55 0 FrameStrobe[7]
rlabel metal2 31510 1279 31510 1279 0 FrameStrobe[8]
rlabel metal2 32246 514 32246 514 0 FrameStrobe[9]
rlabel metal1 32890 8602 32890 8602 0 FrameStrobe_O[0]
rlabel metal1 35788 8330 35788 8330 0 FrameStrobe_O[10]
rlabel metal1 35650 8058 35650 8058 0 FrameStrobe_O[11]
rlabel metal1 36248 8602 36248 8602 0 FrameStrobe_O[12]
rlabel metal1 36202 8058 36202 8058 0 FrameStrobe_O[13]
rlabel metal1 37306 8262 37306 8262 0 FrameStrobe_O[14]
rlabel metal1 36800 8058 36800 8058 0 FrameStrobe_O[15]
rlabel metal1 37352 8602 37352 8602 0 FrameStrobe_O[16]
rlabel metal1 37720 8330 37720 8330 0 FrameStrobe_O[17]
rlabel metal1 38502 8568 38502 8568 0 FrameStrobe_O[18]
rlabel metal1 37904 7990 37904 7990 0 FrameStrobe_O[19]
rlabel metal1 33166 8330 33166 8330 0 FrameStrobe_O[1]
rlabel metal1 33856 8602 33856 8602 0 FrameStrobe_O[2]
rlabel metal1 34270 8364 34270 8364 0 FrameStrobe_O[3]
rlabel metal1 33718 8058 33718 8058 0 FrameStrobe_O[4]
rlabel metal1 34592 8330 34592 8330 0 FrameStrobe_O[5]
rlabel metal1 35190 8364 35190 8364 0 FrameStrobe_O[6]
rlabel metal1 34638 8058 34638 8058 0 FrameStrobe_O[7]
rlabel metal1 35144 8602 35144 8602 0 FrameStrobe_O[8]
rlabel metal1 35558 8262 35558 8262 0 FrameStrobe_O[9]
rlabel metal2 13110 1160 13110 1160 0 I_top0
rlabel metal2 13846 1160 13846 1160 0 I_top1
rlabel metal2 20470 1160 20470 1160 0 I_top10
rlabel metal2 21206 55 21206 55 0 I_top11
rlabel metal2 21942 922 21942 922 0 I_top12
rlabel metal2 22678 1330 22678 1330 0 I_top13
rlabel metal2 23414 1296 23414 1296 0 I_top14
rlabel metal2 24150 1160 24150 1160 0 I_top15
rlabel metal2 14582 1160 14582 1160 0 I_top2
rlabel metal2 15318 599 15318 599 0 I_top3
rlabel metal2 16054 1160 16054 1160 0 I_top4
rlabel metal2 16790 1160 16790 1160 0 I_top5
rlabel metal2 17526 55 17526 55 0 I_top6
rlabel metal2 18262 1160 18262 1160 0 I_top7
rlabel metal2 18998 1160 18998 1160 0 I_top8
rlabel metal2 19734 871 19734 871 0 I_top9
rlabel metal2 19366 4420 19366 4420 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit0.Q
rlabel metal1 20930 4658 20930 4658 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 4738 4250 4738 4250 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 4186 4828 4186 4828 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit11.Q
rlabel metal1 29394 5814 29394 5814 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit12.Q
rlabel metal1 29302 4794 29302 4794 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit13.Q
rlabel metal1 15042 5882 15042 5882 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit14.Q
rlabel metal1 15364 5066 15364 5066 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit15.Q
rlabel metal1 17802 6426 17802 6426 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 18446 6188 18446 6188 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit17.Q
rlabel metal1 8924 3638 8924 3638 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 10166 3927 10166 3927 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit19.Q
rlabel metal1 8924 2890 8924 2890 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit2.Q
rlabel metal1 32154 4658 32154 4658 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit20.Q
rlabel metal1 32430 4250 32430 4250 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit21.Q
rlabel metal1 23000 4250 23000 4250 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 23598 4794 23598 4794 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 20654 8160 20654 8160 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit24.Q
rlabel metal1 21390 7922 21390 7922 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 7038 4148 7038 4148 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 7590 4828 7590 4828 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit27.Q
rlabel metal1 31786 6800 31786 6800 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit28.Q
rlabel metal1 33074 6426 33074 6426 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 19366 1870 19366 1870 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit3.Q
rlabel metal1 12236 4794 12236 4794 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit30.Q
rlabel metal1 13386 5134 13386 5134 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit31.Q
rlabel metal1 31510 3672 31510 3672 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit4.Q
rlabel metal1 30682 3162 30682 3162 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit5.Q
rlabel metal1 23000 2550 23000 2550 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit6.Q
rlabel metal1 23414 7514 23414 7514 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit7.Q
rlabel metal1 9246 7208 9246 7208 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit8.Q
rlabel metal1 8740 6970 8740 6970 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit9.Q
rlabel metal1 13386 5746 13386 5746 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit0.Q
rlabel metal1 22632 5882 22632 5882 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit1.Q
rlabel metal1 3450 4046 3450 4046 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 4922 7208 4922 7208 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 23506 7412 23506 7412 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit12.Q
rlabel metal1 31050 3026 31050 3026 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit13.Q
rlabel metal1 11086 3638 11086 3638 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 19274 4250 19274 4250 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 12006 5916 12006 5916 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit16.Q
rlabel metal1 32706 7344 32706 7344 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit17.Q
rlabel metal1 6348 3162 6348 3162 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit18.Q
rlabel metal1 20884 6834 20884 6834 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 5934 3094 5934 3094 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit2.Q
rlabel metal1 26174 4692 26174 4692 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit20.Q
rlabel metal1 35236 4250 35236 4250 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit21.Q
rlabel metal1 18354 2924 18354 2924 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 17894 7140 17894 7140 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit23.Q
rlabel metal1 11960 7310 11960 7310 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 30130 7038 30130 7038 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 3450 4148 3450 4148 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit26.Q
rlabel metal1 6118 6426 6118 6426 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit27.Q
rlabel metal1 17710 7956 17710 7956 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit28.Q
rlabel metal1 32062 2482 32062 2482 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit29.Q
rlabel metal1 20102 6188 20102 6188 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit3.Q
rlabel metal1 12190 2924 12190 2924 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 18630 3774 18630 3774 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 25622 3604 25622 3604 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit4.Q
rlabel metal1 36202 4250 36202 4250 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit5.Q
rlabel metal1 17710 2550 17710 2550 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit6.Q
rlabel metal1 17204 6834 17204 6834 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit7.Q
rlabel metal1 8970 7752 8970 7752 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit8.Q
rlabel metal1 14030 5712 14030 5712 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit9.Q
rlabel metal1 29486 5338 29486 5338 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit10.Q
rlabel metal1 27462 5576 27462 5576 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 13294 3502 13294 3502 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit12.Q
rlabel metal1 18584 850 18584 850 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit13.Q
rlabel metal1 18170 5066 18170 5066 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 19274 5355 19274 5355 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 12006 6630 12006 6630 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 30774 7514 30774 7514 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit17.Q
rlabel metal1 7590 4692 7590 4692 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 20470 7888 20470 7888 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 23598 6596 23598 6596 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit20.Q
rlabel metal1 30360 4046 30360 4046 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit21.Q
rlabel metal1 11040 2482 11040 2482 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit22.Q
rlabel metal1 20240 4046 20240 4046 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 14398 7310 14398 7310 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 31878 5916 31878 5916 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit25.Q
rlabel metal1 9062 4012 9062 4012 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 8786 6409 8786 6409 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit27.Q
rlabel metal1 26450 6188 26450 6188 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 35466 5916 35466 5916 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit29.Q
rlabel metal1 16100 2958 16100 2958 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 14214 6494 14214 6494 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit31.Q
rlabel metal1 12742 8024 12742 8024 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit8.Q
rlabel metal1 10994 7276 10994 7276 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit9.Q
rlabel metal1 15226 7854 15226 7854 0 Inst_S_CPU_IF_switch_matrix.N1BEG0
rlabel metal2 32338 5440 32338 5440 0 Inst_S_CPU_IF_switch_matrix.N1BEG1
rlabel metal2 11178 4420 11178 4420 0 Inst_S_CPU_IF_switch_matrix.N1BEG2
rlabel metal1 20056 5202 20056 5202 0 Inst_S_CPU_IF_switch_matrix.N1BEG3
rlabel metal1 12926 6766 12926 6766 0 Inst_S_CPU_IF_switch_matrix.N2BEG0
rlabel metal1 30406 6766 30406 6766 0 Inst_S_CPU_IF_switch_matrix.N2BEG1
rlabel metal2 7038 4998 7038 4998 0 Inst_S_CPU_IF_switch_matrix.N2BEG2
rlabel via1 19918 7852 19918 7852 0 Inst_S_CPU_IF_switch_matrix.N2BEG3
rlabel metal1 24380 7514 24380 7514 0 Inst_S_CPU_IF_switch_matrix.N2BEG4
rlabel metal1 31050 4250 31050 4250 0 Inst_S_CPU_IF_switch_matrix.N2BEG5
rlabel metal1 11638 2618 11638 2618 0 Inst_S_CPU_IF_switch_matrix.N2BEG6
rlabel metal1 20700 4114 20700 4114 0 Inst_S_CPU_IF_switch_matrix.N2BEG7
rlabel metal1 14168 7514 14168 7514 0 Inst_S_CPU_IF_switch_matrix.N2BEGb0
rlabel metal1 32522 5882 32522 5882 0 Inst_S_CPU_IF_switch_matrix.N2BEGb1
rlabel metal1 8418 4250 8418 4250 0 Inst_S_CPU_IF_switch_matrix.N2BEGb2
rlabel metal1 18124 6290 18124 6290 0 Inst_S_CPU_IF_switch_matrix.N2BEGb3
rlabel metal1 25944 6086 25944 6086 0 Inst_S_CPU_IF_switch_matrix.N2BEGb4
rlabel metal2 36018 6086 36018 6086 0 Inst_S_CPU_IF_switch_matrix.N2BEGb5
rlabel metal1 15686 2924 15686 2924 0 Inst_S_CPU_IF_switch_matrix.N2BEGb6
rlabel metal1 15364 6970 15364 6970 0 Inst_S_CPU_IF_switch_matrix.N2BEGb7
rlabel metal1 11868 5202 11868 5202 0 Inst_S_CPU_IF_switch_matrix.N4BEG0
rlabel metal2 31142 6596 31142 6596 0 Inst_S_CPU_IF_switch_matrix.N4BEG1
rlabel metal1 2576 4114 2576 4114 0 Inst_S_CPU_IF_switch_matrix.N4BEG10
rlabel metal2 5566 6970 5566 6970 0 Inst_S_CPU_IF_switch_matrix.N4BEG11
rlabel metal1 22172 7854 22172 7854 0 Inst_S_CPU_IF_switch_matrix.N4BEG12
rlabel metal2 30498 2618 30498 2618 0 Inst_S_CPU_IF_switch_matrix.N4BEG13
rlabel metal1 12006 3468 12006 3468 0 Inst_S_CPU_IF_switch_matrix.N4BEG14
rlabel metal1 18676 4114 18676 4114 0 Inst_S_CPU_IF_switch_matrix.N4BEG15
rlabel metal1 4646 3060 4646 3060 0 Inst_S_CPU_IF_switch_matrix.N4BEG2
rlabel metal1 21206 6256 21206 6256 0 Inst_S_CPU_IF_switch_matrix.N4BEG3
rlabel metal1 24932 4114 24932 4114 0 Inst_S_CPU_IF_switch_matrix.N4BEG4
rlabel metal2 35926 4998 35926 4998 0 Inst_S_CPU_IF_switch_matrix.N4BEG5
rlabel metal1 17250 2618 17250 2618 0 Inst_S_CPU_IF_switch_matrix.N4BEG6
rlabel metal1 16376 6766 16376 6766 0 Inst_S_CPU_IF_switch_matrix.N4BEG7
rlabel metal2 11454 6970 11454 6970 0 Inst_S_CPU_IF_switch_matrix.N4BEG8
rlabel metal2 28658 6086 28658 6086 0 Inst_S_CPU_IF_switch_matrix.N4BEG9
rlabel metal1 11316 5678 11316 5678 0 Inst_S_CPU_IF_switch_matrix.NN4BEG0
rlabel metal1 32292 7514 32292 7514 0 Inst_S_CPU_IF_switch_matrix.NN4BEG1
rlabel metal2 2530 3876 2530 3876 0 Inst_S_CPU_IF_switch_matrix.NN4BEG10
rlabel metal1 5198 7310 5198 7310 0 Inst_S_CPU_IF_switch_matrix.NN4BEG11
rlabel metal2 17250 7548 17250 7548 0 Inst_S_CPU_IF_switch_matrix.NN4BEG12
rlabel metal1 31602 2618 31602 2618 0 Inst_S_CPU_IF_switch_matrix.NN4BEG13
rlabel metal1 9246 3094 9246 3094 0 Inst_S_CPU_IF_switch_matrix.NN4BEG14
rlabel viali 20378 3500 20378 3500 0 Inst_S_CPU_IF_switch_matrix.NN4BEG15
rlabel metal1 5290 3502 5290 3502 0 Inst_S_CPU_IF_switch_matrix.NN4BEG2
rlabel metal2 20930 6460 20930 6460 0 Inst_S_CPU_IF_switch_matrix.NN4BEG3
rlabel metal2 25622 4998 25622 4998 0 Inst_S_CPU_IF_switch_matrix.NN4BEG4
rlabel metal2 35006 4658 35006 4658 0 Inst_S_CPU_IF_switch_matrix.NN4BEG5
rlabel metal2 17802 3332 17802 3332 0 Inst_S_CPU_IF_switch_matrix.NN4BEG6
rlabel metal1 16974 7412 16974 7412 0 Inst_S_CPU_IF_switch_matrix.NN4BEG7
rlabel metal2 11546 6970 11546 6970 0 Inst_S_CPU_IF_switch_matrix.NN4BEG8
rlabel metal1 29578 6698 29578 6698 0 Inst_S_CPU_IF_switch_matrix.NN4BEG9
rlabel metal2 3450 8755 3450 8755 0 N1BEG[0]
rlabel metal1 3726 8058 3726 8058 0 N1BEG[1]
rlabel metal1 3634 8602 3634 8602 0 N1BEG[2]
rlabel metal1 4186 8058 4186 8058 0 N1BEG[3]
rlabel metal1 4278 8602 4278 8602 0 N2BEG[0]
rlabel metal1 4738 8058 4738 8058 0 N2BEG[1]
rlabel metal1 4738 8602 4738 8602 0 N2BEG[2]
rlabel metal1 5290 8058 5290 8058 0 N2BEG[3]
rlabel metal1 5198 8330 5198 8330 0 N2BEG[4]
rlabel metal1 5796 8058 5796 8058 0 N2BEG[5]
rlabel metal1 5290 8568 5290 8568 0 N2BEG[6]
rlabel metal1 5980 8602 5980 8602 0 N2BEG[7]
rlabel metal1 6394 8058 6394 8058 0 N2BEGb[0]
rlabel metal1 6026 8364 6026 8364 0 N2BEGb[1]
rlabel metal1 7222 7514 7222 7514 0 N2BEGb[2]
rlabel metal1 6808 8058 6808 8058 0 N2BEGb[3]
rlabel metal1 7406 7990 7406 7990 0 N2BEGb[4]
rlabel metal1 6486 8568 6486 8568 0 N2BEGb[5]
rlabel metal2 7498 8160 7498 8160 0 N2BEGb[6]
rlabel metal1 6762 8602 6762 8602 0 N2BEGb[7]
rlabel metal1 8924 6630 8924 6630 0 N4BEG[0]
rlabel metal1 11040 8330 11040 8330 0 N4BEG[10]
rlabel metal2 10902 9180 10902 9180 0 N4BEG[11]
rlabel metal1 11638 8602 11638 8602 0 N4BEG[12]
rlabel metal1 12098 7990 12098 7990 0 N4BEG[13]
rlabel metal1 13018 7514 13018 7514 0 N4BEG[14]
rlabel metal2 12926 10448 12926 10448 0 N4BEG[15]
rlabel metal1 8050 8602 8050 8602 0 N4BEG[1]
rlabel metal2 9338 10433 9338 10433 0 N4BEG[2]
rlabel metal1 9614 6732 9614 6732 0 N4BEG[3]
rlabel metal1 10028 6970 10028 6970 0 N4BEG[4]
rlabel metal2 9706 8687 9706 8687 0 N4BEG[5]
rlabel metal1 10304 8058 10304 8058 0 N4BEG[6]
rlabel metal1 10212 8262 10212 8262 0 N4BEG[7]
rlabel metal1 11132 7242 11132 7242 0 N4BEG[8]
rlabel metal1 10672 9690 10672 9690 0 N4BEG[9]
rlabel metal2 13202 10873 13202 10873 0 NN4BEG[0]
rlabel metal1 16100 7514 16100 7514 0 NN4BEG[10]
rlabel metal1 15778 8602 15778 8602 0 NN4BEG[11]
rlabel metal1 15732 8330 15732 8330 0 NN4BEG[12]
rlabel metal1 16376 8330 16376 8330 0 NN4BEG[13]
rlabel metal2 16422 9163 16422 9163 0 NN4BEG[14]
rlabel metal1 17204 8602 17204 8602 0 NN4BEG[15]
rlabel metal1 13570 7514 13570 7514 0 NN4BEG[1]
rlabel metal1 13156 8330 13156 8330 0 NN4BEG[2]
rlabel metal2 12834 9299 12834 9299 0 NN4BEG[3]
rlabel metal2 13202 9163 13202 9163 0 NN4BEG[4]
rlabel metal1 14214 8602 14214 8602 0 NN4BEG[5]
rlabel metal1 14950 7514 14950 7514 0 NN4BEG[6]
rlabel metal1 14628 8330 14628 8330 0 NN4BEG[7]
rlabel metal2 14950 9163 14950 9163 0 NN4BEG[8]
rlabel metal1 15640 8058 15640 8058 0 NN4BEG[9]
rlabel metal2 1334 1228 1334 1228 0 O_top0
rlabel metal2 2070 55 2070 55 0 O_top1
rlabel metal2 8694 1194 8694 1194 0 O_top10
rlabel metal2 9430 1228 9430 1228 0 O_top11
rlabel metal2 10166 1228 10166 1228 0 O_top12
rlabel metal2 10902 1228 10902 1228 0 O_top13
rlabel metal2 11638 1194 11638 1194 0 O_top14
rlabel metal2 12374 1228 12374 1228 0 O_top15
rlabel metal1 2898 3026 2898 3026 0 O_top2
rlabel metal2 3542 1228 3542 1228 0 O_top3
rlabel metal2 4278 1262 4278 1262 0 O_top4
rlabel metal2 4922 3060 4922 3060 0 O_top5
rlabel metal2 5750 1296 5750 1296 0 O_top6
rlabel metal2 6486 599 6486 599 0 O_top7
rlabel metal2 7222 599 7222 599 0 O_top8
rlabel metal2 7958 1228 7958 1228 0 O_top9
rlabel metal2 17894 10142 17894 10142 0 S1END[0]
rlabel metal2 18170 9836 18170 9836 0 S1END[1]
rlabel metal1 18354 7922 18354 7922 0 S1END[2]
rlabel metal1 18906 8466 18906 8466 0 S1END[3]
rlabel metal2 21206 10533 21206 10533 0 S2END[0]
rlabel metal2 21482 9836 21482 9836 0 S2END[1]
rlabel metal2 21758 9870 21758 9870 0 S2END[2]
rlabel metal2 22034 9904 22034 9904 0 S2END[3]
rlabel metal2 22310 9870 22310 9870 0 S2END[4]
rlabel metal2 22586 9904 22586 9904 0 S2END[5]
rlabel metal2 22862 10397 22862 10397 0 S2END[6]
rlabel metal2 23138 10601 23138 10601 0 S2END[7]
rlabel metal2 18998 9598 18998 9598 0 S2MID[0]
rlabel metal1 19136 7854 19136 7854 0 S2MID[1]
rlabel metal2 19550 10465 19550 10465 0 S2MID[2]
rlabel metal2 19826 10601 19826 10601 0 S2MID[3]
rlabel metal2 20102 10433 20102 10433 0 S2MID[4]
rlabel metal2 20378 10448 20378 10448 0 S2MID[5]
rlabel metal2 20654 10465 20654 10465 0 S2MID[6]
rlabel metal2 20930 9904 20930 9904 0 S2MID[7]
rlabel metal2 23414 10737 23414 10737 0 S4END[0]
rlabel metal2 26174 9870 26174 9870 0 S4END[10]
rlabel metal2 26450 9768 26450 9768 0 S4END[11]
rlabel metal2 26726 10397 26726 10397 0 S4END[12]
rlabel metal2 27002 10006 27002 10006 0 S4END[13]
rlabel metal2 27278 10941 27278 10941 0 S4END[14]
rlabel metal2 27554 9904 27554 9904 0 S4END[15]
rlabel metal2 23690 9802 23690 9802 0 S4END[1]
rlabel metal2 23966 10397 23966 10397 0 S4END[2]
rlabel metal1 24242 7752 24242 7752 0 S4END[3]
rlabel metal2 24518 9870 24518 9870 0 S4END[4]
rlabel metal2 24794 10533 24794 10533 0 S4END[5]
rlabel metal2 25070 10397 25070 10397 0 S4END[6]
rlabel metal2 25346 10193 25346 10193 0 S4END[7]
rlabel metal2 25622 10720 25622 10720 0 S4END[8]
rlabel metal2 25898 10482 25898 10482 0 S4END[9]
rlabel metal2 27830 9802 27830 9802 0 SS4END[0]
rlabel metal2 30590 9360 30590 9360 0 SS4END[10]
rlabel metal1 31786 7344 31786 7344 0 SS4END[11]
rlabel metal1 32338 7820 32338 7820 0 SS4END[12]
rlabel metal2 31418 9802 31418 9802 0 SS4END[13]
rlabel via1 31878 9605 31878 9605 0 SS4END[14]
rlabel metal2 31970 10346 31970 10346 0 SS4END[15]
rlabel metal2 28106 10414 28106 10414 0 SS4END[1]
rlabel metal2 28382 9292 28382 9292 0 SS4END[2]
rlabel metal2 28658 10006 28658 10006 0 SS4END[3]
rlabel metal2 28934 10533 28934 10533 0 SS4END[4]
rlabel metal2 29210 9802 29210 9802 0 SS4END[5]
rlabel metal2 29486 9870 29486 9870 0 SS4END[6]
rlabel metal1 30636 8602 30636 8602 0 SS4END[7]
rlabel metal2 30038 10414 30038 10414 0 SS4END[8]
rlabel metal2 31786 9775 31786 9775 0 SS4END[9]
rlabel metal2 37582 4063 37582 4063 0 UserCLK
rlabel metal1 32798 8058 32798 8058 0 UserCLKo
rlabel metal1 3864 3162 3864 3162 0 net1
rlabel metal2 6210 5338 6210 5338 0 net10
rlabel metal2 17250 9996 17250 9996 0 net100
rlabel metal1 32614 7514 32614 7514 0 net101
rlabel metal2 19734 8415 19734 8415 0 net102
rlabel metal1 11868 3162 11868 3162 0 net103
rlabel metal2 31326 2329 31326 2329 0 net104
rlabel metal1 17710 7854 17710 7854 0 net105
rlabel metal2 8924 7378 8924 7378 0 net106
rlabel metal2 4462 5015 4462 5015 0 net107
rlabel metal2 29946 7548 29946 7548 0 net108
rlabel metal2 15226 5950 15226 5950 0 net109
rlabel metal1 14766 5814 14766 5814 0 net11
rlabel metal1 17894 7514 17894 7514 0 net110
rlabel metal2 18170 3247 18170 3247 0 net111
rlabel metal2 38502 2465 38502 2465 0 net112
rlabel metal1 39238 3468 39238 3468 0 net113
rlabel metal1 38088 4522 38088 4522 0 net114
rlabel metal2 38962 3876 38962 3876 0 net115
rlabel metal1 38870 5168 38870 5168 0 net116
rlabel metal1 25300 918 25300 918 0 net117
rlabel metal1 16928 5338 16928 5338 0 net118
rlabel metal1 39468 5202 39468 5202 0 net119
rlabel metal1 2622 2550 2622 2550 0 net12
rlabel metal1 33258 6902 33258 6902 0 net120
rlabel metal2 38226 1581 38226 1581 0 net121
rlabel metal2 36478 8160 36478 8160 0 net122
rlabel metal2 38134 1972 38134 1972 0 net123
rlabel metal2 29210 4845 29210 4845 0 net124
rlabel metal1 33948 4726 33948 4726 0 net125
rlabel metal3 32476 6936 32476 6936 0 net126
rlabel metal2 37490 7514 37490 7514 0 net127
rlabel metal2 17434 10404 17434 10404 0 net128
rlabel metal2 34914 7786 34914 7786 0 net129
rlabel metal1 3680 7446 3680 7446 0 net13
rlabel metal2 2346 7735 2346 7735 0 net130
rlabel metal2 37582 8721 37582 8721 0 net131
rlabel metal1 33442 6664 33442 6664 0 net132
rlabel metal1 36800 3366 36800 3366 0 net133
rlabel metal2 33442 1564 33442 1564 0 net134
rlabel metal1 23644 1326 23644 1326 0 net135
rlabel metal2 17250 10574 17250 10574 0 net136
rlabel metal2 38594 2176 38594 2176 0 net137
rlabel metal1 38502 3060 38502 3060 0 net138
rlabel metal1 38778 3026 38778 3026 0 net139
rlabel metal2 34086 4182 34086 4182 0 net14
rlabel metal1 24058 2550 24058 2550 0 net140
rlabel via2 38870 3485 38870 3485 0 net141
rlabel metal1 39100 3026 39100 3026 0 net142
rlabel metal2 35190 3468 35190 3468 0 net143
rlabel metal2 31234 7922 31234 7922 0 net144
rlabel metal1 37674 4726 37674 4726 0 net145
rlabel metal2 36018 4675 36018 4675 0 net146
rlabel metal1 37582 4794 37582 4794 0 net147
rlabel metal1 36432 7854 36432 7854 0 net148
rlabel metal2 37306 8262 37306 8262 0 net149
rlabel metal1 17710 3026 17710 3026 0 net15
rlabel metal1 36708 7854 36708 7854 0 net150
rlabel metal1 38042 8058 38042 8058 0 net151
rlabel metal1 35604 7718 35604 7718 0 net152
rlabel metal2 38594 6902 38594 6902 0 net153
rlabel metal2 37858 7412 37858 7412 0 net154
rlabel metal1 33948 3162 33948 3162 0 net155
rlabel metal1 34638 3706 34638 3706 0 net156
rlabel metal1 38226 6664 38226 6664 0 net157
rlabel metal1 37352 6426 37352 6426 0 net158
rlabel metal1 37306 7514 37306 7514 0 net159
rlabel metal3 16468 4080 16468 4080 0 net16
rlabel metal1 37398 3162 37398 3162 0 net160
rlabel metal1 35006 7922 35006 7922 0 net161
rlabel metal1 36892 5542 36892 5542 0 net162
rlabel metal1 35696 7514 35696 7514 0 net163
rlabel metal1 16790 2380 16790 2380 0 net164
rlabel metal1 14122 2448 14122 2448 0 net165
rlabel metal1 23506 2312 23506 2312 0 net166
rlabel metal1 21528 2414 21528 2414 0 net167
rlabel metal2 22218 2414 22218 2414 0 net168
rlabel metal2 23506 1530 23506 1530 0 net169
rlabel metal2 1702 8806 1702 8806 0 net17
rlabel metal1 24150 2482 24150 2482 0 net170
rlabel metal2 24426 2074 24426 2074 0 net171
rlabel metal2 14950 2040 14950 2040 0 net172
rlabel metal2 24334 2193 24334 2193 0 net173
rlabel metal2 15778 2465 15778 2465 0 net174
rlabel viali 16698 2409 16698 2409 0 net175
rlabel metal2 18170 2006 18170 2006 0 net176
rlabel metal1 17756 2346 17756 2346 0 net177
rlabel metal1 18952 2414 18952 2414 0 net178
rlabel metal2 20930 2244 20930 2244 0 net179
rlabel metal2 2622 8976 2622 8976 0 net18
rlabel metal3 13892 7684 13892 7684 0 net180
rlabel metal2 12558 10200 12558 10200 0 net181
rlabel metal2 8510 8840 8510 8840 0 net182
rlabel via2 20010 5083 20010 5083 0 net183
rlabel metal1 13064 6630 13064 6630 0 net184
rlabel metal3 13708 6664 13708 6664 0 net185
rlabel metal1 5612 5338 5612 5338 0 net186
rlabel metal3 13708 7888 13708 7888 0 net187
rlabel metal2 5106 8823 5106 8823 0 net188
rlabel metal2 13754 4777 13754 4777 0 net189
rlabel metal1 2484 5202 2484 5202 0 net19
rlabel metal1 11638 3638 11638 3638 0 net190
rlabel metal1 16238 9690 16238 9690 0 net191
rlabel metal2 14122 8874 14122 8874 0 net192
rlabel metal1 32292 6426 32292 6426 0 net193
rlabel metal1 7820 4794 7820 4794 0 net194
rlabel metal2 17894 5933 17894 5933 0 net195
rlabel metal3 13524 6800 13524 6800 0 net196
rlabel metal1 35604 6426 35604 6426 0 net197
rlabel metal2 7406 7565 7406 7565 0 net198
rlabel metal1 15410 7514 15410 7514 0 net199
rlabel metal1 1978 3978 1978 3978 0 net2
rlabel metal2 4462 7038 4462 7038 0 net20
rlabel metal1 11500 5338 11500 5338 0 net200
rlabel metal2 2622 5439 2622 5439 0 net201
rlabel metal1 5842 6630 5842 6630 0 net202
rlabel metal2 11362 8874 11362 8874 0 net203
rlabel metal2 30314 1921 30314 1921 0 net204
rlabel metal2 12834 5474 12834 5474 0 net205
rlabel metal1 17526 3910 17526 3910 0 net206
rlabel metal2 7406 8687 7406 8687 0 net207
rlabel metal1 5336 3162 5336 3162 0 net208
rlabel metal2 14674 6596 14674 6596 0 net209
rlabel via2 6854 7939 6854 7939 0 net21
rlabel metal2 19550 1836 19550 1836 0 net210
rlabel metal2 9522 8891 9522 8891 0 net211
rlabel metal1 15410 3706 15410 3706 0 net212
rlabel metal1 16100 6970 16100 6970 0 net213
rlabel metal1 11316 6970 11316 6970 0 net214
rlabel metal2 12742 9180 12742 9180 0 net215
rlabel metal1 11316 5542 11316 5542 0 net216
rlabel via2 2346 3995 2346 3995 0 net217
rlabel metal2 5382 8296 5382 8296 0 net218
rlabel metal1 16744 7514 16744 7514 0 net219
rlabel metal3 14812 6392 14812 6392 0 net22
rlabel metal2 31326 3111 31326 3111 0 net220
rlabel metal2 9798 3264 9798 3264 0 net221
rlabel metal1 18998 3706 18998 3706 0 net222
rlabel metal2 13846 8126 13846 8126 0 net223
rlabel metal2 5198 5525 5198 5525 0 net224
rlabel metal2 13294 8636 13294 8636 0 net225
rlabel metal2 13386 8840 13386 8840 0 net226
rlabel metal2 13662 8415 13662 8415 0 net227
rlabel metal1 17066 3366 17066 3366 0 net228
rlabel metal1 16100 7174 16100 7174 0 net229
rlabel metal1 4968 2414 4968 2414 0 net23
rlabel metal2 13570 8704 13570 8704 0 net230
rlabel metal1 28106 6630 28106 6630 0 net231
rlabel metal1 36708 3978 36708 3978 0 net232
rlabel metal1 17250 8398 17250 8398 0 net233
rlabel metal2 12926 5882 12926 5882 0 net24
rlabel metal2 9522 5491 9522 5491 0 net25
rlabel metal1 19780 2414 19780 2414 0 net26
rlabel metal2 2714 1972 2714 1972 0 net27
rlabel metal2 2530 1972 2530 1972 0 net28
rlabel metal1 5290 3706 5290 3706 0 net29
rlabel metal2 1886 5508 1886 5508 0 net3
rlabel metal1 2300 3570 2300 3570 0 net30
rlabel metal1 7774 7344 7774 7344 0 net31
rlabel metal1 10442 7378 10442 7378 0 net32
rlabel metal2 1702 2176 1702 2176 0 net33
rlabel metal1 10626 2278 10626 2278 0 net34
rlabel metal1 17710 3570 17710 3570 0 net35
rlabel metal1 29716 4658 29716 4658 0 net36
rlabel metal1 34132 3502 34132 3502 0 net37
rlabel metal2 4922 2720 4922 2720 0 net38
rlabel metal4 20516 7956 20516 7956 0 net39
rlabel metal2 13110 4352 13110 4352 0 net4
rlabel metal1 17526 4590 17526 4590 0 net40
rlabel metal1 33396 2618 33396 2618 0 net41
rlabel metal2 14398 5236 14398 5236 0 net42
rlabel metal1 7866 6766 7866 6766 0 net43
rlabel metal1 19274 8330 19274 8330 0 net44
rlabel metal2 31786 7157 31786 7157 0 net45
rlabel metal1 35236 4454 35236 4454 0 net46
rlabel metal2 9706 2142 9706 2142 0 net47
rlabel metal2 16882 3400 16882 3400 0 net48
rlabel metal1 10304 2618 10304 2618 0 net49
rlabel metal2 1610 4896 1610 4896 0 net5
rlabel metal2 12006 2091 12006 2091 0 net50
rlabel metal1 12742 2618 12742 2618 0 net51
rlabel metal1 31004 2278 31004 2278 0 net52
rlabel metal2 17618 7633 17618 7633 0 net53
rlabel metal1 5888 7310 5888 7310 0 net54
rlabel metal3 5658 2652 5658 2652 0 net55
rlabel metal2 9798 1955 9798 1955 0 net56
rlabel metal2 12466 5729 12466 5729 0 net57
rlabel metal2 14766 2213 14766 2213 0 net58
rlabel metal1 17066 2550 17066 2550 0 net59
rlabel metal1 14582 5678 14582 5678 0 net6
rlabel metal2 17434 6902 17434 6902 0 net60
rlabel metal2 12650 3570 12650 3570 0 net61
rlabel metal2 18538 6698 18538 6698 0 net62
rlabel metal1 22586 7956 22586 7956 0 net63
rlabel metal2 14858 7055 14858 7055 0 net64
rlabel metal2 16054 2907 16054 2907 0 net65
rlabel metal1 32062 5576 32062 5576 0 net66
rlabel via1 21114 6069 21114 6069 0 net67
rlabel metal2 17250 6528 17250 6528 0 net68
rlabel metal2 13018 9996 13018 9996 0 net69
rlabel metal1 1886 5576 1886 5576 0 net7
rlabel metal2 24886 8942 24886 8942 0 net70
rlabel metal1 23920 8330 23920 8330 0 net71
rlabel viali 19366 4585 19366 4585 0 net72
rlabel metal1 11362 2414 11362 2414 0 net73
rlabel metal2 32246 4233 32246 4233 0 net74
rlabel metal1 22448 7922 22448 7922 0 net75
rlabel metal1 20056 7922 20056 7922 0 net76
rlabel metal3 14444 4488 14444 4488 0 net77
rlabel metal1 30268 7378 30268 7378 0 net78
rlabel metal2 13754 5440 13754 5440 0 net79
rlabel metal2 1610 6256 1610 6256 0 net8
rlabel metal1 19182 4182 19182 4182 0 net80
rlabel metal2 27738 8211 27738 8211 0 net81
rlabel metal1 26634 4182 26634 4182 0 net82
rlabel metal1 20712 7922 20712 7922 0 net83
rlabel metal2 20562 3604 20562 3604 0 net84
rlabel metal1 31418 6290 31418 6290 0 net85
rlabel metal1 28704 8262 28704 8262 0 net86
rlabel metal1 11270 3536 11270 3536 0 net87
rlabel metal1 28658 6936 28658 6936 0 net88
rlabel metal1 23713 7922 23713 7922 0 net89
rlabel via2 1702 6205 1702 6205 0 net9
rlabel metal2 25806 8874 25806 8874 0 net90
rlabel metal3 14628 5100 14628 5100 0 net91
rlabel metal1 28290 5542 28290 5542 0 net92
rlabel metal1 15847 6222 15847 6222 0 net93
rlabel metal1 26864 8262 26864 8262 0 net94
rlabel metal1 17572 2278 17572 2278 0 net95
rlabel metal2 20286 4420 20286 4420 0 net96
rlabel metal2 32706 4896 32706 4896 0 net97
rlabel metal1 26220 4590 26220 4590 0 net98
rlabel metal2 21022 6817 21022 6817 0 net99
<< properties >>
string FIXED_BBOX 0 0 41000 11250
<< end >>
