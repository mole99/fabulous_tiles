magic
tech sky130A
magscale 1 2
timestamp 1740383593
<< viali >>
rect 3525 8585 3559 8619
rect 4261 8585 4295 8619
rect 4629 8585 4663 8619
rect 4905 8585 4939 8619
rect 5273 8585 5307 8619
rect 5641 8585 5675 8619
rect 6009 8585 6043 8619
rect 6745 8585 6779 8619
rect 7113 8585 7147 8619
rect 7481 8585 7515 8619
rect 7849 8585 7883 8619
rect 8217 8585 8251 8619
rect 8585 8585 8619 8619
rect 9321 8585 9355 8619
rect 9781 8585 9815 8619
rect 10149 8585 10183 8619
rect 10425 8585 10459 8619
rect 10793 8585 10827 8619
rect 11161 8585 11195 8619
rect 11897 8585 11931 8619
rect 12265 8585 12299 8619
rect 12633 8585 12667 8619
rect 13001 8585 13035 8619
rect 13369 8585 13403 8619
rect 13737 8585 13771 8619
rect 14473 8585 14507 8619
rect 14841 8585 14875 8619
rect 15209 8585 15243 8619
rect 15577 8585 15611 8619
rect 15945 8585 15979 8619
rect 16313 8585 16347 8619
rect 16957 8585 16991 8619
rect 17601 8585 17635 8619
rect 17877 8585 17911 8619
rect 32321 8585 32355 8619
rect 32781 8585 32815 8619
rect 33149 8585 33183 8619
rect 33517 8585 33551 8619
rect 33885 8585 33919 8619
rect 34253 8585 34287 8619
rect 35541 8585 35575 8619
rect 36737 8585 36771 8619
rect 37841 8585 37875 8619
rect 38577 8585 38611 8619
rect 2973 8449 3007 8483
rect 3341 8449 3375 8483
rect 4077 8449 4111 8483
rect 4445 8449 4479 8483
rect 5089 8449 5123 8483
rect 5457 8449 5491 8483
rect 5825 8449 5859 8483
rect 6193 8449 6227 8483
rect 6929 8449 6963 8483
rect 7297 8449 7331 8483
rect 7665 8449 7699 8483
rect 8033 8449 8067 8483
rect 8401 8449 8435 8483
rect 8769 8449 8803 8483
rect 9505 8449 9539 8483
rect 9597 8449 9631 8483
rect 9965 8449 9999 8483
rect 10609 8449 10643 8483
rect 10977 8449 11011 8483
rect 11345 8449 11379 8483
rect 12081 8449 12115 8483
rect 12449 8449 12483 8483
rect 12817 8449 12851 8483
rect 13185 8449 13219 8483
rect 13553 8449 13587 8483
rect 13921 8449 13955 8483
rect 14657 8449 14691 8483
rect 15025 8449 15059 8483
rect 15393 8449 15427 8483
rect 15761 8449 15795 8483
rect 16129 8449 16163 8483
rect 16497 8449 16531 8483
rect 17141 8449 17175 8483
rect 17417 8449 17451 8483
rect 18061 8449 18095 8483
rect 32505 8449 32539 8483
rect 32597 8449 32631 8483
rect 32965 8449 32999 8483
rect 33333 8449 33367 8483
rect 33701 8449 33735 8483
rect 34069 8449 34103 8483
rect 34713 8449 34747 8483
rect 35081 8449 35115 8483
rect 35725 8449 35759 8483
rect 35817 8449 35851 8483
rect 36185 8449 36219 8483
rect 36553 8449 36587 8483
rect 37289 8449 37323 8483
rect 37657 8449 37691 8483
rect 38025 8449 38059 8483
rect 38393 8449 38427 8483
rect 38853 8449 38887 8483
rect 39221 8449 39255 8483
rect 18153 8381 18187 8415
rect 3157 8313 3191 8347
rect 34897 8313 34931 8347
rect 36001 8313 36035 8347
rect 38209 8313 38243 8347
rect 39037 8313 39071 8347
rect 39405 8313 39439 8347
rect 35265 8245 35299 8279
rect 36369 8245 36403 8279
rect 37473 8245 37507 8279
rect 3525 8041 3559 8075
rect 4353 8041 4387 8075
rect 5181 8041 5215 8075
rect 6193 8041 6227 8075
rect 6837 8041 6871 8075
rect 7297 8041 7331 8075
rect 8401 8041 8435 8075
rect 9045 8041 9079 8075
rect 9505 8041 9539 8075
rect 10609 8041 10643 8075
rect 11437 8041 11471 8075
rect 11805 8041 11839 8075
rect 12817 8041 12851 8075
rect 13645 8041 13679 8075
rect 14105 8041 14139 8075
rect 14473 8041 14507 8075
rect 15669 8041 15703 8075
rect 16129 8041 16163 8075
rect 19717 8041 19751 8075
rect 21005 8041 21039 8075
rect 21833 8041 21867 8075
rect 23121 8041 23155 8075
rect 23489 8041 23523 8075
rect 31033 8041 31067 8075
rect 34805 8041 34839 8075
rect 35817 8041 35851 8075
rect 36369 8041 36403 8075
rect 36921 8041 36955 8075
rect 37933 8041 37967 8075
rect 38669 8041 38703 8075
rect 8125 7973 8159 8007
rect 12265 7973 12299 8007
rect 13277 7973 13311 8007
rect 15209 7973 15243 8007
rect 22201 7973 22235 8007
rect 4077 7905 4111 7939
rect 3341 7837 3375 7871
rect 4169 7837 4203 7871
rect 4997 7837 5031 7871
rect 6377 7837 6411 7871
rect 6653 7837 6687 7871
rect 7481 7837 7515 7871
rect 7849 7837 7883 7871
rect 7941 7837 7975 7871
rect 8585 7837 8619 7871
rect 9229 7837 9263 7871
rect 9689 7837 9723 7871
rect 9781 7837 9815 7871
rect 10793 7837 10827 7871
rect 11621 7837 11655 7871
rect 11989 7837 12023 7871
rect 12173 7837 12207 7871
rect 12449 7837 12483 7871
rect 13001 7837 13035 7871
rect 13461 7837 13495 7871
rect 13829 7837 13863 7871
rect 14289 7837 14323 7871
rect 14657 7837 14691 7871
rect 15209 7837 15243 7871
rect 15301 7837 15335 7871
rect 15853 7837 15887 7871
rect 16313 7837 16347 7871
rect 17785 7837 17819 7871
rect 19257 7837 19291 7871
rect 19533 7837 19567 7871
rect 19901 7837 19935 7871
rect 21097 7837 21131 7871
rect 21189 7837 21223 7871
rect 21925 7837 21959 7871
rect 22017 7837 22051 7871
rect 23305 7837 23339 7871
rect 23673 7837 23707 7871
rect 27721 7837 27755 7871
rect 31217 7837 31251 7871
rect 33241 7837 33275 7871
rect 34989 7837 35023 7871
rect 35515 7837 35549 7871
rect 35633 7837 35667 7871
rect 36185 7837 36219 7871
rect 36737 7837 36771 7871
rect 38117 7837 38151 7871
rect 38485 7837 38519 7871
rect 38853 7837 38887 7871
rect 39221 7837 39255 7871
rect 3893 7769 3927 7803
rect 7849 7701 7883 7735
rect 9965 7701 9999 7735
rect 15485 7701 15519 7735
rect 17601 7701 17635 7735
rect 19441 7701 19475 7735
rect 21373 7701 21407 7735
rect 27629 7701 27663 7735
rect 27905 7701 27939 7735
rect 33057 7701 33091 7735
rect 35357 7701 35391 7735
rect 39037 7701 39071 7735
rect 39405 7701 39439 7735
rect 2789 7497 2823 7531
rect 9597 7497 9631 7531
rect 14197 7497 14231 7531
rect 21189 7497 21223 7531
rect 23765 7497 23799 7531
rect 38301 7497 38335 7531
rect 38669 7497 38703 7531
rect 39037 7497 39071 7531
rect 14841 7429 14875 7463
rect 2605 7361 2639 7395
rect 7665 7361 7699 7395
rect 9321 7361 9355 7395
rect 9781 7361 9815 7395
rect 14105 7361 14139 7395
rect 14381 7361 14415 7395
rect 14657 7361 14691 7395
rect 14749 7361 14783 7395
rect 16037 7361 16071 7395
rect 17702 7361 17736 7395
rect 21373 7361 21407 7395
rect 23949 7361 23983 7395
rect 31217 7361 31251 7395
rect 37749 7361 37783 7395
rect 38117 7361 38151 7395
rect 38485 7361 38519 7395
rect 38853 7361 38887 7395
rect 39221 7361 39255 7395
rect 17601 7293 17635 7327
rect 9505 7225 9539 7259
rect 14473 7225 14507 7259
rect 15853 7225 15887 7259
rect 17877 7225 17911 7259
rect 7849 7157 7883 7191
rect 14105 7157 14139 7191
rect 31033 7157 31067 7191
rect 37933 7157 37967 7191
rect 39405 7157 39439 7191
rect 22661 6885 22695 6919
rect 2605 6749 2639 6783
rect 2697 6749 2731 6783
rect 9321 6749 9355 6783
rect 9597 6749 9631 6783
rect 22477 6749 22511 6783
rect 25605 6749 25639 6783
rect 30021 6749 30055 6783
rect 34253 6749 34287 6783
rect 38485 6749 38519 6783
rect 38853 6749 38887 6783
rect 39221 6749 39255 6783
rect 2881 6613 2915 6647
rect 9413 6613 9447 6647
rect 25421 6613 25455 6647
rect 29837 6613 29871 6647
rect 34069 6613 34103 6647
rect 38669 6613 38703 6647
rect 39037 6613 39071 6647
rect 39405 6613 39439 6647
rect 3249 6409 3283 6443
rect 3617 6409 3651 6443
rect 4445 6409 4479 6443
rect 7665 6409 7699 6443
rect 8309 6409 8343 6443
rect 10609 6409 10643 6443
rect 11621 6409 11655 6443
rect 26433 6409 26467 6443
rect 29285 6409 29319 6443
rect 39405 6409 39439 6443
rect 2973 6341 3007 6375
rect 3801 6341 3835 6375
rect 3065 6273 3099 6307
rect 3433 6273 3467 6307
rect 3709 6273 3743 6307
rect 4629 6273 4663 6307
rect 7849 6273 7883 6307
rect 8125 6273 8159 6307
rect 8493 6273 8527 6307
rect 8769 6273 8803 6307
rect 10793 6273 10827 6307
rect 11805 6273 11839 6307
rect 19165 6273 19199 6307
rect 19349 6273 19383 6307
rect 24225 6273 24259 6307
rect 26617 6273 26651 6307
rect 29469 6273 29503 6307
rect 38853 6273 38887 6307
rect 39221 6273 39255 6307
rect 8585 6137 8619 6171
rect 19533 6137 19567 6171
rect 24409 6137 24443 6171
rect 39037 6069 39071 6103
rect 3985 5865 4019 5899
rect 4905 5865 4939 5899
rect 5549 5865 5583 5899
rect 6653 5865 6687 5899
rect 7113 5865 7147 5899
rect 11621 5865 11655 5899
rect 26065 5865 26099 5899
rect 35449 5865 35483 5899
rect 37013 5865 37047 5899
rect 38117 5865 38151 5899
rect 39405 5797 39439 5831
rect 4169 5729 4203 5763
rect 3801 5661 3835 5695
rect 4077 5661 4111 5695
rect 5089 5661 5123 5695
rect 5733 5661 5767 5695
rect 6837 5661 6871 5695
rect 7297 5661 7331 5695
rect 11805 5661 11839 5695
rect 18429 5661 18463 5695
rect 18521 5661 18555 5695
rect 25881 5661 25915 5695
rect 28273 5661 28307 5695
rect 35265 5661 35299 5695
rect 35633 5661 35667 5695
rect 37197 5661 37231 5695
rect 38301 5661 38335 5695
rect 38853 5661 38887 5695
rect 39221 5661 39255 5695
rect 18337 5525 18371 5559
rect 18705 5525 18739 5559
rect 28089 5525 28123 5559
rect 35817 5525 35851 5559
rect 39037 5525 39071 5559
rect 5365 5321 5399 5355
rect 5825 5321 5859 5355
rect 13001 5321 13035 5355
rect 15853 5321 15887 5355
rect 16865 5321 16899 5355
rect 39405 5321 39439 5355
rect 5549 5185 5583 5219
rect 5641 5185 5675 5219
rect 13185 5185 13219 5219
rect 16037 5185 16071 5219
rect 16681 5185 16715 5219
rect 16957 5185 16991 5219
rect 17325 5185 17359 5219
rect 17877 5185 17911 5219
rect 22017 5185 22051 5219
rect 27169 5185 27203 5219
rect 38853 5185 38887 5219
rect 39221 5185 39255 5219
rect 17141 5049 17175 5083
rect 18061 5049 18095 5083
rect 21833 4981 21867 5015
rect 26985 4981 27019 5015
rect 39037 4981 39071 5015
rect 14657 4777 14691 4811
rect 16313 4777 16347 4811
rect 16681 4777 16715 4811
rect 18705 4777 18739 4811
rect 33793 4777 33827 4811
rect 11069 4709 11103 4743
rect 23765 4709 23799 4743
rect 24133 4709 24167 4743
rect 39405 4709 39439 4743
rect 11069 4573 11103 4607
rect 11253 4573 11287 4607
rect 14841 4573 14875 4607
rect 16405 4573 16439 4607
rect 16497 4573 16531 4607
rect 18797 4573 18831 4607
rect 18889 4573 18923 4607
rect 20361 4573 20395 4607
rect 23581 4573 23615 4607
rect 23949 4573 23983 4607
rect 28181 4573 28215 4607
rect 31861 4573 31895 4607
rect 33609 4573 33643 4607
rect 38853 4573 38887 4607
rect 39221 4573 39255 4607
rect 11437 4505 11471 4539
rect 19073 4437 19107 4471
rect 20545 4437 20579 4471
rect 28365 4437 28399 4471
rect 32045 4437 32079 4471
rect 39037 4437 39071 4471
rect 13829 4233 13863 4267
rect 5733 4165 5767 4199
rect 9781 4165 9815 4199
rect 13645 4097 13679 4131
rect 23029 4097 23063 4131
rect 23213 4097 23247 4131
rect 30297 4097 30331 4131
rect 36461 4097 36495 4131
rect 38853 4097 38887 4131
rect 39221 4097 39255 4131
rect 9965 3961 9999 3995
rect 39405 3961 39439 3995
rect 5825 3893 5859 3927
rect 23397 3893 23431 3927
rect 30481 3893 30515 3927
rect 36277 3893 36311 3927
rect 39037 3893 39071 3927
rect 14749 3621 14783 3655
rect 20269 3621 20303 3655
rect 39405 3621 39439 3655
rect 11161 3553 11195 3587
rect 10977 3485 11011 3519
rect 14841 3485 14875 3519
rect 14933 3485 14967 3519
rect 17601 3485 17635 3519
rect 20361 3485 20395 3519
rect 20453 3485 20487 3519
rect 29929 3485 29963 3519
rect 38853 3485 38887 3519
rect 39221 3485 39255 3519
rect 15117 3349 15151 3383
rect 17417 3349 17451 3383
rect 20637 3349 20671 3383
rect 30113 3349 30147 3383
rect 39037 3349 39071 3383
rect 18061 3145 18095 3179
rect 18429 3145 18463 3179
rect 20729 3145 20763 3179
rect 21557 3145 21591 3179
rect 33333 3145 33367 3179
rect 33701 3145 33735 3179
rect 39405 3145 39439 3179
rect 8861 3009 8895 3043
rect 13093 3009 13127 3043
rect 13185 3009 13219 3043
rect 15945 3009 15979 3043
rect 16037 3009 16071 3043
rect 16773 3009 16807 3043
rect 18153 3009 18187 3043
rect 18245 3009 18279 3043
rect 20729 3009 20763 3043
rect 20821 3009 20855 3043
rect 21373 3009 21407 3043
rect 23765 3009 23799 3043
rect 23949 3009 23983 3043
rect 24225 3009 24259 3043
rect 24685 3009 24719 3043
rect 24777 3009 24811 3043
rect 26985 3009 27019 3043
rect 28089 3009 28123 3043
rect 28549 3009 28583 3043
rect 28641 3009 28675 3043
rect 30113 3009 30147 3043
rect 30205 3009 30239 3043
rect 33425 3009 33459 3043
rect 33517 3009 33551 3043
rect 38853 3009 38887 3043
rect 39221 3009 39255 3043
rect 17049 2941 17083 2975
rect 9045 2873 9079 2907
rect 15853 2873 15887 2907
rect 16957 2873 16991 2907
rect 21005 2873 21039 2907
rect 24133 2873 24167 2907
rect 13001 2805 13035 2839
rect 13369 2805 13403 2839
rect 16221 2805 16255 2839
rect 24409 2805 24443 2839
rect 24593 2805 24627 2839
rect 24961 2805 24995 2839
rect 27169 2805 27203 2839
rect 28273 2805 28307 2839
rect 28457 2805 28491 2839
rect 28825 2805 28859 2839
rect 30021 2805 30055 2839
rect 30389 2805 30423 2839
rect 39037 2805 39071 2839
rect 39405 2533 39439 2567
rect 37737 2397 37771 2431
rect 38117 2397 38151 2431
rect 38485 2397 38519 2431
rect 38853 2397 38887 2431
rect 39221 2397 39255 2431
rect 37933 2261 37967 2295
rect 38301 2261 38335 2295
rect 38669 2261 38703 2295
rect 39037 2261 39071 2295
<< metal1 >>
rect 7282 11160 7288 11212
rect 7340 11200 7346 11212
rect 27798 11200 27804 11212
rect 7340 11172 27804 11200
rect 7340 11160 7346 11172
rect 27798 11160 27804 11172
rect 27856 11160 27862 11212
rect 6362 11092 6368 11144
rect 6420 11132 6426 11144
rect 18414 11132 18420 11144
rect 6420 11104 18420 11132
rect 6420 11092 6426 11104
rect 18414 11092 18420 11104
rect 18472 11092 18478 11144
rect 16390 10956 16396 11008
rect 16448 10996 16454 11008
rect 22278 10996 22284 11008
rect 16448 10968 22284 10996
rect 16448 10956 16454 10968
rect 22278 10956 22284 10968
rect 22336 10956 22342 11008
rect 16942 10004 16948 10056
rect 17000 10044 17006 10056
rect 23934 10044 23940 10056
rect 17000 10016 23940 10044
rect 17000 10004 17006 10016
rect 23934 10004 23940 10016
rect 23992 10004 23998 10056
rect 13814 9868 13820 9920
rect 13872 9908 13878 9920
rect 18690 9908 18696 9920
rect 13872 9880 18696 9908
rect 13872 9868 13878 9880
rect 18690 9868 18696 9880
rect 18748 9868 18754 9920
rect 19334 9596 19340 9648
rect 19392 9636 19398 9648
rect 24762 9636 24768 9648
rect 19392 9608 24768 9636
rect 19392 9596 19398 9608
rect 24762 9596 24768 9608
rect 24820 9596 24826 9648
rect 1118 9528 1124 9580
rect 1176 9568 1182 9580
rect 23842 9568 23848 9580
rect 1176 9540 23848 9568
rect 1176 9528 1182 9540
rect 23842 9528 23848 9540
rect 23900 9528 23906 9580
rect 17954 9460 17960 9512
rect 18012 9500 18018 9512
rect 24210 9500 24216 9512
rect 18012 9472 24216 9500
rect 18012 9460 18018 9472
rect 24210 9460 24216 9472
rect 24268 9460 24274 9512
rect 1302 9392 1308 9444
rect 1360 9432 1366 9444
rect 26510 9432 26516 9444
rect 1360 9404 26516 9432
rect 1360 9392 1366 9404
rect 26510 9392 26516 9404
rect 26568 9392 26574 9444
rect 13354 9324 13360 9376
rect 13412 9364 13418 9376
rect 17862 9364 17868 9376
rect 13412 9336 17868 9364
rect 13412 9324 13418 9336
rect 17862 9324 17868 9336
rect 17920 9324 17926 9376
rect 22738 9324 22744 9376
rect 22796 9364 22802 9376
rect 36538 9364 36544 9376
rect 22796 9336 36544 9364
rect 22796 9324 22802 9336
rect 36538 9324 36544 9336
rect 36596 9324 36602 9376
rect 15746 9256 15752 9308
rect 15804 9296 15810 9308
rect 26418 9296 26424 9308
rect 15804 9268 26424 9296
rect 15804 9256 15810 9268
rect 26418 9256 26424 9268
rect 26476 9256 26482 9308
rect 8386 9188 8392 9240
rect 8444 9228 8450 9240
rect 17218 9228 17224 9240
rect 8444 9200 17224 9228
rect 8444 9188 8450 9200
rect 17218 9188 17224 9200
rect 17276 9188 17282 9240
rect 24026 9188 24032 9240
rect 24084 9228 24090 9240
rect 38930 9228 38936 9240
rect 24084 9200 38936 9228
rect 24084 9188 24090 9200
rect 38930 9188 38936 9200
rect 38988 9188 38994 9240
rect 198 9120 204 9172
rect 256 9160 262 9172
rect 23934 9160 23940 9172
rect 256 9132 23940 9160
rect 256 9120 262 9132
rect 23934 9120 23940 9132
rect 23992 9120 23998 9172
rect 19242 9092 19248 9104
rect 12406 9064 19248 9092
rect 10778 8984 10784 9036
rect 10836 9024 10842 9036
rect 12406 9024 12434 9064
rect 19242 9052 19248 9064
rect 19300 9052 19306 9104
rect 19610 9052 19616 9104
rect 19668 9092 19674 9104
rect 20622 9092 20628 9104
rect 19668 9064 20628 9092
rect 19668 9052 19674 9064
rect 20622 9052 20628 9064
rect 20680 9052 20686 9104
rect 21726 9052 21732 9104
rect 21784 9092 21790 9104
rect 28074 9092 28080 9104
rect 21784 9064 28080 9092
rect 21784 9052 21790 9064
rect 28074 9052 28080 9064
rect 28132 9052 28138 9104
rect 10836 8996 12434 9024
rect 10836 8984 10842 8996
rect 15562 8984 15568 9036
rect 15620 9024 15626 9036
rect 22922 9024 22928 9036
rect 15620 8996 22928 9024
rect 15620 8984 15626 8996
rect 22922 8984 22928 8996
rect 22980 8984 22986 9036
rect 33594 8984 33600 9036
rect 33652 9024 33658 9036
rect 34238 9024 34244 9036
rect 33652 8996 34244 9024
rect 33652 8984 33658 8996
rect 34238 8984 34244 8996
rect 34296 8984 34302 9036
rect 8662 8916 8668 8968
rect 8720 8956 8726 8968
rect 8720 8928 12434 8956
rect 8720 8916 8726 8928
rect 12406 8888 12434 8928
rect 12802 8916 12808 8968
rect 12860 8956 12866 8968
rect 19702 8956 19708 8968
rect 12860 8928 19708 8956
rect 12860 8916 12866 8928
rect 19702 8916 19708 8928
rect 19760 8916 19766 8968
rect 19794 8916 19800 8968
rect 19852 8956 19858 8968
rect 32582 8956 32588 8968
rect 19852 8928 32588 8956
rect 19852 8916 19858 8928
rect 32582 8916 32588 8928
rect 32640 8916 32646 8968
rect 37274 8956 37280 8968
rect 32876 8928 37280 8956
rect 15838 8888 15844 8900
rect 12406 8860 15844 8888
rect 15838 8848 15844 8860
rect 15896 8848 15902 8900
rect 17034 8848 17040 8900
rect 17092 8888 17098 8900
rect 17862 8888 17868 8900
rect 17092 8860 17868 8888
rect 17092 8848 17098 8860
rect 17862 8848 17868 8860
rect 17920 8848 17926 8900
rect 30742 8848 30748 8900
rect 30800 8888 30806 8900
rect 32876 8888 32904 8928
rect 37274 8916 37280 8928
rect 37332 8916 37338 8968
rect 36170 8888 36176 8900
rect 30800 8860 32904 8888
rect 32968 8860 36176 8888
rect 30800 8848 30806 8860
rect 11330 8780 11336 8832
rect 11388 8820 11394 8832
rect 16022 8820 16028 8832
rect 11388 8792 16028 8820
rect 11388 8780 11394 8792
rect 16022 8780 16028 8792
rect 16080 8780 16086 8832
rect 16114 8780 16120 8832
rect 16172 8820 16178 8832
rect 23474 8820 23480 8832
rect 16172 8792 23480 8820
rect 16172 8780 16178 8792
rect 23474 8780 23480 8792
rect 23532 8780 23538 8832
rect 24578 8780 24584 8832
rect 24636 8820 24642 8832
rect 27246 8820 27252 8832
rect 24636 8792 27252 8820
rect 24636 8780 24642 8792
rect 27246 8780 27252 8792
rect 27304 8780 27310 8832
rect 29914 8780 29920 8832
rect 29972 8820 29978 8832
rect 32968 8820 32996 8860
rect 36170 8848 36176 8860
rect 36228 8848 36234 8900
rect 29972 8792 32996 8820
rect 29972 8780 29978 8792
rect 33042 8780 33048 8832
rect 33100 8820 33106 8832
rect 33502 8820 33508 8832
rect 33100 8792 33508 8820
rect 33100 8780 33106 8792
rect 33502 8780 33508 8792
rect 33560 8780 33566 8832
rect 33778 8780 33784 8832
rect 33836 8820 33842 8832
rect 38010 8820 38016 8832
rect 33836 8792 38016 8820
rect 33836 8780 33842 8792
rect 38010 8780 38016 8792
rect 38068 8780 38074 8832
rect 1104 8730 39836 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 39010 8730
rect 39062 8678 39074 8730
rect 39126 8678 39138 8730
rect 39190 8678 39202 8730
rect 39254 8678 39266 8730
rect 39318 8678 39836 8730
rect 1104 8656 39836 8678
rect 3513 8619 3571 8625
rect 3513 8585 3525 8619
rect 3559 8616 3571 8619
rect 3786 8616 3792 8628
rect 3559 8588 3792 8616
rect 3559 8585 3571 8588
rect 3513 8579 3571 8585
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8616 4307 8619
rect 4338 8616 4344 8628
rect 4295 8588 4344 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 4614 8576 4620 8628
rect 4672 8576 4678 8628
rect 4893 8619 4951 8625
rect 4893 8585 4905 8619
rect 4939 8616 4951 8619
rect 5166 8616 5172 8628
rect 4939 8588 5172 8616
rect 4939 8585 4951 8588
rect 4893 8579 4951 8585
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5261 8619 5319 8625
rect 5261 8585 5273 8619
rect 5307 8616 5319 8619
rect 5442 8616 5448 8628
rect 5307 8588 5448 8616
rect 5307 8585 5319 8588
rect 5261 8579 5319 8585
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8616 5687 8619
rect 5718 8616 5724 8628
rect 5675 8588 5724 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 5718 8576 5724 8588
rect 5776 8576 5782 8628
rect 5997 8619 6055 8625
rect 5997 8585 6009 8619
rect 6043 8616 6055 8619
rect 6270 8616 6276 8628
rect 6043 8588 6276 8616
rect 6043 8585 6055 8588
rect 5997 8579 6055 8585
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 6733 8619 6791 8625
rect 6733 8585 6745 8619
rect 6779 8616 6791 8619
rect 6822 8616 6828 8628
rect 6779 8588 6828 8616
rect 6779 8585 6791 8588
rect 6733 8579 6791 8585
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 7101 8619 7159 8625
rect 7101 8585 7113 8619
rect 7147 8616 7159 8619
rect 7374 8616 7380 8628
rect 7147 8588 7380 8616
rect 7147 8585 7159 8588
rect 7101 8579 7159 8585
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 7469 8619 7527 8625
rect 7469 8585 7481 8619
rect 7515 8616 7527 8619
rect 7650 8616 7656 8628
rect 7515 8588 7656 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 7650 8576 7656 8588
rect 7708 8576 7714 8628
rect 7837 8619 7895 8625
rect 7837 8585 7849 8619
rect 7883 8616 7895 8619
rect 7926 8616 7932 8628
rect 7883 8588 7932 8616
rect 7883 8585 7895 8588
rect 7837 8579 7895 8585
rect 7926 8576 7932 8588
rect 7984 8576 7990 8628
rect 8205 8619 8263 8625
rect 8205 8585 8217 8619
rect 8251 8616 8263 8619
rect 8478 8616 8484 8628
rect 8251 8588 8484 8616
rect 8251 8585 8263 8588
rect 8205 8579 8263 8585
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 8573 8619 8631 8625
rect 8573 8585 8585 8619
rect 8619 8616 8631 8619
rect 8846 8616 8852 8628
rect 8619 8588 8852 8616
rect 8619 8585 8631 8588
rect 8573 8579 8631 8585
rect 8846 8576 8852 8588
rect 8904 8576 8910 8628
rect 9309 8619 9367 8625
rect 9309 8585 9321 8619
rect 9355 8616 9367 8619
rect 9582 8616 9588 8628
rect 9355 8588 9588 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 9769 8619 9827 8625
rect 9769 8585 9781 8619
rect 9815 8616 9827 8619
rect 9858 8616 9864 8628
rect 9815 8588 9864 8616
rect 9815 8585 9827 8588
rect 9769 8579 9827 8585
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 10134 8576 10140 8628
rect 10192 8576 10198 8628
rect 10413 8619 10471 8625
rect 10413 8585 10425 8619
rect 10459 8616 10471 8619
rect 10686 8616 10692 8628
rect 10459 8588 10692 8616
rect 10459 8585 10471 8588
rect 10413 8579 10471 8585
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 10781 8619 10839 8625
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 10962 8616 10968 8628
rect 10827 8588 10968 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11149 8619 11207 8625
rect 11149 8585 11161 8619
rect 11195 8616 11207 8619
rect 11514 8616 11520 8628
rect 11195 8588 11520 8616
rect 11195 8585 11207 8588
rect 11149 8579 11207 8585
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 11885 8619 11943 8625
rect 11885 8585 11897 8619
rect 11931 8616 11943 8619
rect 12066 8616 12072 8628
rect 11931 8588 12072 8616
rect 11931 8585 11943 8588
rect 11885 8579 11943 8585
rect 12066 8576 12072 8588
rect 12124 8576 12130 8628
rect 12253 8619 12311 8625
rect 12253 8585 12265 8619
rect 12299 8616 12311 8619
rect 12342 8616 12348 8628
rect 12299 8588 12348 8616
rect 12299 8585 12311 8588
rect 12253 8579 12311 8585
rect 12342 8576 12348 8588
rect 12400 8576 12406 8628
rect 12621 8619 12679 8625
rect 12621 8585 12633 8619
rect 12667 8616 12679 8619
rect 12894 8616 12900 8628
rect 12667 8588 12900 8616
rect 12667 8585 12679 8588
rect 12621 8579 12679 8585
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 12989 8619 13047 8625
rect 12989 8585 13001 8619
rect 13035 8616 13047 8619
rect 13170 8616 13176 8628
rect 13035 8588 13176 8616
rect 13035 8585 13047 8588
rect 12989 8579 13047 8585
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 13357 8619 13415 8625
rect 13357 8585 13369 8619
rect 13403 8616 13415 8619
rect 13630 8616 13636 8628
rect 13403 8588 13636 8616
rect 13403 8585 13415 8588
rect 13357 8579 13415 8585
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 13725 8619 13783 8625
rect 13725 8585 13737 8619
rect 13771 8616 13783 8619
rect 13998 8616 14004 8628
rect 13771 8588 14004 8616
rect 13771 8585 13783 8588
rect 13725 8579 13783 8585
rect 13998 8576 14004 8588
rect 14056 8576 14062 8628
rect 14461 8619 14519 8625
rect 14461 8585 14473 8619
rect 14507 8616 14519 8619
rect 14550 8616 14556 8628
rect 14507 8588 14556 8616
rect 14507 8585 14519 8588
rect 14461 8579 14519 8585
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 14829 8619 14887 8625
rect 14829 8585 14841 8619
rect 14875 8616 14887 8619
rect 14918 8616 14924 8628
rect 14875 8588 14924 8616
rect 14875 8585 14887 8588
rect 14829 8579 14887 8585
rect 14918 8576 14924 8588
rect 14976 8576 14982 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 15378 8616 15384 8628
rect 15243 8588 15384 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15565 8619 15623 8625
rect 15565 8585 15577 8619
rect 15611 8616 15623 8619
rect 15654 8616 15660 8628
rect 15611 8588 15660 8616
rect 15611 8585 15623 8588
rect 15565 8579 15623 8585
rect 15654 8576 15660 8588
rect 15712 8576 15718 8628
rect 15933 8619 15991 8625
rect 15933 8585 15945 8619
rect 15979 8616 15991 8619
rect 16206 8616 16212 8628
rect 15979 8588 16212 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 16301 8619 16359 8625
rect 16301 8585 16313 8619
rect 16347 8616 16359 8619
rect 16482 8616 16488 8628
rect 16347 8588 16488 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 16482 8576 16488 8588
rect 16540 8576 16546 8628
rect 16758 8576 16764 8628
rect 16816 8616 16822 8628
rect 16945 8619 17003 8625
rect 16945 8616 16957 8619
rect 16816 8588 16957 8616
rect 16816 8576 16822 8588
rect 16945 8585 16957 8588
rect 16991 8585 17003 8619
rect 16945 8579 17003 8585
rect 17310 8576 17316 8628
rect 17368 8616 17374 8628
rect 17589 8619 17647 8625
rect 17589 8616 17601 8619
rect 17368 8588 17601 8616
rect 17368 8576 17374 8588
rect 17589 8585 17601 8588
rect 17635 8585 17647 8619
rect 17589 8579 17647 8585
rect 17862 8576 17868 8628
rect 17920 8576 17926 8628
rect 18230 8616 18236 8628
rect 17972 8588 18236 8616
rect 14734 8548 14740 8560
rect 6196 8520 11192 8548
rect 2866 8440 2872 8492
rect 2924 8480 2930 8492
rect 2961 8483 3019 8489
rect 2961 8480 2973 8483
rect 2924 8452 2973 8480
rect 2924 8440 2930 8452
rect 2961 8449 2973 8452
rect 3007 8449 3019 8483
rect 2961 8443 3019 8449
rect 3329 8483 3387 8489
rect 3329 8449 3341 8483
rect 3375 8480 3387 8483
rect 3418 8480 3424 8492
rect 3375 8452 3424 8480
rect 3375 8449 3387 8452
rect 3329 8443 3387 8449
rect 3418 8440 3424 8452
rect 3476 8440 3482 8492
rect 4062 8440 4068 8492
rect 4120 8440 4126 8492
rect 4430 8440 4436 8492
rect 4488 8440 4494 8492
rect 5074 8440 5080 8492
rect 5132 8440 5138 8492
rect 5442 8440 5448 8492
rect 5500 8440 5506 8492
rect 5810 8440 5816 8492
rect 5868 8440 5874 8492
rect 6196 8489 6224 8520
rect 11164 8492 11192 8520
rect 13556 8520 14740 8548
rect 6181 8483 6239 8489
rect 6181 8449 6193 8483
rect 6227 8449 6239 8483
rect 6181 8443 6239 8449
rect 6914 8440 6920 8492
rect 6972 8440 6978 8492
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 7300 8412 7328 8443
rect 7558 8440 7564 8492
rect 7616 8480 7622 8492
rect 7653 8483 7711 8489
rect 7653 8480 7665 8483
rect 7616 8452 7665 8480
rect 7616 8440 7622 8452
rect 7653 8449 7665 8452
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 7834 8440 7840 8492
rect 7892 8480 7898 8492
rect 8021 8483 8079 8489
rect 8021 8480 8033 8483
rect 7892 8452 8033 8480
rect 7892 8440 7898 8452
rect 8021 8449 8033 8452
rect 8067 8449 8079 8483
rect 8021 8443 8079 8449
rect 8386 8440 8392 8492
rect 8444 8440 8450 8492
rect 8662 8440 8668 8492
rect 8720 8480 8726 8492
rect 8757 8483 8815 8489
rect 8757 8480 8769 8483
rect 8720 8452 8769 8480
rect 8720 8440 8726 8452
rect 8757 8449 8769 8452
rect 8803 8449 8815 8483
rect 8757 8443 8815 8449
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 9585 8483 9643 8489
rect 9585 8449 9597 8483
rect 9631 8449 9643 8483
rect 9585 8443 9643 8449
rect 7742 8412 7748 8424
rect 7300 8384 7748 8412
rect 7742 8372 7748 8384
rect 7800 8372 7806 8424
rect 8478 8372 8484 8424
rect 8536 8412 8542 8424
rect 9600 8412 9628 8443
rect 9950 8440 9956 8492
rect 10008 8440 10014 8492
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8480 10655 8483
rect 10870 8480 10876 8492
rect 10643 8452 10876 8480
rect 10643 8449 10655 8452
rect 10597 8443 10655 8449
rect 10870 8440 10876 8452
rect 10928 8440 10934 8492
rect 10962 8440 10968 8492
rect 11020 8440 11026 8492
rect 11146 8440 11152 8492
rect 11204 8440 11210 8492
rect 11330 8440 11336 8492
rect 11388 8440 11394 8492
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 8536 8384 9628 8412
rect 8536 8372 8542 8384
rect 3145 8347 3203 8353
rect 3145 8313 3157 8347
rect 3191 8344 3203 8347
rect 3602 8344 3608 8356
rect 3191 8316 3608 8344
rect 3191 8313 3203 8316
rect 3145 8307 3203 8313
rect 3602 8304 3608 8316
rect 3660 8304 3666 8356
rect 12084 8344 12112 8443
rect 12452 8412 12480 8443
rect 12802 8440 12808 8492
rect 12860 8440 12866 8492
rect 13170 8440 13176 8492
rect 13228 8440 13234 8492
rect 13556 8489 13584 8520
rect 14734 8508 14740 8520
rect 14792 8508 14798 8560
rect 16574 8548 16580 8560
rect 15672 8520 16580 8548
rect 15672 8492 15700 8520
rect 16574 8508 16580 8520
rect 16632 8508 16638 8560
rect 17972 8548 18000 8588
rect 18230 8576 18236 8588
rect 18288 8576 18294 8628
rect 32214 8576 32220 8628
rect 32272 8616 32278 8628
rect 32309 8619 32367 8625
rect 32309 8616 32321 8619
rect 32272 8588 32321 8616
rect 32272 8576 32278 8588
rect 32309 8585 32321 8588
rect 32355 8585 32367 8619
rect 32309 8579 32367 8585
rect 32490 8576 32496 8628
rect 32548 8616 32554 8628
rect 32769 8619 32827 8625
rect 32769 8616 32781 8619
rect 32548 8588 32781 8616
rect 32548 8576 32554 8588
rect 32769 8585 32781 8588
rect 32815 8585 32827 8619
rect 32769 8579 32827 8585
rect 32858 8576 32864 8628
rect 32916 8616 32922 8628
rect 33137 8619 33195 8625
rect 33137 8616 33149 8619
rect 32916 8588 33149 8616
rect 32916 8576 32922 8588
rect 33137 8585 33149 8588
rect 33183 8585 33195 8619
rect 33137 8579 33195 8585
rect 33502 8576 33508 8628
rect 33560 8576 33566 8628
rect 33873 8619 33931 8625
rect 33873 8585 33885 8619
rect 33919 8585 33931 8619
rect 33873 8579 33931 8585
rect 17052 8520 18000 8548
rect 18064 8520 19334 8548
rect 13541 8483 13599 8489
rect 13541 8449 13553 8483
rect 13587 8449 13599 8483
rect 13541 8443 13599 8449
rect 13909 8483 13967 8489
rect 13909 8449 13921 8483
rect 13955 8449 13967 8483
rect 13909 8443 13967 8449
rect 14645 8483 14703 8489
rect 14645 8449 14657 8483
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8480 15071 8483
rect 15286 8480 15292 8492
rect 15059 8452 15292 8480
rect 15059 8449 15071 8452
rect 15013 8443 15071 8449
rect 13814 8412 13820 8424
rect 12452 8384 13820 8412
rect 13814 8372 13820 8384
rect 13872 8372 13878 8424
rect 13924 8344 13952 8443
rect 14660 8412 14688 8443
rect 15286 8440 15292 8452
rect 15344 8440 15350 8492
rect 15381 8483 15439 8489
rect 15381 8449 15393 8483
rect 15427 8480 15439 8483
rect 15562 8480 15568 8492
rect 15427 8452 15568 8480
rect 15427 8449 15439 8452
rect 15381 8443 15439 8449
rect 15562 8440 15568 8452
rect 15620 8440 15626 8492
rect 15654 8440 15660 8492
rect 15712 8440 15718 8492
rect 15746 8440 15752 8492
rect 15804 8440 15810 8492
rect 16114 8440 16120 8492
rect 16172 8440 16178 8492
rect 16485 8483 16543 8489
rect 16485 8449 16497 8483
rect 16531 8480 16543 8483
rect 17052 8480 17080 8520
rect 16531 8452 17080 8480
rect 17129 8483 17187 8489
rect 16531 8449 16543 8452
rect 16485 8443 16543 8449
rect 17129 8449 17141 8483
rect 17175 8449 17187 8483
rect 17129 8443 17187 8449
rect 16390 8412 16396 8424
rect 14660 8384 16396 8412
rect 16390 8372 16396 8384
rect 16448 8372 16454 8424
rect 17144 8344 17172 8443
rect 17402 8440 17408 8492
rect 17460 8440 17466 8492
rect 17678 8440 17684 8492
rect 17736 8480 17742 8492
rect 18064 8489 18092 8520
rect 18049 8483 18107 8489
rect 17736 8452 18000 8480
rect 17736 8440 17742 8452
rect 17972 8412 18000 8452
rect 18049 8449 18061 8483
rect 18095 8449 18107 8483
rect 19306 8480 19334 8520
rect 23382 8508 23388 8560
rect 23440 8548 23446 8560
rect 23440 8520 33364 8548
rect 23440 8508 23446 8520
rect 20714 8480 20720 8492
rect 19306 8452 20720 8480
rect 18049 8443 18107 8449
rect 20714 8440 20720 8452
rect 20772 8440 20778 8492
rect 30374 8440 30380 8492
rect 30432 8480 30438 8492
rect 32493 8483 32551 8489
rect 32493 8480 32505 8483
rect 30432 8452 32505 8480
rect 30432 8440 30438 8452
rect 32493 8449 32505 8452
rect 32539 8449 32551 8483
rect 32493 8443 32551 8449
rect 32582 8440 32588 8492
rect 32640 8440 32646 8492
rect 32674 8440 32680 8492
rect 32732 8480 32738 8492
rect 33336 8489 33364 8520
rect 33410 8508 33416 8560
rect 33468 8548 33474 8560
rect 33888 8548 33916 8579
rect 34238 8576 34244 8628
rect 34296 8576 34302 8628
rect 34698 8576 34704 8628
rect 34756 8616 34762 8628
rect 35529 8619 35587 8625
rect 35529 8616 35541 8619
rect 34756 8588 35541 8616
rect 34756 8576 34762 8588
rect 35529 8585 35541 8588
rect 35575 8585 35587 8619
rect 35529 8579 35587 8585
rect 35802 8576 35808 8628
rect 35860 8616 35866 8628
rect 36725 8619 36783 8625
rect 36725 8616 36737 8619
rect 35860 8588 36737 8616
rect 35860 8576 35866 8588
rect 36725 8585 36737 8588
rect 36771 8585 36783 8619
rect 36725 8579 36783 8585
rect 36906 8576 36912 8628
rect 36964 8616 36970 8628
rect 37829 8619 37887 8625
rect 37829 8616 37841 8619
rect 36964 8588 37841 8616
rect 36964 8576 36970 8588
rect 37829 8585 37841 8588
rect 37875 8585 37887 8619
rect 37829 8579 37887 8585
rect 38565 8619 38623 8625
rect 38565 8585 38577 8619
rect 38611 8585 38623 8619
rect 38565 8579 38623 8585
rect 33468 8520 33916 8548
rect 33468 8508 33474 8520
rect 34146 8508 34152 8560
rect 34204 8548 34210 8560
rect 34204 8520 34836 8548
rect 34204 8508 34210 8520
rect 32953 8483 33011 8489
rect 32953 8480 32965 8483
rect 32732 8452 32965 8480
rect 32732 8440 32738 8452
rect 32953 8449 32965 8452
rect 32999 8449 33011 8483
rect 32953 8443 33011 8449
rect 33321 8483 33379 8489
rect 33321 8449 33333 8483
rect 33367 8449 33379 8483
rect 33689 8483 33747 8489
rect 33689 8480 33701 8483
rect 33321 8443 33379 8449
rect 33428 8452 33701 8480
rect 18141 8415 18199 8421
rect 18141 8412 18153 8415
rect 17972 8384 18153 8412
rect 18141 8381 18153 8384
rect 18187 8381 18199 8415
rect 18141 8375 18199 8381
rect 18230 8372 18236 8424
rect 18288 8412 18294 8424
rect 23106 8412 23112 8424
rect 18288 8384 23112 8412
rect 18288 8372 18294 8384
rect 23106 8372 23112 8384
rect 23164 8372 23170 8424
rect 24946 8372 24952 8424
rect 25004 8412 25010 8424
rect 33428 8412 33456 8452
rect 33689 8449 33701 8452
rect 33735 8449 33747 8483
rect 33689 8443 33747 8449
rect 34054 8440 34060 8492
rect 34112 8440 34118 8492
rect 34701 8483 34759 8489
rect 34701 8449 34713 8483
rect 34747 8449 34759 8483
rect 34701 8443 34759 8449
rect 34716 8412 34744 8443
rect 25004 8384 33456 8412
rect 33704 8384 34744 8412
rect 34808 8412 34836 8520
rect 35618 8508 35624 8560
rect 35676 8548 35682 8560
rect 35676 8520 37228 8548
rect 35676 8508 35682 8520
rect 34882 8440 34888 8492
rect 34940 8480 34946 8492
rect 35069 8483 35127 8489
rect 35069 8480 35081 8483
rect 34940 8452 35081 8480
rect 34940 8440 34946 8452
rect 35069 8449 35081 8452
rect 35115 8449 35127 8483
rect 35069 8443 35127 8449
rect 35250 8440 35256 8492
rect 35308 8480 35314 8492
rect 35308 8452 35664 8480
rect 35308 8440 35314 8452
rect 35636 8412 35664 8452
rect 35710 8440 35716 8492
rect 35768 8440 35774 8492
rect 35802 8440 35808 8492
rect 35860 8440 35866 8492
rect 36170 8440 36176 8492
rect 36228 8440 36234 8492
rect 36538 8440 36544 8492
rect 36596 8440 36602 8492
rect 34808 8384 35296 8412
rect 35636 8384 36124 8412
rect 25004 8372 25010 8384
rect 23750 8344 23756 8356
rect 12084 8316 13860 8344
rect 13924 8316 17080 8344
rect 17144 8316 23756 8344
rect 7190 8236 7196 8288
rect 7248 8276 7254 8288
rect 13722 8276 13728 8288
rect 7248 8248 13728 8276
rect 7248 8236 7254 8248
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 13832 8276 13860 8316
rect 14366 8276 14372 8288
rect 13832 8248 14372 8276
rect 14366 8236 14372 8248
rect 14424 8236 14430 8288
rect 14458 8236 14464 8288
rect 14516 8276 14522 8288
rect 16942 8276 16948 8288
rect 14516 8248 16948 8276
rect 14516 8236 14522 8248
rect 16942 8236 16948 8248
rect 17000 8236 17006 8288
rect 17052 8276 17080 8316
rect 23750 8304 23756 8316
rect 23808 8304 23814 8356
rect 30926 8304 30932 8356
rect 30984 8344 30990 8356
rect 33704 8344 33732 8384
rect 30984 8316 33732 8344
rect 30984 8304 30990 8316
rect 33962 8304 33968 8356
rect 34020 8344 34026 8356
rect 34885 8347 34943 8353
rect 34885 8344 34897 8347
rect 34020 8316 34897 8344
rect 34020 8304 34026 8316
rect 34885 8313 34897 8316
rect 34931 8313 34943 8347
rect 34885 8307 34943 8313
rect 31018 8276 31024 8288
rect 17052 8248 31024 8276
rect 31018 8236 31024 8248
rect 31076 8236 31082 8288
rect 35268 8285 35296 8384
rect 35342 8304 35348 8356
rect 35400 8344 35406 8356
rect 35989 8347 36047 8353
rect 35989 8344 36001 8347
rect 35400 8316 36001 8344
rect 35400 8304 35406 8316
rect 35989 8313 36001 8316
rect 36035 8313 36047 8347
rect 36096 8344 36124 8384
rect 36354 8372 36360 8424
rect 36412 8412 36418 8424
rect 37200 8412 37228 8520
rect 37458 8508 37464 8560
rect 37516 8548 37522 8560
rect 38580 8548 38608 8579
rect 37516 8520 38608 8548
rect 37516 8508 37522 8520
rect 37274 8440 37280 8492
rect 37332 8440 37338 8492
rect 37366 8440 37372 8492
rect 37424 8480 37430 8492
rect 37645 8483 37703 8489
rect 37645 8480 37657 8483
rect 37424 8452 37657 8480
rect 37424 8440 37430 8452
rect 37645 8449 37657 8452
rect 37691 8449 37703 8483
rect 37645 8443 37703 8449
rect 38010 8440 38016 8492
rect 38068 8440 38074 8492
rect 38381 8483 38439 8489
rect 38381 8449 38393 8483
rect 38427 8449 38439 8483
rect 38381 8443 38439 8449
rect 38396 8412 38424 8443
rect 38562 8440 38568 8492
rect 38620 8480 38626 8492
rect 38841 8483 38899 8489
rect 38841 8480 38853 8483
rect 38620 8452 38853 8480
rect 38620 8440 38626 8452
rect 38841 8449 38853 8452
rect 38887 8449 38899 8483
rect 38841 8443 38899 8449
rect 38930 8440 38936 8492
rect 38988 8480 38994 8492
rect 39209 8483 39267 8489
rect 39209 8480 39221 8483
rect 38988 8452 39221 8480
rect 38988 8440 38994 8452
rect 39209 8449 39221 8452
rect 39255 8449 39267 8483
rect 39209 8443 39267 8449
rect 36412 8384 37136 8412
rect 37200 8384 38424 8412
rect 36412 8372 36418 8384
rect 36096 8316 36400 8344
rect 35989 8307 36047 8313
rect 36372 8285 36400 8316
rect 35253 8279 35311 8285
rect 35253 8245 35265 8279
rect 35299 8245 35311 8279
rect 35253 8239 35311 8245
rect 36357 8279 36415 8285
rect 36357 8245 36369 8279
rect 36403 8245 36415 8279
rect 37108 8276 37136 8384
rect 37182 8304 37188 8356
rect 37240 8344 37246 8356
rect 38197 8347 38255 8353
rect 38197 8344 38209 8347
rect 37240 8316 38209 8344
rect 37240 8304 37246 8316
rect 38197 8313 38209 8316
rect 38243 8313 38255 8347
rect 38197 8307 38255 8313
rect 39022 8304 39028 8356
rect 39080 8304 39086 8356
rect 39390 8304 39396 8356
rect 39448 8304 39454 8356
rect 37461 8279 37519 8285
rect 37461 8276 37473 8279
rect 37108 8248 37473 8276
rect 36357 8239 36415 8245
rect 37461 8245 37473 8248
rect 37507 8245 37519 8279
rect 37461 8239 37519 8245
rect 1104 8186 39836 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 37950 8186
rect 38002 8134 38014 8186
rect 38066 8134 38078 8186
rect 38130 8134 38142 8186
rect 38194 8134 38206 8186
rect 38258 8134 39836 8186
rect 1104 8112 39836 8134
rect 3510 8032 3516 8084
rect 3568 8032 3574 8084
rect 3970 8032 3976 8084
rect 4028 8072 4034 8084
rect 4341 8075 4399 8081
rect 4341 8072 4353 8075
rect 4028 8044 4353 8072
rect 4028 8032 4034 8044
rect 4341 8041 4353 8044
rect 4387 8041 4399 8075
rect 4341 8035 4399 8041
rect 4890 8032 4896 8084
rect 4948 8072 4954 8084
rect 5169 8075 5227 8081
rect 5169 8072 5181 8075
rect 4948 8044 5181 8072
rect 4948 8032 4954 8044
rect 5169 8041 5181 8044
rect 5215 8041 5227 8075
rect 5169 8035 5227 8041
rect 5994 8032 6000 8084
rect 6052 8072 6058 8084
rect 6181 8075 6239 8081
rect 6181 8072 6193 8075
rect 6052 8044 6193 8072
rect 6052 8032 6058 8044
rect 6181 8041 6193 8044
rect 6227 8041 6239 8075
rect 6181 8035 6239 8041
rect 6546 8032 6552 8084
rect 6604 8072 6610 8084
rect 6825 8075 6883 8081
rect 6825 8072 6837 8075
rect 6604 8044 6837 8072
rect 6604 8032 6610 8044
rect 6825 8041 6837 8044
rect 6871 8041 6883 8075
rect 6825 8035 6883 8041
rect 7098 8032 7104 8084
rect 7156 8072 7162 8084
rect 7285 8075 7343 8081
rect 7285 8072 7297 8075
rect 7156 8044 7297 8072
rect 7156 8032 7162 8044
rect 7285 8041 7297 8044
rect 7331 8041 7343 8075
rect 7285 8035 7343 8041
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 8389 8075 8447 8081
rect 8389 8072 8401 8075
rect 8352 8044 8401 8072
rect 8352 8032 8358 8044
rect 8389 8041 8401 8044
rect 8435 8041 8447 8075
rect 8389 8035 8447 8041
rect 8754 8032 8760 8084
rect 8812 8072 8818 8084
rect 9033 8075 9091 8081
rect 9033 8072 9045 8075
rect 8812 8044 9045 8072
rect 8812 8032 8818 8044
rect 9033 8041 9045 8044
rect 9079 8041 9091 8075
rect 9033 8035 9091 8041
rect 9398 8032 9404 8084
rect 9456 8072 9462 8084
rect 9493 8075 9551 8081
rect 9493 8072 9505 8075
rect 9456 8044 9505 8072
rect 9456 8032 9462 8044
rect 9493 8041 9505 8044
rect 9539 8041 9551 8075
rect 9493 8035 9551 8041
rect 10410 8032 10416 8084
rect 10468 8072 10474 8084
rect 10597 8075 10655 8081
rect 10597 8072 10609 8075
rect 10468 8044 10609 8072
rect 10468 8032 10474 8044
rect 10597 8041 10609 8044
rect 10643 8041 10655 8075
rect 10597 8035 10655 8041
rect 11238 8032 11244 8084
rect 11296 8072 11302 8084
rect 11425 8075 11483 8081
rect 11425 8072 11437 8075
rect 11296 8044 11437 8072
rect 11296 8032 11302 8044
rect 11425 8041 11437 8044
rect 11471 8041 11483 8075
rect 11425 8035 11483 8041
rect 11790 8032 11796 8084
rect 11848 8032 11854 8084
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 12805 8075 12863 8081
rect 12805 8072 12817 8075
rect 12676 8044 12817 8072
rect 12676 8032 12682 8044
rect 12805 8041 12817 8044
rect 12851 8041 12863 8075
rect 12805 8035 12863 8041
rect 13446 8032 13452 8084
rect 13504 8072 13510 8084
rect 13633 8075 13691 8081
rect 13633 8072 13645 8075
rect 13504 8044 13645 8072
rect 13504 8032 13510 8044
rect 13633 8041 13645 8044
rect 13679 8041 13691 8075
rect 13633 8035 13691 8041
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 14093 8075 14151 8081
rect 14093 8072 14105 8075
rect 13872 8044 14105 8072
rect 13872 8032 13878 8044
rect 14093 8041 14105 8044
rect 14139 8041 14151 8075
rect 14093 8035 14151 8041
rect 14274 8032 14280 8084
rect 14332 8072 14338 8084
rect 14461 8075 14519 8081
rect 14461 8072 14473 8075
rect 14332 8044 14473 8072
rect 14332 8032 14338 8044
rect 14461 8041 14473 8044
rect 14507 8041 14519 8075
rect 14461 8035 14519 8041
rect 14550 8032 14556 8084
rect 14608 8032 14614 8084
rect 14826 8032 14832 8084
rect 14884 8072 14890 8084
rect 15657 8075 15715 8081
rect 15657 8072 15669 8075
rect 14884 8044 15669 8072
rect 14884 8032 14890 8044
rect 15657 8041 15669 8044
rect 15703 8041 15715 8075
rect 15657 8035 15715 8041
rect 15930 8032 15936 8084
rect 15988 8072 15994 8084
rect 16117 8075 16175 8081
rect 16117 8072 16129 8075
rect 15988 8044 16129 8072
rect 15988 8032 15994 8044
rect 16117 8041 16129 8044
rect 16163 8041 16175 8075
rect 16117 8035 16175 8041
rect 19702 8032 19708 8084
rect 19760 8032 19766 8084
rect 20622 8032 20628 8084
rect 20680 8072 20686 8084
rect 20993 8075 21051 8081
rect 20993 8072 21005 8075
rect 20680 8044 21005 8072
rect 20680 8032 20686 8044
rect 20993 8041 21005 8044
rect 21039 8041 21051 8075
rect 20993 8035 21051 8041
rect 21818 8032 21824 8084
rect 21876 8032 21882 8084
rect 23106 8032 23112 8084
rect 23164 8032 23170 8084
rect 23474 8032 23480 8084
rect 23532 8032 23538 8084
rect 27614 8032 27620 8084
rect 27672 8072 27678 8084
rect 28902 8072 28908 8084
rect 27672 8044 28908 8072
rect 27672 8032 27678 8044
rect 28902 8032 28908 8044
rect 28960 8032 28966 8084
rect 31018 8032 31024 8084
rect 31076 8032 31082 8084
rect 34422 8032 34428 8084
rect 34480 8072 34486 8084
rect 34793 8075 34851 8081
rect 34793 8072 34805 8075
rect 34480 8044 34805 8072
rect 34480 8032 34486 8044
rect 34793 8041 34805 8044
rect 34839 8041 34851 8075
rect 34793 8035 34851 8041
rect 35526 8032 35532 8084
rect 35584 8072 35590 8084
rect 35805 8075 35863 8081
rect 35805 8072 35817 8075
rect 35584 8044 35817 8072
rect 35584 8032 35590 8044
rect 35805 8041 35817 8044
rect 35851 8041 35863 8075
rect 35805 8035 35863 8041
rect 36078 8032 36084 8084
rect 36136 8072 36142 8084
rect 36357 8075 36415 8081
rect 36357 8072 36369 8075
rect 36136 8044 36369 8072
rect 36136 8032 36142 8044
rect 36357 8041 36369 8044
rect 36403 8041 36415 8075
rect 36357 8035 36415 8041
rect 36630 8032 36636 8084
rect 36688 8072 36694 8084
rect 36909 8075 36967 8081
rect 36909 8072 36921 8075
rect 36688 8044 36921 8072
rect 36688 8032 36694 8044
rect 36909 8041 36921 8044
rect 36955 8041 36967 8075
rect 36909 8035 36967 8041
rect 37734 8032 37740 8084
rect 37792 8072 37798 8084
rect 37921 8075 37979 8081
rect 37921 8072 37933 8075
rect 37792 8044 37933 8072
rect 37792 8032 37798 8044
rect 37921 8041 37933 8044
rect 37967 8041 37979 8075
rect 37921 8035 37979 8041
rect 38654 8032 38660 8084
rect 38712 8032 38718 8084
rect 8113 8007 8171 8013
rect 8113 7973 8125 8007
rect 8159 8004 8171 8007
rect 8478 8004 8484 8016
rect 8159 7976 8484 8004
rect 8159 7973 8171 7976
rect 8113 7967 8171 7973
rect 8478 7964 8484 7976
rect 8536 7964 8542 8016
rect 12253 8007 12311 8013
rect 12253 8004 12265 8007
rect 9232 7976 12265 8004
rect 3970 7896 3976 7948
rect 4028 7936 4034 7948
rect 4065 7939 4123 7945
rect 4065 7936 4077 7939
rect 4028 7908 4077 7936
rect 4028 7896 4034 7908
rect 4065 7905 4077 7908
rect 4111 7905 4123 7939
rect 4065 7899 4123 7905
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 3329 7871 3387 7877
rect 3329 7868 3341 7871
rect 2832 7840 3341 7868
rect 2832 7828 2838 7840
rect 3329 7837 3341 7840
rect 3375 7837 3387 7871
rect 3329 7831 3387 7837
rect 4154 7828 4160 7880
rect 4212 7828 4218 7880
rect 4982 7828 4988 7880
rect 5040 7828 5046 7880
rect 6365 7871 6423 7877
rect 6365 7837 6377 7871
rect 6411 7837 6423 7871
rect 6365 7831 6423 7837
rect 3881 7803 3939 7809
rect 3881 7769 3893 7803
rect 3927 7800 3939 7803
rect 6380 7800 6408 7831
rect 6638 7828 6644 7880
rect 6696 7828 6702 7880
rect 7466 7828 7472 7880
rect 7524 7828 7530 7880
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7868 7895 7871
rect 7929 7871 7987 7877
rect 7929 7868 7941 7871
rect 7883 7840 7941 7868
rect 7883 7837 7895 7840
rect 7837 7831 7895 7837
rect 7929 7837 7941 7840
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 8570 7828 8576 7880
rect 8628 7828 8634 7880
rect 9232 7877 9260 7976
rect 12253 7973 12265 7976
rect 12299 7973 12311 8007
rect 13265 8007 13323 8013
rect 13265 8004 13277 8007
rect 12253 7967 12311 7973
rect 12406 7976 13277 8004
rect 11882 7936 11888 7948
rect 9692 7908 11888 7936
rect 9692 7877 9720 7908
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 12406 7936 12434 7976
rect 13265 7973 13277 7976
rect 13311 7973 13323 8007
rect 14568 8004 14596 8032
rect 14918 8004 14924 8016
rect 14568 7976 14924 8004
rect 13265 7967 13323 7973
rect 14918 7964 14924 7976
rect 14976 7964 14982 8016
rect 15197 8007 15255 8013
rect 15197 7973 15209 8007
rect 15243 8004 15255 8007
rect 15470 8004 15476 8016
rect 15243 7976 15476 8004
rect 15243 7973 15255 7976
rect 15197 7967 15255 7973
rect 15470 7964 15476 7976
rect 15528 7964 15534 8016
rect 22189 8007 22247 8013
rect 22189 7973 22201 8007
rect 22235 8004 22247 8007
rect 31570 8004 31576 8016
rect 22235 7976 31576 8004
rect 22235 7973 22247 7976
rect 22189 7967 22247 7973
rect 31570 7964 31576 7976
rect 31628 7964 31634 8016
rect 31726 7976 38516 8004
rect 14550 7936 14556 7948
rect 11992 7908 12434 7936
rect 12912 7908 14556 7936
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7837 9275 7871
rect 9217 7831 9275 7837
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 9769 7871 9827 7877
rect 9769 7837 9781 7871
rect 9815 7837 9827 7871
rect 9769 7831 9827 7837
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7868 10839 7871
rect 11514 7868 11520 7880
rect 10827 7840 11520 7868
rect 10827 7837 10839 7840
rect 10781 7831 10839 7837
rect 7650 7800 7656 7812
rect 3927 7772 5396 7800
rect 6380 7772 7656 7800
rect 3927 7769 3939 7772
rect 3881 7763 3939 7769
rect 5368 7732 5396 7772
rect 7650 7760 7656 7772
rect 7708 7760 7714 7812
rect 8294 7760 8300 7812
rect 8352 7800 8358 7812
rect 9784 7800 9812 7831
rect 11514 7828 11520 7840
rect 11572 7828 11578 7880
rect 11606 7828 11612 7880
rect 11664 7828 11670 7880
rect 11992 7877 12020 7908
rect 11977 7871 12035 7877
rect 11977 7837 11989 7871
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 12161 7871 12219 7877
rect 12161 7837 12173 7871
rect 12207 7868 12219 7871
rect 12437 7871 12495 7877
rect 12437 7868 12449 7871
rect 12207 7840 12449 7868
rect 12207 7837 12219 7840
rect 12161 7831 12219 7837
rect 12437 7837 12449 7840
rect 12483 7868 12495 7871
rect 12912 7868 12940 7908
rect 14550 7896 14556 7908
rect 14608 7896 14614 7948
rect 19794 7936 19800 7948
rect 14660 7908 19800 7936
rect 12483 7840 12940 7868
rect 12989 7871 13047 7877
rect 12483 7837 12495 7840
rect 12437 7831 12495 7837
rect 12989 7837 13001 7871
rect 13035 7837 13047 7871
rect 12989 7831 13047 7837
rect 13004 7800 13032 7831
rect 13446 7828 13452 7880
rect 13504 7828 13510 7880
rect 13814 7828 13820 7880
rect 13872 7828 13878 7880
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7868 14335 7871
rect 14458 7868 14464 7880
rect 14323 7840 14464 7868
rect 14323 7837 14335 7840
rect 14277 7831 14335 7837
rect 14458 7828 14464 7840
rect 14516 7828 14522 7880
rect 14660 7877 14688 7908
rect 19794 7896 19800 7908
rect 19852 7896 19858 7948
rect 19904 7908 22600 7936
rect 14645 7871 14703 7877
rect 14645 7837 14657 7871
rect 14691 7837 14703 7871
rect 14645 7831 14703 7837
rect 15197 7871 15255 7877
rect 15197 7837 15209 7871
rect 15243 7868 15255 7871
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 15243 7840 15301 7868
rect 15243 7837 15255 7840
rect 15197 7831 15255 7837
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 15838 7828 15844 7880
rect 15896 7828 15902 7880
rect 16301 7871 16359 7877
rect 16301 7837 16313 7871
rect 16347 7868 16359 7871
rect 17773 7871 17831 7877
rect 16347 7840 17724 7868
rect 16347 7837 16359 7840
rect 16301 7831 16359 7837
rect 8352 7772 9812 7800
rect 9876 7772 10916 7800
rect 13004 7772 17632 7800
rect 8352 7760 8358 7772
rect 7098 7732 7104 7744
rect 5368 7704 7104 7732
rect 7098 7692 7104 7704
rect 7156 7692 7162 7744
rect 7837 7735 7895 7741
rect 7837 7701 7849 7735
rect 7883 7732 7895 7735
rect 9876 7732 9904 7772
rect 7883 7704 9904 7732
rect 9953 7735 10011 7741
rect 7883 7701 7895 7704
rect 7837 7695 7895 7701
rect 9953 7701 9965 7735
rect 9999 7732 10011 7735
rect 10778 7732 10784 7744
rect 9999 7704 10784 7732
rect 9999 7701 10011 7704
rect 9953 7695 10011 7701
rect 10778 7692 10784 7704
rect 10836 7692 10842 7744
rect 10888 7732 10916 7772
rect 12710 7732 12716 7744
rect 10888 7704 12716 7732
rect 12710 7692 12716 7704
rect 12768 7692 12774 7744
rect 15470 7692 15476 7744
rect 15528 7692 15534 7744
rect 16114 7692 16120 7744
rect 16172 7732 16178 7744
rect 16482 7732 16488 7744
rect 16172 7704 16488 7732
rect 16172 7692 16178 7704
rect 16482 7692 16488 7704
rect 16540 7692 16546 7744
rect 17604 7741 17632 7772
rect 17589 7735 17647 7741
rect 17589 7701 17601 7735
rect 17635 7701 17647 7735
rect 17696 7732 17724 7840
rect 17773 7837 17785 7871
rect 17819 7837 17831 7871
rect 17773 7831 17831 7837
rect 17788 7800 17816 7831
rect 19150 7828 19156 7880
rect 19208 7868 19214 7880
rect 19904 7877 19932 7908
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 19208 7840 19257 7868
rect 19208 7828 19214 7840
rect 19245 7837 19257 7840
rect 19291 7868 19303 7871
rect 19521 7871 19579 7877
rect 19521 7868 19533 7871
rect 19291 7840 19533 7868
rect 19291 7837 19303 7840
rect 19245 7831 19303 7837
rect 19521 7837 19533 7840
rect 19567 7837 19579 7871
rect 19521 7831 19579 7837
rect 19889 7871 19947 7877
rect 19889 7837 19901 7871
rect 19935 7837 19947 7871
rect 19889 7831 19947 7837
rect 21085 7871 21143 7877
rect 21085 7837 21097 7871
rect 21131 7868 21143 7871
rect 21177 7871 21235 7877
rect 21177 7868 21189 7871
rect 21131 7840 21189 7868
rect 21131 7837 21143 7840
rect 21085 7831 21143 7837
rect 21177 7837 21189 7840
rect 21223 7837 21235 7871
rect 21177 7831 21235 7837
rect 21913 7871 21971 7877
rect 21913 7837 21925 7871
rect 21959 7868 21971 7871
rect 22005 7871 22063 7877
rect 22005 7868 22017 7871
rect 21959 7840 22017 7868
rect 21959 7837 21971 7840
rect 21913 7831 21971 7837
rect 22005 7837 22017 7840
rect 22051 7837 22063 7871
rect 22572 7868 22600 7908
rect 22646 7896 22652 7948
rect 22704 7936 22710 7948
rect 31726 7936 31754 7976
rect 22704 7908 31754 7936
rect 22704 7896 22710 7908
rect 31846 7896 31852 7948
rect 31904 7936 31910 7948
rect 31904 7908 35112 7936
rect 31904 7896 31910 7908
rect 23198 7868 23204 7880
rect 22572 7840 23204 7868
rect 22005 7831 22063 7837
rect 23198 7828 23204 7840
rect 23256 7828 23262 7880
rect 23293 7871 23351 7877
rect 23293 7837 23305 7871
rect 23339 7868 23351 7871
rect 23566 7868 23572 7880
rect 23339 7840 23572 7868
rect 23339 7837 23351 7840
rect 23293 7831 23351 7837
rect 23566 7828 23572 7840
rect 23624 7828 23630 7880
rect 23661 7871 23719 7877
rect 23661 7837 23673 7871
rect 23707 7868 23719 7871
rect 27614 7868 27620 7880
rect 23707 7840 27620 7868
rect 23707 7837 23719 7840
rect 23661 7831 23719 7837
rect 27614 7828 27620 7840
rect 27672 7828 27678 7880
rect 27706 7828 27712 7880
rect 27764 7828 27770 7880
rect 31110 7828 31116 7880
rect 31168 7868 31174 7880
rect 31205 7871 31263 7877
rect 31205 7868 31217 7871
rect 31168 7840 31217 7868
rect 31168 7828 31174 7840
rect 31205 7837 31217 7840
rect 31251 7837 31263 7871
rect 31205 7831 31263 7837
rect 31386 7828 31392 7880
rect 31444 7868 31450 7880
rect 33229 7871 33287 7877
rect 33229 7868 33241 7871
rect 31444 7840 33241 7868
rect 31444 7828 31450 7840
rect 33229 7837 33241 7840
rect 33275 7837 33287 7871
rect 33229 7831 33287 7837
rect 34977 7871 35035 7877
rect 34977 7837 34989 7871
rect 35023 7837 35035 7871
rect 35084 7868 35112 7908
rect 35503 7871 35561 7877
rect 35503 7868 35515 7871
rect 35084 7840 35515 7868
rect 34977 7831 35035 7837
rect 35503 7837 35515 7840
rect 35549 7837 35561 7871
rect 35503 7831 35561 7837
rect 35621 7871 35679 7877
rect 35621 7837 35633 7871
rect 35667 7868 35679 7871
rect 35894 7868 35900 7880
rect 35667 7840 35900 7868
rect 35667 7837 35679 7840
rect 35621 7831 35679 7837
rect 20346 7800 20352 7812
rect 17788 7772 20352 7800
rect 20346 7760 20352 7772
rect 20404 7760 20410 7812
rect 20438 7760 20444 7812
rect 20496 7800 20502 7812
rect 34992 7800 35020 7831
rect 35894 7828 35900 7840
rect 35952 7828 35958 7880
rect 36170 7828 36176 7880
rect 36228 7828 36234 7880
rect 36446 7828 36452 7880
rect 36504 7868 36510 7880
rect 36725 7871 36783 7877
rect 36725 7868 36737 7871
rect 36504 7840 36737 7868
rect 36504 7828 36510 7840
rect 36725 7837 36737 7840
rect 36771 7837 36783 7871
rect 36725 7831 36783 7837
rect 38105 7871 38163 7877
rect 38105 7837 38117 7871
rect 38151 7868 38163 7871
rect 38286 7868 38292 7880
rect 38151 7840 38292 7868
rect 38151 7837 38163 7840
rect 38105 7831 38163 7837
rect 38286 7828 38292 7840
rect 38344 7828 38350 7880
rect 38488 7877 38516 7976
rect 38473 7871 38531 7877
rect 38473 7837 38485 7871
rect 38519 7837 38531 7871
rect 38473 7831 38531 7837
rect 38838 7828 38844 7880
rect 38896 7828 38902 7880
rect 39209 7871 39267 7877
rect 39209 7837 39221 7871
rect 39255 7837 39267 7871
rect 39209 7831 39267 7837
rect 20496 7772 31754 7800
rect 34992 7772 35572 7800
rect 20496 7760 20502 7772
rect 19150 7732 19156 7744
rect 17696 7704 19156 7732
rect 17589 7695 17647 7701
rect 19150 7692 19156 7704
rect 19208 7692 19214 7744
rect 19426 7692 19432 7744
rect 19484 7692 19490 7744
rect 21358 7692 21364 7744
rect 21416 7692 21422 7744
rect 27617 7735 27675 7741
rect 27617 7701 27629 7735
rect 27663 7732 27675 7735
rect 27706 7732 27712 7744
rect 27663 7704 27712 7732
rect 27663 7701 27675 7704
rect 27617 7695 27675 7701
rect 27706 7692 27712 7704
rect 27764 7692 27770 7744
rect 27890 7692 27896 7744
rect 27948 7692 27954 7744
rect 31726 7732 31754 7772
rect 33045 7735 33103 7741
rect 33045 7732 33057 7735
rect 31726 7704 33057 7732
rect 33045 7701 33057 7704
rect 33091 7701 33103 7735
rect 33045 7695 33103 7701
rect 35342 7692 35348 7744
rect 35400 7692 35406 7744
rect 35544 7732 35572 7772
rect 36354 7760 36360 7812
rect 36412 7800 36418 7812
rect 39224 7800 39252 7831
rect 36412 7772 39252 7800
rect 36412 7760 36418 7772
rect 36262 7732 36268 7744
rect 35544 7704 36268 7732
rect 36262 7692 36268 7704
rect 36320 7692 36326 7744
rect 38930 7692 38936 7744
rect 38988 7732 38994 7744
rect 39025 7735 39083 7741
rect 39025 7732 39037 7735
rect 38988 7704 39037 7732
rect 38988 7692 38994 7704
rect 39025 7701 39037 7704
rect 39071 7701 39083 7735
rect 39025 7695 39083 7701
rect 39390 7692 39396 7744
rect 39448 7692 39454 7744
rect 1104 7642 39836 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 39010 7642
rect 39062 7590 39074 7642
rect 39126 7590 39138 7642
rect 39190 7590 39202 7642
rect 39254 7590 39266 7642
rect 39318 7590 39836 7642
rect 1104 7568 39836 7590
rect 2774 7488 2780 7540
rect 2832 7488 2838 7540
rect 9490 7488 9496 7540
rect 9548 7528 9554 7540
rect 9585 7531 9643 7537
rect 9585 7528 9597 7531
rect 9548 7500 9597 7528
rect 9548 7488 9554 7500
rect 9585 7497 9597 7500
rect 9631 7497 9643 7531
rect 14185 7531 14243 7537
rect 9585 7491 9643 7497
rect 9692 7500 12388 7528
rect 9692 7460 9720 7500
rect 9324 7432 9720 7460
rect 12360 7460 12388 7500
rect 14185 7497 14197 7531
rect 14231 7528 14243 7531
rect 14366 7528 14372 7540
rect 14231 7500 14372 7528
rect 14231 7497 14243 7500
rect 14185 7491 14243 7497
rect 14366 7488 14372 7500
rect 14424 7488 14430 7540
rect 14734 7488 14740 7540
rect 14792 7528 14798 7540
rect 20438 7528 20444 7540
rect 14792 7500 20444 7528
rect 14792 7488 14798 7500
rect 20438 7488 20444 7500
rect 20496 7488 20502 7540
rect 20714 7488 20720 7540
rect 20772 7528 20778 7540
rect 21177 7531 21235 7537
rect 21177 7528 21189 7531
rect 20772 7500 21189 7528
rect 20772 7488 20778 7500
rect 21177 7497 21189 7500
rect 21223 7497 21235 7531
rect 21177 7491 21235 7497
rect 21358 7488 21364 7540
rect 21416 7528 21422 7540
rect 22646 7528 22652 7540
rect 21416 7500 22652 7528
rect 21416 7488 21422 7500
rect 22646 7488 22652 7500
rect 22704 7488 22710 7540
rect 23750 7488 23756 7540
rect 23808 7488 23814 7540
rect 27890 7488 27896 7540
rect 27948 7528 27954 7540
rect 34146 7528 34152 7540
rect 27948 7500 34152 7528
rect 27948 7488 27954 7500
rect 34146 7488 34152 7500
rect 34204 7488 34210 7540
rect 36446 7528 36452 7540
rect 34256 7500 36452 7528
rect 13078 7460 13084 7472
rect 12360 7432 13084 7460
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7392 2651 7395
rect 7190 7392 7196 7404
rect 2639 7364 7196 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 7282 7352 7288 7404
rect 7340 7392 7346 7404
rect 9324 7401 9352 7432
rect 13078 7420 13084 7432
rect 13136 7420 13142 7472
rect 14829 7463 14887 7469
rect 14829 7429 14841 7463
rect 14875 7460 14887 7463
rect 14918 7460 14924 7472
rect 14875 7432 14924 7460
rect 14875 7429 14887 7432
rect 14829 7423 14887 7429
rect 14918 7420 14924 7432
rect 14976 7420 14982 7472
rect 18046 7460 18052 7472
rect 17788 7432 18052 7460
rect 7653 7395 7711 7401
rect 7653 7392 7665 7395
rect 7340 7364 7665 7392
rect 7340 7352 7346 7364
rect 7653 7361 7665 7364
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7361 9367 7395
rect 9309 7355 9367 7361
rect 9766 7352 9772 7404
rect 9824 7352 9830 7404
rect 14093 7395 14151 7401
rect 14093 7361 14105 7395
rect 14139 7392 14151 7395
rect 14369 7395 14427 7401
rect 14369 7392 14381 7395
rect 14139 7364 14381 7392
rect 14139 7361 14151 7364
rect 14093 7355 14151 7361
rect 14369 7361 14381 7364
rect 14415 7361 14427 7395
rect 14369 7355 14427 7361
rect 14645 7395 14703 7401
rect 14645 7361 14657 7395
rect 14691 7392 14703 7395
rect 14737 7395 14795 7401
rect 14737 7392 14749 7395
rect 14691 7364 14749 7392
rect 14691 7361 14703 7364
rect 14645 7355 14703 7361
rect 14737 7361 14749 7364
rect 14783 7361 14795 7395
rect 14737 7355 14795 7361
rect 16025 7395 16083 7401
rect 16025 7361 16037 7395
rect 16071 7392 16083 7395
rect 17494 7392 17500 7404
rect 16071 7364 17500 7392
rect 16071 7361 16083 7364
rect 16025 7355 16083 7361
rect 17494 7352 17500 7364
rect 17552 7352 17558 7404
rect 17690 7395 17748 7401
rect 17690 7361 17702 7395
rect 17736 7392 17748 7395
rect 17788 7392 17816 7432
rect 18046 7420 18052 7432
rect 18104 7420 18110 7472
rect 19150 7420 19156 7472
rect 19208 7460 19214 7472
rect 24762 7460 24768 7472
rect 19208 7432 24768 7460
rect 19208 7420 19214 7432
rect 24762 7420 24768 7432
rect 24820 7420 24826 7472
rect 30650 7420 30656 7472
rect 30708 7460 30714 7472
rect 34256 7460 34284 7500
rect 36446 7488 36452 7500
rect 36504 7488 36510 7540
rect 38289 7531 38347 7537
rect 38289 7497 38301 7531
rect 38335 7497 38347 7531
rect 38289 7491 38347 7497
rect 38657 7531 38715 7537
rect 38657 7497 38669 7531
rect 38703 7528 38715 7531
rect 38746 7528 38752 7540
rect 38703 7500 38752 7528
rect 38703 7497 38715 7500
rect 38657 7491 38715 7497
rect 30708 7432 34284 7460
rect 30708 7420 30714 7432
rect 17736 7364 17816 7392
rect 17736 7361 17748 7364
rect 17690 7355 17748 7361
rect 3602 7284 3608 7336
rect 3660 7324 3666 7336
rect 8294 7324 8300 7336
rect 3660 7296 8300 7324
rect 3660 7284 3666 7296
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 8570 7284 8576 7336
rect 8628 7324 8634 7336
rect 12250 7324 12256 7336
rect 8628 7296 12256 7324
rect 8628 7284 8634 7296
rect 12250 7284 12256 7296
rect 12308 7284 12314 7336
rect 13446 7284 13452 7336
rect 13504 7324 13510 7336
rect 17589 7327 17647 7333
rect 13504 7296 17540 7324
rect 13504 7284 13510 7296
rect 9493 7259 9551 7265
rect 9493 7225 9505 7259
rect 9539 7256 9551 7259
rect 9950 7256 9956 7268
rect 9539 7228 9956 7256
rect 9539 7225 9551 7228
rect 9493 7219 9551 7225
rect 9950 7216 9956 7228
rect 10008 7216 10014 7268
rect 11882 7216 11888 7268
rect 11940 7256 11946 7268
rect 14461 7259 14519 7265
rect 14461 7256 14473 7259
rect 11940 7228 14473 7256
rect 11940 7216 11946 7228
rect 14461 7225 14473 7228
rect 14507 7225 14519 7259
rect 14461 7219 14519 7225
rect 15841 7259 15899 7265
rect 15841 7225 15853 7259
rect 15887 7256 15899 7259
rect 16022 7256 16028 7268
rect 15887 7228 16028 7256
rect 15887 7225 15899 7228
rect 15841 7219 15899 7225
rect 16022 7216 16028 7228
rect 16080 7216 16086 7268
rect 17512 7256 17540 7296
rect 17589 7293 17601 7327
rect 17635 7324 17647 7327
rect 17696 7324 17724 7355
rect 17862 7352 17868 7404
rect 17920 7392 17926 7404
rect 19334 7392 19340 7404
rect 17920 7364 19340 7392
rect 17920 7352 17926 7364
rect 19334 7352 19340 7364
rect 19392 7352 19398 7404
rect 21361 7395 21419 7401
rect 21361 7361 21373 7395
rect 21407 7392 21419 7395
rect 21726 7392 21732 7404
rect 21407 7364 21732 7392
rect 21407 7361 21419 7364
rect 21361 7355 21419 7361
rect 21726 7352 21732 7364
rect 21784 7352 21790 7404
rect 23937 7395 23995 7401
rect 23937 7361 23949 7395
rect 23983 7392 23995 7395
rect 28350 7392 28356 7404
rect 23983 7364 28356 7392
rect 23983 7361 23995 7364
rect 23937 7355 23995 7361
rect 28350 7352 28356 7364
rect 28408 7352 28414 7404
rect 30834 7352 30840 7404
rect 30892 7392 30898 7404
rect 31205 7395 31263 7401
rect 31205 7392 31217 7395
rect 30892 7364 31217 7392
rect 30892 7352 30898 7364
rect 31205 7361 31217 7364
rect 31251 7361 31263 7395
rect 31205 7355 31263 7361
rect 37734 7352 37740 7404
rect 37792 7352 37798 7404
rect 38105 7395 38163 7401
rect 38105 7361 38117 7395
rect 38151 7361 38163 7395
rect 38304 7392 38332 7491
rect 38746 7488 38752 7500
rect 38804 7488 38810 7540
rect 39025 7531 39083 7537
rect 39025 7497 39037 7531
rect 39071 7528 39083 7531
rect 39482 7528 39488 7540
rect 39071 7500 39488 7528
rect 39071 7497 39083 7500
rect 39025 7491 39083 7497
rect 39482 7488 39488 7500
rect 39540 7488 39546 7540
rect 38562 7420 38568 7472
rect 38620 7460 38626 7472
rect 38620 7432 39252 7460
rect 38620 7420 38626 7432
rect 38378 7392 38384 7404
rect 38304 7364 38384 7392
rect 38105 7355 38163 7361
rect 24486 7324 24492 7336
rect 17635 7296 17724 7324
rect 17788 7296 24492 7324
rect 17635 7293 17647 7296
rect 17589 7287 17647 7293
rect 17788 7256 17816 7296
rect 24486 7284 24492 7296
rect 24544 7284 24550 7336
rect 26878 7284 26884 7336
rect 26936 7324 26942 7336
rect 38120 7324 38148 7355
rect 38378 7352 38384 7364
rect 38436 7352 38442 7404
rect 38470 7352 38476 7404
rect 38528 7352 38534 7404
rect 39224 7401 39252 7432
rect 38841 7395 38899 7401
rect 38841 7361 38853 7395
rect 38887 7361 38899 7395
rect 38841 7355 38899 7361
rect 39209 7395 39267 7401
rect 39209 7361 39221 7395
rect 39255 7361 39267 7395
rect 39209 7355 39267 7361
rect 26936 7296 35296 7324
rect 26936 7284 26942 7296
rect 17512 7228 17816 7256
rect 17865 7259 17923 7265
rect 17865 7225 17877 7259
rect 17911 7256 17923 7259
rect 33686 7256 33692 7268
rect 17911 7228 33692 7256
rect 17911 7225 17923 7228
rect 17865 7219 17923 7225
rect 33686 7216 33692 7228
rect 33744 7216 33750 7268
rect 35268 7256 35296 7296
rect 37108 7296 38148 7324
rect 37108 7256 37136 7296
rect 38194 7284 38200 7336
rect 38252 7324 38258 7336
rect 38856 7324 38884 7355
rect 38252 7296 38884 7324
rect 38252 7284 38258 7296
rect 39482 7256 39488 7268
rect 35268 7228 37136 7256
rect 38304 7228 39488 7256
rect 7837 7191 7895 7197
rect 7837 7157 7849 7191
rect 7883 7188 7895 7191
rect 12158 7188 12164 7200
rect 7883 7160 12164 7188
rect 7883 7157 7895 7160
rect 7837 7151 7895 7157
rect 12158 7148 12164 7160
rect 12216 7148 12222 7200
rect 14093 7191 14151 7197
rect 14093 7157 14105 7191
rect 14139 7188 14151 7191
rect 17954 7188 17960 7200
rect 14139 7160 17960 7188
rect 14139 7157 14151 7160
rect 14093 7151 14151 7157
rect 17954 7148 17960 7160
rect 18012 7148 18018 7200
rect 19794 7148 19800 7200
rect 19852 7188 19858 7200
rect 31021 7191 31079 7197
rect 31021 7188 31033 7191
rect 19852 7160 31033 7188
rect 19852 7148 19858 7160
rect 31021 7157 31033 7160
rect 31067 7157 31079 7191
rect 31021 7151 31079 7157
rect 37921 7191 37979 7197
rect 37921 7157 37933 7191
rect 37967 7188 37979 7191
rect 38304 7188 38332 7228
rect 39482 7216 39488 7228
rect 39540 7216 39546 7268
rect 37967 7160 38332 7188
rect 37967 7157 37979 7160
rect 37921 7151 37979 7157
rect 39390 7148 39396 7200
rect 39448 7148 39454 7200
rect 1104 7098 39836 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 37950 7098
rect 38002 7046 38014 7098
rect 38066 7046 38078 7098
rect 38130 7046 38142 7098
rect 38194 7046 38206 7098
rect 38258 7046 39836 7098
rect 1104 7024 39836 7046
rect 12158 6944 12164 6996
rect 12216 6984 12222 6996
rect 17402 6984 17408 6996
rect 12216 6956 17408 6984
rect 12216 6944 12222 6956
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 19426 6944 19432 6996
rect 19484 6984 19490 6996
rect 26878 6984 26884 6996
rect 19484 6956 26884 6984
rect 19484 6944 19490 6956
rect 26878 6944 26884 6956
rect 26936 6944 26942 6996
rect 32858 6944 32864 6996
rect 32916 6984 32922 6996
rect 38838 6984 38844 6996
rect 32916 6956 38844 6984
rect 32916 6944 32922 6956
rect 38838 6944 38844 6956
rect 38896 6944 38902 6996
rect 9582 6876 9588 6928
rect 9640 6916 9646 6928
rect 22649 6919 22707 6925
rect 9640 6888 11744 6916
rect 9640 6876 9646 6888
rect 4614 6808 4620 6860
rect 4672 6848 4678 6860
rect 11716 6848 11744 6888
rect 22649 6885 22661 6919
rect 22695 6885 22707 6919
rect 22649 6879 22707 6885
rect 20530 6848 20536 6860
rect 4672 6820 11652 6848
rect 11716 6820 20536 6848
rect 4672 6808 4678 6820
rect 2593 6783 2651 6789
rect 2593 6749 2605 6783
rect 2639 6780 2651 6783
rect 2685 6783 2743 6789
rect 2685 6780 2697 6783
rect 2639 6752 2697 6780
rect 2639 6749 2651 6752
rect 2593 6743 2651 6749
rect 2685 6749 2697 6752
rect 2731 6780 2743 6783
rect 6270 6780 6276 6792
rect 2731 6752 6276 6780
rect 2731 6749 2743 6752
rect 2685 6743 2743 6749
rect 6270 6740 6276 6752
rect 6328 6740 6334 6792
rect 9309 6783 9367 6789
rect 9309 6749 9321 6783
rect 9355 6780 9367 6783
rect 9585 6783 9643 6789
rect 9585 6780 9597 6783
rect 9355 6752 9597 6780
rect 9355 6749 9367 6752
rect 9309 6743 9367 6749
rect 9585 6749 9597 6752
rect 9631 6780 9643 6783
rect 11054 6780 11060 6792
rect 9631 6752 11060 6780
rect 9631 6749 9643 6752
rect 9585 6743 9643 6749
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11624 6780 11652 6820
rect 20530 6808 20536 6820
rect 20588 6808 20594 6860
rect 22664 6848 22692 6879
rect 34146 6876 34152 6928
rect 34204 6916 34210 6928
rect 34204 6888 38884 6916
rect 34204 6876 34210 6888
rect 22664 6820 29960 6848
rect 19610 6780 19616 6792
rect 11624 6752 19616 6780
rect 19610 6740 19616 6752
rect 19668 6740 19674 6792
rect 22462 6740 22468 6792
rect 22520 6740 22526 6792
rect 25593 6783 25651 6789
rect 25593 6749 25605 6783
rect 25639 6780 25651 6783
rect 29086 6780 29092 6792
rect 25639 6752 29092 6780
rect 25639 6749 25651 6752
rect 25593 6743 25651 6749
rect 29086 6740 29092 6752
rect 29144 6740 29150 6792
rect 3786 6672 3792 6724
rect 3844 6712 3850 6724
rect 20806 6712 20812 6724
rect 3844 6684 9536 6712
rect 3844 6672 3850 6684
rect 2866 6604 2872 6656
rect 2924 6604 2930 6656
rect 7558 6604 7564 6656
rect 7616 6644 7622 6656
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 7616 6616 9413 6644
rect 7616 6604 7622 6616
rect 9401 6613 9413 6616
rect 9447 6613 9459 6647
rect 9508 6644 9536 6684
rect 9646 6684 20812 6712
rect 9646 6644 9674 6684
rect 20806 6672 20812 6684
rect 20864 6672 20870 6724
rect 29932 6712 29960 6820
rect 30009 6783 30067 6789
rect 30009 6749 30021 6783
rect 30055 6780 30067 6783
rect 30558 6780 30564 6792
rect 30055 6752 30564 6780
rect 30055 6749 30067 6752
rect 30009 6743 30067 6749
rect 30558 6740 30564 6752
rect 30616 6740 30622 6792
rect 31662 6740 31668 6792
rect 31720 6780 31726 6792
rect 34241 6783 34299 6789
rect 34241 6780 34253 6783
rect 31720 6752 34253 6780
rect 31720 6740 31726 6752
rect 34241 6749 34253 6752
rect 34287 6749 34299 6783
rect 34241 6743 34299 6749
rect 38470 6740 38476 6792
rect 38528 6740 38534 6792
rect 38856 6789 38884 6888
rect 38841 6783 38899 6789
rect 38841 6749 38853 6783
rect 38887 6749 38899 6783
rect 38841 6743 38899 6749
rect 38930 6740 38936 6792
rect 38988 6780 38994 6792
rect 39209 6783 39267 6789
rect 39209 6780 39221 6783
rect 38988 6752 39221 6780
rect 38988 6740 38994 6752
rect 39209 6749 39221 6752
rect 39255 6749 39267 6783
rect 39209 6743 39267 6749
rect 32674 6712 32680 6724
rect 22066 6684 29868 6712
rect 29932 6684 32680 6712
rect 9508 6616 9674 6644
rect 9401 6607 9459 6613
rect 11054 6604 11060 6656
rect 11112 6644 11118 6656
rect 12342 6644 12348 6656
rect 11112 6616 12348 6644
rect 11112 6604 11118 6616
rect 12342 6604 12348 6616
rect 12400 6604 12406 6656
rect 16390 6604 16396 6656
rect 16448 6644 16454 6656
rect 22066 6644 22094 6684
rect 16448 6616 22094 6644
rect 16448 6604 16454 6616
rect 24762 6604 24768 6656
rect 24820 6644 24826 6656
rect 29840 6653 29868 6684
rect 32674 6672 32680 6684
rect 32732 6672 32738 6724
rect 39666 6712 39672 6724
rect 39040 6684 39672 6712
rect 25409 6647 25467 6653
rect 25409 6644 25421 6647
rect 24820 6616 25421 6644
rect 24820 6604 24826 6616
rect 25409 6613 25421 6616
rect 25455 6613 25467 6647
rect 25409 6607 25467 6613
rect 29825 6647 29883 6653
rect 29825 6613 29837 6647
rect 29871 6613 29883 6647
rect 29825 6607 29883 6613
rect 30466 6604 30472 6656
rect 30524 6644 30530 6656
rect 34057 6647 34115 6653
rect 34057 6644 34069 6647
rect 30524 6616 34069 6644
rect 30524 6604 30530 6616
rect 34057 6613 34069 6616
rect 34103 6613 34115 6647
rect 34057 6607 34115 6613
rect 38654 6604 38660 6656
rect 38712 6604 38718 6656
rect 39040 6653 39068 6684
rect 39666 6672 39672 6684
rect 39724 6672 39730 6724
rect 39025 6647 39083 6653
rect 39025 6613 39037 6647
rect 39071 6613 39083 6647
rect 39025 6607 39083 6613
rect 39393 6647 39451 6653
rect 39393 6613 39405 6647
rect 39439 6644 39451 6647
rect 39574 6644 39580 6656
rect 39439 6616 39580 6644
rect 39439 6613 39451 6616
rect 39393 6607 39451 6613
rect 39574 6604 39580 6616
rect 39632 6604 39638 6656
rect 1104 6554 39836 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 39010 6554
rect 39062 6502 39074 6554
rect 39126 6502 39138 6554
rect 39190 6502 39202 6554
rect 39254 6502 39266 6554
rect 39318 6502 39836 6554
rect 1104 6480 39836 6502
rect 3237 6443 3295 6449
rect 3237 6409 3249 6443
rect 3283 6440 3295 6443
rect 3418 6440 3424 6452
rect 3283 6412 3424 6440
rect 3283 6409 3295 6412
rect 3237 6403 3295 6409
rect 3418 6400 3424 6412
rect 3476 6400 3482 6452
rect 3605 6443 3663 6449
rect 3605 6409 3617 6443
rect 3651 6440 3663 6443
rect 4062 6440 4068 6452
rect 3651 6412 4068 6440
rect 3651 6409 3663 6412
rect 3605 6403 3663 6409
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 4430 6400 4436 6452
rect 4488 6400 4494 6452
rect 7466 6400 7472 6452
rect 7524 6440 7530 6452
rect 7653 6443 7711 6449
rect 7653 6440 7665 6443
rect 7524 6412 7665 6440
rect 7524 6400 7530 6412
rect 7653 6409 7665 6412
rect 7699 6409 7711 6443
rect 7653 6403 7711 6409
rect 7742 6400 7748 6452
rect 7800 6440 7806 6452
rect 8297 6443 8355 6449
rect 8297 6440 8309 6443
rect 7800 6412 8309 6440
rect 7800 6400 7806 6412
rect 8297 6409 8309 6412
rect 8343 6409 8355 6443
rect 8297 6403 8355 6409
rect 10597 6443 10655 6449
rect 10597 6409 10609 6443
rect 10643 6409 10655 6443
rect 10597 6403 10655 6409
rect 2961 6375 3019 6381
rect 2961 6341 2973 6375
rect 3007 6372 3019 6375
rect 3510 6372 3516 6384
rect 3007 6344 3516 6372
rect 3007 6341 3019 6344
rect 2961 6335 3019 6341
rect 3068 6313 3096 6344
rect 3510 6332 3516 6344
rect 3568 6332 3574 6384
rect 3786 6332 3792 6384
rect 3844 6332 3850 6384
rect 8202 6332 8208 6384
rect 8260 6372 8266 6384
rect 10612 6372 10640 6403
rect 11514 6400 11520 6452
rect 11572 6440 11578 6452
rect 11609 6443 11667 6449
rect 11609 6440 11621 6443
rect 11572 6412 11621 6440
rect 11572 6400 11578 6412
rect 11609 6409 11621 6412
rect 11655 6409 11667 6443
rect 21634 6440 21640 6452
rect 11609 6403 11667 6409
rect 11716 6412 21640 6440
rect 8260 6344 10640 6372
rect 8260 6332 8266 6344
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6304 3111 6307
rect 3421 6307 3479 6313
rect 3099 6276 3133 6304
rect 3099 6273 3111 6276
rect 3053 6267 3111 6273
rect 3421 6273 3433 6307
rect 3467 6304 3479 6307
rect 3697 6307 3755 6313
rect 3697 6304 3709 6307
rect 3467 6276 3709 6304
rect 3467 6273 3479 6276
rect 3421 6267 3479 6273
rect 3697 6273 3709 6276
rect 3743 6273 3755 6307
rect 3697 6267 3755 6273
rect 4614 6264 4620 6316
rect 4672 6264 4678 6316
rect 7374 6264 7380 6316
rect 7432 6304 7438 6316
rect 7837 6307 7895 6313
rect 7837 6304 7849 6307
rect 7432 6276 7849 6304
rect 7432 6264 7438 6276
rect 7837 6273 7849 6276
rect 7883 6273 7895 6307
rect 7837 6267 7895 6273
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6304 8171 6307
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 8159 6276 8493 6304
rect 8159 6273 8171 6276
rect 8113 6267 8171 6273
rect 8481 6273 8493 6276
rect 8527 6304 8539 6307
rect 8757 6307 8815 6313
rect 8527 6276 8708 6304
rect 8527 6273 8539 6276
rect 8481 6267 8539 6273
rect 7650 6128 7656 6180
rect 7708 6168 7714 6180
rect 8573 6171 8631 6177
rect 8573 6168 8585 6171
rect 7708 6140 8585 6168
rect 7708 6128 7714 6140
rect 8573 6137 8585 6140
rect 8619 6137 8631 6171
rect 8680 6168 8708 6276
rect 8757 6273 8769 6307
rect 8803 6304 8815 6307
rect 10686 6304 10692 6316
rect 8803 6276 10692 6304
rect 8803 6273 8815 6276
rect 8757 6267 8815 6273
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6304 10839 6307
rect 11716 6304 11744 6412
rect 21634 6400 21640 6412
rect 21692 6400 21698 6452
rect 26418 6400 26424 6452
rect 26476 6400 26482 6452
rect 29273 6443 29331 6449
rect 29273 6409 29285 6443
rect 29319 6409 29331 6443
rect 29273 6403 29331 6409
rect 25866 6372 25872 6384
rect 11808 6344 25872 6372
rect 11808 6313 11836 6344
rect 25866 6332 25872 6344
rect 25924 6332 25930 6384
rect 10827 6276 11744 6304
rect 11793 6307 11851 6313
rect 10827 6273 10839 6276
rect 10781 6267 10839 6273
rect 11793 6273 11805 6307
rect 11839 6273 11851 6307
rect 11793 6267 11851 6273
rect 11882 6264 11888 6316
rect 11940 6304 11946 6316
rect 18874 6304 18880 6316
rect 11940 6276 18880 6304
rect 11940 6264 11946 6276
rect 18874 6264 18880 6276
rect 18932 6264 18938 6316
rect 19150 6264 19156 6316
rect 19208 6304 19214 6316
rect 19337 6307 19395 6313
rect 19337 6304 19349 6307
rect 19208 6276 19349 6304
rect 19208 6264 19214 6276
rect 19337 6273 19349 6276
rect 19383 6273 19395 6307
rect 19337 6267 19395 6273
rect 23842 6264 23848 6316
rect 23900 6304 23906 6316
rect 24213 6307 24271 6313
rect 24213 6304 24225 6307
rect 23900 6276 24225 6304
rect 23900 6264 23906 6276
rect 24213 6273 24225 6276
rect 24259 6273 24271 6307
rect 24213 6267 24271 6273
rect 26605 6307 26663 6313
rect 26605 6273 26617 6307
rect 26651 6304 26663 6307
rect 29178 6304 29184 6316
rect 26651 6276 29184 6304
rect 26651 6273 26663 6276
rect 26605 6267 26663 6273
rect 29178 6264 29184 6276
rect 29236 6264 29242 6316
rect 15838 6196 15844 6248
rect 15896 6236 15902 6248
rect 29288 6236 29316 6403
rect 39390 6400 39396 6452
rect 39448 6400 39454 6452
rect 31018 6332 31024 6384
rect 31076 6372 31082 6384
rect 35894 6372 35900 6384
rect 31076 6344 35900 6372
rect 31076 6332 31082 6344
rect 35894 6332 35900 6344
rect 35952 6332 35958 6384
rect 29457 6307 29515 6313
rect 29457 6273 29469 6307
rect 29503 6304 29515 6307
rect 30282 6304 30288 6316
rect 29503 6276 30288 6304
rect 29503 6273 29515 6276
rect 29457 6267 29515 6273
rect 30282 6264 30288 6276
rect 30340 6264 30346 6316
rect 34330 6264 34336 6316
rect 34388 6304 34394 6316
rect 38841 6307 38899 6313
rect 38841 6304 38853 6307
rect 34388 6276 38853 6304
rect 34388 6264 34394 6276
rect 38841 6273 38853 6276
rect 38887 6273 38899 6307
rect 38841 6267 38899 6273
rect 39206 6264 39212 6316
rect 39264 6264 39270 6316
rect 15896 6208 29316 6236
rect 15896 6196 15902 6208
rect 29362 6196 29368 6248
rect 29420 6236 29426 6248
rect 37734 6236 37740 6248
rect 29420 6208 37740 6236
rect 29420 6196 29426 6208
rect 37734 6196 37740 6208
rect 37792 6196 37798 6248
rect 16114 6168 16120 6180
rect 8680 6140 16120 6168
rect 8573 6131 8631 6137
rect 16114 6128 16120 6140
rect 16172 6128 16178 6180
rect 19521 6171 19579 6177
rect 19521 6137 19533 6171
rect 19567 6168 19579 6171
rect 24397 6171 24455 6177
rect 19567 6140 22094 6168
rect 19567 6137 19579 6140
rect 19521 6131 19579 6137
rect 11606 6060 11612 6112
rect 11664 6100 11670 6112
rect 17126 6100 17132 6112
rect 11664 6072 17132 6100
rect 11664 6060 11670 6072
rect 17126 6060 17132 6072
rect 17184 6060 17190 6112
rect 22066 6100 22094 6140
rect 24397 6137 24409 6171
rect 24443 6168 24455 6171
rect 38746 6168 38752 6180
rect 24443 6140 38752 6168
rect 24443 6137 24455 6140
rect 24397 6131 24455 6137
rect 38746 6128 38752 6140
rect 38804 6128 38810 6180
rect 38470 6100 38476 6112
rect 22066 6072 38476 6100
rect 38470 6060 38476 6072
rect 38528 6060 38534 6112
rect 39022 6060 39028 6112
rect 39080 6060 39086 6112
rect 1104 6010 39836 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 37950 6010
rect 38002 5958 38014 6010
rect 38066 5958 38078 6010
rect 38130 5958 38142 6010
rect 38194 5958 38206 6010
rect 38258 5958 39836 6010
rect 1104 5936 39836 5958
rect 3973 5899 4031 5905
rect 3973 5865 3985 5899
rect 4019 5896 4031 5899
rect 4154 5896 4160 5908
rect 4019 5868 4160 5896
rect 4019 5865 4031 5868
rect 3973 5859 4031 5865
rect 4154 5856 4160 5868
rect 4212 5856 4218 5908
rect 4893 5899 4951 5905
rect 4893 5865 4905 5899
rect 4939 5896 4951 5899
rect 4982 5896 4988 5908
rect 4939 5868 4988 5896
rect 4939 5865 4951 5868
rect 4893 5859 4951 5865
rect 4982 5856 4988 5868
rect 5040 5856 5046 5908
rect 5442 5856 5448 5908
rect 5500 5896 5506 5908
rect 5537 5899 5595 5905
rect 5537 5896 5549 5899
rect 5500 5868 5549 5896
rect 5500 5856 5506 5868
rect 5537 5865 5549 5868
rect 5583 5865 5595 5899
rect 5537 5859 5595 5865
rect 5810 5856 5816 5908
rect 5868 5896 5874 5908
rect 6641 5899 6699 5905
rect 6641 5896 6653 5899
rect 5868 5868 6653 5896
rect 5868 5856 5874 5868
rect 6641 5865 6653 5868
rect 6687 5865 6699 5899
rect 6641 5859 6699 5865
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7101 5899 7159 5905
rect 7101 5896 7113 5899
rect 6972 5868 7113 5896
rect 6972 5856 6978 5868
rect 7101 5865 7113 5868
rect 7147 5865 7159 5899
rect 7101 5859 7159 5865
rect 11238 5856 11244 5908
rect 11296 5896 11302 5908
rect 11609 5899 11667 5905
rect 11609 5896 11621 5899
rect 11296 5868 11621 5896
rect 11296 5856 11302 5868
rect 11609 5865 11621 5868
rect 11655 5865 11667 5899
rect 11609 5859 11667 5865
rect 26053 5899 26111 5905
rect 26053 5865 26065 5899
rect 26099 5896 26111 5899
rect 30374 5896 30380 5908
rect 26099 5868 30380 5896
rect 26099 5865 26111 5868
rect 26053 5859 26111 5865
rect 30374 5856 30380 5868
rect 30432 5856 30438 5908
rect 35437 5899 35495 5905
rect 35437 5865 35449 5899
rect 35483 5896 35495 5899
rect 35802 5896 35808 5908
rect 35483 5868 35808 5896
rect 35483 5865 35495 5868
rect 35437 5859 35495 5865
rect 35802 5856 35808 5868
rect 35860 5856 35866 5908
rect 35894 5856 35900 5908
rect 35952 5896 35958 5908
rect 37001 5899 37059 5905
rect 37001 5896 37013 5899
rect 35952 5868 37013 5896
rect 35952 5856 35958 5868
rect 37001 5865 37013 5868
rect 37047 5865 37059 5899
rect 37001 5859 37059 5865
rect 38105 5899 38163 5905
rect 38105 5865 38117 5899
rect 38151 5896 38163 5899
rect 38286 5896 38292 5908
rect 38151 5868 38292 5896
rect 38151 5865 38163 5868
rect 38105 5859 38163 5865
rect 38286 5856 38292 5868
rect 38344 5856 38350 5908
rect 38746 5856 38752 5908
rect 38804 5896 38810 5908
rect 39758 5896 39764 5908
rect 38804 5868 39764 5896
rect 38804 5856 38810 5868
rect 39758 5856 39764 5868
rect 39816 5856 39822 5908
rect 11882 5828 11888 5840
rect 5736 5800 11888 5828
rect 4157 5763 4215 5769
rect 4157 5729 4169 5763
rect 4203 5760 4215 5763
rect 5534 5760 5540 5772
rect 4203 5732 5540 5760
rect 4203 5729 4215 5732
rect 4157 5723 4215 5729
rect 5534 5720 5540 5732
rect 5592 5720 5598 5772
rect 5736 5701 5764 5800
rect 11882 5788 11888 5800
rect 11940 5788 11946 5840
rect 19518 5828 19524 5840
rect 12406 5800 19524 5828
rect 12406 5760 12434 5800
rect 19518 5788 19524 5800
rect 19576 5788 19582 5840
rect 27614 5788 27620 5840
rect 27672 5828 27678 5840
rect 39206 5828 39212 5840
rect 27672 5800 39212 5828
rect 27672 5788 27678 5800
rect 39206 5788 39212 5800
rect 39264 5788 39270 5840
rect 39390 5788 39396 5840
rect 39448 5788 39454 5840
rect 16206 5760 16212 5772
rect 6840 5732 12434 5760
rect 15304 5732 16212 5760
rect 6840 5701 6868 5732
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5692 3847 5695
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 3835 5664 4077 5692
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 4065 5661 4077 5664
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5661 5135 5695
rect 5077 5655 5135 5661
rect 5721 5695 5779 5701
rect 5721 5661 5733 5695
rect 5767 5661 5779 5695
rect 5721 5655 5779 5661
rect 6825 5695 6883 5701
rect 6825 5661 6837 5695
rect 6871 5661 6883 5695
rect 6825 5655 6883 5661
rect 7285 5695 7343 5701
rect 7285 5661 7297 5695
rect 7331 5692 7343 5695
rect 11793 5695 11851 5701
rect 7331 5664 11744 5692
rect 7331 5661 7343 5664
rect 7285 5655 7343 5661
rect 5092 5624 5120 5655
rect 9582 5624 9588 5636
rect 5092 5596 9588 5624
rect 9582 5584 9588 5596
rect 9640 5584 9646 5636
rect 11716 5624 11744 5664
rect 11793 5661 11805 5695
rect 11839 5692 11851 5695
rect 15304 5692 15332 5732
rect 16206 5720 16212 5732
rect 16264 5720 16270 5772
rect 20438 5720 20444 5772
rect 20496 5760 20502 5772
rect 20496 5732 31754 5760
rect 20496 5720 20502 5732
rect 11839 5664 15332 5692
rect 11839 5661 11851 5664
rect 11793 5655 11851 5661
rect 15378 5652 15384 5704
rect 15436 5692 15442 5704
rect 18417 5695 18475 5701
rect 15436 5664 18368 5692
rect 15436 5652 15442 5664
rect 16482 5624 16488 5636
rect 11716 5596 16488 5624
rect 16482 5584 16488 5596
rect 16540 5584 16546 5636
rect 18340 5624 18368 5664
rect 18417 5661 18429 5695
rect 18463 5692 18475 5695
rect 18509 5695 18567 5701
rect 18509 5692 18521 5695
rect 18463 5664 18521 5692
rect 18463 5661 18475 5664
rect 18417 5655 18475 5661
rect 18509 5661 18521 5664
rect 18555 5661 18567 5695
rect 18509 5655 18567 5661
rect 25866 5652 25872 5704
rect 25924 5652 25930 5704
rect 28261 5695 28319 5701
rect 28261 5661 28273 5695
rect 28307 5692 28319 5695
rect 30006 5692 30012 5704
rect 28307 5664 30012 5692
rect 28307 5661 28319 5664
rect 28261 5655 28319 5661
rect 30006 5652 30012 5664
rect 30064 5652 30070 5704
rect 31726 5692 31754 5732
rect 35360 5732 38884 5760
rect 35253 5695 35311 5701
rect 35253 5692 35265 5695
rect 31726 5664 35265 5692
rect 35253 5661 35265 5664
rect 35299 5661 35311 5695
rect 35253 5655 35311 5661
rect 18340 5596 28120 5624
rect 14918 5516 14924 5568
rect 14976 5556 14982 5568
rect 18325 5559 18383 5565
rect 18325 5556 18337 5559
rect 14976 5528 18337 5556
rect 14976 5516 14982 5528
rect 18325 5525 18337 5528
rect 18371 5525 18383 5559
rect 18325 5519 18383 5525
rect 18693 5559 18751 5565
rect 18693 5525 18705 5559
rect 18739 5556 18751 5559
rect 26142 5556 26148 5568
rect 18739 5528 26148 5556
rect 18739 5525 18751 5528
rect 18693 5519 18751 5525
rect 26142 5516 26148 5528
rect 26200 5516 26206 5568
rect 28092 5565 28120 5596
rect 28077 5559 28135 5565
rect 28077 5525 28089 5559
rect 28123 5525 28135 5559
rect 28077 5519 28135 5525
rect 28994 5516 29000 5568
rect 29052 5556 29058 5568
rect 35360 5556 35388 5732
rect 35621 5695 35679 5701
rect 35621 5661 35633 5695
rect 35667 5661 35679 5695
rect 35621 5655 35679 5661
rect 35636 5624 35664 5655
rect 37090 5652 37096 5704
rect 37148 5692 37154 5704
rect 37185 5695 37243 5701
rect 37185 5692 37197 5695
rect 37148 5664 37197 5692
rect 37148 5652 37154 5664
rect 37185 5661 37197 5664
rect 37231 5661 37243 5695
rect 37185 5655 37243 5661
rect 38289 5695 38347 5701
rect 38289 5661 38301 5695
rect 38335 5692 38347 5695
rect 38746 5692 38752 5704
rect 38335 5664 38752 5692
rect 38335 5661 38347 5664
rect 38289 5655 38347 5661
rect 38746 5652 38752 5664
rect 38804 5652 38810 5704
rect 38856 5701 38884 5732
rect 38841 5695 38899 5701
rect 38841 5661 38853 5695
rect 38887 5661 38899 5695
rect 39209 5695 39267 5701
rect 39209 5692 39221 5695
rect 38841 5655 38899 5661
rect 38948 5664 39221 5692
rect 37826 5624 37832 5636
rect 35636 5596 37832 5624
rect 37826 5584 37832 5596
rect 37884 5584 37890 5636
rect 29052 5528 35388 5556
rect 29052 5516 29058 5528
rect 35618 5516 35624 5568
rect 35676 5556 35682 5568
rect 35805 5559 35863 5565
rect 35805 5556 35817 5559
rect 35676 5528 35817 5556
rect 35676 5516 35682 5528
rect 35805 5525 35817 5528
rect 35851 5525 35863 5559
rect 35805 5519 35863 5525
rect 36078 5516 36084 5568
rect 36136 5556 36142 5568
rect 38948 5556 38976 5664
rect 39209 5661 39221 5664
rect 39255 5661 39267 5695
rect 39209 5655 39267 5661
rect 36136 5528 38976 5556
rect 39025 5559 39083 5565
rect 36136 5516 36142 5528
rect 39025 5525 39037 5559
rect 39071 5556 39083 5559
rect 39942 5556 39948 5568
rect 39071 5528 39948 5556
rect 39071 5525 39083 5528
rect 39025 5519 39083 5525
rect 39942 5516 39948 5528
rect 40000 5516 40006 5568
rect 1104 5466 39836 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 39010 5466
rect 39062 5414 39074 5466
rect 39126 5414 39138 5466
rect 39190 5414 39202 5466
rect 39254 5414 39266 5466
rect 39318 5414 39836 5466
rect 1104 5392 39836 5414
rect 5074 5312 5080 5364
rect 5132 5352 5138 5364
rect 5353 5355 5411 5361
rect 5353 5352 5365 5355
rect 5132 5324 5365 5352
rect 5132 5312 5138 5324
rect 5353 5321 5365 5324
rect 5399 5321 5411 5355
rect 5353 5315 5411 5321
rect 5813 5355 5871 5361
rect 5813 5321 5825 5355
rect 5859 5352 5871 5355
rect 6638 5352 6644 5364
rect 5859 5324 6644 5352
rect 5859 5321 5871 5324
rect 5813 5315 5871 5321
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 12250 5312 12256 5364
rect 12308 5352 12314 5364
rect 12989 5355 13047 5361
rect 12989 5352 13001 5355
rect 12308 5324 13001 5352
rect 12308 5312 12314 5324
rect 12989 5321 13001 5324
rect 13035 5321 13047 5355
rect 12989 5315 13047 5321
rect 15841 5355 15899 5361
rect 15841 5321 15853 5355
rect 15887 5321 15899 5355
rect 15841 5315 15899 5321
rect 16853 5355 16911 5361
rect 16853 5321 16865 5355
rect 16899 5352 16911 5355
rect 27614 5352 27620 5364
rect 16899 5324 27620 5352
rect 16899 5321 16911 5324
rect 16853 5315 16911 5321
rect 10962 5244 10968 5296
rect 11020 5284 11026 5296
rect 15856 5284 15884 5315
rect 27614 5312 27620 5324
rect 27672 5312 27678 5364
rect 39390 5312 39396 5364
rect 39448 5312 39454 5364
rect 19058 5284 19064 5296
rect 11020 5256 15884 5284
rect 16040 5256 19064 5284
rect 11020 5244 11026 5256
rect 5534 5176 5540 5228
rect 5592 5176 5598 5228
rect 5629 5219 5687 5225
rect 5629 5185 5641 5219
rect 5675 5216 5687 5219
rect 13173 5219 13231 5225
rect 5675 5188 6914 5216
rect 5675 5185 5687 5188
rect 5629 5179 5687 5185
rect 6886 5080 6914 5188
rect 13173 5185 13185 5219
rect 13219 5216 13231 5219
rect 13538 5216 13544 5228
rect 13219 5188 13544 5216
rect 13219 5185 13231 5188
rect 13173 5179 13231 5185
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 16040 5225 16068 5256
rect 19058 5244 19064 5256
rect 19116 5244 19122 5296
rect 16025 5219 16083 5225
rect 16025 5185 16037 5219
rect 16071 5185 16083 5219
rect 16025 5179 16083 5185
rect 16666 5176 16672 5228
rect 16724 5216 16730 5228
rect 16945 5219 17003 5225
rect 16945 5216 16957 5219
rect 16724 5188 16957 5216
rect 16724 5176 16730 5188
rect 16945 5185 16957 5188
rect 16991 5185 17003 5219
rect 16945 5179 17003 5185
rect 17310 5176 17316 5228
rect 17368 5176 17374 5228
rect 17865 5219 17923 5225
rect 17865 5185 17877 5219
rect 17911 5216 17923 5219
rect 19794 5216 19800 5228
rect 17911 5188 19800 5216
rect 17911 5185 17923 5188
rect 17865 5179 17923 5185
rect 19794 5176 19800 5188
rect 19852 5176 19858 5228
rect 22005 5219 22063 5225
rect 22005 5185 22017 5219
rect 22051 5216 22063 5219
rect 24578 5216 24584 5228
rect 22051 5188 24584 5216
rect 22051 5185 22063 5188
rect 22005 5179 22063 5185
rect 24578 5176 24584 5188
rect 24636 5176 24642 5228
rect 27157 5219 27215 5225
rect 27157 5185 27169 5219
rect 27203 5216 27215 5219
rect 27522 5216 27528 5228
rect 27203 5188 27528 5216
rect 27203 5185 27215 5188
rect 27157 5179 27215 5185
rect 27522 5176 27528 5188
rect 27580 5176 27586 5228
rect 37274 5176 37280 5228
rect 37332 5216 37338 5228
rect 38841 5219 38899 5225
rect 38841 5216 38853 5219
rect 37332 5188 38853 5216
rect 37332 5176 37338 5188
rect 38841 5185 38853 5188
rect 38887 5185 38899 5219
rect 38841 5179 38899 5185
rect 39209 5219 39267 5225
rect 39209 5185 39221 5219
rect 39255 5185 39267 5219
rect 39209 5179 39267 5185
rect 15654 5148 15660 5160
rect 12406 5120 15660 5148
rect 12406 5080 12434 5120
rect 15654 5108 15660 5120
rect 15712 5108 15718 5160
rect 16758 5108 16764 5160
rect 16816 5148 16822 5160
rect 29362 5148 29368 5160
rect 16816 5120 29368 5148
rect 16816 5108 16822 5120
rect 29362 5108 29368 5120
rect 29420 5108 29426 5160
rect 35986 5108 35992 5160
rect 36044 5148 36050 5160
rect 39224 5148 39252 5179
rect 36044 5120 39252 5148
rect 36044 5108 36050 5120
rect 6886 5052 12434 5080
rect 17126 5040 17132 5092
rect 17184 5040 17190 5092
rect 18049 5083 18107 5089
rect 18049 5049 18061 5083
rect 18095 5080 18107 5083
rect 22738 5080 22744 5092
rect 18095 5052 22744 5080
rect 18095 5049 18107 5052
rect 18049 5043 18107 5049
rect 22738 5040 22744 5052
rect 22796 5040 22802 5092
rect 26142 5040 26148 5092
rect 26200 5080 26206 5092
rect 38654 5080 38660 5092
rect 26200 5052 38660 5080
rect 26200 5040 26206 5052
rect 38654 5040 38660 5052
rect 38712 5040 38718 5092
rect 21818 4972 21824 5024
rect 21876 4972 21882 5024
rect 22922 4972 22928 5024
rect 22980 5012 22986 5024
rect 26973 5015 27031 5021
rect 26973 5012 26985 5015
rect 22980 4984 26985 5012
rect 22980 4972 22986 4984
rect 26973 4981 26985 4984
rect 27019 4981 27031 5015
rect 26973 4975 27031 4981
rect 39022 4972 39028 5024
rect 39080 4972 39086 5024
rect 1104 4922 39836 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 37950 4922
rect 38002 4870 38014 4922
rect 38066 4870 38078 4922
rect 38130 4870 38142 4922
rect 38194 4870 38206 4922
rect 38258 4870 39836 4922
rect 1104 4848 39836 4870
rect 10870 4768 10876 4820
rect 10928 4808 10934 4820
rect 14645 4811 14703 4817
rect 14645 4808 14657 4811
rect 10928 4780 14657 4808
rect 10928 4768 10934 4780
rect 14645 4777 14657 4780
rect 14691 4777 14703 4811
rect 14645 4771 14703 4777
rect 16298 4768 16304 4820
rect 16356 4768 16362 4820
rect 16669 4811 16727 4817
rect 16669 4777 16681 4811
rect 16715 4808 16727 4811
rect 16758 4808 16764 4820
rect 16715 4780 16764 4808
rect 16715 4777 16727 4780
rect 16669 4771 16727 4777
rect 16758 4768 16764 4780
rect 16816 4768 16822 4820
rect 17862 4768 17868 4820
rect 17920 4808 17926 4820
rect 18693 4811 18751 4817
rect 18693 4808 18705 4811
rect 17920 4780 18705 4808
rect 17920 4768 17926 4780
rect 18693 4777 18705 4780
rect 18739 4777 18751 4811
rect 32858 4808 32864 4820
rect 18693 4771 18751 4777
rect 22066 4780 32864 4808
rect 11057 4743 11115 4749
rect 11057 4709 11069 4743
rect 11103 4740 11115 4743
rect 11146 4740 11152 4752
rect 11103 4712 11152 4740
rect 11103 4709 11115 4712
rect 11057 4703 11115 4709
rect 11146 4700 11152 4712
rect 11204 4700 11210 4752
rect 18414 4700 18420 4752
rect 18472 4740 18478 4752
rect 22066 4740 22094 4780
rect 32858 4768 32864 4780
rect 32916 4768 32922 4820
rect 33778 4768 33784 4820
rect 33836 4768 33842 4820
rect 18472 4712 22094 4740
rect 23753 4743 23811 4749
rect 18472 4700 18478 4712
rect 23753 4709 23765 4743
rect 23799 4740 23811 4743
rect 24026 4740 24032 4752
rect 23799 4712 24032 4740
rect 23799 4709 23811 4712
rect 23753 4703 23811 4709
rect 24026 4700 24032 4712
rect 24084 4700 24090 4752
rect 24121 4743 24179 4749
rect 24121 4709 24133 4743
rect 24167 4740 24179 4743
rect 24167 4712 31754 4740
rect 24167 4709 24179 4712
rect 24121 4703 24179 4709
rect 5534 4632 5540 4684
rect 5592 4672 5598 4684
rect 5592 4644 11744 4672
rect 5592 4632 5598 4644
rect 11057 4607 11115 4613
rect 11057 4573 11069 4607
rect 11103 4604 11115 4607
rect 11241 4607 11299 4613
rect 11241 4604 11253 4607
rect 11103 4576 11253 4604
rect 11103 4573 11115 4576
rect 11057 4567 11115 4573
rect 11241 4573 11253 4576
rect 11287 4573 11299 4607
rect 11241 4567 11299 4573
rect 11422 4496 11428 4548
rect 11480 4496 11486 4548
rect 11716 4536 11744 4644
rect 15930 4632 15936 4684
rect 15988 4672 15994 4684
rect 21818 4672 21824 4684
rect 15988 4644 21824 4672
rect 15988 4632 15994 4644
rect 21818 4632 21824 4644
rect 21876 4632 21882 4684
rect 24302 4672 24308 4684
rect 22066 4644 24308 4672
rect 14826 4564 14832 4616
rect 14884 4564 14890 4616
rect 16393 4607 16451 4613
rect 16393 4573 16405 4607
rect 16439 4604 16451 4607
rect 16485 4607 16543 4613
rect 16485 4604 16497 4607
rect 16439 4576 16497 4604
rect 16439 4573 16451 4576
rect 16393 4567 16451 4573
rect 16485 4573 16497 4576
rect 16531 4573 16543 4607
rect 16485 4567 16543 4573
rect 18785 4607 18843 4613
rect 18785 4573 18797 4607
rect 18831 4604 18843 4607
rect 18877 4607 18935 4613
rect 18877 4604 18889 4607
rect 18831 4576 18889 4604
rect 18831 4573 18843 4576
rect 18785 4567 18843 4573
rect 18877 4573 18889 4576
rect 18923 4573 18935 4607
rect 18877 4567 18935 4573
rect 20349 4607 20407 4613
rect 20349 4573 20361 4607
rect 20395 4604 20407 4607
rect 22066 4604 22094 4644
rect 24302 4632 24308 4644
rect 24360 4632 24366 4684
rect 31726 4672 31754 4712
rect 39390 4700 39396 4752
rect 39448 4700 39454 4752
rect 36170 4672 36176 4684
rect 31726 4644 36176 4672
rect 36170 4632 36176 4644
rect 36228 4632 36234 4684
rect 20395 4576 22094 4604
rect 23569 4607 23627 4613
rect 20395 4573 20407 4576
rect 20349 4567 20407 4573
rect 23569 4573 23581 4607
rect 23615 4604 23627 4607
rect 23842 4604 23848 4616
rect 23615 4576 23848 4604
rect 23615 4573 23627 4576
rect 23569 4567 23627 4573
rect 23842 4564 23848 4576
rect 23900 4564 23906 4616
rect 23937 4607 23995 4613
rect 23937 4573 23949 4607
rect 23983 4604 23995 4607
rect 28074 4604 28080 4616
rect 23983 4576 28080 4604
rect 23983 4573 23995 4576
rect 23937 4567 23995 4573
rect 28074 4564 28080 4576
rect 28132 4564 28138 4616
rect 28169 4607 28227 4613
rect 28169 4573 28181 4607
rect 28215 4604 28227 4607
rect 30098 4604 30104 4616
rect 28215 4576 30104 4604
rect 28215 4573 28227 4576
rect 28169 4567 28227 4573
rect 30098 4564 30104 4576
rect 30156 4564 30162 4616
rect 31849 4607 31907 4613
rect 31849 4573 31861 4607
rect 31895 4573 31907 4607
rect 31849 4567 31907 4573
rect 33597 4607 33655 4613
rect 33597 4573 33609 4607
rect 33643 4604 33655 4607
rect 35894 4604 35900 4616
rect 33643 4576 35900 4604
rect 33643 4573 33655 4576
rect 33597 4567 33655 4573
rect 19702 4536 19708 4548
rect 11716 4508 19708 4536
rect 19702 4496 19708 4508
rect 19760 4496 19766 4548
rect 31018 4536 31024 4548
rect 22066 4508 31024 4536
rect 19058 4428 19064 4480
rect 19116 4428 19122 4480
rect 20533 4471 20591 4477
rect 20533 4437 20545 4471
rect 20579 4468 20591 4471
rect 22066 4468 22094 4508
rect 31018 4496 31024 4508
rect 31076 4496 31082 4548
rect 31864 4536 31892 4567
rect 35894 4564 35900 4576
rect 35952 4564 35958 4616
rect 38838 4564 38844 4616
rect 38896 4564 38902 4616
rect 38930 4564 38936 4616
rect 38988 4604 38994 4616
rect 39209 4607 39267 4613
rect 39209 4604 39221 4607
rect 38988 4576 39221 4604
rect 38988 4564 38994 4576
rect 39209 4573 39221 4576
rect 39255 4573 39267 4607
rect 39209 4567 39267 4573
rect 33962 4536 33968 4548
rect 31864 4508 33968 4536
rect 33962 4496 33968 4508
rect 34020 4496 34026 4548
rect 20579 4440 22094 4468
rect 28353 4471 28411 4477
rect 20579 4437 20591 4440
rect 20533 4431 20591 4437
rect 28353 4437 28365 4471
rect 28399 4468 28411 4471
rect 30742 4468 30748 4480
rect 28399 4440 30748 4468
rect 28399 4437 28411 4440
rect 28353 4431 28411 4437
rect 30742 4428 30748 4440
rect 30800 4428 30806 4480
rect 32033 4471 32091 4477
rect 32033 4437 32045 4471
rect 32079 4468 32091 4471
rect 37182 4468 37188 4480
rect 32079 4440 37188 4468
rect 32079 4437 32091 4440
rect 32033 4431 32091 4437
rect 37182 4428 37188 4440
rect 37240 4428 37246 4480
rect 39025 4471 39083 4477
rect 39025 4437 39037 4471
rect 39071 4468 39083 4471
rect 39942 4468 39948 4480
rect 39071 4440 39948 4468
rect 39071 4437 39083 4440
rect 39025 4431 39083 4437
rect 39942 4428 39948 4440
rect 40000 4428 40006 4480
rect 1104 4378 39836 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 39010 4378
rect 39062 4326 39074 4378
rect 39126 4326 39138 4378
rect 39190 4326 39202 4378
rect 39254 4326 39266 4378
rect 39318 4326 39836 4378
rect 1104 4304 39836 4326
rect 13817 4267 13875 4273
rect 13817 4233 13829 4267
rect 13863 4233 13875 4267
rect 13817 4227 13875 4233
rect 5718 4156 5724 4208
rect 5776 4156 5782 4208
rect 8294 4156 8300 4208
rect 8352 4196 8358 4208
rect 9769 4199 9827 4205
rect 9769 4196 9781 4199
rect 8352 4168 9781 4196
rect 8352 4156 8358 4168
rect 9769 4165 9781 4168
rect 9815 4165 9827 4199
rect 9769 4159 9827 4165
rect 8202 4088 8208 4140
rect 8260 4128 8266 4140
rect 13633 4131 13691 4137
rect 13633 4128 13645 4131
rect 8260 4100 13645 4128
rect 8260 4088 8266 4100
rect 13633 4097 13645 4100
rect 13679 4097 13691 4131
rect 13633 4091 13691 4097
rect 13832 4060 13860 4227
rect 19058 4224 19064 4276
rect 19116 4264 19122 4276
rect 38838 4264 38844 4276
rect 19116 4236 38844 4264
rect 19116 4224 19122 4236
rect 38838 4224 38844 4236
rect 38896 4224 38902 4276
rect 14826 4156 14832 4208
rect 14884 4196 14890 4208
rect 25590 4196 25596 4208
rect 14884 4168 25596 4196
rect 14884 4156 14890 4168
rect 25590 4156 25596 4168
rect 25648 4156 25654 4208
rect 38930 4196 38936 4208
rect 27632 4168 38936 4196
rect 20714 4088 20720 4140
rect 20772 4128 20778 4140
rect 23017 4131 23075 4137
rect 23017 4128 23029 4131
rect 20772 4100 23029 4128
rect 20772 4088 20778 4100
rect 23017 4097 23029 4100
rect 23063 4128 23075 4131
rect 23201 4131 23259 4137
rect 23201 4128 23213 4131
rect 23063 4100 23213 4128
rect 23063 4097 23075 4100
rect 23017 4091 23075 4097
rect 23201 4097 23213 4100
rect 23247 4097 23259 4131
rect 27632 4128 27660 4168
rect 38930 4156 38936 4168
rect 38988 4156 38994 4208
rect 23201 4091 23259 4097
rect 23308 4100 27660 4128
rect 30285 4131 30343 4137
rect 23308 4060 23336 4100
rect 30285 4097 30297 4131
rect 30331 4128 30343 4131
rect 31754 4128 31760 4140
rect 30331 4100 31760 4128
rect 30331 4097 30343 4100
rect 30285 4091 30343 4097
rect 31754 4088 31760 4100
rect 31812 4088 31818 4140
rect 33410 4088 33416 4140
rect 33468 4128 33474 4140
rect 36449 4131 36507 4137
rect 36449 4128 36461 4131
rect 33468 4100 36461 4128
rect 33468 4088 33474 4100
rect 36449 4097 36461 4100
rect 36495 4097 36507 4131
rect 36449 4091 36507 4097
rect 38838 4088 38844 4140
rect 38896 4088 38902 4140
rect 39209 4131 39267 4137
rect 39209 4097 39221 4131
rect 39255 4097 39267 4131
rect 39209 4091 39267 4097
rect 13832 4032 23336 4060
rect 23400 4032 26924 4060
rect 9953 3995 10011 4001
rect 9953 3961 9965 3995
rect 9999 3992 10011 3995
rect 23400 3992 23428 4032
rect 9999 3964 23428 3992
rect 26896 3992 26924 4032
rect 26970 4020 26976 4072
rect 27028 4060 27034 4072
rect 35250 4060 35256 4072
rect 27028 4032 35256 4060
rect 27028 4020 27034 4032
rect 35250 4020 35256 4032
rect 35308 4020 35314 4072
rect 38654 4020 38660 4072
rect 38712 4060 38718 4072
rect 39224 4060 39252 4091
rect 38712 4032 39252 4060
rect 38712 4020 38718 4032
rect 39206 3992 39212 4004
rect 26896 3964 39212 3992
rect 9999 3961 10011 3964
rect 9953 3955 10011 3961
rect 39206 3952 39212 3964
rect 39264 3952 39270 4004
rect 39390 3952 39396 4004
rect 39448 3952 39454 4004
rect 5810 3884 5816 3936
rect 5868 3884 5874 3936
rect 17586 3884 17592 3936
rect 17644 3924 17650 3936
rect 20898 3924 20904 3936
rect 17644 3896 20904 3924
rect 17644 3884 17650 3896
rect 20898 3884 20904 3896
rect 20956 3884 20962 3936
rect 23385 3927 23443 3933
rect 23385 3893 23397 3927
rect 23431 3924 23443 3927
rect 26786 3924 26792 3936
rect 23431 3896 26792 3924
rect 23431 3893 23443 3896
rect 23385 3887 23443 3893
rect 26786 3884 26792 3896
rect 26844 3884 26850 3936
rect 26878 3884 26884 3936
rect 26936 3924 26942 3936
rect 28994 3924 29000 3936
rect 26936 3896 29000 3924
rect 26936 3884 26942 3896
rect 28994 3884 29000 3896
rect 29052 3884 29058 3936
rect 30469 3927 30527 3933
rect 30469 3893 30481 3927
rect 30515 3924 30527 3927
rect 30650 3924 30656 3936
rect 30515 3896 30656 3924
rect 30515 3893 30527 3896
rect 30469 3887 30527 3893
rect 30650 3884 30656 3896
rect 30708 3884 30714 3936
rect 36262 3884 36268 3936
rect 36320 3884 36326 3936
rect 39022 3884 39028 3936
rect 39080 3884 39086 3936
rect 1104 3834 39836 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 37950 3834
rect 38002 3782 38014 3834
rect 38066 3782 38078 3834
rect 38130 3782 38142 3834
rect 38194 3782 38206 3834
rect 38258 3782 39836 3834
rect 1104 3760 39836 3782
rect 5810 3680 5816 3732
rect 5868 3720 5874 3732
rect 37274 3720 37280 3732
rect 5868 3692 37280 3720
rect 5868 3680 5874 3692
rect 37274 3680 37280 3692
rect 37332 3680 37338 3732
rect 14734 3612 14740 3664
rect 14792 3612 14798 3664
rect 16482 3612 16488 3664
rect 16540 3652 16546 3664
rect 20257 3655 20315 3661
rect 20257 3652 20269 3655
rect 16540 3624 20269 3652
rect 16540 3612 16546 3624
rect 20257 3621 20269 3624
rect 20303 3621 20315 3655
rect 20257 3615 20315 3621
rect 28258 3612 28264 3664
rect 28316 3652 28322 3664
rect 28316 3624 31754 3652
rect 28316 3612 28322 3624
rect 11149 3587 11207 3593
rect 11149 3553 11161 3587
rect 11195 3584 11207 3587
rect 11195 3556 30328 3584
rect 11195 3553 11207 3556
rect 11149 3547 11207 3553
rect 7558 3476 7564 3528
rect 7616 3516 7622 3528
rect 10965 3519 11023 3525
rect 10965 3516 10977 3519
rect 7616 3488 10977 3516
rect 7616 3476 7622 3488
rect 10965 3485 10977 3488
rect 11011 3485 11023 3519
rect 10965 3479 11023 3485
rect 14829 3519 14887 3525
rect 14829 3485 14841 3519
rect 14875 3516 14887 3519
rect 14921 3519 14979 3525
rect 14921 3516 14933 3519
rect 14875 3488 14933 3516
rect 14875 3485 14887 3488
rect 14829 3479 14887 3485
rect 14921 3485 14933 3488
rect 14967 3485 14979 3519
rect 14921 3479 14979 3485
rect 17586 3476 17592 3528
rect 17644 3476 17650 3528
rect 20349 3519 20407 3525
rect 20349 3485 20361 3519
rect 20395 3512 20407 3519
rect 20441 3519 20499 3525
rect 20441 3512 20453 3519
rect 20395 3485 20453 3512
rect 20487 3485 20499 3519
rect 26878 3516 26884 3528
rect 20349 3484 20499 3485
rect 20349 3479 20407 3484
rect 20441 3479 20499 3484
rect 21928 3488 26884 3516
rect 21928 3448 21956 3488
rect 26878 3476 26884 3488
rect 26936 3476 26942 3528
rect 28994 3476 29000 3528
rect 29052 3516 29058 3528
rect 29917 3519 29975 3525
rect 29917 3516 29929 3519
rect 29052 3488 29929 3516
rect 29052 3476 29058 3488
rect 29917 3485 29929 3488
rect 29963 3485 29975 3519
rect 29917 3479 29975 3485
rect 30300 3448 30328 3556
rect 31726 3516 31754 3624
rect 39390 3612 39396 3664
rect 39448 3612 39454 3664
rect 34054 3516 34060 3528
rect 31726 3488 34060 3516
rect 34054 3476 34060 3488
rect 34112 3476 34118 3528
rect 35250 3476 35256 3528
rect 35308 3516 35314 3528
rect 38841 3519 38899 3525
rect 38841 3516 38853 3519
rect 35308 3488 38853 3516
rect 35308 3476 35314 3488
rect 38841 3485 38853 3488
rect 38887 3485 38899 3519
rect 38841 3479 38899 3485
rect 39206 3476 39212 3528
rect 39264 3476 39270 3528
rect 35986 3448 35992 3460
rect 15120 3420 19334 3448
rect 15120 3389 15148 3420
rect 15105 3383 15163 3389
rect 15105 3349 15117 3383
rect 15151 3349 15163 3383
rect 15105 3343 15163 3349
rect 17218 3340 17224 3392
rect 17276 3380 17282 3392
rect 17405 3383 17463 3389
rect 17405 3380 17417 3383
rect 17276 3352 17417 3380
rect 17276 3340 17282 3352
rect 17405 3349 17417 3352
rect 17451 3349 17463 3383
rect 19306 3380 19334 3420
rect 20548 3420 21956 3448
rect 22066 3420 30236 3448
rect 30300 3420 35992 3448
rect 20548 3380 20576 3420
rect 19306 3352 20576 3380
rect 20625 3383 20683 3389
rect 17405 3343 17463 3349
rect 20625 3349 20637 3383
rect 20671 3380 20683 3383
rect 22066 3380 22094 3420
rect 20671 3352 22094 3380
rect 20671 3349 20683 3352
rect 20625 3343 20683 3349
rect 29914 3340 29920 3392
rect 29972 3380 29978 3392
rect 30101 3383 30159 3389
rect 30101 3380 30113 3383
rect 29972 3352 30113 3380
rect 29972 3340 29978 3352
rect 30101 3349 30113 3352
rect 30147 3349 30159 3383
rect 30208 3380 30236 3420
rect 35986 3408 35992 3420
rect 36044 3408 36050 3460
rect 38838 3380 38844 3392
rect 30208 3352 38844 3380
rect 30101 3343 30159 3349
rect 38838 3340 38844 3352
rect 38896 3340 38902 3392
rect 39025 3383 39083 3389
rect 39025 3349 39037 3383
rect 39071 3380 39083 3383
rect 39942 3380 39948 3392
rect 39071 3352 39948 3380
rect 39071 3349 39083 3352
rect 39025 3343 39083 3349
rect 39942 3340 39948 3352
rect 40000 3340 40006 3392
rect 1104 3290 39836 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 39010 3290
rect 39062 3238 39074 3290
rect 39126 3238 39138 3290
rect 39190 3238 39202 3290
rect 39254 3238 39266 3290
rect 39318 3238 39836 3290
rect 1104 3216 39836 3238
rect 13722 3136 13728 3188
rect 13780 3176 13786 3188
rect 18049 3179 18107 3185
rect 18049 3176 18061 3179
rect 13780 3148 18061 3176
rect 13780 3136 13786 3148
rect 18049 3145 18061 3148
rect 18095 3145 18107 3179
rect 18049 3139 18107 3145
rect 18414 3136 18420 3188
rect 18472 3136 18478 3188
rect 20714 3136 20720 3188
rect 20772 3136 20778 3188
rect 21545 3179 21603 3185
rect 21545 3145 21557 3179
rect 21591 3176 21603 3179
rect 21591 3148 31754 3176
rect 21591 3145 21603 3148
rect 21545 3139 21603 3145
rect 658 3068 664 3120
rect 716 3108 722 3120
rect 31726 3108 31754 3148
rect 32858 3136 32864 3188
rect 32916 3176 32922 3188
rect 33321 3179 33379 3185
rect 33321 3176 33333 3179
rect 32916 3148 33333 3176
rect 32916 3136 32922 3148
rect 33321 3145 33333 3148
rect 33367 3145 33379 3179
rect 33321 3139 33379 3145
rect 33689 3179 33747 3185
rect 33689 3145 33701 3179
rect 33735 3176 33747 3179
rect 34882 3176 34888 3188
rect 33735 3148 34888 3176
rect 33735 3145 33747 3148
rect 33689 3139 33747 3145
rect 34882 3136 34888 3148
rect 34940 3136 34946 3188
rect 39390 3136 39396 3188
rect 39448 3136 39454 3188
rect 36078 3108 36084 3120
rect 716 3080 24256 3108
rect 31726 3080 36084 3108
rect 716 3068 722 3080
rect 8846 3000 8852 3052
rect 8904 3000 8910 3052
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3040 13139 3043
rect 13173 3043 13231 3049
rect 13173 3040 13185 3043
rect 13127 3012 13185 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 13173 3009 13185 3012
rect 13219 3009 13231 3043
rect 13173 3003 13231 3009
rect 15933 3043 15991 3049
rect 15933 3009 15945 3043
rect 15979 3040 15991 3043
rect 16025 3043 16083 3049
rect 16025 3040 16037 3043
rect 15979 3012 16037 3040
rect 15979 3009 15991 3012
rect 15933 3003 15991 3009
rect 16025 3009 16037 3012
rect 16071 3009 16083 3043
rect 16025 3003 16083 3009
rect 16761 3043 16819 3049
rect 16761 3009 16773 3043
rect 16807 3009 16819 3043
rect 16761 3003 16819 3009
rect 18141 3043 18199 3049
rect 18141 3009 18153 3043
rect 18187 3040 18199 3043
rect 18233 3043 18291 3049
rect 18233 3040 18245 3043
rect 18187 3012 18245 3040
rect 18187 3009 18199 3012
rect 18141 3003 18199 3009
rect 18233 3009 18245 3012
rect 18279 3009 18291 3043
rect 18233 3003 18291 3009
rect 20717 3043 20775 3049
rect 20717 3009 20729 3043
rect 20763 3040 20775 3043
rect 20809 3043 20867 3049
rect 20809 3040 20821 3043
rect 20763 3012 20821 3040
rect 20763 3009 20775 3012
rect 20717 3003 20775 3009
rect 20809 3009 20821 3012
rect 20855 3009 20867 3043
rect 20809 3003 20867 3009
rect 9398 2932 9404 2984
rect 9456 2972 9462 2984
rect 16776 2972 16804 3003
rect 21358 3000 21364 3052
rect 21416 3000 21422 3052
rect 23750 3000 23756 3052
rect 23808 3040 23814 3052
rect 24228 3049 24256 3080
rect 36078 3068 36084 3080
rect 36136 3068 36142 3120
rect 36188 3080 39252 3108
rect 23937 3043 23995 3049
rect 23937 3040 23949 3043
rect 23808 3012 23949 3040
rect 23808 3000 23814 3012
rect 23937 3009 23949 3012
rect 23983 3009 23995 3043
rect 23937 3003 23995 3009
rect 24213 3043 24271 3049
rect 24213 3009 24225 3043
rect 24259 3009 24271 3043
rect 24213 3003 24271 3009
rect 24673 3043 24731 3049
rect 24673 3009 24685 3043
rect 24719 3040 24731 3043
rect 24765 3043 24823 3049
rect 24765 3040 24777 3043
rect 24719 3012 24777 3040
rect 24719 3009 24731 3012
rect 24673 3003 24731 3009
rect 24765 3009 24777 3012
rect 24811 3009 24823 3043
rect 24765 3003 24823 3009
rect 26510 3000 26516 3052
rect 26568 3040 26574 3052
rect 26973 3043 27031 3049
rect 26973 3040 26985 3043
rect 26568 3012 26985 3040
rect 26568 3000 26574 3012
rect 26973 3009 26985 3012
rect 27019 3009 27031 3043
rect 26973 3003 27031 3009
rect 28074 3000 28080 3052
rect 28132 3000 28138 3052
rect 28537 3043 28595 3049
rect 28537 3009 28549 3043
rect 28583 3040 28595 3043
rect 28629 3043 28687 3049
rect 28629 3040 28641 3043
rect 28583 3012 28641 3040
rect 28583 3009 28595 3012
rect 28537 3003 28595 3009
rect 28629 3009 28641 3012
rect 28675 3009 28687 3043
rect 28629 3003 28687 3009
rect 30101 3043 30159 3049
rect 30101 3009 30113 3043
rect 30147 3040 30159 3043
rect 30193 3043 30251 3049
rect 30193 3040 30205 3043
rect 30147 3012 30205 3040
rect 30147 3009 30159 3012
rect 30101 3003 30159 3009
rect 30193 3009 30205 3012
rect 30239 3009 30251 3043
rect 30193 3003 30251 3009
rect 33413 3043 33471 3049
rect 33413 3009 33425 3043
rect 33459 3040 33471 3043
rect 33505 3043 33563 3049
rect 33505 3040 33517 3043
rect 33459 3012 33517 3040
rect 33459 3009 33471 3012
rect 33413 3003 33471 3009
rect 33505 3009 33517 3012
rect 33551 3009 33563 3043
rect 33505 3003 33563 3009
rect 17037 2975 17095 2981
rect 17037 2972 17049 2975
rect 9456 2944 17049 2972
rect 9456 2932 9462 2944
rect 17037 2941 17049 2944
rect 17083 2941 17095 2975
rect 36188 2972 36216 3080
rect 39224 3049 39252 3080
rect 38841 3043 38899 3049
rect 38841 3009 38853 3043
rect 38887 3009 38899 3043
rect 38841 3003 38899 3009
rect 39209 3043 39267 3049
rect 39209 3009 39221 3043
rect 39255 3009 39267 3043
rect 39209 3003 39267 3009
rect 17037 2935 17095 2941
rect 22066 2944 36216 2972
rect 9030 2864 9036 2916
rect 9088 2864 9094 2916
rect 9490 2864 9496 2916
rect 9548 2904 9554 2916
rect 15841 2907 15899 2913
rect 15841 2904 15853 2907
rect 9548 2876 15853 2904
rect 9548 2864 9554 2876
rect 15841 2873 15853 2876
rect 15887 2873 15899 2907
rect 15841 2867 15899 2873
rect 16945 2907 17003 2913
rect 16945 2873 16957 2907
rect 16991 2904 17003 2907
rect 20993 2907 21051 2913
rect 16991 2876 19334 2904
rect 16991 2873 17003 2876
rect 16945 2867 17003 2873
rect 9582 2796 9588 2848
rect 9640 2836 9646 2848
rect 12989 2839 13047 2845
rect 12989 2836 13001 2839
rect 9640 2808 13001 2836
rect 9640 2796 9646 2808
rect 12989 2805 13001 2808
rect 13035 2805 13047 2839
rect 12989 2799 13047 2805
rect 13354 2796 13360 2848
rect 13412 2796 13418 2848
rect 16206 2796 16212 2848
rect 16264 2796 16270 2848
rect 19306 2836 19334 2876
rect 20993 2873 21005 2907
rect 21039 2904 21051 2907
rect 22066 2904 22094 2944
rect 21039 2876 22094 2904
rect 24121 2907 24179 2913
rect 21039 2873 21051 2876
rect 20993 2867 21051 2873
rect 24121 2873 24133 2907
rect 24167 2904 24179 2907
rect 38856 2904 38884 3003
rect 24167 2876 38884 2904
rect 24167 2873 24179 2876
rect 24121 2867 24179 2873
rect 24026 2836 24032 2848
rect 19306 2808 24032 2836
rect 24026 2796 24032 2808
rect 24084 2796 24090 2848
rect 24394 2796 24400 2848
rect 24452 2796 24458 2848
rect 24578 2796 24584 2848
rect 24636 2796 24642 2848
rect 24946 2796 24952 2848
rect 25004 2796 25010 2848
rect 27157 2839 27215 2845
rect 27157 2805 27169 2839
rect 27203 2836 27215 2839
rect 27338 2836 27344 2848
rect 27203 2808 27344 2836
rect 27203 2805 27215 2808
rect 27157 2799 27215 2805
rect 27338 2796 27344 2808
rect 27396 2796 27402 2848
rect 28258 2796 28264 2848
rect 28316 2796 28322 2848
rect 28442 2796 28448 2848
rect 28500 2796 28506 2848
rect 28810 2796 28816 2848
rect 28868 2796 28874 2848
rect 30006 2796 30012 2848
rect 30064 2796 30070 2848
rect 30377 2839 30435 2845
rect 30377 2805 30389 2839
rect 30423 2836 30435 2839
rect 30926 2836 30932 2848
rect 30423 2808 30932 2836
rect 30423 2805 30435 2808
rect 30377 2799 30435 2805
rect 30926 2796 30932 2808
rect 30984 2796 30990 2848
rect 39022 2796 39028 2848
rect 39080 2796 39086 2848
rect 1104 2746 39836 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 37950 2746
rect 38002 2694 38014 2746
rect 38066 2694 38078 2746
rect 38130 2694 38142 2746
rect 38194 2694 38206 2746
rect 38258 2694 39836 2746
rect 1104 2672 39836 2694
rect 38102 2632 38108 2644
rect 26528 2604 38108 2632
rect 16206 2524 16212 2576
rect 16264 2564 16270 2576
rect 26528 2564 26556 2604
rect 38102 2592 38108 2604
rect 38160 2592 38166 2644
rect 16264 2536 26556 2564
rect 16264 2524 16270 2536
rect 38562 2524 38568 2576
rect 38620 2564 38626 2576
rect 38620 2536 38884 2564
rect 38620 2524 38626 2536
rect 13354 2456 13360 2508
rect 13412 2496 13418 2508
rect 26510 2496 26516 2508
rect 13412 2468 26516 2496
rect 13412 2456 13418 2468
rect 26510 2456 26516 2468
rect 26568 2456 26574 2508
rect 26694 2456 26700 2508
rect 26752 2496 26758 2508
rect 31570 2496 31576 2508
rect 26752 2468 31576 2496
rect 26752 2456 26758 2468
rect 31570 2456 31576 2468
rect 31628 2456 31634 2508
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 26418 2428 26424 2440
rect 9088 2400 26424 2428
rect 9088 2388 9094 2400
rect 26418 2388 26424 2400
rect 26476 2388 26482 2440
rect 26786 2388 26792 2440
rect 26844 2428 26850 2440
rect 32582 2428 32588 2440
rect 26844 2400 32588 2428
rect 26844 2388 26850 2400
rect 32582 2388 32588 2400
rect 32640 2388 32646 2440
rect 32674 2388 32680 2440
rect 32732 2428 32738 2440
rect 37725 2431 37783 2437
rect 37725 2428 37737 2431
rect 32732 2400 37737 2428
rect 32732 2388 32738 2400
rect 37725 2397 37737 2400
rect 37771 2397 37783 2431
rect 37725 2391 37783 2397
rect 38102 2388 38108 2440
rect 38160 2388 38166 2440
rect 38470 2388 38476 2440
rect 38528 2388 38534 2440
rect 38856 2437 38884 2536
rect 39390 2524 39396 2576
rect 39448 2524 39454 2576
rect 38841 2431 38899 2437
rect 38841 2397 38853 2431
rect 38887 2397 38899 2431
rect 38841 2391 38899 2397
rect 39209 2431 39267 2437
rect 39209 2397 39221 2431
rect 39255 2397 39267 2431
rect 39209 2391 39267 2397
rect 3418 2320 3424 2372
rect 3476 2360 3482 2372
rect 21358 2360 21364 2372
rect 3476 2332 21364 2360
rect 3476 2320 3482 2332
rect 21358 2320 21364 2332
rect 21416 2320 21422 2372
rect 24026 2320 24032 2372
rect 24084 2360 24090 2372
rect 24084 2332 27016 2360
rect 24084 2320 24090 2332
rect 16574 2252 16580 2304
rect 16632 2292 16638 2304
rect 26878 2292 26884 2304
rect 16632 2264 26884 2292
rect 16632 2252 16638 2264
rect 26878 2252 26884 2264
rect 26936 2252 26942 2304
rect 26988 2292 27016 2332
rect 28810 2320 28816 2372
rect 28868 2360 28874 2372
rect 39224 2360 39252 2391
rect 28868 2332 33088 2360
rect 28868 2320 28874 2332
rect 32674 2292 32680 2304
rect 26988 2264 32680 2292
rect 32674 2252 32680 2264
rect 32732 2252 32738 2304
rect 33060 2292 33088 2332
rect 33244 2332 39252 2360
rect 33244 2292 33272 2332
rect 33060 2264 33272 2292
rect 37918 2252 37924 2304
rect 37976 2252 37982 2304
rect 38286 2252 38292 2304
rect 38344 2252 38350 2304
rect 38654 2252 38660 2304
rect 38712 2252 38718 2304
rect 39025 2295 39083 2301
rect 39025 2261 39037 2295
rect 39071 2292 39083 2295
rect 39942 2292 39948 2304
rect 39071 2264 39948 2292
rect 39071 2261 39083 2264
rect 39025 2255 39083 2261
rect 39942 2252 39948 2264
rect 40000 2252 40006 2304
rect 1104 2202 39836 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 39010 2202
rect 39062 2150 39074 2202
rect 39126 2150 39138 2202
rect 39190 2150 39202 2202
rect 39254 2150 39266 2202
rect 39318 2150 39836 2202
rect 1104 2128 39836 2150
rect 12710 2048 12716 2100
rect 12768 2088 12774 2100
rect 30006 2088 30012 2100
rect 12768 2060 30012 2088
rect 12768 2048 12774 2060
rect 30006 2048 30012 2060
rect 30064 2048 30070 2100
rect 26878 1912 26884 1964
rect 26936 1952 26942 1964
rect 33410 1952 33416 1964
rect 26936 1924 33416 1952
rect 26936 1912 26942 1924
rect 33410 1912 33416 1924
rect 33468 1912 33474 1964
rect 22370 1368 22376 1420
rect 22428 1408 22434 1420
rect 28994 1408 29000 1420
rect 22428 1380 29000 1408
rect 22428 1368 22434 1380
rect 28994 1368 29000 1380
rect 29052 1368 29058 1420
rect 4982 144 4988 196
rect 5040 184 5046 196
rect 22462 184 22468 196
rect 5040 156 22468 184
rect 5040 144 5046 156
rect 22462 144 22468 156
rect 22520 144 22526 196
rect 18598 76 18604 128
rect 18656 116 18662 128
rect 37090 116 37096 128
rect 18656 88 37096 116
rect 18656 76 18662 88
rect 37090 76 37096 88
rect 37148 76 37154 128
rect 1210 8 1216 60
rect 1268 48 1274 60
rect 25866 48 25872 60
rect 1268 20 25872 48
rect 1268 8 1274 20
rect 25866 8 25872 20
rect 25924 8 25930 60
<< via1 >>
rect 7288 11160 7340 11212
rect 27804 11160 27856 11212
rect 6368 11092 6420 11144
rect 18420 11092 18472 11144
rect 16396 10956 16448 11008
rect 22284 10956 22336 11008
rect 16948 10004 17000 10056
rect 23940 10004 23992 10056
rect 13820 9868 13872 9920
rect 18696 9868 18748 9920
rect 19340 9596 19392 9648
rect 24768 9596 24820 9648
rect 1124 9528 1176 9580
rect 23848 9528 23900 9580
rect 17960 9460 18012 9512
rect 24216 9460 24268 9512
rect 1308 9392 1360 9444
rect 26516 9392 26568 9444
rect 13360 9324 13412 9376
rect 17868 9324 17920 9376
rect 22744 9324 22796 9376
rect 36544 9324 36596 9376
rect 15752 9256 15804 9308
rect 26424 9256 26476 9308
rect 8392 9188 8444 9240
rect 17224 9188 17276 9240
rect 24032 9188 24084 9240
rect 38936 9188 38988 9240
rect 204 9120 256 9172
rect 23940 9120 23992 9172
rect 10784 8984 10836 9036
rect 19248 9052 19300 9104
rect 19616 9052 19668 9104
rect 20628 9052 20680 9104
rect 21732 9052 21784 9104
rect 28080 9052 28132 9104
rect 15568 8984 15620 9036
rect 22928 8984 22980 9036
rect 33600 8984 33652 9036
rect 34244 8984 34296 9036
rect 8668 8916 8720 8968
rect 12808 8916 12860 8968
rect 19708 8916 19760 8968
rect 19800 8916 19852 8968
rect 32588 8916 32640 8968
rect 15844 8848 15896 8900
rect 17040 8848 17092 8900
rect 17868 8848 17920 8900
rect 30748 8848 30800 8900
rect 37280 8916 37332 8968
rect 11336 8780 11388 8832
rect 16028 8780 16080 8832
rect 16120 8780 16172 8832
rect 23480 8780 23532 8832
rect 24584 8780 24636 8832
rect 27252 8780 27304 8832
rect 29920 8780 29972 8832
rect 36176 8848 36228 8900
rect 33048 8780 33100 8832
rect 33508 8780 33560 8832
rect 33784 8780 33836 8832
rect 38016 8780 38068 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 39010 8678 39062 8730
rect 39074 8678 39126 8730
rect 39138 8678 39190 8730
rect 39202 8678 39254 8730
rect 39266 8678 39318 8730
rect 3792 8576 3844 8628
rect 4344 8576 4396 8628
rect 4620 8619 4672 8628
rect 4620 8585 4629 8619
rect 4629 8585 4663 8619
rect 4663 8585 4672 8619
rect 4620 8576 4672 8585
rect 5172 8576 5224 8628
rect 5448 8576 5500 8628
rect 5724 8576 5776 8628
rect 6276 8576 6328 8628
rect 6828 8576 6880 8628
rect 7380 8576 7432 8628
rect 7656 8576 7708 8628
rect 7932 8576 7984 8628
rect 8484 8576 8536 8628
rect 8852 8576 8904 8628
rect 9588 8576 9640 8628
rect 9864 8576 9916 8628
rect 10140 8619 10192 8628
rect 10140 8585 10149 8619
rect 10149 8585 10183 8619
rect 10183 8585 10192 8619
rect 10140 8576 10192 8585
rect 10692 8576 10744 8628
rect 10968 8576 11020 8628
rect 11520 8576 11572 8628
rect 12072 8576 12124 8628
rect 12348 8576 12400 8628
rect 12900 8576 12952 8628
rect 13176 8576 13228 8628
rect 13636 8576 13688 8628
rect 14004 8576 14056 8628
rect 14556 8576 14608 8628
rect 14924 8576 14976 8628
rect 15384 8576 15436 8628
rect 15660 8576 15712 8628
rect 16212 8576 16264 8628
rect 16488 8576 16540 8628
rect 16764 8576 16816 8628
rect 17316 8576 17368 8628
rect 17868 8619 17920 8628
rect 17868 8585 17877 8619
rect 17877 8585 17911 8619
rect 17911 8585 17920 8619
rect 17868 8576 17920 8585
rect 2872 8440 2924 8492
rect 3424 8440 3476 8492
rect 4068 8483 4120 8492
rect 4068 8449 4077 8483
rect 4077 8449 4111 8483
rect 4111 8449 4120 8483
rect 4068 8440 4120 8449
rect 4436 8483 4488 8492
rect 4436 8449 4445 8483
rect 4445 8449 4479 8483
rect 4479 8449 4488 8483
rect 4436 8440 4488 8449
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 5448 8483 5500 8492
rect 5448 8449 5457 8483
rect 5457 8449 5491 8483
rect 5491 8449 5500 8483
rect 5448 8440 5500 8449
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 7564 8440 7616 8492
rect 7840 8440 7892 8492
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 8668 8440 8720 8492
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 7748 8372 7800 8424
rect 8484 8372 8536 8424
rect 9956 8483 10008 8492
rect 9956 8449 9965 8483
rect 9965 8449 9999 8483
rect 9999 8449 10008 8483
rect 9956 8440 10008 8449
rect 10876 8440 10928 8492
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 11152 8440 11204 8492
rect 11336 8483 11388 8492
rect 11336 8449 11345 8483
rect 11345 8449 11379 8483
rect 11379 8449 11388 8483
rect 11336 8440 11388 8449
rect 3608 8304 3660 8356
rect 12808 8483 12860 8492
rect 12808 8449 12817 8483
rect 12817 8449 12851 8483
rect 12851 8449 12860 8483
rect 12808 8440 12860 8449
rect 13176 8483 13228 8492
rect 13176 8449 13185 8483
rect 13185 8449 13219 8483
rect 13219 8449 13228 8483
rect 13176 8440 13228 8449
rect 14740 8508 14792 8560
rect 16580 8508 16632 8560
rect 18236 8576 18288 8628
rect 32220 8576 32272 8628
rect 32496 8576 32548 8628
rect 32864 8576 32916 8628
rect 33508 8619 33560 8628
rect 33508 8585 33517 8619
rect 33517 8585 33551 8619
rect 33551 8585 33560 8619
rect 33508 8576 33560 8585
rect 13820 8372 13872 8424
rect 15292 8440 15344 8492
rect 15568 8440 15620 8492
rect 15660 8440 15712 8492
rect 15752 8483 15804 8492
rect 15752 8449 15761 8483
rect 15761 8449 15795 8483
rect 15795 8449 15804 8483
rect 15752 8440 15804 8449
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 16396 8372 16448 8424
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 17684 8440 17736 8492
rect 23388 8508 23440 8560
rect 20720 8440 20772 8492
rect 30380 8440 30432 8492
rect 32588 8483 32640 8492
rect 32588 8449 32597 8483
rect 32597 8449 32631 8483
rect 32631 8449 32640 8483
rect 32588 8440 32640 8449
rect 32680 8440 32732 8492
rect 33416 8508 33468 8560
rect 34244 8619 34296 8628
rect 34244 8585 34253 8619
rect 34253 8585 34287 8619
rect 34287 8585 34296 8619
rect 34244 8576 34296 8585
rect 34704 8576 34756 8628
rect 35808 8576 35860 8628
rect 36912 8576 36964 8628
rect 34152 8508 34204 8560
rect 18236 8372 18288 8424
rect 23112 8372 23164 8424
rect 24952 8372 25004 8424
rect 34060 8483 34112 8492
rect 34060 8449 34069 8483
rect 34069 8449 34103 8483
rect 34103 8449 34112 8483
rect 34060 8440 34112 8449
rect 35624 8508 35676 8560
rect 34888 8440 34940 8492
rect 35256 8440 35308 8492
rect 35716 8483 35768 8492
rect 35716 8449 35725 8483
rect 35725 8449 35759 8483
rect 35759 8449 35768 8483
rect 35716 8440 35768 8449
rect 35808 8483 35860 8492
rect 35808 8449 35817 8483
rect 35817 8449 35851 8483
rect 35851 8449 35860 8483
rect 35808 8440 35860 8449
rect 36176 8483 36228 8492
rect 36176 8449 36185 8483
rect 36185 8449 36219 8483
rect 36219 8449 36228 8483
rect 36176 8440 36228 8449
rect 36544 8483 36596 8492
rect 36544 8449 36553 8483
rect 36553 8449 36587 8483
rect 36587 8449 36596 8483
rect 36544 8440 36596 8449
rect 7196 8236 7248 8288
rect 13728 8236 13780 8288
rect 14372 8236 14424 8288
rect 14464 8236 14516 8288
rect 16948 8236 17000 8288
rect 23756 8304 23808 8356
rect 30932 8304 30984 8356
rect 33968 8304 34020 8356
rect 31024 8236 31076 8288
rect 35348 8304 35400 8356
rect 36360 8372 36412 8424
rect 37464 8508 37516 8560
rect 37280 8483 37332 8492
rect 37280 8449 37289 8483
rect 37289 8449 37323 8483
rect 37323 8449 37332 8483
rect 37280 8440 37332 8449
rect 37372 8440 37424 8492
rect 38016 8483 38068 8492
rect 38016 8449 38025 8483
rect 38025 8449 38059 8483
rect 38059 8449 38068 8483
rect 38016 8440 38068 8449
rect 38568 8440 38620 8492
rect 38936 8440 38988 8492
rect 37188 8304 37240 8356
rect 39028 8347 39080 8356
rect 39028 8313 39037 8347
rect 39037 8313 39071 8347
rect 39071 8313 39080 8347
rect 39028 8304 39080 8313
rect 39396 8347 39448 8356
rect 39396 8313 39405 8347
rect 39405 8313 39439 8347
rect 39439 8313 39448 8347
rect 39396 8304 39448 8313
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 37950 8134 38002 8186
rect 38014 8134 38066 8186
rect 38078 8134 38130 8186
rect 38142 8134 38194 8186
rect 38206 8134 38258 8186
rect 3516 8075 3568 8084
rect 3516 8041 3525 8075
rect 3525 8041 3559 8075
rect 3559 8041 3568 8075
rect 3516 8032 3568 8041
rect 3976 8032 4028 8084
rect 4896 8032 4948 8084
rect 6000 8032 6052 8084
rect 6552 8032 6604 8084
rect 7104 8032 7156 8084
rect 8300 8032 8352 8084
rect 8760 8032 8812 8084
rect 9404 8032 9456 8084
rect 10416 8032 10468 8084
rect 11244 8032 11296 8084
rect 11796 8075 11848 8084
rect 11796 8041 11805 8075
rect 11805 8041 11839 8075
rect 11839 8041 11848 8075
rect 11796 8032 11848 8041
rect 12624 8032 12676 8084
rect 13452 8032 13504 8084
rect 13820 8032 13872 8084
rect 14280 8032 14332 8084
rect 14556 8032 14608 8084
rect 14832 8032 14884 8084
rect 15936 8032 15988 8084
rect 19708 8075 19760 8084
rect 19708 8041 19717 8075
rect 19717 8041 19751 8075
rect 19751 8041 19760 8075
rect 19708 8032 19760 8041
rect 20628 8032 20680 8084
rect 21824 8075 21876 8084
rect 21824 8041 21833 8075
rect 21833 8041 21867 8075
rect 21867 8041 21876 8075
rect 21824 8032 21876 8041
rect 23112 8075 23164 8084
rect 23112 8041 23121 8075
rect 23121 8041 23155 8075
rect 23155 8041 23164 8075
rect 23112 8032 23164 8041
rect 23480 8075 23532 8084
rect 23480 8041 23489 8075
rect 23489 8041 23523 8075
rect 23523 8041 23532 8075
rect 23480 8032 23532 8041
rect 27620 8032 27672 8084
rect 28908 8032 28960 8084
rect 31024 8075 31076 8084
rect 31024 8041 31033 8075
rect 31033 8041 31067 8075
rect 31067 8041 31076 8075
rect 31024 8032 31076 8041
rect 34428 8032 34480 8084
rect 35532 8032 35584 8084
rect 36084 8032 36136 8084
rect 36636 8032 36688 8084
rect 37740 8032 37792 8084
rect 38660 8075 38712 8084
rect 38660 8041 38669 8075
rect 38669 8041 38703 8075
rect 38703 8041 38712 8075
rect 38660 8032 38712 8041
rect 8484 7964 8536 8016
rect 3976 7896 4028 7948
rect 2780 7828 2832 7880
rect 4160 7871 4212 7880
rect 4160 7837 4169 7871
rect 4169 7837 4203 7871
rect 4203 7837 4212 7871
rect 4160 7828 4212 7837
rect 4988 7871 5040 7880
rect 4988 7837 4997 7871
rect 4997 7837 5031 7871
rect 5031 7837 5040 7871
rect 4988 7828 5040 7837
rect 6644 7871 6696 7880
rect 6644 7837 6653 7871
rect 6653 7837 6687 7871
rect 6687 7837 6696 7871
rect 6644 7828 6696 7837
rect 7472 7871 7524 7880
rect 7472 7837 7481 7871
rect 7481 7837 7515 7871
rect 7515 7837 7524 7871
rect 7472 7828 7524 7837
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 11888 7896 11940 7948
rect 14924 7964 14976 8016
rect 15476 7964 15528 8016
rect 31576 7964 31628 8016
rect 7656 7760 7708 7812
rect 8300 7760 8352 7812
rect 11520 7828 11572 7880
rect 11612 7871 11664 7880
rect 11612 7837 11621 7871
rect 11621 7837 11655 7871
rect 11655 7837 11664 7871
rect 11612 7828 11664 7837
rect 14556 7896 14608 7948
rect 13452 7871 13504 7880
rect 13452 7837 13461 7871
rect 13461 7837 13495 7871
rect 13495 7837 13504 7871
rect 13452 7828 13504 7837
rect 13820 7871 13872 7880
rect 13820 7837 13829 7871
rect 13829 7837 13863 7871
rect 13863 7837 13872 7871
rect 13820 7828 13872 7837
rect 14464 7828 14516 7880
rect 19800 7896 19852 7948
rect 15844 7871 15896 7880
rect 15844 7837 15853 7871
rect 15853 7837 15887 7871
rect 15887 7837 15896 7871
rect 15844 7828 15896 7837
rect 7104 7692 7156 7744
rect 10784 7692 10836 7744
rect 12716 7692 12768 7744
rect 15476 7735 15528 7744
rect 15476 7701 15485 7735
rect 15485 7701 15519 7735
rect 15519 7701 15528 7735
rect 15476 7692 15528 7701
rect 16120 7692 16172 7744
rect 16488 7692 16540 7744
rect 19156 7828 19208 7880
rect 22652 7896 22704 7948
rect 31852 7896 31904 7948
rect 23204 7828 23256 7880
rect 23572 7828 23624 7880
rect 27620 7828 27672 7880
rect 27712 7871 27764 7880
rect 27712 7837 27721 7871
rect 27721 7837 27755 7871
rect 27755 7837 27764 7871
rect 27712 7828 27764 7837
rect 31116 7828 31168 7880
rect 31392 7828 31444 7880
rect 20352 7760 20404 7812
rect 20444 7760 20496 7812
rect 35900 7828 35952 7880
rect 36176 7871 36228 7880
rect 36176 7837 36185 7871
rect 36185 7837 36219 7871
rect 36219 7837 36228 7871
rect 36176 7828 36228 7837
rect 36452 7828 36504 7880
rect 38292 7828 38344 7880
rect 38844 7871 38896 7880
rect 38844 7837 38853 7871
rect 38853 7837 38887 7871
rect 38887 7837 38896 7871
rect 38844 7828 38896 7837
rect 19156 7692 19208 7744
rect 19432 7735 19484 7744
rect 19432 7701 19441 7735
rect 19441 7701 19475 7735
rect 19475 7701 19484 7735
rect 19432 7692 19484 7701
rect 21364 7735 21416 7744
rect 21364 7701 21373 7735
rect 21373 7701 21407 7735
rect 21407 7701 21416 7735
rect 21364 7692 21416 7701
rect 27712 7692 27764 7744
rect 27896 7735 27948 7744
rect 27896 7701 27905 7735
rect 27905 7701 27939 7735
rect 27939 7701 27948 7735
rect 27896 7692 27948 7701
rect 35348 7735 35400 7744
rect 35348 7701 35357 7735
rect 35357 7701 35391 7735
rect 35391 7701 35400 7735
rect 35348 7692 35400 7701
rect 36360 7760 36412 7812
rect 36268 7692 36320 7744
rect 38936 7692 38988 7744
rect 39396 7735 39448 7744
rect 39396 7701 39405 7735
rect 39405 7701 39439 7735
rect 39439 7701 39448 7735
rect 39396 7692 39448 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 39010 7590 39062 7642
rect 39074 7590 39126 7642
rect 39138 7590 39190 7642
rect 39202 7590 39254 7642
rect 39266 7590 39318 7642
rect 2780 7531 2832 7540
rect 2780 7497 2789 7531
rect 2789 7497 2823 7531
rect 2823 7497 2832 7531
rect 2780 7488 2832 7497
rect 9496 7488 9548 7540
rect 14372 7488 14424 7540
rect 14740 7488 14792 7540
rect 20444 7488 20496 7540
rect 20720 7488 20772 7540
rect 21364 7488 21416 7540
rect 22652 7488 22704 7540
rect 23756 7531 23808 7540
rect 23756 7497 23765 7531
rect 23765 7497 23799 7531
rect 23799 7497 23808 7531
rect 23756 7488 23808 7497
rect 27896 7488 27948 7540
rect 34152 7488 34204 7540
rect 7196 7352 7248 7404
rect 7288 7352 7340 7404
rect 13084 7420 13136 7472
rect 14924 7420 14976 7472
rect 9772 7395 9824 7404
rect 9772 7361 9781 7395
rect 9781 7361 9815 7395
rect 9815 7361 9824 7395
rect 9772 7352 9824 7361
rect 17500 7352 17552 7404
rect 18052 7420 18104 7472
rect 19156 7420 19208 7472
rect 24768 7420 24820 7472
rect 30656 7420 30708 7472
rect 36452 7488 36504 7540
rect 3608 7284 3660 7336
rect 8300 7284 8352 7336
rect 8576 7284 8628 7336
rect 12256 7284 12308 7336
rect 13452 7284 13504 7336
rect 9956 7216 10008 7268
rect 11888 7216 11940 7268
rect 16028 7216 16080 7268
rect 17868 7352 17920 7404
rect 19340 7352 19392 7404
rect 21732 7352 21784 7404
rect 28356 7352 28408 7404
rect 30840 7352 30892 7404
rect 37740 7395 37792 7404
rect 37740 7361 37749 7395
rect 37749 7361 37783 7395
rect 37783 7361 37792 7395
rect 37740 7352 37792 7361
rect 38752 7488 38804 7540
rect 39488 7488 39540 7540
rect 38568 7420 38620 7472
rect 24492 7284 24544 7336
rect 26884 7284 26936 7336
rect 38384 7352 38436 7404
rect 38476 7395 38528 7404
rect 38476 7361 38485 7395
rect 38485 7361 38519 7395
rect 38519 7361 38528 7395
rect 38476 7352 38528 7361
rect 33692 7216 33744 7268
rect 38200 7284 38252 7336
rect 12164 7148 12216 7200
rect 17960 7148 18012 7200
rect 19800 7148 19852 7200
rect 39488 7216 39540 7268
rect 39396 7191 39448 7200
rect 39396 7157 39405 7191
rect 39405 7157 39439 7191
rect 39439 7157 39448 7191
rect 39396 7148 39448 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 37950 7046 38002 7098
rect 38014 7046 38066 7098
rect 38078 7046 38130 7098
rect 38142 7046 38194 7098
rect 38206 7046 38258 7098
rect 12164 6944 12216 6996
rect 17408 6944 17460 6996
rect 19432 6944 19484 6996
rect 26884 6944 26936 6996
rect 32864 6944 32916 6996
rect 38844 6944 38896 6996
rect 9588 6876 9640 6928
rect 4620 6808 4672 6860
rect 6276 6740 6328 6792
rect 11060 6740 11112 6792
rect 20536 6808 20588 6860
rect 34152 6876 34204 6928
rect 19616 6740 19668 6792
rect 22468 6783 22520 6792
rect 22468 6749 22477 6783
rect 22477 6749 22511 6783
rect 22511 6749 22520 6783
rect 22468 6740 22520 6749
rect 29092 6740 29144 6792
rect 3792 6672 3844 6724
rect 2872 6647 2924 6656
rect 2872 6613 2881 6647
rect 2881 6613 2915 6647
rect 2915 6613 2924 6647
rect 2872 6604 2924 6613
rect 7564 6604 7616 6656
rect 20812 6672 20864 6724
rect 30564 6740 30616 6792
rect 31668 6740 31720 6792
rect 38476 6783 38528 6792
rect 38476 6749 38485 6783
rect 38485 6749 38519 6783
rect 38519 6749 38528 6783
rect 38476 6740 38528 6749
rect 38936 6740 38988 6792
rect 11060 6604 11112 6656
rect 12348 6604 12400 6656
rect 16396 6604 16448 6656
rect 24768 6604 24820 6656
rect 32680 6672 32732 6724
rect 30472 6604 30524 6656
rect 38660 6647 38712 6656
rect 38660 6613 38669 6647
rect 38669 6613 38703 6647
rect 38703 6613 38712 6647
rect 38660 6604 38712 6613
rect 39672 6672 39724 6724
rect 39580 6604 39632 6656
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 39010 6502 39062 6554
rect 39074 6502 39126 6554
rect 39138 6502 39190 6554
rect 39202 6502 39254 6554
rect 39266 6502 39318 6554
rect 3424 6400 3476 6452
rect 4068 6400 4120 6452
rect 4436 6443 4488 6452
rect 4436 6409 4445 6443
rect 4445 6409 4479 6443
rect 4479 6409 4488 6443
rect 4436 6400 4488 6409
rect 7472 6400 7524 6452
rect 7748 6400 7800 6452
rect 3516 6332 3568 6384
rect 3792 6375 3844 6384
rect 3792 6341 3801 6375
rect 3801 6341 3835 6375
rect 3835 6341 3844 6375
rect 3792 6332 3844 6341
rect 8208 6332 8260 6384
rect 11520 6400 11572 6452
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 7380 6264 7432 6316
rect 7656 6128 7708 6180
rect 10692 6264 10744 6316
rect 21640 6400 21692 6452
rect 26424 6443 26476 6452
rect 26424 6409 26433 6443
rect 26433 6409 26467 6443
rect 26467 6409 26476 6443
rect 26424 6400 26476 6409
rect 25872 6332 25924 6384
rect 11888 6264 11940 6316
rect 18880 6264 18932 6316
rect 19156 6307 19208 6316
rect 19156 6273 19165 6307
rect 19165 6273 19199 6307
rect 19199 6273 19208 6307
rect 19156 6264 19208 6273
rect 23848 6264 23900 6316
rect 29184 6264 29236 6316
rect 15844 6196 15896 6248
rect 39396 6443 39448 6452
rect 39396 6409 39405 6443
rect 39405 6409 39439 6443
rect 39439 6409 39448 6443
rect 39396 6400 39448 6409
rect 31024 6332 31076 6384
rect 35900 6332 35952 6384
rect 30288 6264 30340 6316
rect 34336 6264 34388 6316
rect 39212 6307 39264 6316
rect 39212 6273 39221 6307
rect 39221 6273 39255 6307
rect 39255 6273 39264 6307
rect 39212 6264 39264 6273
rect 29368 6196 29420 6248
rect 37740 6196 37792 6248
rect 16120 6128 16172 6180
rect 11612 6060 11664 6112
rect 17132 6060 17184 6112
rect 38752 6128 38804 6180
rect 38476 6060 38528 6112
rect 39028 6103 39080 6112
rect 39028 6069 39037 6103
rect 39037 6069 39071 6103
rect 39071 6069 39080 6103
rect 39028 6060 39080 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 37950 5958 38002 6010
rect 38014 5958 38066 6010
rect 38078 5958 38130 6010
rect 38142 5958 38194 6010
rect 38206 5958 38258 6010
rect 4160 5856 4212 5908
rect 4988 5856 5040 5908
rect 5448 5856 5500 5908
rect 5816 5856 5868 5908
rect 6920 5856 6972 5908
rect 11244 5856 11296 5908
rect 30380 5856 30432 5908
rect 35808 5856 35860 5908
rect 35900 5856 35952 5908
rect 38292 5856 38344 5908
rect 38752 5856 38804 5908
rect 39764 5856 39816 5908
rect 5540 5720 5592 5772
rect 11888 5788 11940 5840
rect 19524 5788 19576 5840
rect 27620 5788 27672 5840
rect 39212 5788 39264 5840
rect 39396 5831 39448 5840
rect 39396 5797 39405 5831
rect 39405 5797 39439 5831
rect 39439 5797 39448 5831
rect 39396 5788 39448 5797
rect 9588 5584 9640 5636
rect 16212 5720 16264 5772
rect 20444 5720 20496 5772
rect 15384 5652 15436 5704
rect 16488 5584 16540 5636
rect 25872 5695 25924 5704
rect 25872 5661 25881 5695
rect 25881 5661 25915 5695
rect 25915 5661 25924 5695
rect 25872 5652 25924 5661
rect 30012 5652 30064 5704
rect 14924 5516 14976 5568
rect 26148 5516 26200 5568
rect 29000 5516 29052 5568
rect 37096 5652 37148 5704
rect 38752 5652 38804 5704
rect 37832 5584 37884 5636
rect 35624 5516 35676 5568
rect 36084 5516 36136 5568
rect 39948 5516 40000 5568
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 39010 5414 39062 5466
rect 39074 5414 39126 5466
rect 39138 5414 39190 5466
rect 39202 5414 39254 5466
rect 39266 5414 39318 5466
rect 5080 5312 5132 5364
rect 6644 5312 6696 5364
rect 12256 5312 12308 5364
rect 10968 5244 11020 5296
rect 27620 5312 27672 5364
rect 39396 5355 39448 5364
rect 39396 5321 39405 5355
rect 39405 5321 39439 5355
rect 39439 5321 39448 5355
rect 39396 5312 39448 5321
rect 5540 5219 5592 5228
rect 5540 5185 5549 5219
rect 5549 5185 5583 5219
rect 5583 5185 5592 5219
rect 5540 5176 5592 5185
rect 13544 5176 13596 5228
rect 19064 5244 19116 5296
rect 16672 5219 16724 5228
rect 16672 5185 16681 5219
rect 16681 5185 16715 5219
rect 16715 5185 16724 5219
rect 16672 5176 16724 5185
rect 17316 5219 17368 5228
rect 17316 5185 17325 5219
rect 17325 5185 17359 5219
rect 17359 5185 17368 5219
rect 17316 5176 17368 5185
rect 19800 5176 19852 5228
rect 24584 5176 24636 5228
rect 27528 5176 27580 5228
rect 37280 5176 37332 5228
rect 15660 5108 15712 5160
rect 16764 5108 16816 5160
rect 29368 5108 29420 5160
rect 35992 5108 36044 5160
rect 17132 5083 17184 5092
rect 17132 5049 17141 5083
rect 17141 5049 17175 5083
rect 17175 5049 17184 5083
rect 17132 5040 17184 5049
rect 22744 5040 22796 5092
rect 26148 5040 26200 5092
rect 38660 5040 38712 5092
rect 21824 5015 21876 5024
rect 21824 4981 21833 5015
rect 21833 4981 21867 5015
rect 21867 4981 21876 5015
rect 21824 4972 21876 4981
rect 22928 4972 22980 5024
rect 39028 5015 39080 5024
rect 39028 4981 39037 5015
rect 39037 4981 39071 5015
rect 39071 4981 39080 5015
rect 39028 4972 39080 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 37950 4870 38002 4922
rect 38014 4870 38066 4922
rect 38078 4870 38130 4922
rect 38142 4870 38194 4922
rect 38206 4870 38258 4922
rect 10876 4768 10928 4820
rect 16304 4811 16356 4820
rect 16304 4777 16313 4811
rect 16313 4777 16347 4811
rect 16347 4777 16356 4811
rect 16304 4768 16356 4777
rect 16764 4768 16816 4820
rect 17868 4768 17920 4820
rect 11152 4700 11204 4752
rect 18420 4700 18472 4752
rect 32864 4768 32916 4820
rect 33784 4811 33836 4820
rect 33784 4777 33793 4811
rect 33793 4777 33827 4811
rect 33827 4777 33836 4811
rect 33784 4768 33836 4777
rect 24032 4700 24084 4752
rect 5540 4632 5592 4684
rect 11428 4539 11480 4548
rect 11428 4505 11437 4539
rect 11437 4505 11471 4539
rect 11471 4505 11480 4539
rect 11428 4496 11480 4505
rect 15936 4632 15988 4684
rect 21824 4632 21876 4684
rect 14832 4607 14884 4616
rect 14832 4573 14841 4607
rect 14841 4573 14875 4607
rect 14875 4573 14884 4607
rect 14832 4564 14884 4573
rect 24308 4632 24360 4684
rect 39396 4743 39448 4752
rect 39396 4709 39405 4743
rect 39405 4709 39439 4743
rect 39439 4709 39448 4743
rect 39396 4700 39448 4709
rect 36176 4632 36228 4684
rect 23848 4564 23900 4616
rect 28080 4564 28132 4616
rect 30104 4564 30156 4616
rect 19708 4496 19760 4548
rect 19064 4471 19116 4480
rect 19064 4437 19073 4471
rect 19073 4437 19107 4471
rect 19107 4437 19116 4471
rect 19064 4428 19116 4437
rect 31024 4496 31076 4548
rect 35900 4564 35952 4616
rect 38844 4607 38896 4616
rect 38844 4573 38853 4607
rect 38853 4573 38887 4607
rect 38887 4573 38896 4607
rect 38844 4564 38896 4573
rect 38936 4564 38988 4616
rect 33968 4496 34020 4548
rect 30748 4428 30800 4480
rect 37188 4428 37240 4480
rect 39948 4428 40000 4480
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 39010 4326 39062 4378
rect 39074 4326 39126 4378
rect 39138 4326 39190 4378
rect 39202 4326 39254 4378
rect 39266 4326 39318 4378
rect 5724 4199 5776 4208
rect 5724 4165 5733 4199
rect 5733 4165 5767 4199
rect 5767 4165 5776 4199
rect 5724 4156 5776 4165
rect 8300 4156 8352 4208
rect 8208 4088 8260 4140
rect 19064 4224 19116 4276
rect 38844 4224 38896 4276
rect 14832 4156 14884 4208
rect 25596 4156 25648 4208
rect 20720 4088 20772 4140
rect 38936 4156 38988 4208
rect 31760 4088 31812 4140
rect 33416 4088 33468 4140
rect 38844 4131 38896 4140
rect 38844 4097 38853 4131
rect 38853 4097 38887 4131
rect 38887 4097 38896 4131
rect 38844 4088 38896 4097
rect 26976 4020 27028 4072
rect 35256 4020 35308 4072
rect 38660 4020 38712 4072
rect 39212 3952 39264 4004
rect 39396 3995 39448 4004
rect 39396 3961 39405 3995
rect 39405 3961 39439 3995
rect 39439 3961 39448 3995
rect 39396 3952 39448 3961
rect 5816 3927 5868 3936
rect 5816 3893 5825 3927
rect 5825 3893 5859 3927
rect 5859 3893 5868 3927
rect 5816 3884 5868 3893
rect 17592 3884 17644 3936
rect 20904 3884 20956 3936
rect 26792 3884 26844 3936
rect 26884 3884 26936 3936
rect 29000 3884 29052 3936
rect 30656 3884 30708 3936
rect 36268 3927 36320 3936
rect 36268 3893 36277 3927
rect 36277 3893 36311 3927
rect 36311 3893 36320 3927
rect 36268 3884 36320 3893
rect 39028 3927 39080 3936
rect 39028 3893 39037 3927
rect 39037 3893 39071 3927
rect 39071 3893 39080 3927
rect 39028 3884 39080 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 37950 3782 38002 3834
rect 38014 3782 38066 3834
rect 38078 3782 38130 3834
rect 38142 3782 38194 3834
rect 38206 3782 38258 3834
rect 5816 3680 5868 3732
rect 37280 3680 37332 3732
rect 14740 3655 14792 3664
rect 14740 3621 14749 3655
rect 14749 3621 14783 3655
rect 14783 3621 14792 3655
rect 14740 3612 14792 3621
rect 16488 3612 16540 3664
rect 28264 3612 28316 3664
rect 7564 3476 7616 3528
rect 17592 3519 17644 3528
rect 17592 3485 17601 3519
rect 17601 3485 17635 3519
rect 17635 3485 17644 3519
rect 17592 3476 17644 3485
rect 26884 3476 26936 3528
rect 29000 3476 29052 3528
rect 39396 3655 39448 3664
rect 39396 3621 39405 3655
rect 39405 3621 39439 3655
rect 39439 3621 39448 3655
rect 39396 3612 39448 3621
rect 34060 3476 34112 3528
rect 35256 3476 35308 3528
rect 39212 3519 39264 3528
rect 39212 3485 39221 3519
rect 39221 3485 39255 3519
rect 39255 3485 39264 3519
rect 39212 3476 39264 3485
rect 17224 3340 17276 3392
rect 29920 3340 29972 3392
rect 35992 3408 36044 3460
rect 38844 3340 38896 3392
rect 39948 3340 40000 3392
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 39010 3238 39062 3290
rect 39074 3238 39126 3290
rect 39138 3238 39190 3290
rect 39202 3238 39254 3290
rect 39266 3238 39318 3290
rect 13728 3136 13780 3188
rect 18420 3179 18472 3188
rect 18420 3145 18429 3179
rect 18429 3145 18463 3179
rect 18463 3145 18472 3179
rect 18420 3136 18472 3145
rect 20720 3179 20772 3188
rect 20720 3145 20729 3179
rect 20729 3145 20763 3179
rect 20763 3145 20772 3179
rect 20720 3136 20772 3145
rect 664 3068 716 3120
rect 32864 3136 32916 3188
rect 34888 3136 34940 3188
rect 39396 3179 39448 3188
rect 39396 3145 39405 3179
rect 39405 3145 39439 3179
rect 39439 3145 39448 3179
rect 39396 3136 39448 3145
rect 8852 3043 8904 3052
rect 8852 3009 8861 3043
rect 8861 3009 8895 3043
rect 8895 3009 8904 3043
rect 8852 3000 8904 3009
rect 9404 2932 9456 2984
rect 21364 3043 21416 3052
rect 21364 3009 21373 3043
rect 21373 3009 21407 3043
rect 21407 3009 21416 3043
rect 21364 3000 21416 3009
rect 23756 3043 23808 3052
rect 23756 3009 23765 3043
rect 23765 3009 23799 3043
rect 23799 3009 23808 3043
rect 36084 3068 36136 3120
rect 23756 3000 23808 3009
rect 26516 3000 26568 3052
rect 28080 3043 28132 3052
rect 28080 3009 28089 3043
rect 28089 3009 28123 3043
rect 28123 3009 28132 3043
rect 28080 3000 28132 3009
rect 9036 2907 9088 2916
rect 9036 2873 9045 2907
rect 9045 2873 9079 2907
rect 9079 2873 9088 2907
rect 9036 2864 9088 2873
rect 9496 2864 9548 2916
rect 9588 2796 9640 2848
rect 13360 2839 13412 2848
rect 13360 2805 13369 2839
rect 13369 2805 13403 2839
rect 13403 2805 13412 2839
rect 13360 2796 13412 2805
rect 16212 2839 16264 2848
rect 16212 2805 16221 2839
rect 16221 2805 16255 2839
rect 16255 2805 16264 2839
rect 16212 2796 16264 2805
rect 24032 2796 24084 2848
rect 24400 2839 24452 2848
rect 24400 2805 24409 2839
rect 24409 2805 24443 2839
rect 24443 2805 24452 2839
rect 24400 2796 24452 2805
rect 24584 2839 24636 2848
rect 24584 2805 24593 2839
rect 24593 2805 24627 2839
rect 24627 2805 24636 2839
rect 24584 2796 24636 2805
rect 24952 2839 25004 2848
rect 24952 2805 24961 2839
rect 24961 2805 24995 2839
rect 24995 2805 25004 2839
rect 24952 2796 25004 2805
rect 27344 2796 27396 2848
rect 28264 2839 28316 2848
rect 28264 2805 28273 2839
rect 28273 2805 28307 2839
rect 28307 2805 28316 2839
rect 28264 2796 28316 2805
rect 28448 2839 28500 2848
rect 28448 2805 28457 2839
rect 28457 2805 28491 2839
rect 28491 2805 28500 2839
rect 28448 2796 28500 2805
rect 28816 2839 28868 2848
rect 28816 2805 28825 2839
rect 28825 2805 28859 2839
rect 28859 2805 28868 2839
rect 28816 2796 28868 2805
rect 30012 2839 30064 2848
rect 30012 2805 30021 2839
rect 30021 2805 30055 2839
rect 30055 2805 30064 2839
rect 30012 2796 30064 2805
rect 30932 2796 30984 2848
rect 39028 2839 39080 2848
rect 39028 2805 39037 2839
rect 39037 2805 39071 2839
rect 39071 2805 39080 2839
rect 39028 2796 39080 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 37950 2694 38002 2746
rect 38014 2694 38066 2746
rect 38078 2694 38130 2746
rect 38142 2694 38194 2746
rect 38206 2694 38258 2746
rect 16212 2524 16264 2576
rect 38108 2592 38160 2644
rect 38568 2524 38620 2576
rect 13360 2456 13412 2508
rect 26516 2456 26568 2508
rect 26700 2456 26752 2508
rect 31576 2456 31628 2508
rect 9036 2388 9088 2440
rect 26424 2388 26476 2440
rect 26792 2388 26844 2440
rect 32588 2388 32640 2440
rect 32680 2388 32732 2440
rect 38108 2431 38160 2440
rect 38108 2397 38117 2431
rect 38117 2397 38151 2431
rect 38151 2397 38160 2431
rect 38108 2388 38160 2397
rect 38476 2431 38528 2440
rect 38476 2397 38485 2431
rect 38485 2397 38519 2431
rect 38519 2397 38528 2431
rect 38476 2388 38528 2397
rect 39396 2567 39448 2576
rect 39396 2533 39405 2567
rect 39405 2533 39439 2567
rect 39439 2533 39448 2567
rect 39396 2524 39448 2533
rect 3424 2320 3476 2372
rect 21364 2320 21416 2372
rect 24032 2320 24084 2372
rect 16580 2252 16632 2304
rect 26884 2252 26936 2304
rect 28816 2320 28868 2372
rect 32680 2252 32732 2304
rect 37924 2295 37976 2304
rect 37924 2261 37933 2295
rect 37933 2261 37967 2295
rect 37967 2261 37976 2295
rect 37924 2252 37976 2261
rect 38292 2295 38344 2304
rect 38292 2261 38301 2295
rect 38301 2261 38335 2295
rect 38335 2261 38344 2295
rect 38292 2252 38344 2261
rect 38660 2295 38712 2304
rect 38660 2261 38669 2295
rect 38669 2261 38703 2295
rect 38703 2261 38712 2295
rect 38660 2252 38712 2261
rect 39948 2252 40000 2304
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 39010 2150 39062 2202
rect 39074 2150 39126 2202
rect 39138 2150 39190 2202
rect 39202 2150 39254 2202
rect 39266 2150 39318 2202
rect 12716 2048 12768 2100
rect 30012 2048 30064 2100
rect 26884 1912 26936 1964
rect 33416 1912 33468 1964
rect 22376 1368 22428 1420
rect 29000 1368 29052 1420
rect 4988 144 5040 196
rect 22468 144 22520 196
rect 18604 76 18656 128
rect 37096 76 37148 128
rect 1216 8 1268 60
rect 25872 8 25924 60
<< metal2 >>
rect 3238 11194 3294 11250
rect 3514 11194 3570 11250
rect 3790 11194 3846 11250
rect 4066 11194 4122 11250
rect 4342 11194 4398 11250
rect 4618 11194 4674 11250
rect 4894 11194 4950 11250
rect 5170 11194 5226 11250
rect 5446 11194 5502 11250
rect 5722 11194 5778 11250
rect 5998 11194 6054 11250
rect 6274 11194 6330 11250
rect 6550 11194 6606 11250
rect 6826 11194 6882 11250
rect 7102 11194 7158 11250
rect 7288 11212 7340 11218
rect 1124 9580 1176 9586
rect 1124 9522 1176 9528
rect 204 9172 256 9178
rect 204 9114 256 9120
rect 216 7993 244 9114
rect 1136 8265 1164 9522
rect 1308 9444 1360 9450
rect 1308 9386 1360 9392
rect 1122 8256 1178 8265
rect 1122 8191 1178 8200
rect 202 7984 258 7993
rect 202 7919 258 7928
rect 662 7712 718 7721
rect 662 7647 718 7656
rect 676 3126 704 7647
rect 1320 7177 1348 9386
rect 3252 9194 3280 11194
rect 3528 9330 3556 11194
rect 3528 9302 3648 9330
rect 3252 9166 3556 9194
rect 2778 8800 2834 8809
rect 2778 8735 2834 8744
rect 2792 8401 2820 8735
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 2778 8392 2834 8401
rect 2778 8327 2834 8336
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2792 7546 2820 7822
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 1306 7168 1362 7177
rect 1306 7103 1362 7112
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1766 6760 1822 6769
rect 1766 6695 1822 6704
rect 1780 6089 1808 6695
rect 2884 6662 2912 8434
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 2872 6656 2924 6662
rect 2778 6624 2834 6633
rect 2872 6598 2924 6604
rect 2778 6559 2834 6568
rect 1766 6080 1822 6089
rect 1766 6015 1822 6024
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2792 5681 2820 6559
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 3436 6458 3464 8434
rect 3528 8090 3556 9166
rect 3620 8362 3648 9302
rect 3804 8634 3832 11194
rect 4080 8650 4108 11194
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3988 8622 4108 8650
rect 4356 8634 4384 11194
rect 4632 8634 4660 11194
rect 4344 8628 4396 8634
rect 3608 8356 3660 8362
rect 3608 8298 3660 8304
rect 3988 8090 4016 8622
rect 4344 8570 4396 8576
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 3974 7984 4030 7993
rect 3974 7919 3976 7928
rect 4028 7919 4030 7928
rect 3976 7890 4028 7896
rect 3608 7336 3660 7342
rect 3514 7304 3570 7313
rect 3608 7278 3660 7284
rect 3514 7239 3570 7248
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3528 6390 3556 7239
rect 3516 6384 3568 6390
rect 3516 6326 3568 6332
rect 3422 5808 3478 5817
rect 3422 5743 3478 5752
rect 2778 5672 2834 5681
rect 2778 5607 2834 5616
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 2686 5264 2742 5273
rect 2686 5199 2742 5208
rect 2700 5001 2728 5199
rect 2686 4992 2742 5001
rect 1950 4924 2258 4933
rect 2686 4927 2742 4936
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 2870 4040 2926 4049
rect 2870 3975 2926 3984
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2884 3369 2912 3975
rect 2870 3360 2926 3369
rect 2870 3295 2926 3304
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 664 3120 716 3126
rect 664 3062 716 3068
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 3436 2378 3464 5743
rect 3424 2372 3476 2378
rect 3424 2314 3476 2320
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 1136 66 1256 82
rect 1136 60 1268 66
rect 1136 56 1216 60
rect 1122 54 1216 56
rect 1122 0 1178 54
rect 3068 56 3188 82
rect 1216 2 1268 8
rect 3054 54 3188 56
rect 3054 0 3110 54
rect 3160 42 3188 54
rect 3620 42 3648 7278
rect 3792 6724 3844 6730
rect 3792 6666 3844 6672
rect 3804 6390 3832 6666
rect 4080 6458 4108 8434
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 3792 6384 3844 6390
rect 3792 6326 3844 6332
rect 4172 5914 4200 7822
rect 4448 6458 4476 8434
rect 4908 8090 4936 11194
rect 5184 8634 5212 11194
rect 5460 8634 5488 11194
rect 5736 8634 5764 11194
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4436 6452 4488 6458
rect 4436 6394 4488 6400
rect 4632 6322 4660 6802
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 5000 5914 5028 7822
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 5092 5370 5120 8434
rect 5460 5914 5488 8434
rect 5538 6216 5594 6225
rect 5538 6151 5594 6160
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5552 5778 5580 6151
rect 5828 5914 5856 8434
rect 6012 8090 6040 11194
rect 6288 8634 6316 11194
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 6380 6914 6408 11086
rect 6564 8090 6592 11194
rect 6840 8634 6868 11194
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6288 6886 6408 6914
rect 6288 6798 6316 6886
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 6656 5370 6684 7822
rect 6932 5914 6960 8434
rect 7116 8090 7144 11194
rect 7378 11194 7434 11250
rect 7654 11194 7710 11250
rect 7930 11194 7986 11250
rect 8206 11194 8262 11250
rect 8482 11194 8538 11250
rect 8758 11194 8814 11250
rect 9034 11194 9090 11250
rect 9310 11194 9366 11250
rect 9586 11194 9642 11250
rect 9862 11194 9918 11250
rect 10138 11194 10194 11250
rect 10414 11194 10470 11250
rect 10690 11194 10746 11250
rect 10966 11194 11022 11250
rect 11242 11194 11298 11250
rect 11518 11194 11574 11250
rect 11794 11194 11850 11250
rect 12070 11194 12126 11250
rect 12346 11194 12402 11250
rect 12622 11194 12678 11250
rect 12898 11194 12954 11250
rect 13174 11194 13230 11250
rect 13450 11194 13506 11250
rect 13726 11194 13782 11250
rect 14002 11194 14058 11250
rect 14278 11194 14334 11250
rect 14554 11194 14610 11250
rect 14830 11194 14886 11250
rect 15106 11194 15162 11250
rect 15382 11194 15438 11250
rect 15658 11194 15714 11250
rect 15934 11194 15990 11250
rect 16210 11194 16266 11250
rect 16486 11194 16542 11250
rect 16762 11194 16818 11250
rect 17038 11194 17094 11250
rect 17314 11194 17370 11250
rect 17590 11194 17646 11250
rect 17866 11194 17922 11250
rect 18142 11194 18198 11250
rect 18418 11194 18474 11250
rect 18694 11194 18750 11250
rect 18970 11194 19026 11250
rect 19246 11194 19302 11250
rect 19522 11194 19578 11250
rect 19798 11194 19854 11250
rect 20074 11194 20130 11250
rect 20350 11194 20406 11250
rect 20626 11194 20682 11250
rect 20902 11194 20958 11250
rect 21178 11194 21234 11250
rect 21454 11194 21510 11250
rect 21730 11194 21786 11250
rect 22006 11194 22062 11250
rect 22282 11194 22338 11250
rect 22558 11194 22614 11250
rect 22834 11194 22890 11250
rect 23110 11194 23166 11250
rect 23386 11194 23442 11250
rect 23662 11194 23718 11250
rect 23938 11194 23994 11250
rect 24214 11194 24270 11250
rect 24490 11194 24546 11250
rect 24766 11194 24822 11250
rect 25042 11194 25098 11250
rect 25318 11194 25374 11250
rect 25594 11194 25650 11250
rect 25870 11194 25926 11250
rect 26146 11194 26202 11250
rect 26422 11194 26478 11250
rect 26698 11194 26754 11250
rect 26974 11194 27030 11250
rect 27250 11194 27306 11250
rect 27526 11194 27582 11250
rect 27802 11212 27858 11250
rect 27802 11194 27804 11212
rect 7288 11154 7340 11160
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5552 4690 5580 5170
rect 5722 5128 5778 5137
rect 5722 5063 5778 5072
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5736 4214 5764 5063
rect 5724 4208 5776 4214
rect 5724 4150 5776 4156
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5828 3738 5856 3878
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 4988 196 5040 202
rect 4988 138 5040 144
rect 5000 56 5028 138
rect 6932 56 7052 82
rect 3160 14 3648 42
rect 4986 0 5042 56
rect 6918 54 7052 56
rect 6918 0 6974 54
rect 7024 42 7052 54
rect 7116 42 7144 7686
rect 7208 7410 7236 8230
rect 7300 7410 7328 11154
rect 7392 8634 7420 11194
rect 7470 11112 7526 11121
rect 7470 11047 7526 11056
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7484 8514 7512 11047
rect 7668 8634 7696 11194
rect 7944 8634 7972 11194
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7392 8486 7512 8514
rect 7564 8492 7616 8498
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7392 6322 7420 8486
rect 7564 8434 7616 8440
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7484 6458 7512 7822
rect 7576 6662 7604 8434
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7668 6186 7696 7754
rect 7760 6458 7788 8366
rect 7852 6914 7880 8434
rect 8220 8378 8248 11194
rect 8392 9240 8444 9246
rect 8392 9182 8444 9188
rect 8404 8498 8432 9182
rect 8496 8634 8524 11194
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8680 8498 8708 8910
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8484 8424 8536 8430
rect 8220 8350 8340 8378
rect 8484 8366 8536 8372
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 8312 8090 8340 8350
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8496 8022 8524 8366
rect 8772 8090 8800 11194
rect 9048 8820 9076 11194
rect 8864 8792 9076 8820
rect 9324 8820 9352 11194
rect 9324 8792 9444 8820
rect 8864 8634 8892 8792
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 9416 8090 9444 8792
rect 9600 8634 9628 11194
rect 9770 10296 9826 10305
rect 9770 10231 9826 10240
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 8484 8016 8536 8022
rect 8484 7958 8536 7964
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8312 7342 8340 7754
rect 8588 7342 8616 7822
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 9508 7546 9536 8434
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9784 7410 9812 10231
rect 9876 8634 9904 11194
rect 10152 8634 10180 11194
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 9968 7274 9996 8434
rect 10428 8090 10456 11194
rect 10704 8634 10732 11194
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 10796 7970 10824 8978
rect 10980 8634 11008 11194
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 10704 7942 10824 7970
rect 10230 7712 10286 7721
rect 10230 7647 10286 7656
rect 10244 7313 10272 7647
rect 10230 7304 10286 7313
rect 9956 7268 10008 7274
rect 10230 7239 10286 7248
rect 9956 7210 10008 7216
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 9588 6928 9640 6934
rect 7852 6886 8248 6914
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 8220 6390 8248 6886
rect 9588 6870 9640 6876
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 7656 6180 7708 6186
rect 7656 6122 7708 6128
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 9600 5642 9628 6870
rect 10704 6322 10732 7942
rect 10782 7848 10838 7857
rect 10782 7783 10838 7792
rect 10796 7750 10824 7783
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 7562 4992 7618 5001
rect 7562 4927 7618 4936
rect 7576 3534 7604 4927
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 10888 4826 10916 8434
rect 10980 5302 11008 8434
rect 11164 6914 11192 8434
rect 11256 8090 11284 11194
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11348 8498 11376 8774
rect 11532 8634 11560 11194
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11808 8090 11836 11194
rect 12084 8634 12112 11194
rect 12360 8634 12388 11194
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12636 8090 12664 11194
rect 12714 10976 12770 10985
rect 12714 10911 12770 10920
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11164 6886 11284 6914
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11150 6760 11206 6769
rect 11072 6662 11100 6734
rect 11150 6695 11206 6704
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 10968 5296 11020 5302
rect 10968 5238 11020 5244
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 11164 4758 11192 6695
rect 11256 5914 11284 6886
rect 11532 6458 11560 7822
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11624 6118 11652 7822
rect 11900 7274 11928 7890
rect 12728 7750 12756 10911
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12820 8498 12848 8910
rect 12912 8634 12940 11194
rect 13082 10840 13138 10849
rect 13082 10775 13138 10784
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 13096 7478 13124 10775
rect 13188 8634 13216 11194
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13188 7857 13216 8434
rect 13174 7848 13230 7857
rect 13174 7783 13230 7792
rect 13084 7472 13136 7478
rect 12346 7440 12402 7449
rect 13084 7414 13136 7420
rect 12346 7375 12402 7384
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 11888 7268 11940 7274
rect 11888 7210 11940 7216
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12176 7002 12204 7142
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11900 5846 11928 6258
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 12268 5370 12296 7278
rect 12360 6662 12388 7375
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 13372 6225 13400 9318
rect 13464 8090 13492 11194
rect 13542 8936 13598 8945
rect 13542 8871 13598 8880
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13464 7342 13492 7822
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13358 6216 13414 6225
rect 13358 6151 13414 6160
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 13556 5234 13584 8871
rect 13636 8628 13688 8634
rect 13740 8616 13768 11194
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13688 8588 13768 8616
rect 13636 8570 13688 8576
rect 13832 8514 13860 9862
rect 14016 8634 14044 11194
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 13740 8486 13860 8514
rect 13740 8294 13768 8486
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13832 8090 13860 8366
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 14292 8090 14320 11194
rect 14568 8634 14596 11194
rect 14646 10704 14702 10713
rect 14646 10639 14702 10648
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 14464 8288 14516 8294
rect 14660 8242 14688 10639
rect 14740 8560 14792 8566
rect 14740 8502 14792 8508
rect 14464 8230 14516 8236
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13726 7304 13782 7313
rect 13726 7239 13782 7248
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 11152 4752 11204 4758
rect 8206 4720 8262 4729
rect 11152 4694 11204 4700
rect 8206 4655 8262 4664
rect 8220 4146 8248 4655
rect 11426 4584 11482 4593
rect 11426 4519 11428 4528
rect 11480 4519 11482 4528
rect 11428 4490 11480 4496
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 7564 3528 7616 3534
rect 8312 3505 8340 4150
rect 7564 3470 7616 3476
rect 8298 3496 8354 3505
rect 8298 3431 8354 3440
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 10782 3224 10838 3233
rect 13740 3194 13768 7239
rect 13832 6769 13860 7822
rect 14384 7546 14412 8230
rect 14476 7886 14504 8230
rect 14568 8214 14688 8242
rect 14568 8090 14596 8214
rect 14646 8120 14702 8129
rect 14556 8084 14608 8090
rect 14646 8055 14702 8064
rect 14556 8026 14608 8032
rect 14556 7948 14608 7954
rect 14556 7890 14608 7896
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14568 7449 14596 7890
rect 14660 7721 14688 8055
rect 14646 7712 14702 7721
rect 14646 7647 14702 7656
rect 14752 7546 14780 8502
rect 14844 8090 14872 11194
rect 15120 8922 15148 11194
rect 14936 8894 15148 8922
rect 14936 8634 14964 8894
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 15396 8634 15424 11194
rect 15474 9072 15530 9081
rect 15474 9007 15530 9016
rect 15568 9036 15620 9042
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14924 8016 14976 8022
rect 14924 7958 14976 7964
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14936 7478 14964 7958
rect 15304 7732 15332 8434
rect 15488 8022 15516 9007
rect 15568 8978 15620 8984
rect 15580 8498 15608 8978
rect 15672 8634 15700 11194
rect 15752 9308 15804 9314
rect 15752 9250 15804 9256
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15764 8498 15792 9250
rect 15844 8900 15896 8906
rect 15844 8842 15896 8848
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15476 8016 15528 8022
rect 15476 7958 15528 7964
rect 15476 7744 15528 7750
rect 15304 7704 15424 7732
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 14924 7472 14976 7478
rect 14278 7440 14334 7449
rect 14278 7375 14334 7384
rect 14554 7440 14610 7449
rect 14924 7414 14976 7420
rect 14554 7375 14610 7384
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 14292 7018 14320 7375
rect 14370 7032 14426 7041
rect 14292 6990 14370 7018
rect 14370 6967 14426 6976
rect 13818 6760 13874 6769
rect 13818 6695 13874 6704
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 15396 5710 15424 7704
rect 15476 7686 15528 7692
rect 15488 5817 15516 7686
rect 15474 5808 15530 5817
rect 15474 5743 15530 5752
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 14738 5264 14794 5273
rect 14738 5199 14794 5208
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 14752 3670 14780 5199
rect 14832 4616 14884 4622
rect 14832 4558 14884 4564
rect 14844 4214 14872 4558
rect 14832 4208 14884 4214
rect 14936 4185 14964 5510
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 15672 5166 15700 8434
rect 15856 7970 15884 8842
rect 15948 8090 15976 11194
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 15856 7942 15976 7970
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15856 6254 15884 7822
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 15948 4690 15976 7942
rect 16040 7274 16068 8774
rect 16132 8498 16160 8774
rect 16224 8634 16252 11194
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16302 9752 16358 9761
rect 16302 9687 16358 9696
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16316 8514 16344 9687
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16224 8486 16344 8514
rect 16408 8514 16436 10950
rect 16500 8634 16528 11194
rect 16578 9072 16634 9081
rect 16578 9007 16634 9016
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16592 8566 16620 9007
rect 16776 8634 16804 11194
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16580 8560 16632 8566
rect 16408 8486 16528 8514
rect 16580 8502 16632 8508
rect 16120 7744 16172 7750
rect 16120 7686 16172 7692
rect 16028 7268 16080 7274
rect 16028 7210 16080 7216
rect 16132 6186 16160 7686
rect 16120 6180 16172 6186
rect 16120 6122 16172 6128
rect 16224 5778 16252 8486
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16302 6896 16358 6905
rect 16302 6831 16358 6840
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 16316 4826 16344 6831
rect 16408 6662 16436 8366
rect 16500 7750 16528 8486
rect 16960 8294 16988 9998
rect 17052 8906 17080 11194
rect 17224 9240 17276 9246
rect 17224 9182 17276 9188
rect 17040 8900 17092 8906
rect 17040 8842 17092 8848
rect 16948 8288 17000 8294
rect 16948 8230 17000 8236
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16486 7304 16542 7313
rect 16486 7239 16542 7248
rect 16396 6656 16448 6662
rect 16396 6598 16448 6604
rect 16500 5642 16528 7239
rect 17132 6112 17184 6118
rect 17132 6054 17184 6060
rect 16670 5672 16726 5681
rect 16488 5636 16540 5642
rect 16670 5607 16726 5616
rect 16488 5578 16540 5584
rect 16684 5234 16712 5607
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16776 4826 16804 5102
rect 17144 5098 17172 6054
rect 17132 5092 17184 5098
rect 17132 5034 17184 5040
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 14832 4150 14884 4156
rect 14922 4176 14978 4185
rect 14922 4111 14978 4120
rect 14740 3664 14792 3670
rect 16488 3664 16540 3670
rect 14740 3606 14792 3612
rect 16486 3632 16488 3641
rect 16540 3632 16542 3641
rect 16486 3567 16542 3576
rect 14646 3496 14702 3505
rect 14646 3431 14702 3440
rect 10782 3159 10838 3168
rect 13728 3188 13780 3194
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 8864 2417 8892 2994
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 9048 2446 9076 2858
rect 9036 2440 9088 2446
rect 8850 2408 8906 2417
rect 9036 2382 9088 2388
rect 8850 2343 8906 2352
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 9416 2009 9444 2926
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 9402 2000 9458 2009
rect 9402 1935 9458 1944
rect 9508 1737 9536 2858
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9494 1728 9550 1737
rect 9494 1663 9550 1672
rect 9600 1465 9628 2790
rect 9586 1456 9642 1465
rect 9586 1391 9642 1400
rect 7024 14 7144 42
rect 8850 96 8906 105
rect 10796 56 10824 3159
rect 13728 3130 13780 3136
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 13372 2514 13400 2790
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 12716 2100 12768 2106
rect 12716 2042 12768 2048
rect 12728 56 12756 2042
rect 14660 56 14688 3431
rect 17236 3398 17264 9182
rect 17328 8634 17356 11194
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17408 8492 17460 8498
rect 17604 8480 17632 11194
rect 17880 9382 17908 11194
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17868 8900 17920 8906
rect 17868 8842 17920 8848
rect 17880 8634 17908 8842
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17684 8492 17736 8498
rect 17604 8452 17684 8480
rect 17408 8434 17460 8440
rect 17684 8434 17736 8440
rect 17420 7002 17448 8434
rect 17500 7404 17552 7410
rect 17868 7404 17920 7410
rect 17552 7364 17868 7392
rect 17500 7346 17552 7352
rect 17868 7346 17920 7352
rect 17972 7206 18000 9454
rect 18050 9344 18106 9353
rect 18050 9279 18106 9288
rect 18064 7478 18092 9279
rect 18052 7472 18104 7478
rect 18052 7414 18104 7420
rect 17960 7200 18012 7206
rect 18156 7177 18184 11194
rect 18432 11150 18460 11194
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18708 9926 18736 11194
rect 18878 10160 18934 10169
rect 18878 10095 18934 10104
rect 18696 9920 18748 9926
rect 18696 9862 18748 9868
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18248 8430 18276 8570
rect 18236 8424 18288 8430
rect 18236 8366 18288 8372
rect 17960 7142 18012 7148
rect 18142 7168 18198 7177
rect 18142 7103 18198 7112
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 18892 6322 18920 10095
rect 18984 9761 19012 11194
rect 19062 10024 19118 10033
rect 19062 9959 19118 9968
rect 18970 9752 19026 9761
rect 18970 9687 19026 9696
rect 18880 6316 18932 6322
rect 18880 6258 18932 6264
rect 19076 5302 19104 9959
rect 19154 9888 19210 9897
rect 19154 9823 19210 9832
rect 19168 7886 19196 9823
rect 19260 9110 19288 11194
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19248 9104 19300 9110
rect 19248 9046 19300 9052
rect 19156 7880 19208 7886
rect 19156 7822 19208 7828
rect 19156 7744 19208 7750
rect 19156 7686 19208 7692
rect 19168 7478 19196 7686
rect 19156 7472 19208 7478
rect 19156 7414 19208 7420
rect 19352 7410 19380 9590
rect 19432 7744 19484 7750
rect 19432 7686 19484 7692
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 19444 7002 19472 7686
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19154 6352 19210 6361
rect 19154 6287 19156 6296
rect 19208 6287 19210 6296
rect 19156 6258 19208 6264
rect 19536 5846 19564 11194
rect 19812 10169 19840 11194
rect 19798 10160 19854 10169
rect 19798 10095 19854 10104
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 19628 6798 19656 9046
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19800 8968 19852 8974
rect 19800 8910 19852 8916
rect 19720 8090 19748 8910
rect 19812 8129 19840 8910
rect 20088 8673 20116 11194
rect 20364 9058 20392 11194
rect 20640 9110 20668 11194
rect 20628 9104 20680 9110
rect 20364 9030 20576 9058
rect 20916 9058 20944 11194
rect 20628 9046 20680 9052
rect 20074 8664 20130 8673
rect 20074 8599 20130 8608
rect 20350 8256 20406 8265
rect 19950 8188 20258 8197
rect 20350 8191 20406 8200
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19798 8120 19854 8129
rect 19950 8123 20258 8132
rect 19708 8084 19760 8090
rect 19798 8055 19854 8064
rect 19708 8026 19760 8032
rect 19800 7948 19852 7954
rect 19800 7890 19852 7896
rect 19812 7206 19840 7890
rect 20364 7818 20392 8191
rect 20352 7812 20404 7818
rect 20352 7754 20404 7760
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 20456 7546 20484 7754
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 19800 7200 19852 7206
rect 19800 7142 19852 7148
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 20548 6866 20576 9030
rect 20824 9030 20944 9058
rect 20626 8528 20682 8537
rect 20626 8463 20682 8472
rect 20720 8492 20772 8498
rect 20640 8090 20668 8463
rect 20720 8434 20772 8440
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20732 7546 20760 8434
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20536 6860 20588 6866
rect 20536 6802 20588 6808
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 20824 6730 20852 9030
rect 21192 8922 21220 11194
rect 21468 8945 21496 11194
rect 21744 9194 21772 11194
rect 21652 9166 21772 9194
rect 20916 8894 21220 8922
rect 21454 8936 21510 8945
rect 20812 6724 20864 6730
rect 20812 6666 20864 6672
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 19524 5840 19576 5846
rect 19524 5782 19576 5788
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 19706 5536 19762 5545
rect 19706 5471 19762 5480
rect 19064 5296 19116 5302
rect 17314 5264 17370 5273
rect 19064 5238 19116 5244
rect 17314 5199 17316 5208
rect 17368 5199 17370 5208
rect 17316 5170 17368 5176
rect 17866 5128 17922 5137
rect 17866 5063 17922 5072
rect 17880 4826 17908 5063
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 18420 4752 18472 4758
rect 18420 4694 18472 4700
rect 17592 3936 17644 3942
rect 17592 3878 17644 3884
rect 17604 3534 17632 3878
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 14830 3224 14886 3233
rect 15010 3227 15318 3236
rect 18432 3194 18460 4694
rect 19720 4554 19748 5471
rect 19800 5228 19852 5234
rect 19800 5170 19852 5176
rect 19708 4548 19760 4554
rect 19708 4490 19760 4496
rect 19064 4480 19116 4486
rect 19064 4422 19116 4428
rect 19076 4282 19104 4422
rect 19064 4276 19116 4282
rect 19064 4218 19116 4224
rect 19812 4185 19840 5170
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 19798 4176 19854 4185
rect 19798 4111 19854 4120
rect 19950 3836 20258 3845
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 14830 3159 14886 3168
rect 18420 3188 18472 3194
rect 14844 2825 14872 3159
rect 18420 3130 18472 3136
rect 16212 2848 16264 2854
rect 14830 2816 14886 2825
rect 16212 2790 16264 2796
rect 14830 2751 14886 2760
rect 16224 2582 16252 2790
rect 19950 2748 20258 2757
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 16580 2304 16632 2310
rect 16580 2246 16632 2252
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 16592 56 16620 2246
rect 18604 128 18656 134
rect 18524 76 18604 82
rect 18524 70 18656 76
rect 18524 56 18644 70
rect 20456 56 20484 5714
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 20732 4049 20760 4082
rect 20718 4040 20774 4049
rect 20718 3975 20774 3984
rect 20916 3942 20944 8894
rect 21454 8871 21510 8880
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 21364 7744 21416 7750
rect 21364 7686 21416 7692
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 21376 7546 21404 7686
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 21652 6458 21680 9166
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 21744 7410 21772 9046
rect 21822 8392 21878 8401
rect 21822 8327 21878 8336
rect 21836 8090 21864 8327
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21732 7404 21784 7410
rect 21732 7346 21784 7352
rect 22020 7041 22048 11194
rect 22296 11014 22324 11194
rect 22572 11121 22600 11194
rect 22558 11112 22614 11121
rect 22558 11047 22614 11056
rect 22284 11008 22336 11014
rect 22284 10950 22336 10956
rect 22744 9376 22796 9382
rect 22744 9318 22796 9324
rect 22652 7948 22704 7954
rect 22652 7890 22704 7896
rect 22664 7546 22692 7890
rect 22652 7540 22704 7546
rect 22652 7482 22704 7488
rect 22006 7032 22062 7041
rect 22006 6967 22062 6976
rect 22468 6792 22520 6798
rect 22468 6734 22520 6740
rect 21640 6452 21692 6458
rect 21640 6394 21692 6400
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 21824 5024 21876 5030
rect 21824 4966 21876 4972
rect 21836 4690 21864 4966
rect 21824 4684 21876 4690
rect 21824 4626 21876 4632
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 20718 3224 20774 3233
rect 21010 3227 21318 3236
rect 20718 3159 20720 3168
rect 20772 3159 20774 3168
rect 20720 3130 20772 3136
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 21376 2378 21404 2994
rect 21364 2372 21416 2378
rect 21364 2314 21416 2320
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 22376 1420 22428 1426
rect 22376 1362 22428 1368
rect 22388 56 22416 1362
rect 22480 202 22508 6734
rect 22756 5098 22784 9318
rect 22848 7313 22876 11194
rect 23124 9081 23152 11194
rect 23400 9674 23428 11194
rect 23570 9888 23626 9897
rect 23570 9823 23626 9832
rect 23216 9646 23428 9674
rect 23110 9072 23166 9081
rect 22928 9036 22980 9042
rect 23110 9007 23166 9016
rect 22928 8978 22980 8984
rect 22834 7304 22890 7313
rect 22834 7239 22890 7248
rect 22744 5092 22796 5098
rect 22744 5034 22796 5040
rect 22940 5030 22968 8978
rect 23112 8424 23164 8430
rect 23112 8366 23164 8372
rect 23124 8090 23152 8366
rect 23112 8084 23164 8090
rect 23112 8026 23164 8032
rect 23216 7886 23244 9646
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23388 8560 23440 8566
rect 23388 8502 23440 8508
rect 23400 7993 23428 8502
rect 23492 8090 23520 8774
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 23386 7984 23442 7993
rect 23386 7919 23442 7928
rect 23584 7886 23612 9823
rect 23676 8265 23704 11194
rect 23952 10062 23980 11194
rect 23940 10056 23992 10062
rect 23940 9998 23992 10004
rect 23848 9580 23900 9586
rect 23848 9522 23900 9528
rect 23756 8356 23808 8362
rect 23756 8298 23808 8304
rect 23662 8256 23718 8265
rect 23662 8191 23718 8200
rect 23204 7880 23256 7886
rect 23204 7822 23256 7828
rect 23572 7880 23624 7886
rect 23572 7822 23624 7828
rect 23768 7546 23796 8298
rect 23756 7540 23808 7546
rect 23756 7482 23808 7488
rect 23860 6322 23888 9522
rect 24228 9518 24256 11194
rect 24216 9512 24268 9518
rect 24216 9454 24268 9460
rect 24032 9240 24084 9246
rect 24032 9182 24084 9188
rect 23940 9172 23992 9178
rect 23940 9114 23992 9120
rect 23848 6316 23900 6322
rect 23848 6258 23900 6264
rect 23952 6202 23980 9114
rect 23860 6174 23980 6202
rect 22928 5024 22980 5030
rect 22928 4966 22980 4972
rect 23860 4622 23888 6174
rect 24044 4758 24072 9182
rect 24504 7342 24532 11194
rect 24780 9654 24808 11194
rect 24768 9648 24820 9654
rect 24768 9590 24820 9596
rect 24584 8832 24636 8838
rect 24584 8774 24636 8780
rect 24492 7336 24544 7342
rect 24398 7304 24454 7313
rect 24492 7278 24544 7284
rect 24398 7239 24454 7248
rect 24032 4752 24084 4758
rect 24032 4694 24084 4700
rect 24308 4684 24360 4690
rect 24308 4626 24360 4632
rect 23848 4616 23900 4622
rect 23848 4558 23900 4564
rect 23754 3088 23810 3097
rect 23754 3023 23756 3032
rect 23808 3023 23810 3032
rect 23756 2994 23808 3000
rect 24032 2848 24084 2854
rect 24032 2790 24084 2796
rect 24044 2378 24072 2790
rect 24032 2372 24084 2378
rect 24032 2314 24084 2320
rect 22468 196 22520 202
rect 22468 138 22520 144
rect 24320 56 24348 4626
rect 24412 2854 24440 7239
rect 24596 5234 24624 8774
rect 24952 8424 25004 8430
rect 24952 8366 25004 8372
rect 24768 7472 24820 7478
rect 24768 7414 24820 7420
rect 24780 6662 24808 7414
rect 24768 6656 24820 6662
rect 24768 6598 24820 6604
rect 24584 5228 24636 5234
rect 24584 5170 24636 5176
rect 24964 2854 24992 8366
rect 25056 5273 25084 11194
rect 25332 10033 25360 11194
rect 25318 10024 25374 10033
rect 25318 9959 25374 9968
rect 25042 5264 25098 5273
rect 25042 5199 25098 5208
rect 25608 4214 25636 11194
rect 25884 6390 25912 11194
rect 26160 10849 26188 11194
rect 26436 10985 26464 11194
rect 26422 10976 26478 10985
rect 26422 10911 26478 10920
rect 26146 10840 26202 10849
rect 26146 10775 26202 10784
rect 26712 10305 26740 11194
rect 26988 10713 27016 11194
rect 26974 10704 27030 10713
rect 26974 10639 27030 10648
rect 26698 10296 26754 10305
rect 26698 10231 26754 10240
rect 26516 9444 26568 9450
rect 26516 9386 26568 9392
rect 26424 9308 26476 9314
rect 26424 9250 26476 9256
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 26436 6458 26464 9250
rect 26424 6452 26476 6458
rect 26424 6394 26476 6400
rect 25872 6384 25924 6390
rect 25872 6326 25924 6332
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 25872 5704 25924 5710
rect 25872 5646 25924 5652
rect 25596 4208 25648 4214
rect 25596 4150 25648 4156
rect 24400 2848 24452 2854
rect 24400 2790 24452 2796
rect 24584 2848 24636 2854
rect 24584 2790 24636 2796
rect 24952 2848 25004 2854
rect 24952 2790 25004 2796
rect 24596 105 24624 2790
rect 24582 96 24638 105
rect 8850 0 8906 40
rect 10782 0 10838 56
rect 12714 0 12770 56
rect 14646 0 14702 56
rect 16578 0 16634 56
rect 18510 54 18644 56
rect 18510 0 18566 54
rect 20442 0 20498 56
rect 22374 0 22430 56
rect 24306 0 24362 56
rect 25884 66 25912 5646
rect 26148 5568 26200 5574
rect 26148 5510 26200 5516
rect 26160 5098 26188 5510
rect 26148 5092 26200 5098
rect 26148 5034 26200 5040
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 26330 4176 26386 4185
rect 26330 4111 26386 4120
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 26344 1442 26372 4111
rect 26528 3058 26556 9386
rect 27264 8838 27292 11194
rect 27540 9874 27568 11194
rect 27856 11194 27858 11212
rect 28078 11194 28134 11250
rect 28354 11194 28410 11250
rect 28630 11194 28686 11250
rect 28906 11194 28962 11250
rect 29182 11194 29238 11250
rect 29458 11194 29514 11250
rect 29734 11194 29790 11250
rect 30010 11194 30066 11250
rect 30286 11194 30342 11250
rect 30562 11194 30618 11250
rect 30838 11194 30894 11250
rect 31114 11194 31170 11250
rect 31390 11194 31446 11250
rect 31666 11194 31722 11250
rect 31942 11194 31998 11250
rect 32218 11194 32274 11250
rect 32494 11194 32550 11250
rect 32770 11194 32826 11250
rect 33046 11194 33102 11250
rect 33322 11194 33378 11250
rect 33598 11194 33654 11250
rect 33874 11194 33930 11250
rect 34150 11194 34206 11250
rect 34426 11194 34482 11250
rect 34702 11194 34758 11250
rect 34978 11194 35034 11250
rect 35254 11194 35310 11250
rect 35530 11194 35586 11250
rect 35806 11194 35862 11250
rect 36082 11194 36138 11250
rect 36358 11194 36414 11250
rect 36634 11194 36690 11250
rect 36910 11194 36966 11250
rect 37186 11194 37242 11250
rect 37462 11194 37518 11250
rect 37738 11194 37794 11250
rect 27804 11154 27856 11160
rect 27448 9846 27568 9874
rect 27252 8832 27304 8838
rect 27252 8774 27304 8780
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 27448 7449 27476 9846
rect 27526 9752 27582 9761
rect 27526 9687 27582 9696
rect 27434 7440 27490 7449
rect 27434 7375 27490 7384
rect 26884 7336 26936 7342
rect 26884 7278 26936 7284
rect 26896 7002 26924 7278
rect 26884 6996 26936 7002
rect 26884 6938 26936 6944
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 27540 5234 27568 9687
rect 27710 9616 27766 9625
rect 27710 9551 27766 9560
rect 27620 8084 27672 8090
rect 27620 8026 27672 8032
rect 27632 7886 27660 8026
rect 27724 7886 27752 9551
rect 28092 9110 28120 11194
rect 28080 9104 28132 9110
rect 28080 9046 28132 9052
rect 27620 7880 27672 7886
rect 27620 7822 27672 7828
rect 27712 7880 27764 7886
rect 27712 7822 27764 7828
rect 27724 7750 27752 7822
rect 27712 7744 27764 7750
rect 27712 7686 27764 7692
rect 27896 7744 27948 7750
rect 27896 7686 27948 7692
rect 27908 7546 27936 7686
rect 27896 7540 27948 7546
rect 27896 7482 27948 7488
rect 28368 7410 28396 11194
rect 28644 9897 28672 11194
rect 28630 9888 28686 9897
rect 28630 9823 28686 9832
rect 28920 8090 28948 11194
rect 29196 9058 29224 11194
rect 29104 9030 29224 9058
rect 28908 8084 28960 8090
rect 28908 8026 28960 8032
rect 28356 7404 28408 7410
rect 28356 7346 28408 7352
rect 29104 6798 29132 9030
rect 29472 8786 29500 11194
rect 29748 9761 29776 11194
rect 29734 9752 29790 9761
rect 29734 9687 29790 9696
rect 29196 8758 29500 8786
rect 29920 8832 29972 8838
rect 29920 8774 29972 8780
rect 29092 6792 29144 6798
rect 29092 6734 29144 6740
rect 29196 6322 29224 8758
rect 29184 6316 29236 6322
rect 29184 6258 29236 6264
rect 29368 6248 29420 6254
rect 29368 6190 29420 6196
rect 27620 5840 27672 5846
rect 27620 5782 27672 5788
rect 27632 5370 27660 5782
rect 29000 5568 29052 5574
rect 29000 5510 29052 5516
rect 27620 5364 27672 5370
rect 27620 5306 27672 5312
rect 27528 5228 27580 5234
rect 27528 5170 27580 5176
rect 28080 4616 28132 4622
rect 28080 4558 28132 4564
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 26976 4072 27028 4078
rect 26804 4020 26976 4026
rect 26804 4014 27028 4020
rect 26804 3998 27016 4014
rect 26804 3942 26832 3998
rect 26792 3936 26844 3942
rect 26792 3878 26844 3884
rect 26884 3936 26936 3942
rect 26884 3878 26936 3884
rect 26896 3534 26924 3878
rect 28092 3754 28120 4558
rect 29012 3942 29040 5510
rect 29380 5166 29408 6190
rect 29368 5160 29420 5166
rect 29368 5102 29420 5108
rect 29000 3936 29052 3942
rect 29000 3878 29052 3884
rect 28092 3726 28212 3754
rect 26884 3528 26936 3534
rect 26884 3470 26936 3476
rect 27342 3496 27398 3505
rect 27342 3431 27398 3440
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 26516 3052 26568 3058
rect 26516 2994 26568 3000
rect 27356 2854 27384 3431
rect 28080 3052 28132 3058
rect 28080 2994 28132 3000
rect 28092 2961 28120 2994
rect 28078 2952 28134 2961
rect 28078 2887 28134 2896
rect 27344 2848 27396 2854
rect 27344 2790 27396 2796
rect 26528 2514 26740 2530
rect 26516 2508 26752 2514
rect 26568 2502 26700 2508
rect 26516 2450 26568 2456
rect 26700 2450 26752 2456
rect 26424 2440 26476 2446
rect 26792 2440 26844 2446
rect 26476 2388 26792 2394
rect 26424 2382 26844 2388
rect 26436 2366 26832 2382
rect 26884 2304 26936 2310
rect 26884 2246 26936 2252
rect 26896 1970 26924 2246
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 26884 1964 26936 1970
rect 26884 1906 26936 1912
rect 26252 1414 26372 1442
rect 24582 31 24638 40
rect 25872 60 25924 66
rect 26252 56 26280 1414
rect 28184 56 28212 3726
rect 28264 3664 28316 3670
rect 28264 3606 28316 3612
rect 28276 2854 28304 3606
rect 29000 3528 29052 3534
rect 29000 3470 29052 3476
rect 28264 2848 28316 2854
rect 28264 2790 28316 2796
rect 28448 2848 28500 2854
rect 28448 2790 28500 2796
rect 28816 2848 28868 2854
rect 28816 2790 28868 2796
rect 28460 2553 28488 2790
rect 28446 2544 28502 2553
rect 28446 2479 28502 2488
rect 28828 2378 28856 2790
rect 28816 2372 28868 2378
rect 28816 2314 28868 2320
rect 29012 1426 29040 3470
rect 29932 3398 29960 8774
rect 30024 5710 30052 11194
rect 30300 6322 30328 11194
rect 30380 8492 30432 8498
rect 30380 8434 30432 8440
rect 30288 6316 30340 6322
rect 30288 6258 30340 6264
rect 30392 5914 30420 8434
rect 30576 6798 30604 11194
rect 30748 8900 30800 8906
rect 30748 8842 30800 8848
rect 30656 7472 30708 7478
rect 30656 7414 30708 7420
rect 30564 6792 30616 6798
rect 30470 6760 30526 6769
rect 30564 6734 30616 6740
rect 30470 6695 30526 6704
rect 30484 6662 30512 6695
rect 30472 6656 30524 6662
rect 30472 6598 30524 6604
rect 30380 5908 30432 5914
rect 30380 5850 30432 5856
rect 30012 5704 30064 5710
rect 30012 5646 30064 5652
rect 30104 4616 30156 4622
rect 30104 4558 30156 4564
rect 29920 3392 29972 3398
rect 29920 3334 29972 3340
rect 30012 2848 30064 2854
rect 30012 2790 30064 2796
rect 30024 2106 30052 2790
rect 30012 2100 30064 2106
rect 30012 2042 30064 2048
rect 29000 1420 29052 1426
rect 29000 1362 29052 1368
rect 30116 56 30144 4558
rect 30668 3942 30696 7414
rect 30760 4486 30788 8842
rect 30852 7410 30880 11194
rect 30932 8356 30984 8362
rect 30932 8298 30984 8304
rect 30840 7404 30892 7410
rect 30840 7346 30892 7352
rect 30748 4480 30800 4486
rect 30748 4422 30800 4428
rect 30656 3936 30708 3942
rect 30656 3878 30708 3884
rect 30944 2854 30972 8298
rect 31024 8288 31076 8294
rect 31024 8230 31076 8236
rect 31036 8090 31064 8230
rect 31024 8084 31076 8090
rect 31024 8026 31076 8032
rect 31128 7886 31156 11194
rect 31404 7886 31432 11194
rect 31576 8016 31628 8022
rect 31574 7984 31576 7993
rect 31628 7984 31630 7993
rect 31574 7919 31630 7928
rect 31116 7880 31168 7886
rect 31116 7822 31168 7828
rect 31392 7880 31444 7886
rect 31392 7822 31444 7828
rect 31680 6798 31708 11194
rect 31956 9674 31984 11194
rect 31864 9646 31984 9674
rect 31864 7954 31892 9646
rect 32232 8634 32260 11194
rect 32508 8634 32536 11194
rect 32784 9602 32812 11194
rect 32784 9574 32904 9602
rect 32588 8968 32640 8974
rect 32588 8910 32640 8916
rect 32220 8628 32272 8634
rect 32220 8570 32272 8576
rect 32496 8628 32548 8634
rect 32496 8570 32548 8576
rect 32600 8498 32628 8910
rect 32876 8634 32904 9574
rect 33060 8838 33088 11194
rect 33336 9058 33364 11194
rect 33336 9030 33456 9058
rect 33612 9042 33640 11194
rect 33048 8832 33100 8838
rect 33048 8774 33100 8780
rect 33010 8732 33318 8741
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 33010 8667 33318 8676
rect 32864 8628 32916 8634
rect 32864 8570 32916 8576
rect 33428 8566 33456 9030
rect 33600 9036 33652 9042
rect 33600 8978 33652 8984
rect 33508 8832 33560 8838
rect 33508 8774 33560 8780
rect 33784 8832 33836 8838
rect 33784 8774 33836 8780
rect 33520 8634 33548 8774
rect 33508 8628 33560 8634
rect 33508 8570 33560 8576
rect 33416 8560 33468 8566
rect 33416 8502 33468 8508
rect 32588 8492 32640 8498
rect 32588 8434 32640 8440
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 31852 7948 31904 7954
rect 31852 7890 31904 7896
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 31668 6792 31720 6798
rect 31668 6734 31720 6740
rect 32692 6730 32720 8434
rect 33010 7644 33318 7653
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 33690 7440 33746 7449
rect 33690 7375 33746 7384
rect 33704 7274 33732 7375
rect 33692 7268 33744 7274
rect 33692 7210 33744 7216
rect 32864 6996 32916 7002
rect 32864 6938 32916 6944
rect 32680 6724 32732 6730
rect 32680 6666 32732 6672
rect 31024 6384 31076 6390
rect 31024 6326 31076 6332
rect 31036 4554 31064 6326
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 32876 4826 32904 6938
rect 33010 6556 33318 6565
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 33010 5468 33318 5477
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 33010 5403 33318 5412
rect 33796 4826 33824 8774
rect 33888 8378 33916 11194
rect 34164 8566 34192 11194
rect 34244 9036 34296 9042
rect 34244 8978 34296 8984
rect 34256 8634 34284 8978
rect 34244 8628 34296 8634
rect 34244 8570 34296 8576
rect 34152 8560 34204 8566
rect 34152 8502 34204 8508
rect 34060 8492 34112 8498
rect 34060 8434 34112 8440
rect 33888 8362 34008 8378
rect 33888 8356 34020 8362
rect 33888 8350 33968 8356
rect 33968 8298 34020 8304
rect 32864 4820 32916 4826
rect 32864 4762 32916 4768
rect 33784 4820 33836 4826
rect 33784 4762 33836 4768
rect 31024 4548 31076 4554
rect 31024 4490 31076 4496
rect 33968 4548 34020 4554
rect 33968 4490 34020 4496
rect 33010 4380 33318 4389
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 31760 4140 31812 4146
rect 31760 4082 31812 4088
rect 33416 4140 33468 4146
rect 33416 4082 33468 4088
rect 30932 2848 30984 2854
rect 30932 2790 30984 2796
rect 31574 2544 31630 2553
rect 31574 2479 31576 2488
rect 31628 2479 31630 2488
rect 31576 2450 31628 2456
rect 25872 2 25924 8
rect 26238 0 26294 56
rect 28170 0 28226 56
rect 30102 0 30158 56
rect 31772 42 31800 4082
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 32862 3632 32918 3641
rect 32862 3567 32918 3576
rect 32876 3194 32904 3567
rect 33010 3292 33318 3301
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 32864 3188 32916 3194
rect 32864 3130 32916 3136
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 32588 2440 32640 2446
rect 32586 2408 32588 2417
rect 32680 2440 32732 2446
rect 32640 2408 32642 2417
rect 32680 2382 32732 2388
rect 32586 2343 32642 2352
rect 32692 2310 32720 2382
rect 32680 2304 32732 2310
rect 32680 2246 32732 2252
rect 33010 2204 33318 2213
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 33428 1970 33456 4082
rect 33416 1964 33468 1970
rect 33416 1906 33468 1912
rect 31956 56 32076 82
rect 33980 56 34008 4490
rect 34072 3534 34100 8434
rect 34440 8090 34468 11194
rect 34716 8634 34744 11194
rect 34704 8628 34756 8634
rect 34704 8570 34756 8576
rect 34888 8492 34940 8498
rect 34888 8434 34940 8440
rect 34428 8084 34480 8090
rect 34428 8026 34480 8032
rect 34152 7540 34204 7546
rect 34152 7482 34204 7488
rect 34164 6934 34192 7482
rect 34152 6928 34204 6934
rect 34152 6870 34204 6876
rect 34336 6316 34388 6322
rect 34336 6258 34388 6264
rect 34348 4593 34376 6258
rect 34334 4584 34390 4593
rect 34334 4519 34390 4528
rect 34060 3528 34112 3534
rect 34060 3470 34112 3476
rect 34900 3194 34928 8434
rect 34992 8378 35020 11194
rect 35268 8498 35296 11194
rect 35256 8492 35308 8498
rect 35256 8434 35308 8440
rect 34992 8362 35388 8378
rect 34992 8356 35400 8362
rect 34992 8350 35348 8356
rect 35348 8298 35400 8304
rect 35544 8090 35572 11194
rect 35820 8634 35848 11194
rect 35808 8628 35860 8634
rect 35808 8570 35860 8576
rect 35624 8560 35676 8566
rect 35624 8502 35676 8508
rect 35532 8084 35584 8090
rect 35532 8026 35584 8032
rect 35346 7848 35402 7857
rect 35346 7783 35402 7792
rect 35360 7750 35388 7783
rect 35348 7744 35400 7750
rect 35348 7686 35400 7692
rect 35636 5574 35664 8502
rect 35716 8492 35768 8498
rect 35716 8434 35768 8440
rect 35808 8492 35860 8498
rect 35808 8434 35860 8440
rect 35728 5794 35756 8434
rect 35820 5914 35848 8434
rect 36096 8090 36124 11194
rect 36176 8900 36228 8906
rect 36176 8842 36228 8848
rect 36188 8498 36216 8842
rect 36176 8492 36228 8498
rect 36176 8434 36228 8440
rect 36372 8430 36400 11194
rect 36544 9376 36596 9382
rect 36544 9318 36596 9324
rect 36556 8498 36584 9318
rect 36544 8492 36596 8498
rect 36544 8434 36596 8440
rect 36360 8424 36412 8430
rect 36360 8366 36412 8372
rect 36648 8090 36676 11194
rect 36924 8634 36952 11194
rect 36912 8628 36964 8634
rect 36912 8570 36964 8576
rect 37200 8362 37228 11194
rect 37280 8968 37332 8974
rect 37280 8910 37332 8916
rect 37292 8498 37320 8910
rect 37476 8566 37504 11194
rect 37464 8560 37516 8566
rect 37464 8502 37516 8508
rect 37280 8492 37332 8498
rect 37280 8434 37332 8440
rect 37372 8492 37424 8498
rect 37372 8434 37424 8440
rect 37384 8378 37412 8434
rect 37188 8356 37240 8362
rect 37188 8298 37240 8304
rect 37292 8350 37412 8378
rect 37292 8242 37320 8350
rect 37200 8214 37320 8242
rect 36084 8084 36136 8090
rect 36084 8026 36136 8032
rect 36636 8084 36688 8090
rect 36636 8026 36688 8032
rect 35900 7880 35952 7886
rect 35900 7822 35952 7828
rect 36176 7880 36228 7886
rect 36176 7822 36228 7828
rect 36452 7880 36504 7886
rect 36452 7822 36504 7828
rect 35912 6390 35940 7822
rect 35900 6384 35952 6390
rect 35900 6326 35952 6332
rect 35808 5908 35860 5914
rect 35808 5850 35860 5856
rect 35900 5908 35952 5914
rect 35900 5850 35952 5856
rect 35912 5794 35940 5850
rect 35728 5766 35940 5794
rect 35624 5568 35676 5574
rect 35624 5510 35676 5516
rect 36084 5568 36136 5574
rect 36084 5510 36136 5516
rect 35992 5160 36044 5166
rect 35992 5102 36044 5108
rect 35900 4616 35952 4622
rect 35900 4558 35952 4564
rect 35256 4072 35308 4078
rect 35256 4014 35308 4020
rect 35268 3534 35296 4014
rect 35256 3528 35308 3534
rect 35256 3470 35308 3476
rect 34888 3188 34940 3194
rect 34888 3130 34940 3136
rect 35912 56 35940 4558
rect 36004 3466 36032 5102
rect 35992 3460 36044 3466
rect 35992 3402 36044 3408
rect 36096 3126 36124 5510
rect 36188 4690 36216 7822
rect 36360 7812 36412 7818
rect 36360 7754 36412 7760
rect 36268 7744 36320 7750
rect 36268 7686 36320 7692
rect 36176 4684 36228 4690
rect 36176 4626 36228 4632
rect 36280 3942 36308 7686
rect 36372 7313 36400 7754
rect 36464 7546 36492 7822
rect 36452 7540 36504 7546
rect 36452 7482 36504 7488
rect 36358 7304 36414 7313
rect 36358 7239 36414 7248
rect 37096 5704 37148 5710
rect 37096 5646 37148 5652
rect 36268 3936 36320 3942
rect 36268 3878 36320 3884
rect 36084 3120 36136 3126
rect 36084 3062 36136 3068
rect 37108 134 37136 5646
rect 37200 4486 37228 8214
rect 37752 8090 37780 11194
rect 38382 9888 38438 9897
rect 38382 9823 38438 9832
rect 38016 8832 38068 8838
rect 38016 8774 38068 8780
rect 38028 8498 38056 8774
rect 38016 8492 38068 8498
rect 38016 8434 38068 8440
rect 37950 8188 38258 8197
rect 37950 8186 37956 8188
rect 38012 8186 38036 8188
rect 38092 8186 38116 8188
rect 38172 8186 38196 8188
rect 38252 8186 38258 8188
rect 38012 8134 38014 8186
rect 38194 8134 38196 8186
rect 37950 8132 37956 8134
rect 38012 8132 38036 8134
rect 38092 8132 38116 8134
rect 38172 8132 38196 8134
rect 38252 8132 38258 8134
rect 37950 8123 38258 8132
rect 37740 8084 37792 8090
rect 37740 8026 37792 8032
rect 38198 7984 38254 7993
rect 38198 7919 38254 7928
rect 37740 7404 37792 7410
rect 37740 7346 37792 7352
rect 37752 6254 37780 7346
rect 38212 7342 38240 7919
rect 38292 7880 38344 7886
rect 38292 7822 38344 7828
rect 38200 7336 38252 7342
rect 38200 7278 38252 7284
rect 37950 7100 38258 7109
rect 37950 7098 37956 7100
rect 38012 7098 38036 7100
rect 38092 7098 38116 7100
rect 38172 7098 38196 7100
rect 38252 7098 38258 7100
rect 38012 7046 38014 7098
rect 38194 7046 38196 7098
rect 37950 7044 37956 7046
rect 38012 7044 38036 7046
rect 38092 7044 38116 7046
rect 38172 7044 38196 7046
rect 38252 7044 38258 7046
rect 37950 7035 38258 7044
rect 37740 6248 37792 6254
rect 37740 6190 37792 6196
rect 37950 6012 38258 6021
rect 37950 6010 37956 6012
rect 38012 6010 38036 6012
rect 38092 6010 38116 6012
rect 38172 6010 38196 6012
rect 38252 6010 38258 6012
rect 38012 5958 38014 6010
rect 38194 5958 38196 6010
rect 37950 5956 37956 5958
rect 38012 5956 38036 5958
rect 38092 5956 38116 5958
rect 38172 5956 38196 5958
rect 38252 5956 38258 5958
rect 37950 5947 38258 5956
rect 38304 5914 38332 7822
rect 38396 7410 38424 9823
rect 39670 9616 39726 9625
rect 39670 9551 39726 9560
rect 38750 9344 38806 9353
rect 38750 9279 38806 9288
rect 38658 8528 38714 8537
rect 38568 8492 38620 8498
rect 38658 8463 38714 8472
rect 38568 8434 38620 8440
rect 38580 7970 38608 8434
rect 38672 8090 38700 8463
rect 38660 8084 38712 8090
rect 38660 8026 38712 8032
rect 38580 7942 38700 7970
rect 38568 7472 38620 7478
rect 38474 7440 38530 7449
rect 38384 7404 38436 7410
rect 38568 7414 38620 7420
rect 38474 7375 38476 7384
rect 38384 7346 38436 7352
rect 38528 7375 38530 7384
rect 38476 7346 38528 7352
rect 38476 6792 38528 6798
rect 38476 6734 38528 6740
rect 38488 6118 38516 6734
rect 38476 6112 38528 6118
rect 38476 6054 38528 6060
rect 38292 5908 38344 5914
rect 38292 5850 38344 5856
rect 37832 5636 37884 5642
rect 37832 5578 37884 5584
rect 37280 5228 37332 5234
rect 37280 5170 37332 5176
rect 37188 4480 37240 4486
rect 37188 4422 37240 4428
rect 37292 3738 37320 5170
rect 37280 3732 37332 3738
rect 37280 3674 37332 3680
rect 37096 128 37148 134
rect 37096 70 37148 76
rect 37844 56 37872 5578
rect 37950 4924 38258 4933
rect 37950 4922 37956 4924
rect 38012 4922 38036 4924
rect 38092 4922 38116 4924
rect 38172 4922 38196 4924
rect 38252 4922 38258 4924
rect 38012 4870 38014 4922
rect 38194 4870 38196 4922
rect 37950 4868 37956 4870
rect 38012 4868 38036 4870
rect 38092 4868 38116 4870
rect 38172 4868 38196 4870
rect 38252 4868 38258 4870
rect 37950 4859 38258 4868
rect 37950 3836 38258 3845
rect 37950 3834 37956 3836
rect 38012 3834 38036 3836
rect 38092 3834 38116 3836
rect 38172 3834 38196 3836
rect 38252 3834 38258 3836
rect 38012 3782 38014 3834
rect 38194 3782 38196 3834
rect 37950 3780 37956 3782
rect 38012 3780 38036 3782
rect 38092 3780 38116 3782
rect 38172 3780 38196 3782
rect 38252 3780 38258 3782
rect 37950 3771 38258 3780
rect 38580 3505 38608 7414
rect 38672 6746 38700 7942
rect 38764 7546 38792 9279
rect 38936 9240 38988 9246
rect 38936 9182 38988 9188
rect 38948 8498 38976 9182
rect 39578 9072 39634 9081
rect 39578 9007 39634 9016
rect 39486 8800 39542 8809
rect 39010 8732 39318 8741
rect 39486 8735 39542 8744
rect 39010 8730 39016 8732
rect 39072 8730 39096 8732
rect 39152 8730 39176 8732
rect 39232 8730 39256 8732
rect 39312 8730 39318 8732
rect 39072 8678 39074 8730
rect 39254 8678 39256 8730
rect 39010 8676 39016 8678
rect 39072 8676 39096 8678
rect 39152 8676 39176 8678
rect 39232 8676 39256 8678
rect 39312 8676 39318 8678
rect 39010 8667 39318 8676
rect 38936 8492 38988 8498
rect 38936 8434 38988 8440
rect 39028 8356 39080 8362
rect 39028 8298 39080 8304
rect 39396 8356 39448 8362
rect 39396 8298 39448 8304
rect 39040 8265 39068 8298
rect 39026 8256 39082 8265
rect 39026 8191 39082 8200
rect 39408 7993 39436 8298
rect 39394 7984 39450 7993
rect 39394 7919 39450 7928
rect 38844 7880 38896 7886
rect 38844 7822 38896 7828
rect 38752 7540 38804 7546
rect 38752 7482 38804 7488
rect 38856 7002 38884 7822
rect 38936 7744 38988 7750
rect 39396 7744 39448 7750
rect 38936 7686 38988 7692
rect 39394 7712 39396 7721
rect 39448 7712 39450 7721
rect 38948 7449 38976 7686
rect 39010 7644 39318 7653
rect 39394 7647 39450 7656
rect 39010 7642 39016 7644
rect 39072 7642 39096 7644
rect 39152 7642 39176 7644
rect 39232 7642 39256 7644
rect 39312 7642 39318 7644
rect 39072 7590 39074 7642
rect 39254 7590 39256 7642
rect 39010 7588 39016 7590
rect 39072 7588 39096 7590
rect 39152 7588 39176 7590
rect 39232 7588 39256 7590
rect 39312 7588 39318 7590
rect 39010 7579 39318 7588
rect 39500 7546 39528 8735
rect 39488 7540 39540 7546
rect 39488 7482 39540 7488
rect 38934 7440 38990 7449
rect 38934 7375 38990 7384
rect 39488 7268 39540 7274
rect 39488 7210 39540 7216
rect 39396 7200 39448 7206
rect 39394 7168 39396 7177
rect 39448 7168 39450 7177
rect 39394 7103 39450 7112
rect 38844 6996 38896 7002
rect 38844 6938 38896 6944
rect 39500 6905 39528 7210
rect 39486 6896 39542 6905
rect 39486 6831 39542 6840
rect 38936 6792 38988 6798
rect 38672 6718 38792 6746
rect 38936 6734 38988 6740
rect 38660 6656 38712 6662
rect 38660 6598 38712 6604
rect 38672 6361 38700 6598
rect 38658 6352 38714 6361
rect 38658 6287 38714 6296
rect 38764 6186 38792 6718
rect 38752 6180 38804 6186
rect 38752 6122 38804 6128
rect 38752 5908 38804 5914
rect 38752 5850 38804 5856
rect 38764 5710 38792 5850
rect 38948 5817 38976 6734
rect 39592 6662 39620 9007
rect 39684 6730 39712 9551
rect 39672 6724 39724 6730
rect 39672 6666 39724 6672
rect 39580 6656 39632 6662
rect 39394 6624 39450 6633
rect 39580 6598 39632 6604
rect 39010 6556 39318 6565
rect 39394 6559 39450 6568
rect 39010 6554 39016 6556
rect 39072 6554 39096 6556
rect 39152 6554 39176 6556
rect 39232 6554 39256 6556
rect 39312 6554 39318 6556
rect 39072 6502 39074 6554
rect 39254 6502 39256 6554
rect 39010 6500 39016 6502
rect 39072 6500 39096 6502
rect 39152 6500 39176 6502
rect 39232 6500 39256 6502
rect 39312 6500 39318 6502
rect 39010 6491 39318 6500
rect 39408 6458 39436 6559
rect 39396 6452 39448 6458
rect 39396 6394 39448 6400
rect 39212 6316 39264 6322
rect 39212 6258 39264 6264
rect 39028 6112 39080 6118
rect 39026 6080 39028 6089
rect 39080 6080 39082 6089
rect 39026 6015 39082 6024
rect 39224 5846 39252 6258
rect 39764 5908 39816 5914
rect 39764 5850 39816 5856
rect 39212 5840 39264 5846
rect 38934 5808 38990 5817
rect 39396 5840 39448 5846
rect 39212 5782 39264 5788
rect 39394 5808 39396 5817
rect 39448 5808 39450 5817
rect 38934 5743 38990 5752
rect 39394 5743 39450 5752
rect 38752 5704 38804 5710
rect 38752 5646 38804 5652
rect 39010 5468 39318 5477
rect 39010 5466 39016 5468
rect 39072 5466 39096 5468
rect 39152 5466 39176 5468
rect 39232 5466 39256 5468
rect 39312 5466 39318 5468
rect 39072 5414 39074 5466
rect 39254 5414 39256 5466
rect 39010 5412 39016 5414
rect 39072 5412 39096 5414
rect 39152 5412 39176 5414
rect 39232 5412 39256 5414
rect 39312 5412 39318 5414
rect 39010 5403 39318 5412
rect 39396 5364 39448 5370
rect 39396 5306 39448 5312
rect 39408 5273 39436 5306
rect 39394 5264 39450 5273
rect 39394 5199 39450 5208
rect 38660 5092 38712 5098
rect 38660 5034 38712 5040
rect 38672 4078 38700 5034
rect 39028 5024 39080 5030
rect 39026 4992 39028 5001
rect 39080 4992 39082 5001
rect 39026 4927 39082 4936
rect 39396 4752 39448 4758
rect 39394 4720 39396 4729
rect 39448 4720 39450 4729
rect 39394 4655 39450 4664
rect 38844 4616 38896 4622
rect 38844 4558 38896 4564
rect 38936 4616 38988 4622
rect 38936 4558 38988 4564
rect 38856 4282 38884 4558
rect 38844 4276 38896 4282
rect 38844 4218 38896 4224
rect 38948 4214 38976 4558
rect 39010 4380 39318 4389
rect 39010 4378 39016 4380
rect 39072 4378 39096 4380
rect 39152 4378 39176 4380
rect 39232 4378 39256 4380
rect 39312 4378 39318 4380
rect 39072 4326 39074 4378
rect 39254 4326 39256 4378
rect 39010 4324 39016 4326
rect 39072 4324 39096 4326
rect 39152 4324 39176 4326
rect 39232 4324 39256 4326
rect 39312 4324 39318 4326
rect 39010 4315 39318 4324
rect 38936 4208 38988 4214
rect 38936 4150 38988 4156
rect 39394 4176 39450 4185
rect 38844 4140 38896 4146
rect 39394 4111 39450 4120
rect 38844 4082 38896 4088
rect 38660 4072 38712 4078
rect 38660 4014 38712 4020
rect 38566 3496 38622 3505
rect 38566 3431 38622 3440
rect 38856 3398 38884 4082
rect 39408 4010 39436 4111
rect 39212 4004 39264 4010
rect 39212 3946 39264 3952
rect 39396 4004 39448 4010
rect 39396 3946 39448 3952
rect 39028 3936 39080 3942
rect 39026 3904 39028 3913
rect 39080 3904 39082 3913
rect 39026 3839 39082 3848
rect 39224 3534 39252 3946
rect 39396 3664 39448 3670
rect 39394 3632 39396 3641
rect 39448 3632 39450 3641
rect 39394 3567 39450 3576
rect 39212 3528 39264 3534
rect 39212 3470 39264 3476
rect 38844 3392 38896 3398
rect 38844 3334 38896 3340
rect 39010 3292 39318 3301
rect 39010 3290 39016 3292
rect 39072 3290 39096 3292
rect 39152 3290 39176 3292
rect 39232 3290 39256 3292
rect 39312 3290 39318 3292
rect 39072 3238 39074 3290
rect 39254 3238 39256 3290
rect 39010 3236 39016 3238
rect 39072 3236 39096 3238
rect 39152 3236 39176 3238
rect 39232 3236 39256 3238
rect 39312 3236 39318 3238
rect 39010 3227 39318 3236
rect 39396 3188 39448 3194
rect 39396 3130 39448 3136
rect 39408 3097 39436 3130
rect 39394 3088 39450 3097
rect 39394 3023 39450 3032
rect 39028 2848 39080 2854
rect 39026 2816 39028 2825
rect 39080 2816 39082 2825
rect 37950 2748 38258 2757
rect 39026 2751 39082 2760
rect 37950 2746 37956 2748
rect 38012 2746 38036 2748
rect 38092 2746 38116 2748
rect 38172 2746 38196 2748
rect 38252 2746 38258 2748
rect 38012 2694 38014 2746
rect 38194 2694 38196 2746
rect 37950 2692 37956 2694
rect 38012 2692 38036 2694
rect 38092 2692 38116 2694
rect 38172 2692 38196 2694
rect 38252 2692 38258 2694
rect 37950 2683 38258 2692
rect 38108 2644 38160 2650
rect 38108 2586 38160 2592
rect 38120 2446 38148 2586
rect 38568 2576 38620 2582
rect 38474 2544 38530 2553
rect 39396 2576 39448 2582
rect 38568 2518 38620 2524
rect 39394 2544 39396 2553
rect 39448 2544 39450 2553
rect 38474 2479 38530 2488
rect 38488 2446 38516 2479
rect 38108 2440 38160 2446
rect 38108 2382 38160 2388
rect 38476 2440 38528 2446
rect 38580 2417 38608 2518
rect 39394 2479 39450 2488
rect 38476 2382 38528 2388
rect 38566 2408 38622 2417
rect 38566 2343 38622 2352
rect 37924 2304 37976 2310
rect 37924 2246 37976 2252
rect 38292 2304 38344 2310
rect 38292 2246 38344 2252
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 37936 2009 37964 2246
rect 37922 2000 37978 2009
rect 37922 1935 37978 1944
rect 38304 1737 38332 2246
rect 38290 1728 38346 1737
rect 38290 1663 38346 1672
rect 38672 1465 38700 2246
rect 39010 2204 39318 2213
rect 39010 2202 39016 2204
rect 39072 2202 39096 2204
rect 39152 2202 39176 2204
rect 39232 2202 39256 2204
rect 39312 2202 39318 2204
rect 39072 2150 39074 2202
rect 39254 2150 39256 2202
rect 39010 2148 39016 2150
rect 39072 2148 39096 2150
rect 39152 2148 39176 2150
rect 39232 2148 39256 2150
rect 39312 2148 39318 2150
rect 39010 2139 39318 2148
rect 38658 1456 38714 1465
rect 38658 1391 38714 1400
rect 39776 56 39804 5850
rect 39948 5568 40000 5574
rect 39946 5536 39948 5545
rect 40000 5536 40002 5545
rect 39946 5471 40002 5480
rect 39948 4480 40000 4486
rect 39946 4448 39948 4457
rect 40000 4448 40002 4457
rect 39946 4383 40002 4392
rect 39948 3392 40000 3398
rect 39946 3360 39948 3369
rect 40000 3360 40002 3369
rect 39946 3295 40002 3304
rect 39948 2304 40000 2310
rect 39946 2272 39948 2281
rect 40000 2272 40002 2281
rect 39946 2207 40002 2216
rect 31956 54 32090 56
rect 31956 42 31984 54
rect 31772 14 31984 42
rect 32034 0 32090 54
rect 33966 0 34022 56
rect 35898 0 35954 56
rect 37830 0 37886 56
rect 39762 0 39818 56
<< via2 >>
rect 1122 8200 1178 8256
rect 202 7928 258 7984
rect 662 7656 718 7712
rect 2778 8744 2834 8800
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 2778 8336 2834 8392
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 1306 7112 1362 7168
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1766 6704 1822 6760
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 2778 6568 2834 6624
rect 1766 6024 1822 6080
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 3974 7948 4030 7984
rect 3974 7928 3976 7948
rect 3976 7928 4028 7948
rect 4028 7928 4030 7948
rect 3514 7248 3570 7304
rect 3422 5752 3478 5808
rect 2778 5616 2834 5672
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 2686 5208 2742 5264
rect 2686 4936 2742 4992
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 2870 3984 2926 4040
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 2870 3304 2926 3360
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 5538 6160 5594 6216
rect 5722 5072 5778 5128
rect 7470 11056 7526 11112
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 9770 10240 9826 10296
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 10230 7656 10286 7712
rect 10230 7248 10286 7304
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 10782 7792 10838 7848
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 7562 4936 7618 4992
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 12714 10920 12770 10976
rect 11150 6704 11206 6760
rect 13082 10784 13138 10840
rect 13174 7792 13230 7848
rect 12346 7384 12402 7440
rect 13542 8880 13598 8936
rect 13358 6160 13414 6216
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 14646 10648 14702 10704
rect 13726 7248 13782 7304
rect 8206 4664 8262 4720
rect 11426 4548 11482 4584
rect 11426 4528 11428 4548
rect 11428 4528 11480 4548
rect 11480 4528 11482 4548
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 8298 3440 8354 3496
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 10782 3168 10838 3224
rect 14646 8064 14702 8120
rect 14646 7656 14702 7712
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 15474 9016 15530 9072
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 14278 7384 14334 7440
rect 14554 7384 14610 7440
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 14370 6976 14426 7032
rect 13818 6704 13874 6760
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 15474 5752 15530 5808
rect 14738 5208 14794 5264
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 16302 9696 16358 9752
rect 16578 9016 16634 9072
rect 16302 6840 16358 6896
rect 16486 7248 16542 7304
rect 16670 5616 16726 5672
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 14922 4120 14978 4176
rect 16486 3612 16488 3632
rect 16488 3612 16540 3632
rect 16540 3612 16542 3632
rect 16486 3576 16542 3612
rect 14646 3440 14702 3496
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 8850 2352 8906 2408
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 9402 1944 9458 2000
rect 9494 1672 9550 1728
rect 9586 1400 9642 1456
rect 8850 40 8906 96
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 18050 9288 18106 9344
rect 18878 10104 18934 10160
rect 18142 7112 18198 7168
rect 19062 9968 19118 10024
rect 18970 9696 19026 9752
rect 19154 9832 19210 9888
rect 19154 6316 19210 6352
rect 19154 6296 19156 6316
rect 19156 6296 19208 6316
rect 19208 6296 19210 6316
rect 19798 10104 19854 10160
rect 20074 8608 20130 8664
rect 20350 8200 20406 8256
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 19798 8064 19854 8120
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 20626 8472 20682 8528
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 19706 5480 19762 5536
rect 17314 5228 17370 5264
rect 17314 5208 17316 5228
rect 17316 5208 17368 5228
rect 17368 5208 17370 5228
rect 17866 5072 17922 5128
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 14830 3168 14886 3224
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 19798 4120 19854 4176
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 14830 2760 14886 2816
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 20718 3984 20774 4040
rect 21454 8880 21510 8936
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 21822 8336 21878 8392
rect 22558 11056 22614 11112
rect 22006 6976 22062 7032
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 20718 3188 20774 3224
rect 20718 3168 20720 3188
rect 20720 3168 20772 3188
rect 20772 3168 20774 3188
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 23570 9832 23626 9888
rect 23110 9016 23166 9072
rect 22834 7248 22890 7304
rect 23386 7928 23442 7984
rect 23662 8200 23718 8256
rect 24398 7248 24454 7304
rect 23754 3052 23810 3088
rect 23754 3032 23756 3052
rect 23756 3032 23808 3052
rect 23808 3032 23810 3052
rect 25318 9968 25374 10024
rect 25042 5208 25098 5264
rect 26422 10920 26478 10976
rect 26146 10784 26202 10840
rect 26974 10648 27030 10704
rect 26698 10240 26754 10296
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 24582 40 24638 96
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 26330 4120 26386 4176
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 27526 9696 27582 9752
rect 27434 7384 27490 7440
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27710 9560 27766 9616
rect 28630 9832 28686 9888
rect 29734 9696 29790 9752
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 27342 3440 27398 3496
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 28078 2896 28134 2952
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 28446 2488 28502 2544
rect 30470 6704 30526 6760
rect 31574 7964 31576 7984
rect 31576 7964 31628 7984
rect 31628 7964 31630 7984
rect 31574 7928 31630 7964
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 33690 7384 33746 7440
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 31574 2508 31630 2544
rect 31574 2488 31576 2508
rect 31576 2488 31628 2508
rect 31628 2488 31630 2508
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 32862 3576 32918 3632
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 32586 2388 32588 2408
rect 32588 2388 32640 2408
rect 32640 2388 32642 2408
rect 32586 2352 32642 2388
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
rect 34334 4528 34390 4584
rect 35346 7792 35402 7848
rect 36358 7248 36414 7304
rect 38382 9832 38438 9888
rect 37956 8186 38012 8188
rect 38036 8186 38092 8188
rect 38116 8186 38172 8188
rect 38196 8186 38252 8188
rect 37956 8134 38002 8186
rect 38002 8134 38012 8186
rect 38036 8134 38066 8186
rect 38066 8134 38078 8186
rect 38078 8134 38092 8186
rect 38116 8134 38130 8186
rect 38130 8134 38142 8186
rect 38142 8134 38172 8186
rect 38196 8134 38206 8186
rect 38206 8134 38252 8186
rect 37956 8132 38012 8134
rect 38036 8132 38092 8134
rect 38116 8132 38172 8134
rect 38196 8132 38252 8134
rect 38198 7928 38254 7984
rect 37956 7098 38012 7100
rect 38036 7098 38092 7100
rect 38116 7098 38172 7100
rect 38196 7098 38252 7100
rect 37956 7046 38002 7098
rect 38002 7046 38012 7098
rect 38036 7046 38066 7098
rect 38066 7046 38078 7098
rect 38078 7046 38092 7098
rect 38116 7046 38130 7098
rect 38130 7046 38142 7098
rect 38142 7046 38172 7098
rect 38196 7046 38206 7098
rect 38206 7046 38252 7098
rect 37956 7044 38012 7046
rect 38036 7044 38092 7046
rect 38116 7044 38172 7046
rect 38196 7044 38252 7046
rect 37956 6010 38012 6012
rect 38036 6010 38092 6012
rect 38116 6010 38172 6012
rect 38196 6010 38252 6012
rect 37956 5958 38002 6010
rect 38002 5958 38012 6010
rect 38036 5958 38066 6010
rect 38066 5958 38078 6010
rect 38078 5958 38092 6010
rect 38116 5958 38130 6010
rect 38130 5958 38142 6010
rect 38142 5958 38172 6010
rect 38196 5958 38206 6010
rect 38206 5958 38252 6010
rect 37956 5956 38012 5958
rect 38036 5956 38092 5958
rect 38116 5956 38172 5958
rect 38196 5956 38252 5958
rect 39670 9560 39726 9616
rect 38750 9288 38806 9344
rect 38658 8472 38714 8528
rect 38474 7404 38530 7440
rect 38474 7384 38476 7404
rect 38476 7384 38528 7404
rect 38528 7384 38530 7404
rect 37956 4922 38012 4924
rect 38036 4922 38092 4924
rect 38116 4922 38172 4924
rect 38196 4922 38252 4924
rect 37956 4870 38002 4922
rect 38002 4870 38012 4922
rect 38036 4870 38066 4922
rect 38066 4870 38078 4922
rect 38078 4870 38092 4922
rect 38116 4870 38130 4922
rect 38130 4870 38142 4922
rect 38142 4870 38172 4922
rect 38196 4870 38206 4922
rect 38206 4870 38252 4922
rect 37956 4868 38012 4870
rect 38036 4868 38092 4870
rect 38116 4868 38172 4870
rect 38196 4868 38252 4870
rect 37956 3834 38012 3836
rect 38036 3834 38092 3836
rect 38116 3834 38172 3836
rect 38196 3834 38252 3836
rect 37956 3782 38002 3834
rect 38002 3782 38012 3834
rect 38036 3782 38066 3834
rect 38066 3782 38078 3834
rect 38078 3782 38092 3834
rect 38116 3782 38130 3834
rect 38130 3782 38142 3834
rect 38142 3782 38172 3834
rect 38196 3782 38206 3834
rect 38206 3782 38252 3834
rect 37956 3780 38012 3782
rect 38036 3780 38092 3782
rect 38116 3780 38172 3782
rect 38196 3780 38252 3782
rect 39578 9016 39634 9072
rect 39486 8744 39542 8800
rect 39016 8730 39072 8732
rect 39096 8730 39152 8732
rect 39176 8730 39232 8732
rect 39256 8730 39312 8732
rect 39016 8678 39062 8730
rect 39062 8678 39072 8730
rect 39096 8678 39126 8730
rect 39126 8678 39138 8730
rect 39138 8678 39152 8730
rect 39176 8678 39190 8730
rect 39190 8678 39202 8730
rect 39202 8678 39232 8730
rect 39256 8678 39266 8730
rect 39266 8678 39312 8730
rect 39016 8676 39072 8678
rect 39096 8676 39152 8678
rect 39176 8676 39232 8678
rect 39256 8676 39312 8678
rect 39026 8200 39082 8256
rect 39394 7928 39450 7984
rect 39394 7692 39396 7712
rect 39396 7692 39448 7712
rect 39448 7692 39450 7712
rect 39394 7656 39450 7692
rect 39016 7642 39072 7644
rect 39096 7642 39152 7644
rect 39176 7642 39232 7644
rect 39256 7642 39312 7644
rect 39016 7590 39062 7642
rect 39062 7590 39072 7642
rect 39096 7590 39126 7642
rect 39126 7590 39138 7642
rect 39138 7590 39152 7642
rect 39176 7590 39190 7642
rect 39190 7590 39202 7642
rect 39202 7590 39232 7642
rect 39256 7590 39266 7642
rect 39266 7590 39312 7642
rect 39016 7588 39072 7590
rect 39096 7588 39152 7590
rect 39176 7588 39232 7590
rect 39256 7588 39312 7590
rect 38934 7384 38990 7440
rect 39394 7148 39396 7168
rect 39396 7148 39448 7168
rect 39448 7148 39450 7168
rect 39394 7112 39450 7148
rect 39486 6840 39542 6896
rect 38658 6296 38714 6352
rect 39394 6568 39450 6624
rect 39016 6554 39072 6556
rect 39096 6554 39152 6556
rect 39176 6554 39232 6556
rect 39256 6554 39312 6556
rect 39016 6502 39062 6554
rect 39062 6502 39072 6554
rect 39096 6502 39126 6554
rect 39126 6502 39138 6554
rect 39138 6502 39152 6554
rect 39176 6502 39190 6554
rect 39190 6502 39202 6554
rect 39202 6502 39232 6554
rect 39256 6502 39266 6554
rect 39266 6502 39312 6554
rect 39016 6500 39072 6502
rect 39096 6500 39152 6502
rect 39176 6500 39232 6502
rect 39256 6500 39312 6502
rect 39026 6060 39028 6080
rect 39028 6060 39080 6080
rect 39080 6060 39082 6080
rect 39026 6024 39082 6060
rect 38934 5752 38990 5808
rect 39394 5788 39396 5808
rect 39396 5788 39448 5808
rect 39448 5788 39450 5808
rect 39394 5752 39450 5788
rect 39016 5466 39072 5468
rect 39096 5466 39152 5468
rect 39176 5466 39232 5468
rect 39256 5466 39312 5468
rect 39016 5414 39062 5466
rect 39062 5414 39072 5466
rect 39096 5414 39126 5466
rect 39126 5414 39138 5466
rect 39138 5414 39152 5466
rect 39176 5414 39190 5466
rect 39190 5414 39202 5466
rect 39202 5414 39232 5466
rect 39256 5414 39266 5466
rect 39266 5414 39312 5466
rect 39016 5412 39072 5414
rect 39096 5412 39152 5414
rect 39176 5412 39232 5414
rect 39256 5412 39312 5414
rect 39394 5208 39450 5264
rect 39026 4972 39028 4992
rect 39028 4972 39080 4992
rect 39080 4972 39082 4992
rect 39026 4936 39082 4972
rect 39394 4700 39396 4720
rect 39396 4700 39448 4720
rect 39448 4700 39450 4720
rect 39394 4664 39450 4700
rect 39016 4378 39072 4380
rect 39096 4378 39152 4380
rect 39176 4378 39232 4380
rect 39256 4378 39312 4380
rect 39016 4326 39062 4378
rect 39062 4326 39072 4378
rect 39096 4326 39126 4378
rect 39126 4326 39138 4378
rect 39138 4326 39152 4378
rect 39176 4326 39190 4378
rect 39190 4326 39202 4378
rect 39202 4326 39232 4378
rect 39256 4326 39266 4378
rect 39266 4326 39312 4378
rect 39016 4324 39072 4326
rect 39096 4324 39152 4326
rect 39176 4324 39232 4326
rect 39256 4324 39312 4326
rect 39394 4120 39450 4176
rect 38566 3440 38622 3496
rect 39026 3884 39028 3904
rect 39028 3884 39080 3904
rect 39080 3884 39082 3904
rect 39026 3848 39082 3884
rect 39394 3612 39396 3632
rect 39396 3612 39448 3632
rect 39448 3612 39450 3632
rect 39394 3576 39450 3612
rect 39016 3290 39072 3292
rect 39096 3290 39152 3292
rect 39176 3290 39232 3292
rect 39256 3290 39312 3292
rect 39016 3238 39062 3290
rect 39062 3238 39072 3290
rect 39096 3238 39126 3290
rect 39126 3238 39138 3290
rect 39138 3238 39152 3290
rect 39176 3238 39190 3290
rect 39190 3238 39202 3290
rect 39202 3238 39232 3290
rect 39256 3238 39266 3290
rect 39266 3238 39312 3290
rect 39016 3236 39072 3238
rect 39096 3236 39152 3238
rect 39176 3236 39232 3238
rect 39256 3236 39312 3238
rect 39394 3032 39450 3088
rect 39026 2796 39028 2816
rect 39028 2796 39080 2816
rect 39080 2796 39082 2816
rect 39026 2760 39082 2796
rect 37956 2746 38012 2748
rect 38036 2746 38092 2748
rect 38116 2746 38172 2748
rect 38196 2746 38252 2748
rect 37956 2694 38002 2746
rect 38002 2694 38012 2746
rect 38036 2694 38066 2746
rect 38066 2694 38078 2746
rect 38078 2694 38092 2746
rect 38116 2694 38130 2746
rect 38130 2694 38142 2746
rect 38142 2694 38172 2746
rect 38196 2694 38206 2746
rect 38206 2694 38252 2746
rect 37956 2692 38012 2694
rect 38036 2692 38092 2694
rect 38116 2692 38172 2694
rect 38196 2692 38252 2694
rect 38474 2488 38530 2544
rect 39394 2524 39396 2544
rect 39396 2524 39448 2544
rect 39448 2524 39450 2544
rect 39394 2488 39450 2524
rect 38566 2352 38622 2408
rect 37922 1944 37978 2000
rect 38290 1672 38346 1728
rect 39016 2202 39072 2204
rect 39096 2202 39152 2204
rect 39176 2202 39232 2204
rect 39256 2202 39312 2204
rect 39016 2150 39062 2202
rect 39062 2150 39072 2202
rect 39096 2150 39126 2202
rect 39126 2150 39138 2202
rect 39138 2150 39152 2202
rect 39176 2150 39190 2202
rect 39190 2150 39202 2202
rect 39202 2150 39232 2202
rect 39256 2150 39266 2202
rect 39266 2150 39312 2202
rect 39016 2148 39072 2150
rect 39096 2148 39152 2150
rect 39176 2148 39232 2150
rect 39256 2148 39312 2150
rect 38658 1400 38714 1456
rect 39946 5516 39948 5536
rect 39948 5516 40000 5536
rect 40000 5516 40002 5536
rect 39946 5480 40002 5516
rect 39946 4428 39948 4448
rect 39948 4428 40000 4448
rect 40000 4428 40002 4448
rect 39946 4392 40002 4428
rect 39946 3340 39948 3360
rect 39948 3340 40000 3360
rect 40000 3340 40002 3360
rect 39946 3304 40002 3340
rect 39946 2252 39948 2272
rect 39948 2252 40000 2272
rect 40000 2252 40002 2272
rect 39946 2216 40002 2252
<< metal3 >>
rect 7465 11114 7531 11117
rect 22553 11114 22619 11117
rect 7465 11112 22619 11114
rect 7465 11056 7470 11112
rect 7526 11056 22558 11112
rect 22614 11056 22619 11112
rect 7465 11054 22619 11056
rect 7465 11051 7531 11054
rect 22553 11051 22619 11054
rect 12709 10978 12775 10981
rect 26417 10978 26483 10981
rect 12709 10976 26483 10978
rect 12709 10920 12714 10976
rect 12770 10920 26422 10976
rect 26478 10920 26483 10976
rect 12709 10918 26483 10920
rect 12709 10915 12775 10918
rect 26417 10915 26483 10918
rect 13077 10842 13143 10845
rect 26141 10842 26207 10845
rect 13077 10840 26207 10842
rect 13077 10784 13082 10840
rect 13138 10784 26146 10840
rect 26202 10784 26207 10840
rect 13077 10782 26207 10784
rect 13077 10779 13143 10782
rect 26141 10779 26207 10782
rect 14641 10706 14707 10709
rect 26969 10706 27035 10709
rect 14641 10704 27035 10706
rect 14641 10648 14646 10704
rect 14702 10648 26974 10704
rect 27030 10648 27035 10704
rect 14641 10646 27035 10648
rect 14641 10643 14707 10646
rect 26969 10643 27035 10646
rect 9765 10298 9831 10301
rect 26693 10298 26759 10301
rect 9765 10296 26759 10298
rect 9765 10240 9770 10296
rect 9826 10240 26698 10296
rect 26754 10240 26759 10296
rect 9765 10238 26759 10240
rect 9765 10235 9831 10238
rect 26693 10235 26759 10238
rect 18873 10162 18939 10165
rect 19793 10162 19859 10165
rect 18873 10160 19859 10162
rect 18873 10104 18878 10160
rect 18934 10104 19798 10160
rect 19854 10104 19859 10160
rect 18873 10102 19859 10104
rect 18873 10099 18939 10102
rect 19793 10099 19859 10102
rect 19057 10026 19123 10029
rect 25313 10026 25379 10029
rect 19057 10024 25379 10026
rect 19057 9968 19062 10024
rect 19118 9968 25318 10024
rect 25374 9968 25379 10024
rect 19057 9966 25379 9968
rect 19057 9963 19123 9966
rect 25313 9963 25379 9966
rect 0 9890 120 9920
rect 19149 9890 19215 9893
rect 0 9888 19215 9890
rect 0 9832 19154 9888
rect 19210 9832 19215 9888
rect 0 9830 19215 9832
rect 0 9800 120 9830
rect 19149 9827 19215 9830
rect 23565 9890 23631 9893
rect 28625 9890 28691 9893
rect 23565 9888 28691 9890
rect 23565 9832 23570 9888
rect 23626 9832 28630 9888
rect 28686 9832 28691 9888
rect 23565 9830 28691 9832
rect 23565 9827 23631 9830
rect 28625 9827 28691 9830
rect 38377 9890 38443 9893
rect 40880 9890 41000 9920
rect 38377 9888 41000 9890
rect 38377 9832 38382 9888
rect 38438 9832 41000 9888
rect 38377 9830 41000 9832
rect 38377 9827 38443 9830
rect 40880 9800 41000 9830
rect 16297 9754 16363 9757
rect 18965 9754 19031 9757
rect 16297 9752 19031 9754
rect 16297 9696 16302 9752
rect 16358 9696 18970 9752
rect 19026 9696 19031 9752
rect 16297 9694 19031 9696
rect 16297 9691 16363 9694
rect 18965 9691 19031 9694
rect 27521 9754 27587 9757
rect 29729 9754 29795 9757
rect 27521 9752 29795 9754
rect 27521 9696 27526 9752
rect 27582 9696 29734 9752
rect 29790 9696 29795 9752
rect 27521 9694 29795 9696
rect 27521 9691 27587 9694
rect 29729 9691 29795 9694
rect 0 9618 120 9648
rect 27705 9618 27771 9621
rect 0 9616 27771 9618
rect 0 9560 27710 9616
rect 27766 9560 27771 9616
rect 0 9558 27771 9560
rect 0 9528 120 9558
rect 27705 9555 27771 9558
rect 39665 9618 39731 9621
rect 40880 9618 41000 9648
rect 39665 9616 41000 9618
rect 39665 9560 39670 9616
rect 39726 9560 41000 9616
rect 39665 9558 41000 9560
rect 39665 9555 39731 9558
rect 40880 9528 41000 9558
rect 0 9346 120 9376
rect 18045 9346 18111 9349
rect 0 9344 18111 9346
rect 0 9288 18050 9344
rect 18106 9288 18111 9344
rect 0 9286 18111 9288
rect 0 9256 120 9286
rect 18045 9283 18111 9286
rect 38745 9346 38811 9349
rect 40880 9346 41000 9376
rect 38745 9344 41000 9346
rect 38745 9288 38750 9344
rect 38806 9288 41000 9344
rect 38745 9286 41000 9288
rect 38745 9283 38811 9286
rect 40880 9256 41000 9286
rect 0 9074 120 9104
rect 15469 9074 15535 9077
rect 0 9072 15535 9074
rect 0 9016 15474 9072
rect 15530 9016 15535 9072
rect 0 9014 15535 9016
rect 0 8984 120 9014
rect 15469 9011 15535 9014
rect 16573 9074 16639 9077
rect 23105 9074 23171 9077
rect 16573 9072 23171 9074
rect 16573 9016 16578 9072
rect 16634 9016 23110 9072
rect 23166 9016 23171 9072
rect 16573 9014 23171 9016
rect 16573 9011 16639 9014
rect 23105 9011 23171 9014
rect 39573 9074 39639 9077
rect 40880 9074 41000 9104
rect 39573 9072 41000 9074
rect 39573 9016 39578 9072
rect 39634 9016 41000 9072
rect 39573 9014 41000 9016
rect 39573 9011 39639 9014
rect 40880 8984 41000 9014
rect 13537 8938 13603 8941
rect 21449 8938 21515 8941
rect 13537 8936 21515 8938
rect 13537 8880 13542 8936
rect 13598 8880 21454 8936
rect 21510 8880 21515 8936
rect 13537 8878 21515 8880
rect 13537 8875 13603 8878
rect 21449 8875 21515 8878
rect 0 8802 120 8832
rect 2773 8802 2839 8805
rect 0 8800 2839 8802
rect 0 8744 2778 8800
rect 2834 8744 2839 8800
rect 0 8742 2839 8744
rect 0 8712 120 8742
rect 2773 8739 2839 8742
rect 39481 8802 39547 8805
rect 40880 8802 41000 8832
rect 39481 8800 41000 8802
rect 39481 8744 39486 8800
rect 39542 8744 41000 8800
rect 39481 8742 41000 8744
rect 39481 8739 39547 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 33006 8671 33322 8672
rect 39006 8736 39322 8737
rect 39006 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39322 8736
rect 40880 8712 41000 8742
rect 39006 8671 39322 8672
rect 19742 8604 19748 8668
rect 19812 8666 19818 8668
rect 20069 8666 20135 8669
rect 19812 8664 20135 8666
rect 19812 8608 20074 8664
rect 20130 8608 20135 8664
rect 19812 8606 20135 8608
rect 19812 8604 19818 8606
rect 20069 8603 20135 8606
rect 0 8530 120 8560
rect 20621 8530 20687 8533
rect 0 8528 20687 8530
rect 0 8472 20626 8528
rect 20682 8472 20687 8528
rect 0 8470 20687 8472
rect 0 8440 120 8470
rect 20621 8467 20687 8470
rect 38653 8530 38719 8533
rect 40880 8530 41000 8560
rect 38653 8528 41000 8530
rect 38653 8472 38658 8528
rect 38714 8472 41000 8528
rect 38653 8470 41000 8472
rect 38653 8467 38719 8470
rect 40880 8440 41000 8470
rect 2773 8394 2839 8397
rect 21817 8394 21883 8397
rect 2773 8392 21883 8394
rect 2773 8336 2778 8392
rect 2834 8336 21822 8392
rect 21878 8336 21883 8392
rect 2773 8334 21883 8336
rect 2773 8331 2839 8334
rect 21817 8331 21883 8334
rect 0 8258 120 8288
rect 1117 8258 1183 8261
rect 0 8256 1183 8258
rect 0 8200 1122 8256
rect 1178 8200 1183 8256
rect 0 8198 1183 8200
rect 0 8168 120 8198
rect 1117 8195 1183 8198
rect 20345 8258 20411 8261
rect 23657 8258 23723 8261
rect 20345 8256 23723 8258
rect 20345 8200 20350 8256
rect 20406 8200 23662 8256
rect 23718 8200 23723 8256
rect 20345 8198 23723 8200
rect 20345 8195 20411 8198
rect 23657 8195 23723 8198
rect 39021 8258 39087 8261
rect 40880 8258 41000 8288
rect 39021 8256 41000 8258
rect 39021 8200 39026 8256
rect 39082 8200 41000 8256
rect 39021 8198 41000 8200
rect 39021 8195 39087 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 37946 8192 38262 8193
rect 37946 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38262 8192
rect 40880 8168 41000 8198
rect 37946 8127 38262 8128
rect 14641 8122 14707 8125
rect 19793 8122 19859 8125
rect 14641 8120 19859 8122
rect 14641 8064 14646 8120
rect 14702 8064 19798 8120
rect 19854 8064 19859 8120
rect 14641 8062 19859 8064
rect 14641 8059 14707 8062
rect 19793 8059 19859 8062
rect 0 7986 120 8016
rect 197 7986 263 7989
rect 0 7984 263 7986
rect 0 7928 202 7984
rect 258 7928 263 7984
rect 0 7926 263 7928
rect 0 7896 120 7926
rect 197 7923 263 7926
rect 3969 7986 4035 7989
rect 23381 7986 23447 7989
rect 3969 7984 23447 7986
rect 3969 7928 3974 7984
rect 4030 7928 23386 7984
rect 23442 7928 23447 7984
rect 3969 7926 23447 7928
rect 3969 7923 4035 7926
rect 23381 7923 23447 7926
rect 31569 7986 31635 7989
rect 38193 7986 38259 7989
rect 31569 7984 38259 7986
rect 31569 7928 31574 7984
rect 31630 7928 38198 7984
rect 38254 7928 38259 7984
rect 31569 7926 38259 7928
rect 31569 7923 31635 7926
rect 38193 7923 38259 7926
rect 39389 7986 39455 7989
rect 40880 7986 41000 8016
rect 39389 7984 41000 7986
rect 39389 7928 39394 7984
rect 39450 7928 41000 7984
rect 39389 7926 41000 7928
rect 39389 7923 39455 7926
rect 40880 7896 41000 7926
rect 10777 7850 10843 7853
rect 13169 7850 13235 7853
rect 35341 7850 35407 7853
rect 10777 7848 13002 7850
rect 10777 7792 10782 7848
rect 10838 7792 13002 7848
rect 10777 7790 13002 7792
rect 10777 7787 10843 7790
rect 0 7714 120 7744
rect 657 7714 723 7717
rect 0 7712 723 7714
rect 0 7656 662 7712
rect 718 7656 723 7712
rect 0 7654 723 7656
rect 0 7624 120 7654
rect 657 7651 723 7654
rect 10225 7714 10291 7717
rect 12942 7714 13002 7790
rect 13169 7848 35407 7850
rect 13169 7792 13174 7848
rect 13230 7792 35346 7848
rect 35402 7792 35407 7848
rect 13169 7790 35407 7792
rect 13169 7787 13235 7790
rect 35341 7787 35407 7790
rect 14641 7714 14707 7717
rect 10225 7712 12450 7714
rect 10225 7656 10230 7712
rect 10286 7656 12450 7712
rect 10225 7654 12450 7656
rect 12942 7712 14707 7714
rect 12942 7656 14646 7712
rect 14702 7656 14707 7712
rect 12942 7654 14707 7656
rect 10225 7651 10291 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 12390 7578 12450 7654
rect 14641 7651 14707 7654
rect 39389 7714 39455 7717
rect 40880 7714 41000 7744
rect 39389 7712 41000 7714
rect 39389 7656 39394 7712
rect 39450 7656 41000 7712
rect 39389 7654 41000 7656
rect 39389 7651 39455 7654
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 33006 7583 33322 7584
rect 39006 7648 39322 7649
rect 39006 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39322 7648
rect 40880 7624 41000 7654
rect 39006 7583 39322 7584
rect 12390 7518 14474 7578
rect 0 7442 120 7472
rect 12341 7442 12407 7445
rect 14273 7442 14339 7445
rect 0 7382 10426 7442
rect 0 7352 120 7382
rect 3509 7306 3575 7309
rect 10225 7306 10291 7309
rect 3509 7304 10291 7306
rect 3509 7248 3514 7304
rect 3570 7248 10230 7304
rect 10286 7248 10291 7304
rect 3509 7246 10291 7248
rect 10366 7306 10426 7382
rect 12341 7440 14339 7442
rect 12341 7384 12346 7440
rect 12402 7384 14278 7440
rect 14334 7384 14339 7440
rect 12341 7382 14339 7384
rect 12341 7379 12407 7382
rect 14273 7379 14339 7382
rect 13721 7306 13787 7309
rect 10366 7304 13787 7306
rect 10366 7248 13726 7304
rect 13782 7248 13787 7304
rect 10366 7246 13787 7248
rect 3509 7243 3575 7246
rect 10225 7243 10291 7246
rect 13721 7243 13787 7246
rect 0 7170 120 7200
rect 1301 7170 1367 7173
rect 0 7168 1367 7170
rect 0 7112 1306 7168
rect 1362 7112 1367 7168
rect 0 7110 1367 7112
rect 14414 7170 14474 7518
rect 14549 7442 14615 7445
rect 27429 7442 27495 7445
rect 14549 7440 27495 7442
rect 14549 7384 14554 7440
rect 14610 7384 27434 7440
rect 27490 7384 27495 7440
rect 14549 7382 27495 7384
rect 14549 7379 14615 7382
rect 27429 7379 27495 7382
rect 33685 7442 33751 7445
rect 38469 7442 38535 7445
rect 33685 7440 38535 7442
rect 33685 7384 33690 7440
rect 33746 7384 38474 7440
rect 38530 7384 38535 7440
rect 33685 7382 38535 7384
rect 33685 7379 33751 7382
rect 38469 7379 38535 7382
rect 38929 7442 38995 7445
rect 40880 7442 41000 7472
rect 38929 7440 41000 7442
rect 38929 7384 38934 7440
rect 38990 7384 41000 7440
rect 38929 7382 41000 7384
rect 38929 7379 38995 7382
rect 40880 7352 41000 7382
rect 16481 7306 16547 7309
rect 22829 7306 22895 7309
rect 16481 7304 22895 7306
rect 16481 7248 16486 7304
rect 16542 7248 22834 7304
rect 22890 7248 22895 7304
rect 16481 7246 22895 7248
rect 16481 7243 16547 7246
rect 22829 7243 22895 7246
rect 24393 7306 24459 7309
rect 36353 7306 36419 7309
rect 24393 7304 36419 7306
rect 24393 7248 24398 7304
rect 24454 7248 36358 7304
rect 36414 7248 36419 7304
rect 24393 7246 36419 7248
rect 24393 7243 24459 7246
rect 36353 7243 36419 7246
rect 18137 7170 18203 7173
rect 14414 7168 18203 7170
rect 14414 7112 18142 7168
rect 18198 7112 18203 7168
rect 14414 7110 18203 7112
rect 0 7080 120 7110
rect 1301 7107 1367 7110
rect 18137 7107 18203 7110
rect 39389 7170 39455 7173
rect 40880 7170 41000 7200
rect 39389 7168 41000 7170
rect 39389 7112 39394 7168
rect 39450 7112 41000 7168
rect 39389 7110 41000 7112
rect 39389 7107 39455 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 37946 7104 38262 7105
rect 37946 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38262 7104
rect 40880 7080 41000 7110
rect 37946 7039 38262 7040
rect 14365 7034 14431 7037
rect 22001 7034 22067 7037
rect 14365 7032 19810 7034
rect 14365 6976 14370 7032
rect 14426 6976 19810 7032
rect 14365 6974 19810 6976
rect 14365 6971 14431 6974
rect 0 6898 120 6928
rect 16297 6898 16363 6901
rect 0 6896 16363 6898
rect 0 6840 16302 6896
rect 16358 6840 16363 6896
rect 0 6838 16363 6840
rect 19750 6898 19810 6974
rect 20486 7032 22067 7034
rect 20486 6976 22006 7032
rect 22062 6976 22067 7032
rect 20486 6974 22067 6976
rect 20486 6898 20546 6974
rect 22001 6971 22067 6974
rect 19750 6838 20546 6898
rect 39481 6898 39547 6901
rect 40880 6898 41000 6928
rect 39481 6896 41000 6898
rect 39481 6840 39486 6896
rect 39542 6840 41000 6896
rect 39481 6838 41000 6840
rect 0 6808 120 6838
rect 16297 6835 16363 6838
rect 39481 6835 39547 6838
rect 40880 6808 41000 6838
rect 1761 6762 1827 6765
rect 11145 6762 11211 6765
rect 1761 6760 11211 6762
rect 1761 6704 1766 6760
rect 1822 6704 11150 6760
rect 11206 6704 11211 6760
rect 1761 6702 11211 6704
rect 1761 6699 1827 6702
rect 11145 6699 11211 6702
rect 13813 6762 13879 6765
rect 30465 6762 30531 6765
rect 13813 6760 30531 6762
rect 13813 6704 13818 6760
rect 13874 6704 30470 6760
rect 30526 6704 30531 6760
rect 13813 6702 30531 6704
rect 13813 6699 13879 6702
rect 30465 6699 30531 6702
rect 0 6626 120 6656
rect 2773 6626 2839 6629
rect 0 6624 2839 6626
rect 0 6568 2778 6624
rect 2834 6568 2839 6624
rect 0 6566 2839 6568
rect 0 6536 120 6566
rect 2773 6563 2839 6566
rect 39389 6626 39455 6629
rect 40880 6626 41000 6656
rect 39389 6624 41000 6626
rect 39389 6568 39394 6624
rect 39450 6568 41000 6624
rect 39389 6566 41000 6568
rect 39389 6563 39455 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 33006 6495 33322 6496
rect 39006 6560 39322 6561
rect 39006 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39322 6560
rect 40880 6536 41000 6566
rect 39006 6495 39322 6496
rect 0 6354 120 6384
rect 19149 6354 19215 6357
rect 0 6352 19215 6354
rect 0 6296 19154 6352
rect 19210 6296 19215 6352
rect 0 6294 19215 6296
rect 0 6264 120 6294
rect 19149 6291 19215 6294
rect 38653 6354 38719 6357
rect 40880 6354 41000 6384
rect 38653 6352 41000 6354
rect 38653 6296 38658 6352
rect 38714 6296 41000 6352
rect 38653 6294 41000 6296
rect 38653 6291 38719 6294
rect 40880 6264 41000 6294
rect 5533 6218 5599 6221
rect 13353 6218 13419 6221
rect 5533 6216 13419 6218
rect 5533 6160 5538 6216
rect 5594 6160 13358 6216
rect 13414 6160 13419 6216
rect 5533 6158 13419 6160
rect 5533 6155 5599 6158
rect 13353 6155 13419 6158
rect 0 6082 120 6112
rect 1761 6082 1827 6085
rect 0 6080 1827 6082
rect 0 6024 1766 6080
rect 1822 6024 1827 6080
rect 0 6022 1827 6024
rect 0 5992 120 6022
rect 1761 6019 1827 6022
rect 39021 6082 39087 6085
rect 40880 6082 41000 6112
rect 39021 6080 41000 6082
rect 39021 6024 39026 6080
rect 39082 6024 41000 6080
rect 39021 6022 41000 6024
rect 39021 6019 39087 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 37946 6016 38262 6017
rect 37946 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38262 6016
rect 40880 5992 41000 6022
rect 37946 5951 38262 5952
rect 0 5810 120 5840
rect 3417 5810 3483 5813
rect 0 5808 3483 5810
rect 0 5752 3422 5808
rect 3478 5752 3483 5808
rect 0 5750 3483 5752
rect 0 5720 120 5750
rect 3417 5747 3483 5750
rect 15469 5810 15535 5813
rect 38929 5810 38995 5813
rect 15469 5808 38995 5810
rect 15469 5752 15474 5808
rect 15530 5752 38934 5808
rect 38990 5752 38995 5808
rect 15469 5750 38995 5752
rect 15469 5747 15535 5750
rect 38929 5747 38995 5750
rect 39389 5810 39455 5813
rect 40880 5810 41000 5840
rect 39389 5808 41000 5810
rect 39389 5752 39394 5808
rect 39450 5752 41000 5808
rect 39389 5750 41000 5752
rect 39389 5747 39455 5750
rect 40880 5720 41000 5750
rect 2773 5674 2839 5677
rect 16665 5674 16731 5677
rect 2773 5672 16731 5674
rect 2773 5616 2778 5672
rect 2834 5616 16670 5672
rect 16726 5616 16731 5672
rect 2773 5614 16731 5616
rect 2773 5611 2839 5614
rect 16665 5611 16731 5614
rect 0 5538 120 5568
rect 19701 5540 19767 5541
rect 19701 5538 19748 5540
rect 0 5478 2882 5538
rect 19656 5536 19748 5538
rect 19656 5480 19706 5536
rect 19656 5478 19748 5480
rect 0 5448 120 5478
rect 0 5266 120 5296
rect 2681 5266 2747 5269
rect 0 5264 2747 5266
rect 0 5208 2686 5264
rect 2742 5208 2747 5264
rect 0 5206 2747 5208
rect 2822 5266 2882 5478
rect 19701 5476 19748 5478
rect 19812 5476 19818 5540
rect 39941 5538 40007 5541
rect 40880 5538 41000 5568
rect 39941 5536 41000 5538
rect 39941 5480 39946 5536
rect 40002 5480 41000 5536
rect 39941 5478 41000 5480
rect 19701 5475 19767 5476
rect 39941 5475 40007 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 33006 5407 33322 5408
rect 39006 5472 39322 5473
rect 39006 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39322 5472
rect 40880 5448 41000 5478
rect 39006 5407 39322 5408
rect 14733 5266 14799 5269
rect 2822 5264 14799 5266
rect 2822 5208 14738 5264
rect 14794 5208 14799 5264
rect 2822 5206 14799 5208
rect 0 5176 120 5206
rect 2681 5203 2747 5206
rect 14733 5203 14799 5206
rect 17309 5266 17375 5269
rect 25037 5266 25103 5269
rect 17309 5264 25103 5266
rect 17309 5208 17314 5264
rect 17370 5208 25042 5264
rect 25098 5208 25103 5264
rect 17309 5206 25103 5208
rect 17309 5203 17375 5206
rect 25037 5203 25103 5206
rect 39389 5266 39455 5269
rect 40880 5266 41000 5296
rect 39389 5264 41000 5266
rect 39389 5208 39394 5264
rect 39450 5208 41000 5264
rect 39389 5206 41000 5208
rect 39389 5203 39455 5206
rect 40880 5176 41000 5206
rect 5717 5130 5783 5133
rect 17861 5130 17927 5133
rect 1718 5128 5783 5130
rect 1718 5072 5722 5128
rect 5778 5072 5783 5128
rect 1718 5070 5783 5072
rect 0 4994 120 5024
rect 1718 4994 1778 5070
rect 5717 5067 5783 5070
rect 8342 5128 17927 5130
rect 8342 5072 17866 5128
rect 17922 5072 17927 5128
rect 8342 5070 17927 5072
rect 0 4934 1778 4994
rect 2681 4994 2747 4997
rect 7557 4994 7623 4997
rect 2681 4992 7623 4994
rect 2681 4936 2686 4992
rect 2742 4936 7562 4992
rect 7618 4936 7623 4992
rect 2681 4934 7623 4936
rect 0 4904 120 4934
rect 2681 4931 2747 4934
rect 7557 4931 7623 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 0 4722 120 4752
rect 8201 4722 8267 4725
rect 0 4720 8267 4722
rect 0 4664 8206 4720
rect 8262 4664 8267 4720
rect 0 4662 8267 4664
rect 0 4632 120 4662
rect 8201 4659 8267 4662
rect 8342 4586 8402 5070
rect 17861 5067 17927 5070
rect 39021 4994 39087 4997
rect 40880 4994 41000 5024
rect 39021 4992 41000 4994
rect 39021 4936 39026 4992
rect 39082 4936 41000 4992
rect 39021 4934 41000 4936
rect 39021 4931 39087 4934
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 37946 4928 38262 4929
rect 37946 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38262 4928
rect 40880 4904 41000 4934
rect 37946 4863 38262 4864
rect 39389 4722 39455 4725
rect 40880 4722 41000 4752
rect 39389 4720 41000 4722
rect 39389 4664 39394 4720
rect 39450 4664 41000 4720
rect 39389 4662 41000 4664
rect 39389 4659 39455 4662
rect 40880 4632 41000 4662
rect 2822 4526 8402 4586
rect 11421 4586 11487 4589
rect 34329 4586 34395 4589
rect 11421 4584 34395 4586
rect 11421 4528 11426 4584
rect 11482 4528 34334 4584
rect 34390 4528 34395 4584
rect 11421 4526 34395 4528
rect 0 4450 120 4480
rect 2822 4450 2882 4526
rect 11421 4523 11487 4526
rect 34329 4523 34395 4526
rect 0 4390 2882 4450
rect 39941 4450 40007 4453
rect 40880 4450 41000 4480
rect 39941 4448 41000 4450
rect 39941 4392 39946 4448
rect 40002 4392 41000 4448
rect 39941 4390 41000 4392
rect 0 4360 120 4390
rect 39941 4387 40007 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 33006 4319 33322 4320
rect 39006 4384 39322 4385
rect 39006 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39322 4384
rect 40880 4360 41000 4390
rect 39006 4319 39322 4320
rect 0 4178 120 4208
rect 14917 4178 14983 4181
rect 0 4176 14983 4178
rect 0 4120 14922 4176
rect 14978 4120 14983 4176
rect 0 4118 14983 4120
rect 0 4088 120 4118
rect 14917 4115 14983 4118
rect 19793 4178 19859 4181
rect 26325 4178 26391 4181
rect 19793 4176 26391 4178
rect 19793 4120 19798 4176
rect 19854 4120 26330 4176
rect 26386 4120 26391 4176
rect 19793 4118 26391 4120
rect 19793 4115 19859 4118
rect 26325 4115 26391 4118
rect 39389 4178 39455 4181
rect 40880 4178 41000 4208
rect 39389 4176 41000 4178
rect 39389 4120 39394 4176
rect 39450 4120 41000 4176
rect 39389 4118 41000 4120
rect 39389 4115 39455 4118
rect 40880 4088 41000 4118
rect 2865 4042 2931 4045
rect 20713 4042 20779 4045
rect 1718 3982 2514 4042
rect 0 3906 120 3936
rect 1718 3906 1778 3982
rect 0 3846 1778 3906
rect 2454 3906 2514 3982
rect 2865 4040 20779 4042
rect 2865 3984 2870 4040
rect 2926 3984 20718 4040
rect 20774 3984 20779 4040
rect 2865 3982 20779 3984
rect 2865 3979 2931 3982
rect 20713 3979 20779 3982
rect 39021 3906 39087 3909
rect 40880 3906 41000 3936
rect 2454 3846 6930 3906
rect 0 3816 120 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 0 3634 120 3664
rect 6870 3634 6930 3846
rect 39021 3904 41000 3906
rect 39021 3848 39026 3904
rect 39082 3848 41000 3904
rect 39021 3846 41000 3848
rect 39021 3843 39087 3846
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 37946 3840 38262 3841
rect 37946 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38262 3840
rect 40880 3816 41000 3846
rect 37946 3775 38262 3776
rect 16481 3634 16547 3637
rect 32857 3634 32923 3637
rect 0 3574 3572 3634
rect 6870 3632 16547 3634
rect 6870 3576 16486 3632
rect 16542 3576 16547 3632
rect 6870 3574 16547 3576
rect 0 3544 120 3574
rect 3512 3498 3572 3574
rect 16481 3571 16547 3574
rect 22050 3632 32923 3634
rect 22050 3576 32862 3632
rect 32918 3576 32923 3632
rect 22050 3574 32923 3576
rect 8293 3498 8359 3501
rect 3512 3496 8359 3498
rect 3512 3440 8298 3496
rect 8354 3440 8359 3496
rect 3512 3438 8359 3440
rect 8293 3435 8359 3438
rect 14641 3498 14707 3501
rect 22050 3498 22110 3574
rect 32857 3571 32923 3574
rect 39389 3634 39455 3637
rect 40880 3634 41000 3664
rect 39389 3632 41000 3634
rect 39389 3576 39394 3632
rect 39450 3576 41000 3632
rect 39389 3574 41000 3576
rect 39389 3571 39455 3574
rect 40880 3544 41000 3574
rect 14641 3496 22110 3498
rect 14641 3440 14646 3496
rect 14702 3440 22110 3496
rect 14641 3438 22110 3440
rect 27337 3498 27403 3501
rect 38561 3498 38627 3501
rect 27337 3496 38627 3498
rect 27337 3440 27342 3496
rect 27398 3440 38566 3496
rect 38622 3440 38627 3496
rect 27337 3438 38627 3440
rect 14641 3435 14707 3438
rect 27337 3435 27403 3438
rect 38561 3435 38627 3438
rect 0 3362 120 3392
rect 2865 3362 2931 3365
rect 0 3360 2931 3362
rect 0 3304 2870 3360
rect 2926 3304 2931 3360
rect 0 3302 2931 3304
rect 0 3272 120 3302
rect 2865 3299 2931 3302
rect 39941 3362 40007 3365
rect 40880 3362 41000 3392
rect 39941 3360 41000 3362
rect 39941 3304 39946 3360
rect 40002 3304 41000 3360
rect 39941 3302 41000 3304
rect 39941 3299 40007 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 33006 3231 33322 3232
rect 39006 3296 39322 3297
rect 39006 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39322 3296
rect 40880 3272 41000 3302
rect 39006 3231 39322 3232
rect 10777 3226 10843 3229
rect 14825 3226 14891 3229
rect 20713 3226 20779 3229
rect 10777 3224 14891 3226
rect 10777 3168 10782 3224
rect 10838 3168 14830 3224
rect 14886 3168 14891 3224
rect 10777 3166 14891 3168
rect 10777 3163 10843 3166
rect 14825 3163 14891 3166
rect 16990 3224 20779 3226
rect 16990 3168 20718 3224
rect 20774 3168 20779 3224
rect 16990 3166 20779 3168
rect 0 3090 120 3120
rect 16990 3090 17050 3166
rect 20713 3163 20779 3166
rect 23749 3090 23815 3093
rect 0 3030 17050 3090
rect 17174 3088 23815 3090
rect 17174 3032 23754 3088
rect 23810 3032 23815 3088
rect 17174 3030 23815 3032
rect 0 3000 120 3030
rect 17174 2954 17234 3030
rect 23749 3027 23815 3030
rect 39389 3090 39455 3093
rect 40880 3090 41000 3120
rect 39389 3088 41000 3090
rect 39389 3032 39394 3088
rect 39450 3032 41000 3088
rect 39389 3030 41000 3032
rect 39389 3027 39455 3030
rect 40880 3000 41000 3030
rect 28073 2954 28139 2957
rect 1718 2894 17234 2954
rect 17358 2952 28139 2954
rect 17358 2896 28078 2952
rect 28134 2896 28139 2952
rect 17358 2894 28139 2896
rect 0 2818 120 2848
rect 1718 2818 1778 2894
rect 0 2758 1778 2818
rect 14825 2818 14891 2821
rect 17358 2818 17418 2894
rect 28073 2891 28139 2894
rect 14825 2816 17418 2818
rect 14825 2760 14830 2816
rect 14886 2760 17418 2816
rect 14825 2758 17418 2760
rect 39021 2818 39087 2821
rect 40880 2818 41000 2848
rect 39021 2816 41000 2818
rect 39021 2760 39026 2816
rect 39082 2760 41000 2816
rect 39021 2758 41000 2760
rect 0 2728 120 2758
rect 14825 2755 14891 2758
rect 39021 2755 39087 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 37946 2752 38262 2753
rect 37946 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38262 2752
rect 40880 2728 41000 2758
rect 37946 2687 38262 2688
rect 0 2546 120 2576
rect 28441 2546 28507 2549
rect 0 2544 28507 2546
rect 0 2488 28446 2544
rect 28502 2488 28507 2544
rect 0 2486 28507 2488
rect 0 2456 120 2486
rect 28441 2483 28507 2486
rect 31569 2546 31635 2549
rect 38469 2546 38535 2549
rect 31569 2544 38535 2546
rect 31569 2488 31574 2544
rect 31630 2488 38474 2544
rect 38530 2488 38535 2544
rect 31569 2486 38535 2488
rect 31569 2483 31635 2486
rect 38469 2483 38535 2486
rect 39389 2546 39455 2549
rect 40880 2546 41000 2576
rect 39389 2544 41000 2546
rect 39389 2488 39394 2544
rect 39450 2488 41000 2544
rect 39389 2486 41000 2488
rect 39389 2483 39455 2486
rect 40880 2456 41000 2486
rect 8845 2410 8911 2413
rect 2822 2408 8911 2410
rect 2822 2352 8850 2408
rect 8906 2352 8911 2408
rect 2822 2350 8911 2352
rect 0 2274 120 2304
rect 2822 2274 2882 2350
rect 8845 2347 8911 2350
rect 32581 2410 32647 2413
rect 38561 2410 38627 2413
rect 32581 2408 38627 2410
rect 32581 2352 32586 2408
rect 32642 2352 38566 2408
rect 38622 2352 38627 2408
rect 32581 2350 38627 2352
rect 32581 2347 32647 2350
rect 38561 2347 38627 2350
rect 0 2214 2882 2274
rect 39941 2274 40007 2277
rect 40880 2274 41000 2304
rect 39941 2272 41000 2274
rect 39941 2216 39946 2272
rect 40002 2216 41000 2272
rect 39941 2214 41000 2216
rect 0 2184 120 2214
rect 39941 2211 40007 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 33006 2143 33322 2144
rect 39006 2208 39322 2209
rect 39006 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39322 2208
rect 40880 2184 41000 2214
rect 39006 2143 39322 2144
rect 0 2002 120 2032
rect 9397 2002 9463 2005
rect 0 2000 9463 2002
rect 0 1944 9402 2000
rect 9458 1944 9463 2000
rect 0 1942 9463 1944
rect 0 1912 120 1942
rect 9397 1939 9463 1942
rect 37917 2002 37983 2005
rect 40880 2002 41000 2032
rect 37917 2000 41000 2002
rect 37917 1944 37922 2000
rect 37978 1944 41000 2000
rect 37917 1942 41000 1944
rect 37917 1939 37983 1942
rect 40880 1912 41000 1942
rect 0 1730 120 1760
rect 9489 1730 9555 1733
rect 0 1728 9555 1730
rect 0 1672 9494 1728
rect 9550 1672 9555 1728
rect 0 1670 9555 1672
rect 0 1640 120 1670
rect 9489 1667 9555 1670
rect 38285 1730 38351 1733
rect 40880 1730 41000 1760
rect 38285 1728 41000 1730
rect 38285 1672 38290 1728
rect 38346 1672 41000 1728
rect 38285 1670 41000 1672
rect 38285 1667 38351 1670
rect 40880 1640 41000 1670
rect 0 1458 120 1488
rect 9581 1458 9647 1461
rect 0 1456 9647 1458
rect 0 1400 9586 1456
rect 9642 1400 9647 1456
rect 0 1398 9647 1400
rect 0 1368 120 1398
rect 9581 1395 9647 1398
rect 38653 1458 38719 1461
rect 40880 1458 41000 1488
rect 38653 1456 41000 1458
rect 38653 1400 38658 1456
rect 38714 1400 41000 1456
rect 38653 1398 41000 1400
rect 38653 1395 38719 1398
rect 40880 1368 41000 1398
rect 8845 98 8911 101
rect 24577 98 24643 101
rect 8845 96 24643 98
rect 8845 40 8850 96
rect 8906 40 24582 96
rect 24638 40 24643 96
rect 8845 38 24643 40
rect 8845 35 8911 38
rect 24577 35 24643 38
<< via3 >>
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 39012 8732 39076 8736
rect 39012 8676 39016 8732
rect 39016 8676 39072 8732
rect 39072 8676 39076 8732
rect 39012 8672 39076 8676
rect 39092 8732 39156 8736
rect 39092 8676 39096 8732
rect 39096 8676 39152 8732
rect 39152 8676 39156 8732
rect 39092 8672 39156 8676
rect 39172 8732 39236 8736
rect 39172 8676 39176 8732
rect 39176 8676 39232 8732
rect 39232 8676 39236 8732
rect 39172 8672 39236 8676
rect 39252 8732 39316 8736
rect 39252 8676 39256 8732
rect 39256 8676 39312 8732
rect 39312 8676 39316 8732
rect 39252 8672 39316 8676
rect 19748 8604 19812 8668
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 37952 8188 38016 8192
rect 37952 8132 37956 8188
rect 37956 8132 38012 8188
rect 38012 8132 38016 8188
rect 37952 8128 38016 8132
rect 38032 8188 38096 8192
rect 38032 8132 38036 8188
rect 38036 8132 38092 8188
rect 38092 8132 38096 8188
rect 38032 8128 38096 8132
rect 38112 8188 38176 8192
rect 38112 8132 38116 8188
rect 38116 8132 38172 8188
rect 38172 8132 38176 8188
rect 38112 8128 38176 8132
rect 38192 8188 38256 8192
rect 38192 8132 38196 8188
rect 38196 8132 38252 8188
rect 38252 8132 38256 8188
rect 38192 8128 38256 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 39012 7644 39076 7648
rect 39012 7588 39016 7644
rect 39016 7588 39072 7644
rect 39072 7588 39076 7644
rect 39012 7584 39076 7588
rect 39092 7644 39156 7648
rect 39092 7588 39096 7644
rect 39096 7588 39152 7644
rect 39152 7588 39156 7644
rect 39092 7584 39156 7588
rect 39172 7644 39236 7648
rect 39172 7588 39176 7644
rect 39176 7588 39232 7644
rect 39232 7588 39236 7644
rect 39172 7584 39236 7588
rect 39252 7644 39316 7648
rect 39252 7588 39256 7644
rect 39256 7588 39312 7644
rect 39312 7588 39316 7644
rect 39252 7584 39316 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 37952 7100 38016 7104
rect 37952 7044 37956 7100
rect 37956 7044 38012 7100
rect 38012 7044 38016 7100
rect 37952 7040 38016 7044
rect 38032 7100 38096 7104
rect 38032 7044 38036 7100
rect 38036 7044 38092 7100
rect 38092 7044 38096 7100
rect 38032 7040 38096 7044
rect 38112 7100 38176 7104
rect 38112 7044 38116 7100
rect 38116 7044 38172 7100
rect 38172 7044 38176 7100
rect 38112 7040 38176 7044
rect 38192 7100 38256 7104
rect 38192 7044 38196 7100
rect 38196 7044 38252 7100
rect 38252 7044 38256 7100
rect 38192 7040 38256 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 39012 6556 39076 6560
rect 39012 6500 39016 6556
rect 39016 6500 39072 6556
rect 39072 6500 39076 6556
rect 39012 6496 39076 6500
rect 39092 6556 39156 6560
rect 39092 6500 39096 6556
rect 39096 6500 39152 6556
rect 39152 6500 39156 6556
rect 39092 6496 39156 6500
rect 39172 6556 39236 6560
rect 39172 6500 39176 6556
rect 39176 6500 39232 6556
rect 39232 6500 39236 6556
rect 39172 6496 39236 6500
rect 39252 6556 39316 6560
rect 39252 6500 39256 6556
rect 39256 6500 39312 6556
rect 39312 6500 39316 6556
rect 39252 6496 39316 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 37952 6012 38016 6016
rect 37952 5956 37956 6012
rect 37956 5956 38012 6012
rect 38012 5956 38016 6012
rect 37952 5952 38016 5956
rect 38032 6012 38096 6016
rect 38032 5956 38036 6012
rect 38036 5956 38092 6012
rect 38092 5956 38096 6012
rect 38032 5952 38096 5956
rect 38112 6012 38176 6016
rect 38112 5956 38116 6012
rect 38116 5956 38172 6012
rect 38172 5956 38176 6012
rect 38112 5952 38176 5956
rect 38192 6012 38256 6016
rect 38192 5956 38196 6012
rect 38196 5956 38252 6012
rect 38252 5956 38256 6012
rect 38192 5952 38256 5956
rect 19748 5536 19812 5540
rect 19748 5480 19762 5536
rect 19762 5480 19812 5536
rect 19748 5476 19812 5480
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 39012 5468 39076 5472
rect 39012 5412 39016 5468
rect 39016 5412 39072 5468
rect 39072 5412 39076 5468
rect 39012 5408 39076 5412
rect 39092 5468 39156 5472
rect 39092 5412 39096 5468
rect 39096 5412 39152 5468
rect 39152 5412 39156 5468
rect 39092 5408 39156 5412
rect 39172 5468 39236 5472
rect 39172 5412 39176 5468
rect 39176 5412 39232 5468
rect 39232 5412 39236 5468
rect 39172 5408 39236 5412
rect 39252 5468 39316 5472
rect 39252 5412 39256 5468
rect 39256 5412 39312 5468
rect 39312 5412 39316 5468
rect 39252 5408 39316 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 37952 4924 38016 4928
rect 37952 4868 37956 4924
rect 37956 4868 38012 4924
rect 38012 4868 38016 4924
rect 37952 4864 38016 4868
rect 38032 4924 38096 4928
rect 38032 4868 38036 4924
rect 38036 4868 38092 4924
rect 38092 4868 38096 4924
rect 38032 4864 38096 4868
rect 38112 4924 38176 4928
rect 38112 4868 38116 4924
rect 38116 4868 38172 4924
rect 38172 4868 38176 4924
rect 38112 4864 38176 4868
rect 38192 4924 38256 4928
rect 38192 4868 38196 4924
rect 38196 4868 38252 4924
rect 38252 4868 38256 4924
rect 38192 4864 38256 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 39012 4380 39076 4384
rect 39012 4324 39016 4380
rect 39016 4324 39072 4380
rect 39072 4324 39076 4380
rect 39012 4320 39076 4324
rect 39092 4380 39156 4384
rect 39092 4324 39096 4380
rect 39096 4324 39152 4380
rect 39152 4324 39156 4380
rect 39092 4320 39156 4324
rect 39172 4380 39236 4384
rect 39172 4324 39176 4380
rect 39176 4324 39232 4380
rect 39232 4324 39236 4380
rect 39172 4320 39236 4324
rect 39252 4380 39316 4384
rect 39252 4324 39256 4380
rect 39256 4324 39312 4380
rect 39312 4324 39316 4380
rect 39252 4320 39316 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 37952 3836 38016 3840
rect 37952 3780 37956 3836
rect 37956 3780 38012 3836
rect 38012 3780 38016 3836
rect 37952 3776 38016 3780
rect 38032 3836 38096 3840
rect 38032 3780 38036 3836
rect 38036 3780 38092 3836
rect 38092 3780 38096 3836
rect 38032 3776 38096 3780
rect 38112 3836 38176 3840
rect 38112 3780 38116 3836
rect 38116 3780 38172 3836
rect 38172 3780 38176 3836
rect 38112 3776 38176 3780
rect 38192 3836 38256 3840
rect 38192 3780 38196 3836
rect 38196 3780 38252 3836
rect 38252 3780 38256 3836
rect 38192 3776 38256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 39012 3292 39076 3296
rect 39012 3236 39016 3292
rect 39016 3236 39072 3292
rect 39072 3236 39076 3292
rect 39012 3232 39076 3236
rect 39092 3292 39156 3296
rect 39092 3236 39096 3292
rect 39096 3236 39152 3292
rect 39152 3236 39156 3292
rect 39092 3232 39156 3236
rect 39172 3292 39236 3296
rect 39172 3236 39176 3292
rect 39176 3236 39232 3292
rect 39232 3236 39236 3292
rect 39172 3232 39236 3236
rect 39252 3292 39316 3296
rect 39252 3236 39256 3292
rect 39256 3236 39312 3292
rect 39312 3236 39316 3292
rect 39252 3232 39316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 37952 2748 38016 2752
rect 37952 2692 37956 2748
rect 37956 2692 38012 2748
rect 38012 2692 38016 2748
rect 37952 2688 38016 2692
rect 38032 2748 38096 2752
rect 38032 2692 38036 2748
rect 38036 2692 38092 2748
rect 38092 2692 38096 2748
rect 38032 2688 38096 2692
rect 38112 2748 38176 2752
rect 38112 2692 38116 2748
rect 38116 2692 38172 2748
rect 38172 2692 38176 2748
rect 38112 2688 38176 2692
rect 38192 2748 38256 2752
rect 38192 2692 38196 2748
rect 38196 2692 38252 2748
rect 38252 2692 38256 2748
rect 38192 2688 38256 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
rect 39012 2204 39076 2208
rect 39012 2148 39016 2204
rect 39016 2148 39072 2204
rect 39072 2148 39076 2204
rect 39012 2144 39076 2148
rect 39092 2204 39156 2208
rect 39092 2148 39096 2204
rect 39096 2148 39152 2204
rect 39152 2148 39156 2204
rect 39092 2144 39156 2148
rect 39172 2204 39236 2208
rect 39172 2148 39176 2204
rect 39176 2148 39232 2204
rect 39232 2148 39236 2204
rect 39172 2144 39236 2148
rect 39252 2204 39316 2208
rect 39252 2148 39256 2204
rect 39256 2148 39312 2204
rect 39312 2148 39316 2204
rect 39252 2144 39316 2148
<< metal4 >>
rect 1944 8192 2264 11250
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 8736 3324 11250
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11250
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 8736 9324 11250
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 8192 14264 11250
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13944 0 14264 2688
rect 15004 8736 15324 11250
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 19747 8668 19813 8669
rect 19747 8604 19748 8668
rect 19812 8604 19813 8668
rect 19747 8603 19813 8604
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 19750 5541 19810 8603
rect 19944 8192 20264 11250
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 19747 5540 19813 5541
rect 19747 5476 19748 5540
rect 19812 5476 19813 5540
rect 19747 5475 19813 5476
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19944 0 20264 2688
rect 21004 8736 21324 11250
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 21004 6560 21324 7584
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25944 8192 26264 11250
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25944 0 26264 2688
rect 27004 8736 27324 11250
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 31944 8192 32264 11250
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 0 32264 2688
rect 33004 8736 33324 11250
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
rect 37944 8192 38264 11250
rect 37944 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38264 8192
rect 37944 7104 38264 8128
rect 37944 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38264 7104
rect 37944 6016 38264 7040
rect 37944 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38264 6016
rect 37944 4928 38264 5952
rect 37944 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38264 4928
rect 37944 3840 38264 4864
rect 37944 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38264 3840
rect 37944 2752 38264 3776
rect 37944 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38264 2752
rect 37944 0 38264 2688
rect 39004 8736 39324 11250
rect 39004 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39324 8736
rect 39004 7648 39324 8672
rect 39004 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39324 7648
rect 39004 6560 39324 7584
rect 39004 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39324 6560
rect 39004 5472 39324 6496
rect 39004 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39324 5472
rect 39004 4384 39324 5408
rect 39004 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39324 4384
rect 39004 3296 39324 4320
rect 39004 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39324 3296
rect 39004 2208 39324 3232
rect 39004 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39324 2208
rect 39004 0 39324 2144
use sky130_fd_sc_hd__buf_1  _001_
timestamp -3599
transform 1 0 13156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _002_
timestamp -3599
transform -1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _003_
timestamp -3599
transform 1 0 16744 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _004_
timestamp -3599
transform 1 0 8740 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _005_
timestamp -3599
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _006_
timestamp -3599
transform 1 0 23920 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _007_
timestamp -3599
transform 1 0 20792 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _008_
timestamp -3599
transform 1 0 23184 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _009_
timestamp -3599
transform 1 0 9660 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _010_
timestamp -3599
transform 1 0 20424 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _011_
timestamp -3599
transform 1 0 18492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _012_
timestamp -3599
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _013_
timestamp -3599
transform 1 0 13616 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _014_
timestamp -3599
transform 1 0 5612 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _015_
timestamp -3599
transform 1 0 10856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _016_
timestamp -3599
transform 1 0 14904 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _017_
timestamp -3599
transform 1 0 21344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _018_
timestamp -3599
transform 1 0 11132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _019_
timestamp -3599
transform 1 0 19320 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _020_
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _021_
timestamp -3599
transform 1 0 16468 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _022_
timestamp -3599
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _023_
timestamp -3599
transform 1 0 18216 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _024_
timestamp -3599
transform 1 0 24196 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _025_
timestamp -3599
transform 1 0 23552 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _026_
timestamp -3599
transform 1 0 24196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _027_
timestamp -3599
transform 1 0 21160 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _028_
timestamp -3599
transform 1 0 21988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _029_
timestamp -3599
transform 1 0 15272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _030_
timestamp -3599
transform 1 0 17664 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _031_
timestamp -3599
transform 1 0 27692 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _032_
timestamp -3599
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _033_
timestamp -3599
transform -1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _034_
timestamp -3599
transform 1 0 22448 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _035_
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _036_
timestamp -3599
transform 1 0 24748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp -3599
transform -1 0 28336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _038_
timestamp -3599
transform -1 0 30452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _039_
timestamp -3599
transform -1 0 33764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp -3599
transform 1 0 36248 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp -3599
transform 1 0 36984 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp -3599
transform -1 0 35512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp -3599
transform -1 0 30176 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _044_
timestamp -3599
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _045_
timestamp -3599
transform 1 0 17848 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _046_
timestamp -3599
transform 1 0 23920 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp -3599
transform -1 0 28428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp -3599
transform -1 0 30544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp -3599
transform -1 0 32108 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp -3599
transform -1 0 33856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp -3599
transform -1 0 35880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _052_
timestamp -3599
transform 1 0 38088 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _053_
timestamp -3599
transform -1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _054_
timestamp -3599
transform -1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _055_
timestamp -3599
transform -1 0 3312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp -3599
transform -1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp -3599
transform -1 0 3680 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp -3599
transform 1 0 4416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp -3599
transform 1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp -3599
transform 1 0 5336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp -3599
transform 1 0 5520 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp -3599
transform 1 0 6624 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp -3599
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp -3599
transform 1 0 11592 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp -3599
transform -1 0 5888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp -3599
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp -3599
transform 1 0 7636 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp -3599
transform 1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp -3599
transform 1 0 9384 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp -3599
transform 1 0 10580 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp -3599
transform 1 0 12972 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _072_
timestamp -3599
transform -1 0 17664 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp -3599
transform 1 0 12236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _074_
timestamp -3599
transform -1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp -3599
transform 1 0 14444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp -3599
transform 1 0 9568 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp -3599
transform -1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp -3599
transform -1 0 9568 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp -3599
transform 1 0 11592 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp -3599
transform 1 0 14628 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp -3599
transform 1 0 15824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp -3599
transform 1 0 17112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp -3599
transform 1 0 15824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp -3599
transform 1 0 13248 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp -3599
transform 1 0 14168 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp -3599
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp -3599
transform 1 0 17572 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp -3599
transform 1 0 19688 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _089_
timestamp -3599
transform -1 0 35604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _090_
timestamp -3599
transform -1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _091_
timestamp -3599
transform -1 0 33304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _092_
timestamp -3599
transform -1 0 31280 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _093_
timestamp -3599
transform -1 0 31280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _094_
timestamp -3599
transform -1 0 30084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _095_
timestamp -3599
transform -1 0 29532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _096_
timestamp -3599
transform -1 0 28336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _097_
timestamp -3599
transform -1 0 27232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _098_
timestamp -3599
transform -1 0 26680 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp -3599
transform 1 0 25392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp -3599
transform 1 0 23460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp -3599
transform 1 0 23092 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp -3599
transform 1 0 23736 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp -3599
transform 1 0 21160 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp -3599
transform -1 0 7912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp -3599
transform 1 0 25852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform 1 0 12972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform -1 0 18492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform -1 0 18860 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform 1 0 14720 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform 1 0 10948 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform -1 0 19320 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 17112 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform 1 0 15824 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform 1 0 16284 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform -1 0 18216 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform 1 0 20976 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform 1 0 21804 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform 1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform -1 0 17664 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform -1 0 17204 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform 1 0 27508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp -3599
transform -1 0 19688 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp -3599
transform 1 0 28428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp -3599
transform 1 0 23736 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp -3599
transform -1 0 20792 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp -3599
transform 1 0 23000 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp -3599
transform 1 0 20240 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp -3599
transform 1 0 24564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp -3599
transform 1 0 29992 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp -3599
transform 1 0 33304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp -3599
transform 1 0 4048 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp -3599
transform -1 0 3036 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp -3599
transform -1 0 9384 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp -3599
transform -1 0 8280 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp -3599
transform -1 0 3864 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp -3599
transform -1 0 7912 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp -3599
transform -1 0 14904 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp -3599
transform -1 0 12236 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp -3599
transform -1 0 14168 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp -3599
transform -1 0 2668 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636964856
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636964856
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636964856
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636964856
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636964856
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636964856
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636964856
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636964856
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -3599
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636964856
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636964856
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -3599
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636964856
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636964856
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -3599
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636964856
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636964856
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp -3599
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636964856
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636964856
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -3599
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636964856
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636964856
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -3599
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636964856
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636964856
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -3599
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636964856
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636964856
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -3599
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636964856
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1636964856
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp -3599
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1636964856
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1636964856
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp -3599
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1636964856
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1636964856
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp -3599
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_393
timestamp -3599
transform 1 0 37260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_397
timestamp -3599
transform 1 0 37628 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636964856
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636964856
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636964856
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636964856
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp -3599
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -3599
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636964856
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636964856
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_81
timestamp -3599
transform 1 0 8556 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_87
timestamp 1636964856
transform 1 0 9108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_99
timestamp 1636964856
transform 1 0 10212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -3599
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636964856
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp -3599
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_134
timestamp 1636964856
transform 1 0 13432 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_146
timestamp 1636964856
transform 1 0 14536 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_158
timestamp -3599
transform 1 0 15640 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp -3599
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp -3599
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_175
timestamp -3599
transform 1 0 17204 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_183
timestamp -3599
transform 1 0 17940 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_189
timestamp 1636964856
transform 1 0 18492 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_201
timestamp -3599
transform 1 0 19596 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_209
timestamp -3599
transform 1 0 20332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_217
timestamp -3599
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp -3599
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636964856
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_237
timestamp -3599
transform 1 0 22908 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_245
timestamp -3599
transform 1 0 23644 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_254
timestamp -3599
transform 1 0 24472 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_260
timestamp 1636964856
transform 1 0 25024 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_272
timestamp -3599
transform 1 0 26128 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_284
timestamp -3599
transform 1 0 27232 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_292
timestamp -3599
transform 1 0 27968 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_296
timestamp -3599
transform 1 0 28336 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_302
timestamp 1636964856
transform 1 0 28888 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_319
timestamp 1636964856
transform 1 0 30452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp -3599
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp -3599
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636964856
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_349
timestamp -3599
transform 1 0 33212 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_355
timestamp 1636964856
transform 1 0 33764 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_367
timestamp 1636964856
transform 1 0 34868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_379
timestamp 1636964856
transform 1 0 35972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp -3599
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636964856
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_405
timestamp -3599
transform 1 0 38364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_409
timestamp -3599
transform 1 0 38732 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636964856
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636964856
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636964856
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636964856
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636964856
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636964856
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636964856
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_97
timestamp -3599
transform 1 0 10028 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_105
timestamp -3599
transform 1 0 10764 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_110
timestamp 1636964856
transform 1 0 11224 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_122
timestamp 1636964856
transform 1 0 12328 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_134
timestamp -3599
transform 1 0 13432 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_141
timestamp -3599
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_147
timestamp -3599
transform 1 0 14628 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636964856
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636964856
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_180
timestamp 1636964856
transform 1 0 17664 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp -3599
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_197
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_205
timestamp -3599
transform 1 0 19964 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_213
timestamp 1636964856
transform 1 0 20700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_225
timestamp 1636964856
transform 1 0 21804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_237
timestamp 1636964856
transform 1 0 22908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp -3599
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636964856
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636964856
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636964856
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636964856
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp -3599
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp -3599
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_309
timestamp -3599
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_316
timestamp 1636964856
transform 1 0 30176 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_328
timestamp 1636964856
transform 1 0 31280 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_340
timestamp 1636964856
transform 1 0 32384 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_352
timestamp 1636964856
transform 1 0 33488 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636964856
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636964856
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636964856
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_401
timestamp -3599
transform 1 0 37996 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_409
timestamp -3599
transform 1 0 38732 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636964856
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636964856
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636964856
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_39
timestamp -3599
transform 1 0 4692 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_47
timestamp -3599
transform 1 0 5428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp -3599
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636964856
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636964856
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636964856
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_97
timestamp 1636964856
transform 1 0 10028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp -3599
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636964856
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_125
timestamp -3599
transform 1 0 12604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_133
timestamp -3599
transform 1 0 13340 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_139
timestamp 1636964856
transform 1 0 13892 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_151
timestamp 1636964856
transform 1 0 14996 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp -3599
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -3599
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636964856
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636964856
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636964856
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636964856
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp -3599
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp -3599
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636964856
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_237
timestamp -3599
transform 1 0 22908 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_243
timestamp 1636964856
transform 1 0 23460 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_255
timestamp 1636964856
transform 1 0 24564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_267
timestamp 1636964856
transform 1 0 25668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp -3599
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636964856
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636964856
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636964856
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_320
timestamp 1636964856
transform 1 0 30544 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_332
timestamp -3599
transform 1 0 31648 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636964856
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636964856
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636964856
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_373
timestamp -3599
transform 1 0 35420 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_381
timestamp -3599
transform 1 0 36156 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp -3599
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp -3599
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636964856
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_405
timestamp -3599
transform 1 0 38364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_409
timestamp -3599
transform 1 0 38732 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636964856
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636964856
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636964856
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636964856
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636964856
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636964856
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp -3599
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -3599
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636964856
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_97
timestamp -3599
transform 1 0 10028 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_105
timestamp -3599
transform 1 0 10764 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_113
timestamp 1636964856
transform 1 0 11500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_125
timestamp 1636964856
transform 1 0 12604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp -3599
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_141
timestamp -3599
transform 1 0 14076 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_150
timestamp 1636964856
transform 1 0 14904 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_162
timestamp -3599
transform 1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_170
timestamp 1636964856
transform 1 0 16744 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_182
timestamp -3599
transform 1 0 17848 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_190
timestamp -3599
transform 1 0 18584 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636964856
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_212
timestamp 1636964856
transform 1 0 20608 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_224
timestamp 1636964856
transform 1 0 21712 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_236
timestamp -3599
transform 1 0 22816 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_247
timestamp -3599
transform 1 0 23828 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp -3599
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636964856
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636964856
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636964856
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_289
timestamp -3599
transform 1 0 27692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_293
timestamp -3599
transform 1 0 28060 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_297
timestamp -3599
transform 1 0 28428 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp -3599
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636964856
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636964856
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_333
timestamp -3599
transform 1 0 31740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_337
timestamp 1636964856
transform 1 0 32108 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_349
timestamp -3599
transform 1 0 33212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_356
timestamp -3599
transform 1 0 33856 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636964856
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636964856
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1636964856
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_401
timestamp -3599
transform 1 0 37996 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_409
timestamp -3599
transform 1 0 38732 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636964856
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636964856
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636964856
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_39
timestamp -3599
transform 1 0 4692 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_45
timestamp -3599
transform 1 0 5244 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp -3599
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636964856
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636964856
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636964856
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636964856
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp -3599
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp -3599
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636964856
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_125
timestamp -3599
transform 1 0 12604 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_132
timestamp 1636964856
transform 1 0 13248 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_144
timestamp 1636964856
transform 1 0 14352 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_156
timestamp -3599
transform 1 0 15456 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_163
timestamp -3599
transform 1 0 16100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp -3599
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_177
timestamp -3599
transform 1 0 17388 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_181
timestamp -3599
transform 1 0 17756 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_185
timestamp 1636964856
transform 1 0 18124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_197
timestamp 1636964856
transform 1 0 19228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_209
timestamp 1636964856
transform 1 0 20332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_221
timestamp -3599
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_228
timestamp 1636964856
transform 1 0 22080 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_240
timestamp 1636964856
transform 1 0 23184 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_252
timestamp 1636964856
transform 1 0 24288 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_264
timestamp 1636964856
transform 1 0 25392 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp -3599
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_284
timestamp 1636964856
transform 1 0 27232 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_296
timestamp 1636964856
transform 1 0 28336 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_308
timestamp 1636964856
transform 1 0 29440 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_320
timestamp 1636964856
transform 1 0 30544 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp -3599
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636964856
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636964856
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636964856
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636964856
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp -3599
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp -3599
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636964856
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_405
timestamp -3599
transform 1 0 38364 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_409
timestamp -3599
transform 1 0 38732 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636964856
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636964856
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_34
timestamp -3599
transform 1 0 4232 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_40
timestamp -3599
transform 1 0 4784 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_44
timestamp -3599
transform 1 0 5152 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_51
timestamp -3599
transform 1 0 5796 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_59
timestamp -3599
transform 1 0 6532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_63
timestamp -3599
transform 1 0 6900 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_68
timestamp 1636964856
transform 1 0 7360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp -3599
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636964856
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636964856
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_109
timestamp -3599
transform 1 0 11132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_113
timestamp -3599
transform 1 0 11500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_117
timestamp 1636964856
transform 1 0 11868 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_129
timestamp -3599
transform 1 0 12972 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_137
timestamp -3599
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636964856
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636964856
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636964856
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_177
timestamp -3599
transform 1 0 17388 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_185
timestamp -3599
transform 1 0 18124 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp -3599
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636964856
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636964856
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1636964856
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1636964856
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp -3599
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp -3599
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636964856
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_265
timestamp -3599
transform 1 0 25484 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_273
timestamp 1636964856
transform 1 0 26220 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_285
timestamp -3599
transform 1 0 27324 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_296
timestamp 1636964856
transform 1 0 28336 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636964856
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1636964856
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1636964856
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1636964856
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp -3599
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp -3599
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_365
timestamp -3599
transform 1 0 34684 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_374
timestamp -3599
transform 1 0 35512 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_378
timestamp 1636964856
transform 1 0 35880 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_393
timestamp -3599
transform 1 0 37260 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_401
timestamp -3599
transform 1 0 37996 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_405
timestamp -3599
transform 1 0 38364 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_409
timestamp -3599
transform 1 0 38732 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636964856
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_15
timestamp -3599
transform 1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_24
timestamp -3599
transform 1 0 3312 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_30
timestamp -3599
transform 1 0 3864 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636964856
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp -3599
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -3599
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636964856
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_69
timestamp -3599
transform 1 0 7452 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_74
timestamp -3599
transform 1 0 7912 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_84
timestamp 1636964856
transform 1 0 8832 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_96
timestamp -3599
transform 1 0 9936 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_102
timestamp -3599
transform 1 0 10488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_106
timestamp -3599
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp -3599
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_117
timestamp 1636964856
transform 1 0 11868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_129
timestamp 1636964856
transform 1 0 12972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_141
timestamp 1636964856
transform 1 0 14076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_153
timestamp 1636964856
transform 1 0 15180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp -3599
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636964856
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636964856
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_193
timestamp -3599
transform 1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_201
timestamp 1636964856
transform 1 0 19596 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_213
timestamp -3599
transform 1 0 20700 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_221
timestamp -3599
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636964856
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636964856
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_249
timestamp -3599
transform 1 0 24012 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_254
timestamp 1636964856
transform 1 0 24472 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_266
timestamp -3599
transform 1 0 25576 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_274
timestamp -3599
transform 1 0 26312 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp -3599
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636964856
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1636964856
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_305
timestamp -3599
transform 1 0 29164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_309
timestamp 1636964856
transform 1 0 29532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_321
timestamp 1636964856
transform 1 0 30636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_333
timestamp -3599
transform 1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1636964856
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1636964856
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1636964856
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1636964856
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp -3599
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp -3599
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1636964856
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_405
timestamp -3599
transform 1 0 38364 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_409
timestamp -3599
transform 1 0 38732 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636964856
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp -3599
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636964856
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636964856
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636964856
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636964856
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp -3599
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp -3599
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_93
timestamp 1636964856
transform 1 0 9660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_105
timestamp 1636964856
transform 1 0 10764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_117
timestamp 1636964856
transform 1 0 11868 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_129
timestamp -3599
transform 1 0 12972 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp -3599
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636964856
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636964856
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636964856
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1636964856
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp -3599
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp -3599
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636964856
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636964856
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_221
timestamp -3599
transform 1 0 21436 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_229
timestamp -3599
transform 1 0 22172 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_235
timestamp 1636964856
transform 1 0 22724 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_247
timestamp -3599
transform 1 0 23828 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp -3599
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_253
timestamp -3599
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_261
timestamp -3599
transform 1 0 25116 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_267
timestamp 1636964856
transform 1 0 25668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_279
timestamp 1636964856
transform 1 0 26772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_291
timestamp 1636964856
transform 1 0 27876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_303
timestamp -3599
transform 1 0 28980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp -3599
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_309
timestamp -3599
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_315
timestamp 1636964856
transform 1 0 30084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_327
timestamp 1636964856
transform 1 0 31188 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_339
timestamp 1636964856
transform 1 0 32292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_351
timestamp -3599
transform 1 0 33396 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_357
timestamp -3599
transform 1 0 33948 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_361
timestamp -3599
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1636964856
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1636964856
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1636964856
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_401
timestamp -3599
transform 1 0 37996 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_405
timestamp -3599
transform 1 0 38364 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636964856
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_15
timestamp -3599
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_19
timestamp 1636964856
transform 1 0 2852 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_31
timestamp 1636964856
transform 1 0 3956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_43
timestamp 1636964856
transform 1 0 5060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -3599
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636964856
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_69
timestamp -3599
transform 1 0 7452 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_74
timestamp 1636964856
transform 1 0 7912 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_86
timestamp -3599
transform 1 0 9016 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_95
timestamp 1636964856
transform 1 0 9844 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_107
timestamp -3599
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp -3599
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636964856
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1636964856
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_137
timestamp -3599
transform 1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_150
timestamp -3599
transform 1 0 14904 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_158
timestamp -3599
transform 1 0 15640 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp -3599
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp -3599
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_169
timestamp -3599
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_177
timestamp -3599
transform 1 0 17388 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_183
timestamp 1636964856
transform 1 0 17940 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_195
timestamp 1636964856
transform 1 0 19044 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_207
timestamp -3599
transform 1 0 20148 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_215
timestamp -3599
transform 1 0 20884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp -3599
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1636964856
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_237
timestamp -3599
transform 1 0 22908 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_245
timestamp -3599
transform 1 0 23644 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1636964856
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1636964856
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp -3599
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp -3599
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636964856
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1636964856
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1636964856
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_317
timestamp -3599
transform 1 0 30268 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_328
timestamp -3599
transform 1 0 31280 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1636964856
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1636964856
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1636964856
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1636964856
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp -3599
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp -3599
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_393
timestamp -3599
transform 1 0 37260 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_397
timestamp -3599
transform 1 0 37628 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636964856
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_15
timestamp -3599
transform 1 0 2484 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_23
timestamp -3599
transform 1 0 3220 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_37
timestamp -3599
transform 1 0 4508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_41
timestamp -3599
transform 1 0 4876 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_46
timestamp -3599
transform 1 0 5336 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_58
timestamp -3599
transform 1 0 6440 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_64
timestamp -3599
transform 1 0 6992 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_70
timestamp -3599
transform 1 0 7544 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_77
timestamp -3599
transform 1 0 8188 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp -3599
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_89
timestamp -3599
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_97
timestamp -3599
transform 1 0 10028 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_101
timestamp -3599
transform 1 0 10396 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_106
timestamp -3599
transform 1 0 10856 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_110
timestamp -3599
transform 1 0 11224 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_124
timestamp -3599
transform 1 0 12512 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_130
timestamp -3599
transform 1 0 13064 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp -3599
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_148
timestamp -3599
transform 1 0 14720 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_161
timestamp -3599
transform 1 0 15916 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_166
timestamp 1636964856
transform 1 0 16376 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_178
timestamp -3599
transform 1 0 17480 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_182
timestamp 1636964856
transform 1 0 17848 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp -3599
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_205
timestamp -3599
transform 1 0 19964 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_213
timestamp -3599
transform 1 0 20700 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_221
timestamp -3599
transform 1 0 21436 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_230
timestamp -3599
transform 1 0 22264 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_238
timestamp -3599
transform 1 0 23000 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_242
timestamp -3599
transform 1 0 23368 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_246
timestamp -3599
transform 1 0 23736 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1636964856
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1636964856
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_277
timestamp -3599
transform 1 0 26588 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_285
timestamp -3599
transform 1 0 27324 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_292
timestamp 1636964856
transform 1 0 27968 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp -3599
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1636964856
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_321
timestamp -3599
transform 1 0 30636 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_328
timestamp 1636964856
transform 1 0 31280 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_340
timestamp -3599
transform 1 0 32384 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_346
timestamp -3599
transform 1 0 32936 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_350
timestamp 1636964856
transform 1 0 33304 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp -3599
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_369
timestamp -3599
transform 1 0 35052 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_379
timestamp -3599
transform 1 0 35972 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_385
timestamp -3599
transform 1 0 36524 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_391
timestamp -3599
transform 1 0 37076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_403
timestamp -3599
transform 1 0 38180 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636964856
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp -3599
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_19
timestamp -3599
transform 1 0 2852 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_29
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp -3599
transform 1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_141
timestamp -3599
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp -3599
transform 1 0 17204 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_188
timestamp -3599
transform 1 0 18400 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_197
timestamp 1636964856
transform 1 0 19228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_209
timestamp 1636964856
transform 1 0 20332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp -3599
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1636964856
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1636964856
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_249
timestamp -3599
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_253
timestamp 1636964856
transform 1 0 24380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_265
timestamp 1636964856
transform 1 0 25484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp -3599
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1636964856
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1636964856
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_305
timestamp -3599
transform 1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_309
timestamp 1636964856
transform 1 0 29532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_321
timestamp 1636964856
transform 1 0 30636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp -3599
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp -3599
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_362
timestamp -3599
transform 1 0 34408 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp -3599
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_409
timestamp -3599
transform 1 0 38732 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output1
timestamp -3599
transform 1 0 38456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform 1 0 39192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform 1 0 38824 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform 1 0 39192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform 1 0 38824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform 1 0 39192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 38824 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform 1 0 39192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 38824 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -3599
transform 1 0 38456 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -3599
transform 1 0 39192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -3599
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp -3599
transform 1 0 37720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp -3599
transform 1 0 39192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp -3599
transform 1 0 38824 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp -3599
transform 1 0 39192 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp -3599
transform 1 0 39192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -3599
transform 1 0 38824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp -3599
transform 1 0 38456 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp -3599
transform 1 0 38824 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp -3599
transform 1 0 39192 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp -3599
transform 1 0 38456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp -3599
transform 1 0 37720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp -3599
transform 1 0 38824 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp -3599
transform 1 0 38088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp -3599
transform 1 0 38824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp -3599
transform 1 0 39192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp -3599
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp -3599
transform 1 0 39192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp -3599
transform 1 0 38824 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp -3599
transform 1 0 39192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp -3599
transform 1 0 38824 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp -3599
transform 1 0 32568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp -3599
transform 1 0 36156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp -3599
transform 1 0 35604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp -3599
transform 1 0 36524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp -3599
transform 1 0 36156 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp -3599
transform 1 0 37260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp -3599
transform 1 0 36708 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp -3599
transform 1 0 37628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp -3599
transform 1 0 37996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp -3599
transform 1 0 38364 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp -3599
transform -1 0 38180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp -3599
transform 1 0 32936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp -3599
transform 1 0 33304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp -3599
transform 1 0 33672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp -3599
transform 1 0 34040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp -3599
transform 1 0 34684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp -3599
transform 1 0 35052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp -3599
transform -1 0 35052 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp -3599
transform -1 0 35788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp -3599
transform 1 0 35788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp -3599
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp -3599
transform 1 0 2944 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp -3599
transform 1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp -3599
transform 1 0 4140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp -3599
transform 1 0 4048 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp -3599
transform 1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp -3599
transform 1 0 4968 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp -3599
transform -1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp -3599
transform -1 0 5520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp -3599
transform -1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp -3599
transform -1 0 6440 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp -3599
transform -1 0 6256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp -3599
transform 1 0 6624 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp -3599
transform -1 0 6992 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp -3599
transform -1 0 7544 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp -3599
transform -1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp -3599
transform -1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp -3599
transform -1 0 8096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp -3599
transform -1 0 8648 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp -3599
transform -1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp -3599
transform -1 0 9292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp -3599
transform -1 0 11408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp -3599
transform -1 0 12052 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp -3599
transform -1 0 12144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform -1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform -1 0 13064 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform -1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform -1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform -1 0 9752 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform -1 0 9568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform 1 0 9568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform 1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform -1 0 10856 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform -1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform -1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform -1 0 11684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform -1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform -1 0 16376 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform -1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform -1 0 16560 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform -1 0 17204 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform -1 0 18124 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform 1 0 17388 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform -1 0 13892 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform -1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform -1 0 13984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform -1 0 14720 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform -1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform -1 0 15916 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform -1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform -1 0 15456 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform -1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output105
timestamp -3599
transform -1 0 32568 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 39836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 39836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 39836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 39836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 39836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 39836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 39836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 39836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 39836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 39836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  S_term_single_106
timestamp -3599
transform -1 0 18400 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_38
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -3599
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_45
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_48
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_49
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_50
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -3599
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_52
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_53
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_54
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_55
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_56
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_57
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_58
timestamp -3599
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_59
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_60
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_61
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_62
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_63
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_65
timestamp -3599
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_66
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_67
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_68
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_69
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_70
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_71
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp -3599
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_73
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_74
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_75
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_76
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp -3599
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_83
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_84
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_85
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp -3599
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_87
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_88
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_92
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_93
timestamp -3599
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_95
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_96
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_97
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_98
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_99
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_100
timestamp -3599
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_101
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_102
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_103
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_104
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_105
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp -3599
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_108
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_109
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_110
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_111
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_112
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_113
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_114
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_115
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_116
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_117
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_118
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_119
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp -3599
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_121
timestamp -3599
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 17590 11194 17646 11250 0 FreeSans 224 0 0 0 Co
port 0 nsew signal output
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[0]
port 1 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[10]
port 2 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[11]
port 3 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[12]
port 4 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[13]
port 5 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[14]
port 6 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[15]
port 7 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[16]
port 8 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[17]
port 9 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[18]
port 10 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[19]
port 11 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[1]
port 12 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[20]
port 13 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[21]
port 14 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[22]
port 15 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[23]
port 16 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[24]
port 17 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[25]
port 18 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[26]
port 19 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[27]
port 20 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[28]
port 21 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[29]
port 22 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[2]
port 23 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[30]
port 24 nsew signal input
flabel metal3 s 0 9800 120 9920 0 FreeSans 480 0 0 0 FrameData[31]
port 25 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[3]
port 26 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[4]
port 27 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[5]
port 28 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[6]
port 29 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[7]
port 30 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[8]
port 31 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[9]
port 32 nsew signal input
flabel metal3 s 40880 1368 41000 1488 0 FreeSans 480 0 0 0 FrameData_O[0]
port 33 nsew signal output
flabel metal3 s 40880 4088 41000 4208 0 FreeSans 480 0 0 0 FrameData_O[10]
port 34 nsew signal output
flabel metal3 s 40880 4360 41000 4480 0 FreeSans 480 0 0 0 FrameData_O[11]
port 35 nsew signal output
flabel metal3 s 40880 4632 41000 4752 0 FreeSans 480 0 0 0 FrameData_O[12]
port 36 nsew signal output
flabel metal3 s 40880 4904 41000 5024 0 FreeSans 480 0 0 0 FrameData_O[13]
port 37 nsew signal output
flabel metal3 s 40880 5176 41000 5296 0 FreeSans 480 0 0 0 FrameData_O[14]
port 38 nsew signal output
flabel metal3 s 40880 5448 41000 5568 0 FreeSans 480 0 0 0 FrameData_O[15]
port 39 nsew signal output
flabel metal3 s 40880 5720 41000 5840 0 FreeSans 480 0 0 0 FrameData_O[16]
port 40 nsew signal output
flabel metal3 s 40880 5992 41000 6112 0 FreeSans 480 0 0 0 FrameData_O[17]
port 41 nsew signal output
flabel metal3 s 40880 6264 41000 6384 0 FreeSans 480 0 0 0 FrameData_O[18]
port 42 nsew signal output
flabel metal3 s 40880 6536 41000 6656 0 FreeSans 480 0 0 0 FrameData_O[19]
port 43 nsew signal output
flabel metal3 s 40880 1640 41000 1760 0 FreeSans 480 0 0 0 FrameData_O[1]
port 44 nsew signal output
flabel metal3 s 40880 6808 41000 6928 0 FreeSans 480 0 0 0 FrameData_O[20]
port 45 nsew signal output
flabel metal3 s 40880 7080 41000 7200 0 FreeSans 480 0 0 0 FrameData_O[21]
port 46 nsew signal output
flabel metal3 s 40880 7352 41000 7472 0 FreeSans 480 0 0 0 FrameData_O[22]
port 47 nsew signal output
flabel metal3 s 40880 7624 41000 7744 0 FreeSans 480 0 0 0 FrameData_O[23]
port 48 nsew signal output
flabel metal3 s 40880 7896 41000 8016 0 FreeSans 480 0 0 0 FrameData_O[24]
port 49 nsew signal output
flabel metal3 s 40880 8168 41000 8288 0 FreeSans 480 0 0 0 FrameData_O[25]
port 50 nsew signal output
flabel metal3 s 40880 8440 41000 8560 0 FreeSans 480 0 0 0 FrameData_O[26]
port 51 nsew signal output
flabel metal3 s 40880 8712 41000 8832 0 FreeSans 480 0 0 0 FrameData_O[27]
port 52 nsew signal output
flabel metal3 s 40880 8984 41000 9104 0 FreeSans 480 0 0 0 FrameData_O[28]
port 53 nsew signal output
flabel metal3 s 40880 9256 41000 9376 0 FreeSans 480 0 0 0 FrameData_O[29]
port 54 nsew signal output
flabel metal3 s 40880 1912 41000 2032 0 FreeSans 480 0 0 0 FrameData_O[2]
port 55 nsew signal output
flabel metal3 s 40880 9528 41000 9648 0 FreeSans 480 0 0 0 FrameData_O[30]
port 56 nsew signal output
flabel metal3 s 40880 9800 41000 9920 0 FreeSans 480 0 0 0 FrameData_O[31]
port 57 nsew signal output
flabel metal3 s 40880 2184 41000 2304 0 FreeSans 480 0 0 0 FrameData_O[3]
port 58 nsew signal output
flabel metal3 s 40880 2456 41000 2576 0 FreeSans 480 0 0 0 FrameData_O[4]
port 59 nsew signal output
flabel metal3 s 40880 2728 41000 2848 0 FreeSans 480 0 0 0 FrameData_O[5]
port 60 nsew signal output
flabel metal3 s 40880 3000 41000 3120 0 FreeSans 480 0 0 0 FrameData_O[6]
port 61 nsew signal output
flabel metal3 s 40880 3272 41000 3392 0 FreeSans 480 0 0 0 FrameData_O[7]
port 62 nsew signal output
flabel metal3 s 40880 3544 41000 3664 0 FreeSans 480 0 0 0 FrameData_O[8]
port 63 nsew signal output
flabel metal3 s 40880 3816 41000 3936 0 FreeSans 480 0 0 0 FrameData_O[9]
port 64 nsew signal output
flabel metal2 s 3054 0 3110 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 65 nsew signal input
flabel metal2 s 22374 0 22430 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 66 nsew signal input
flabel metal2 s 24306 0 24362 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 67 nsew signal input
flabel metal2 s 26238 0 26294 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 68 nsew signal input
flabel metal2 s 28170 0 28226 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 69 nsew signal input
flabel metal2 s 30102 0 30158 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 70 nsew signal input
flabel metal2 s 32034 0 32090 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 71 nsew signal input
flabel metal2 s 33966 0 34022 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 72 nsew signal input
flabel metal2 s 35898 0 35954 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 73 nsew signal input
flabel metal2 s 37830 0 37886 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 74 nsew signal input
flabel metal2 s 39762 0 39818 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 75 nsew signal input
flabel metal2 s 4986 0 5042 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 76 nsew signal input
flabel metal2 s 6918 0 6974 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 77 nsew signal input
flabel metal2 s 8850 0 8906 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 78 nsew signal input
flabel metal2 s 10782 0 10838 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 79 nsew signal input
flabel metal2 s 12714 0 12770 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 80 nsew signal input
flabel metal2 s 14646 0 14702 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 81 nsew signal input
flabel metal2 s 16578 0 16634 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 82 nsew signal input
flabel metal2 s 18510 0 18566 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 83 nsew signal input
flabel metal2 s 20442 0 20498 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 84 nsew signal input
flabel metal2 s 32494 11194 32550 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 85 nsew signal output
flabel metal2 s 35254 11194 35310 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 86 nsew signal output
flabel metal2 s 35530 11194 35586 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 87 nsew signal output
flabel metal2 s 35806 11194 35862 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 88 nsew signal output
flabel metal2 s 36082 11194 36138 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 89 nsew signal output
flabel metal2 s 36358 11194 36414 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 90 nsew signal output
flabel metal2 s 36634 11194 36690 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 91 nsew signal output
flabel metal2 s 36910 11194 36966 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 92 nsew signal output
flabel metal2 s 37186 11194 37242 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 93 nsew signal output
flabel metal2 s 37462 11194 37518 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 94 nsew signal output
flabel metal2 s 37738 11194 37794 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 95 nsew signal output
flabel metal2 s 32770 11194 32826 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 96 nsew signal output
flabel metal2 s 33046 11194 33102 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 97 nsew signal output
flabel metal2 s 33322 11194 33378 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 98 nsew signal output
flabel metal2 s 33598 11194 33654 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 99 nsew signal output
flabel metal2 s 33874 11194 33930 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 100 nsew signal output
flabel metal2 s 34150 11194 34206 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 101 nsew signal output
flabel metal2 s 34426 11194 34482 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 102 nsew signal output
flabel metal2 s 34702 11194 34758 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 103 nsew signal output
flabel metal2 s 34978 11194 35034 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 104 nsew signal output
flabel metal2 s 3238 11194 3294 11250 0 FreeSans 224 0 0 0 N1BEG[0]
port 105 nsew signal output
flabel metal2 s 3514 11194 3570 11250 0 FreeSans 224 0 0 0 N1BEG[1]
port 106 nsew signal output
flabel metal2 s 3790 11194 3846 11250 0 FreeSans 224 0 0 0 N1BEG[2]
port 107 nsew signal output
flabel metal2 s 4066 11194 4122 11250 0 FreeSans 224 0 0 0 N1BEG[3]
port 108 nsew signal output
flabel metal2 s 4342 11194 4398 11250 0 FreeSans 224 0 0 0 N2BEG[0]
port 109 nsew signal output
flabel metal2 s 4618 11194 4674 11250 0 FreeSans 224 0 0 0 N2BEG[1]
port 110 nsew signal output
flabel metal2 s 4894 11194 4950 11250 0 FreeSans 224 0 0 0 N2BEG[2]
port 111 nsew signal output
flabel metal2 s 5170 11194 5226 11250 0 FreeSans 224 0 0 0 N2BEG[3]
port 112 nsew signal output
flabel metal2 s 5446 11194 5502 11250 0 FreeSans 224 0 0 0 N2BEG[4]
port 113 nsew signal output
flabel metal2 s 5722 11194 5778 11250 0 FreeSans 224 0 0 0 N2BEG[5]
port 114 nsew signal output
flabel metal2 s 5998 11194 6054 11250 0 FreeSans 224 0 0 0 N2BEG[6]
port 115 nsew signal output
flabel metal2 s 6274 11194 6330 11250 0 FreeSans 224 0 0 0 N2BEG[7]
port 116 nsew signal output
flabel metal2 s 6550 11194 6606 11250 0 FreeSans 224 0 0 0 N2BEGb[0]
port 117 nsew signal output
flabel metal2 s 6826 11194 6882 11250 0 FreeSans 224 0 0 0 N2BEGb[1]
port 118 nsew signal output
flabel metal2 s 7102 11194 7158 11250 0 FreeSans 224 0 0 0 N2BEGb[2]
port 119 nsew signal output
flabel metal2 s 7378 11194 7434 11250 0 FreeSans 224 0 0 0 N2BEGb[3]
port 120 nsew signal output
flabel metal2 s 7654 11194 7710 11250 0 FreeSans 224 0 0 0 N2BEGb[4]
port 121 nsew signal output
flabel metal2 s 7930 11194 7986 11250 0 FreeSans 224 0 0 0 N2BEGb[5]
port 122 nsew signal output
flabel metal2 s 8206 11194 8262 11250 0 FreeSans 224 0 0 0 N2BEGb[6]
port 123 nsew signal output
flabel metal2 s 8482 11194 8538 11250 0 FreeSans 224 0 0 0 N2BEGb[7]
port 124 nsew signal output
flabel metal2 s 8758 11194 8814 11250 0 FreeSans 224 0 0 0 N4BEG[0]
port 125 nsew signal output
flabel metal2 s 11518 11194 11574 11250 0 FreeSans 224 0 0 0 N4BEG[10]
port 126 nsew signal output
flabel metal2 s 11794 11194 11850 11250 0 FreeSans 224 0 0 0 N4BEG[11]
port 127 nsew signal output
flabel metal2 s 12070 11194 12126 11250 0 FreeSans 224 0 0 0 N4BEG[12]
port 128 nsew signal output
flabel metal2 s 12346 11194 12402 11250 0 FreeSans 224 0 0 0 N4BEG[13]
port 129 nsew signal output
flabel metal2 s 12622 11194 12678 11250 0 FreeSans 224 0 0 0 N4BEG[14]
port 130 nsew signal output
flabel metal2 s 12898 11194 12954 11250 0 FreeSans 224 0 0 0 N4BEG[15]
port 131 nsew signal output
flabel metal2 s 9034 11194 9090 11250 0 FreeSans 224 0 0 0 N4BEG[1]
port 132 nsew signal output
flabel metal2 s 9310 11194 9366 11250 0 FreeSans 224 0 0 0 N4BEG[2]
port 133 nsew signal output
flabel metal2 s 9586 11194 9642 11250 0 FreeSans 224 0 0 0 N4BEG[3]
port 134 nsew signal output
flabel metal2 s 9862 11194 9918 11250 0 FreeSans 224 0 0 0 N4BEG[4]
port 135 nsew signal output
flabel metal2 s 10138 11194 10194 11250 0 FreeSans 224 0 0 0 N4BEG[5]
port 136 nsew signal output
flabel metal2 s 10414 11194 10470 11250 0 FreeSans 224 0 0 0 N4BEG[6]
port 137 nsew signal output
flabel metal2 s 10690 11194 10746 11250 0 FreeSans 224 0 0 0 N4BEG[7]
port 138 nsew signal output
flabel metal2 s 10966 11194 11022 11250 0 FreeSans 224 0 0 0 N4BEG[8]
port 139 nsew signal output
flabel metal2 s 11242 11194 11298 11250 0 FreeSans 224 0 0 0 N4BEG[9]
port 140 nsew signal output
flabel metal2 s 13174 11194 13230 11250 0 FreeSans 224 0 0 0 NN4BEG[0]
port 141 nsew signal output
flabel metal2 s 15934 11194 15990 11250 0 FreeSans 224 0 0 0 NN4BEG[10]
port 142 nsew signal output
flabel metal2 s 16210 11194 16266 11250 0 FreeSans 224 0 0 0 NN4BEG[11]
port 143 nsew signal output
flabel metal2 s 16486 11194 16542 11250 0 FreeSans 224 0 0 0 NN4BEG[12]
port 144 nsew signal output
flabel metal2 s 16762 11194 16818 11250 0 FreeSans 224 0 0 0 NN4BEG[13]
port 145 nsew signal output
flabel metal2 s 17038 11194 17094 11250 0 FreeSans 224 0 0 0 NN4BEG[14]
port 146 nsew signal output
flabel metal2 s 17314 11194 17370 11250 0 FreeSans 224 0 0 0 NN4BEG[15]
port 147 nsew signal output
flabel metal2 s 13450 11194 13506 11250 0 FreeSans 224 0 0 0 NN4BEG[1]
port 148 nsew signal output
flabel metal2 s 13726 11194 13782 11250 0 FreeSans 224 0 0 0 NN4BEG[2]
port 149 nsew signal output
flabel metal2 s 14002 11194 14058 11250 0 FreeSans 224 0 0 0 NN4BEG[3]
port 150 nsew signal output
flabel metal2 s 14278 11194 14334 11250 0 FreeSans 224 0 0 0 NN4BEG[4]
port 151 nsew signal output
flabel metal2 s 14554 11194 14610 11250 0 FreeSans 224 0 0 0 NN4BEG[5]
port 152 nsew signal output
flabel metal2 s 14830 11194 14886 11250 0 FreeSans 224 0 0 0 NN4BEG[6]
port 153 nsew signal output
flabel metal2 s 15106 11194 15162 11250 0 FreeSans 224 0 0 0 NN4BEG[7]
port 154 nsew signal output
flabel metal2 s 15382 11194 15438 11250 0 FreeSans 224 0 0 0 NN4BEG[8]
port 155 nsew signal output
flabel metal2 s 15658 11194 15714 11250 0 FreeSans 224 0 0 0 NN4BEG[9]
port 156 nsew signal output
flabel metal2 s 17866 11194 17922 11250 0 FreeSans 224 0 0 0 S1END[0]
port 157 nsew signal input
flabel metal2 s 18142 11194 18198 11250 0 FreeSans 224 0 0 0 S1END[1]
port 158 nsew signal input
flabel metal2 s 18418 11194 18474 11250 0 FreeSans 224 0 0 0 S1END[2]
port 159 nsew signal input
flabel metal2 s 18694 11194 18750 11250 0 FreeSans 224 0 0 0 S1END[3]
port 160 nsew signal input
flabel metal2 s 21178 11194 21234 11250 0 FreeSans 224 0 0 0 S2END[0]
port 161 nsew signal input
flabel metal2 s 21454 11194 21510 11250 0 FreeSans 224 0 0 0 S2END[1]
port 162 nsew signal input
flabel metal2 s 21730 11194 21786 11250 0 FreeSans 224 0 0 0 S2END[2]
port 163 nsew signal input
flabel metal2 s 22006 11194 22062 11250 0 FreeSans 224 0 0 0 S2END[3]
port 164 nsew signal input
flabel metal2 s 22282 11194 22338 11250 0 FreeSans 224 0 0 0 S2END[4]
port 165 nsew signal input
flabel metal2 s 22558 11194 22614 11250 0 FreeSans 224 0 0 0 S2END[5]
port 166 nsew signal input
flabel metal2 s 22834 11194 22890 11250 0 FreeSans 224 0 0 0 S2END[6]
port 167 nsew signal input
flabel metal2 s 23110 11194 23166 11250 0 FreeSans 224 0 0 0 S2END[7]
port 168 nsew signal input
flabel metal2 s 18970 11194 19026 11250 0 FreeSans 224 0 0 0 S2MID[0]
port 169 nsew signal input
flabel metal2 s 19246 11194 19302 11250 0 FreeSans 224 0 0 0 S2MID[1]
port 170 nsew signal input
flabel metal2 s 19522 11194 19578 11250 0 FreeSans 224 0 0 0 S2MID[2]
port 171 nsew signal input
flabel metal2 s 19798 11194 19854 11250 0 FreeSans 224 0 0 0 S2MID[3]
port 172 nsew signal input
flabel metal2 s 20074 11194 20130 11250 0 FreeSans 224 0 0 0 S2MID[4]
port 173 nsew signal input
flabel metal2 s 20350 11194 20406 11250 0 FreeSans 224 0 0 0 S2MID[5]
port 174 nsew signal input
flabel metal2 s 20626 11194 20682 11250 0 FreeSans 224 0 0 0 S2MID[6]
port 175 nsew signal input
flabel metal2 s 20902 11194 20958 11250 0 FreeSans 224 0 0 0 S2MID[7]
port 176 nsew signal input
flabel metal2 s 23386 11194 23442 11250 0 FreeSans 224 0 0 0 S4END[0]
port 177 nsew signal input
flabel metal2 s 26146 11194 26202 11250 0 FreeSans 224 0 0 0 S4END[10]
port 178 nsew signal input
flabel metal2 s 26422 11194 26478 11250 0 FreeSans 224 0 0 0 S4END[11]
port 179 nsew signal input
flabel metal2 s 26698 11194 26754 11250 0 FreeSans 224 0 0 0 S4END[12]
port 180 nsew signal input
flabel metal2 s 26974 11194 27030 11250 0 FreeSans 224 0 0 0 S4END[13]
port 181 nsew signal input
flabel metal2 s 27250 11194 27306 11250 0 FreeSans 224 0 0 0 S4END[14]
port 182 nsew signal input
flabel metal2 s 27526 11194 27582 11250 0 FreeSans 224 0 0 0 S4END[15]
port 183 nsew signal input
flabel metal2 s 23662 11194 23718 11250 0 FreeSans 224 0 0 0 S4END[1]
port 184 nsew signal input
flabel metal2 s 23938 11194 23994 11250 0 FreeSans 224 0 0 0 S4END[2]
port 185 nsew signal input
flabel metal2 s 24214 11194 24270 11250 0 FreeSans 224 0 0 0 S4END[3]
port 186 nsew signal input
flabel metal2 s 24490 11194 24546 11250 0 FreeSans 224 0 0 0 S4END[4]
port 187 nsew signal input
flabel metal2 s 24766 11194 24822 11250 0 FreeSans 224 0 0 0 S4END[5]
port 188 nsew signal input
flabel metal2 s 25042 11194 25098 11250 0 FreeSans 224 0 0 0 S4END[6]
port 189 nsew signal input
flabel metal2 s 25318 11194 25374 11250 0 FreeSans 224 0 0 0 S4END[7]
port 190 nsew signal input
flabel metal2 s 25594 11194 25650 11250 0 FreeSans 224 0 0 0 S4END[8]
port 191 nsew signal input
flabel metal2 s 25870 11194 25926 11250 0 FreeSans 224 0 0 0 S4END[9]
port 192 nsew signal input
flabel metal2 s 27802 11194 27858 11250 0 FreeSans 224 0 0 0 SS4END[0]
port 193 nsew signal input
flabel metal2 s 30562 11194 30618 11250 0 FreeSans 224 0 0 0 SS4END[10]
port 194 nsew signal input
flabel metal2 s 30838 11194 30894 11250 0 FreeSans 224 0 0 0 SS4END[11]
port 195 nsew signal input
flabel metal2 s 31114 11194 31170 11250 0 FreeSans 224 0 0 0 SS4END[12]
port 196 nsew signal input
flabel metal2 s 31390 11194 31446 11250 0 FreeSans 224 0 0 0 SS4END[13]
port 197 nsew signal input
flabel metal2 s 31666 11194 31722 11250 0 FreeSans 224 0 0 0 SS4END[14]
port 198 nsew signal input
flabel metal2 s 31942 11194 31998 11250 0 FreeSans 224 0 0 0 SS4END[15]
port 199 nsew signal input
flabel metal2 s 28078 11194 28134 11250 0 FreeSans 224 0 0 0 SS4END[1]
port 200 nsew signal input
flabel metal2 s 28354 11194 28410 11250 0 FreeSans 224 0 0 0 SS4END[2]
port 201 nsew signal input
flabel metal2 s 28630 11194 28686 11250 0 FreeSans 224 0 0 0 SS4END[3]
port 202 nsew signal input
flabel metal2 s 28906 11194 28962 11250 0 FreeSans 224 0 0 0 SS4END[4]
port 203 nsew signal input
flabel metal2 s 29182 11194 29238 11250 0 FreeSans 224 0 0 0 SS4END[5]
port 204 nsew signal input
flabel metal2 s 29458 11194 29514 11250 0 FreeSans 224 0 0 0 SS4END[6]
port 205 nsew signal input
flabel metal2 s 29734 11194 29790 11250 0 FreeSans 224 0 0 0 SS4END[7]
port 206 nsew signal input
flabel metal2 s 30010 11194 30066 11250 0 FreeSans 224 0 0 0 SS4END[8]
port 207 nsew signal input
flabel metal2 s 30286 11194 30342 11250 0 FreeSans 224 0 0 0 SS4END[9]
port 208 nsew signal input
flabel metal2 s 1122 0 1178 56 0 FreeSans 224 0 0 0 UserCLK
port 209 nsew signal input
flabel metal2 s 32218 11194 32274 11250 0 FreeSans 224 0 0 0 UserCLKo
port 210 nsew signal output
flabel metal4 s 3004 0 3324 11250 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 3004 11190 3324 11250 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11250 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 9004 11190 9324 11250 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11250 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 15004 11190 15324 11250 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11250 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 21004 11190 21324 11250 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11250 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 27004 11190 27324 11250 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11250 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 33004 11190 33324 11250 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 39004 0 39324 11250 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 39004 0 39324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 39004 11190 39324 11250 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11250 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 1944 11190 2264 11250 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 7944 0 8264 11250 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 7944 11190 8264 11250 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 13944 0 14264 11250 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 13944 11190 14264 11250 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 19944 0 20264 11250 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 19944 11190 20264 11250 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 25944 0 26264 11250 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 25944 11190 26264 11250 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 31944 0 32264 11250 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 31944 11190 32264 11250 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 37944 0 38264 11250 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 37944 0 38264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 37944 11190 38264 11250 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
rlabel metal1 20470 8704 20470 8704 0 VGND
rlabel metal1 20470 8160 20470 8160 0 VPWR
rlabel metal2 9614 2125 9614 2125 0 FrameData[0]
rlabel metal1 16652 5542 16652 5542 0 FrameData[10]
rlabel metal3 1471 4420 1471 4420 0 FrameData[11]
rlabel metal2 8234 4403 8234 4403 0 FrameData[12]
rlabel metal3 919 4964 919 4964 0 FrameData[13]
rlabel metal3 1402 5236 1402 5236 0 FrameData[14]
rlabel metal3 1471 5508 1471 5508 0 FrameData[15]
rlabel metal3 1770 5780 1770 5780 0 FrameData[16]
rlabel metal3 942 6052 942 6052 0 FrameData[17]
rlabel via2 19182 6307 19182 6307 0 FrameData[18]
rlabel metal3 1448 6596 1448 6596 0 FrameData[19]
rlabel metal2 9522 2295 9522 2295 0 FrameData[1]
rlabel metal2 16330 5831 16330 5831 0 FrameData[20]
rlabel metal3 712 7140 712 7140 0 FrameData[21]
rlabel metal3 10396 7344 10396 7344 0 FrameData[22]
rlabel metal3 390 7684 390 7684 0 FrameData[23]
rlabel metal3 160 7956 160 7956 0 FrameData[24]
rlabel metal3 620 8228 620 8228 0 FrameData[25]
rlabel metal1 20838 8058 20838 8058 0 FrameData[26]
rlabel metal3 1448 8772 1448 8772 0 FrameData[27]
rlabel metal1 15364 7990 15364 7990 0 FrameData[28]
rlabel metal1 17760 7378 17760 7378 0 FrameData[29]
rlabel metal2 9430 2465 9430 2465 0 FrameData[2]
rlabel metal2 27738 8721 27738 8721 0 FrameData[30]
rlabel metal1 19228 7854 19228 7854 0 FrameData[31]
rlabel metal3 1471 2244 1471 2244 0 FrameData[3]
rlabel metal3 14282 2516 14282 2516 0 FrameData[4]
rlabel metal3 919 2788 919 2788 0 FrameData[5]
rlabel via2 20746 3179 20746 3179 0 FrameData[6]
rlabel metal3 1494 3332 1494 3332 0 FrameData[7]
rlabel metal3 1816 3604 1816 3604 0 FrameData[8]
rlabel metal3 919 3876 919 3876 0 FrameData[9]
rlabel metal3 39798 1428 39798 1428 0 FrameData_O[0]
rlabel metal3 40166 4148 40166 4148 0 FrameData_O[10]
rlabel metal3 40442 4420 40442 4420 0 FrameData_O[11]
rlabel metal3 40166 4692 40166 4692 0 FrameData_O[12]
rlabel metal3 39982 4964 39982 4964 0 FrameData_O[13]
rlabel metal3 40166 5236 40166 5236 0 FrameData_O[14]
rlabel metal3 40442 5508 40442 5508 0 FrameData_O[15]
rlabel metal3 40166 5780 40166 5780 0 FrameData_O[16]
rlabel metal3 39982 6052 39982 6052 0 FrameData_O[17]
rlabel metal3 39798 6324 39798 6324 0 FrameData_O[18]
rlabel metal2 39422 6511 39422 6511 0 FrameData_O[19]
rlabel metal3 39614 1700 39614 1700 0 FrameData_O[1]
rlabel metal3 40212 6868 40212 6868 0 FrameData_O[20]
rlabel metal3 40166 7140 40166 7140 0 FrameData_O[21]
rlabel metal3 39936 7412 39936 7412 0 FrameData_O[22]
rlabel metal3 40166 7684 40166 7684 0 FrameData_O[23]
rlabel metal3 40166 7956 40166 7956 0 FrameData_O[24]
rlabel metal3 39982 8228 39982 8228 0 FrameData_O[25]
rlabel metal2 38686 8279 38686 8279 0 FrameData_O[26]
rlabel metal1 39284 7514 39284 7514 0 FrameData_O[27]
rlabel metal1 39514 6630 39514 6630 0 FrameData_O[28]
rlabel metal1 38732 7514 38732 7514 0 FrameData_O[29]
rlabel metal3 39430 1972 39430 1972 0 FrameData_O[2]
rlabel metal1 39054 6664 39054 6664 0 FrameData_O[30]
rlabel metal3 39660 9860 39660 9860 0 FrameData_O[31]
rlabel metal3 40442 2244 40442 2244 0 FrameData_O[3]
rlabel metal3 40166 2516 40166 2516 0 FrameData_O[4]
rlabel metal3 39982 2788 39982 2788 0 FrameData_O[5]
rlabel metal3 40166 3060 40166 3060 0 FrameData_O[6]
rlabel metal3 40442 3332 40442 3332 0 FrameData_O[7]
rlabel metal3 40166 3604 40166 3604 0 FrameData_O[8]
rlabel metal3 39982 3876 39982 3876 0 FrameData_O[9]
rlabel metal2 3082 55 3082 55 0 FrameStrobe[0]
rlabel metal2 22402 718 22402 718 0 FrameStrobe[10]
rlabel metal1 21229 4590 21229 4590 0 FrameStrobe[11]
rlabel metal2 19826 4675 19826 4675 0 FrameStrobe[12]
rlabel metal2 28152 3740 28152 3740 0 FrameStrobe[13]
rlabel metal1 29164 4590 29164 4590 0 FrameStrobe[14]
rlabel metal2 32062 55 32062 55 0 FrameStrobe[15]
rlabel metal1 32936 4522 32936 4522 0 FrameStrobe[16]
rlabel metal1 34776 4590 34776 4590 0 FrameStrobe[17]
rlabel metal1 36754 5610 36754 5610 0 FrameStrobe[18]
rlabel metal1 39284 5882 39284 5882 0 FrameStrobe[19]
rlabel metal2 5014 106 5014 106 0 FrameStrobe[1]
rlabel metal1 5382 7752 5382 7752 0 FrameStrobe[2]
rlabel via2 8878 55 8878 55 0 FrameStrobe[3]
rlabel metal2 10810 1619 10810 1619 0 FrameStrobe[4]
rlabel metal2 12742 1058 12742 1058 0 FrameStrobe[5]
rlabel metal2 14674 1755 14674 1755 0 FrameStrobe[6]
rlabel metal2 16606 1160 16606 1160 0 FrameStrobe[7]
rlabel metal2 18538 55 18538 55 0 FrameStrobe[8]
rlabel metal2 20470 2894 20470 2894 0 FrameStrobe[9]
rlabel metal1 32660 8602 32660 8602 0 FrameStrobe_O[0]
rlabel metal1 36386 8296 36386 8296 0 FrameStrobe_O[10]
rlabel metal1 35696 8058 35696 8058 0 FrameStrobe_O[11]
rlabel metal1 36294 8602 36294 8602 0 FrameStrobe_O[12]
rlabel metal1 36248 8058 36248 8058 0 FrameStrobe_O[13]
rlabel metal1 37306 8262 37306 8262 0 FrameStrobe_O[14]
rlabel metal1 36800 8058 36800 8058 0 FrameStrobe_O[15]
rlabel metal1 37398 8602 37398 8602 0 FrameStrobe_O[16]
rlabel metal1 37720 8330 37720 8330 0 FrameStrobe_O[17]
rlabel metal1 38594 8568 38594 8568 0 FrameStrobe_O[18]
rlabel metal1 37858 8058 37858 8058 0 FrameStrobe_O[19]
rlabel metal1 33028 8602 33028 8602 0 FrameStrobe_O[1]
rlabel metal2 33534 8704 33534 8704 0 FrameStrobe_O[2]
rlabel metal1 33902 8568 33902 8568 0 FrameStrobe_O[3]
rlabel metal2 34270 8806 34270 8806 0 FrameStrobe_O[4]
rlabel metal1 34454 8330 34454 8330 0 FrameStrobe_O[5]
rlabel metal1 35282 8330 35282 8330 0 FrameStrobe_O[6]
rlabel metal1 34638 8058 34638 8058 0 FrameStrobe_O[7]
rlabel metal1 35144 8602 35144 8602 0 FrameStrobe_O[8]
rlabel metal1 35696 8330 35696 8330 0 FrameStrobe_O[9]
rlabel metal2 3542 8619 3542 8619 0 N1BEG[0]
rlabel metal1 3404 8330 3404 8330 0 N1BEG[1]
rlabel metal1 3680 8602 3680 8602 0 N1BEG[2]
rlabel metal1 4186 8058 4186 8058 0 N1BEG[3]
rlabel metal1 4324 8602 4324 8602 0 N2BEG[0]
rlabel metal2 4646 9904 4646 9904 0 N2BEG[1]
rlabel metal1 5060 8058 5060 8058 0 N2BEG[2]
rlabel metal1 5060 8602 5060 8602 0 N2BEG[3]
rlabel metal1 5382 8602 5382 8602 0 N2BEG[4]
rlabel metal1 5704 8602 5704 8602 0 N2BEG[5]
rlabel metal1 6118 8058 6118 8058 0 N2BEG[6]
rlabel metal1 6164 8602 6164 8602 0 N2BEG[7]
rlabel metal1 6716 8058 6716 8058 0 N2BEGb[0]
rlabel metal1 6808 8602 6808 8602 0 N2BEGb[1]
rlabel metal1 7222 8058 7222 8058 0 N2BEGb[2]
rlabel metal1 7268 8602 7268 8602 0 N2BEGb[3]
rlabel metal1 7590 8602 7590 8602 0 N2BEGb[4]
rlabel metal1 7912 8602 7912 8602 0 N2BEGb[5]
rlabel metal1 8372 8058 8372 8058 0 N2BEGb[6]
rlabel metal1 8372 8602 8372 8602 0 N2BEGb[7]
rlabel metal1 8924 8058 8924 8058 0 N4BEG[0]
rlabel metal1 11362 8602 11362 8602 0 N4BEG[10]
rlabel metal2 11822 9632 11822 9632 0 N4BEG[11]
rlabel metal1 12006 8602 12006 8602 0 N4BEG[12]
rlabel metal1 12328 8602 12328 8602 0 N4BEG[13]
rlabel metal1 12742 8058 12742 8058 0 N4BEG[14]
rlabel metal1 12788 8602 12788 8602 0 N4BEG[15]
rlabel metal1 8740 8602 8740 8602 0 N4BEG[1]
rlabel metal1 9476 8058 9476 8058 0 N4BEG[2]
rlabel metal1 9476 8602 9476 8602 0 N4BEG[3]
rlabel metal1 9844 8602 9844 8602 0 N4BEG[4]
rlabel metal2 10166 9904 10166 9904 0 N4BEG[5]
rlabel metal1 10534 8058 10534 8058 0 N4BEG[6]
rlabel metal1 10580 8602 10580 8602 0 N4BEG[7]
rlabel metal1 10902 8602 10902 8602 0 N4BEG[8]
rlabel metal1 11362 8058 11362 8058 0 N4BEG[9]
rlabel metal1 13110 8602 13110 8602 0 NN4BEG[0]
rlabel metal1 16054 8058 16054 8058 0 NN4BEG[10]
rlabel metal1 16100 8602 16100 8602 0 NN4BEG[11]
rlabel metal1 16422 8602 16422 8602 0 NN4BEG[12]
rlabel metal1 16882 8602 16882 8602 0 NN4BEG[13]
rlabel metal2 17894 8738 17894 8738 0 NN4BEG[14]
rlabel metal1 17480 8602 17480 8602 0 NN4BEG[15]
rlabel metal1 13570 8058 13570 8058 0 NN4BEG[1]
rlabel metal1 13524 8602 13524 8602 0 NN4BEG[2]
rlabel metal1 13892 8602 13892 8602 0 NN4BEG[3]
rlabel metal1 14398 8058 14398 8058 0 NN4BEG[4]
rlabel metal1 14536 8602 14536 8602 0 NN4BEG[5]
rlabel metal1 15272 8058 15272 8058 0 NN4BEG[6]
rlabel metal1 14904 8602 14904 8602 0 NN4BEG[7]
rlabel metal1 15318 8602 15318 8602 0 NN4BEG[8]
rlabel metal1 15640 8602 15640 8602 0 NN4BEG[9]
rlabel metal1 4876 5746 4876 5746 0 S1END[0]
rlabel metal1 3266 6358 3266 6358 0 S1END[1]
rlabel metal1 4508 6766 4508 6766 0 S1END[2]
rlabel metal2 7222 7820 7222 7820 0 S1END[3]
rlabel metal2 21206 10057 21206 10057 0 S2END[0]
rlabel metal2 21482 10057 21482 10057 0 S2END[1]
rlabel metal1 11730 6358 11730 6358 0 S2END[2]
rlabel metal1 10350 6766 10350 6766 0 S2END[3]
rlabel metal1 8602 6290 8602 6290 0 S2END[4]
rlabel metal1 7636 6290 7636 6290 0 S2END[5]
rlabel metal1 11730 5644 11730 5644 0 S2END[6]
rlabel metal1 6279 5202 6279 5202 0 S2END[7]
rlabel metal2 18998 10465 18998 10465 0 S2MID[0]
rlabel metal1 9752 6290 9752 6290 0 S2MID[1]
rlabel metal1 6854 5712 6854 5712 0 S2MID[2]
rlabel metal1 5750 5746 5750 5746 0 S2MID[3]
rlabel metal2 5566 4930 5566 4930 0 S2MID[4]
rlabel metal1 5106 5644 5106 5644 0 S2MID[5]
rlabel metal2 4646 6562 4646 6562 0 S2MID[6]
rlabel metal2 3818 6528 3818 6528 0 S2MID[7]
rlabel metal2 23414 10433 23414 10433 0 S4END[0]
rlabel metal1 12374 7480 12374 7480 0 S4END[10]
rlabel metal1 8878 7718 8878 7718 0 S4END[11]
rlabel metal2 9798 8823 9798 8823 0 S4END[12]
rlabel metal1 14904 7446 14904 7446 0 S4END[13]
rlabel metal2 27278 10006 27278 10006 0 S4END[14]
rlabel metal1 12926 7888 12926 7888 0 S4END[15]
rlabel metal2 20378 8007 20378 8007 0 S4END[1]
rlabel metal2 16974 9146 16974 9146 0 S4END[2]
rlabel metal1 16054 7174 16054 7174 0 S4END[3]
rlabel metal2 24518 9258 24518 9258 0 S4END[4]
rlabel metal2 19366 8500 19366 8500 0 S4END[5]
rlabel via2 17342 5219 17342 5219 0 S4END[6]
rlabel metal2 19090 7633 19090 7633 0 S4END[7]
rlabel metal2 14858 4386 14858 4386 0 S4END[8]
rlabel metal1 11822 6324 11822 6324 0 S4END[9]
rlabel metal2 7314 9282 7314 9282 0 SS4END[0]
rlabel metal2 30590 8986 30590 8986 0 SS4END[10]
rlabel metal2 30866 9292 30866 9292 0 SS4END[11]
rlabel metal2 31142 9530 31142 9530 0 SS4END[12]
rlabel metal2 31418 9530 31418 9530 0 SS4END[13]
rlabel metal2 31694 8986 31694 8986 0 SS4END[14]
rlabel metal2 31970 10433 31970 10433 0 SS4END[15]
rlabel metal2 21758 8228 21758 8228 0 SS4END[1]
rlabel metal2 28382 9292 28382 9292 0 SS4END[2]
rlabel metal2 28658 10533 28658 10533 0 SS4END[3]
rlabel metal2 28934 9632 28934 9632 0 SS4END[4]
rlabel metal2 29210 10125 29210 10125 0 SS4END[5]
rlabel metal2 29486 9989 29486 9989 0 SS4END[6]
rlabel metal2 29762 10465 29762 10465 0 SS4END[7]
rlabel metal2 30038 8442 30038 8442 0 SS4END[8]
rlabel metal2 30314 8748 30314 8748 0 SS4END[9]
rlabel metal2 1150 55 1150 55 0 UserCLK
rlabel metal1 32292 8602 32292 8602 0 UserCLKo
rlabel metal2 13386 2652 13386 2652 0 net1
rlabel metal2 38502 6426 38502 6426 0 net10
rlabel metal2 16422 7514 16422 7514 0 net100
rlabel metal2 15870 7038 15870 7038 0 net101
rlabel metal1 18354 5644 18354 5644 0 net102
rlabel metal2 15594 8738 15594 8738 0 net103
rlabel metal2 15778 8874 15778 8874 0 net104
rlabel metal1 28244 5882 28244 5882 0 net105
rlabel metal1 18078 8398 18078 8398 0 net106
rlabel metal2 39238 6052 39238 6052 0 net11
rlabel metal2 16238 2686 16238 2686 0 net12
rlabel metal1 16744 4794 16744 4794 0 net13
rlabel metal1 39238 7412 39238 7412 0 net14
rlabel metal2 18446 3944 18446 3944 0 net15
rlabel metal2 36386 7531 36386 7531 0 net16
rlabel metal2 38962 8840 38962 8840 0 net17
rlabel metal2 38778 6443 38778 6443 0 net18
rlabel metal2 21390 7616 21390 7616 0 net19
rlabel metal2 38686 4556 38686 4556 0 net2
rlabel metal1 38870 7344 38870 7344 0 net20
rlabel metal2 15502 6749 15502 6749 0 net21
rlabel metal2 33718 7327 33718 7327 0 net22
rlabel metal1 18147 2890 18147 2890 0 net23
rlabel metal2 34178 7208 34178 7208 0 net24
rlabel metal2 19458 7344 19458 7344 0 net25
rlabel metal2 9062 2652 9062 2652 0 net26
rlabel metal1 39238 2380 39238 2380 0 net27
rlabel metal1 38870 2958 38870 2958 0 net28
rlabel metal1 36202 3026 36202 3026 0 net29
rlabel metal2 19090 4352 19090 4352 0 net3
rlabel metal2 35282 3774 35282 3774 0 net30
rlabel metal2 39238 3740 39238 3740 0 net31
rlabel metal2 38870 3740 38870 3740 0 net32
rlabel metal2 10810 7769 10810 7769 0 net33
rlabel metal1 32982 8840 32982 8840 0 net34
rlabel metal1 21321 4454 21321 4454 0 net35
rlabel metal2 36570 8908 36570 8908 0 net36
rlabel metal2 36202 6256 36202 6256 0 net37
rlabel metal1 32890 8908 32890 8908 0 net38
rlabel metal1 34270 7480 34270 7480 0 net39
rlabel metal1 13846 4148 13846 4148 0 net4
rlabel metal1 34638 4454 34638 4454 0 net40
rlabel metal2 33810 6800 33810 6800 0 net41
rlabel metal1 35742 5542 35742 5542 0 net42
rlabel metal1 38226 5882 38226 5882 0 net43
rlabel metal2 32706 7582 32706 7582 0 net44
rlabel via2 4002 7939 4002 7939 0 net45
rlabel metal1 33442 8432 33442 8432 0 net46
rlabel metal2 34086 5984 34086 5984 0 net47
rlabel metal1 33718 8364 33718 8364 0 net48
rlabel metal1 34316 3162 34316 3162 0 net49
rlabel metal2 5842 3808 5842 3808 0 net5
rlabel metal2 36294 5814 36294 5814 0 net50
rlabel metal1 36478 5882 36478 5882 0 net51
rlabel metal1 35650 5882 35650 5882 0 net52
rlabel metal2 2806 7684 2806 7684 0 net53
rlabel metal1 2944 8466 2944 8466 0 net54
rlabel metal1 3358 6426 3358 6426 0 net55
rlabel metal1 4094 5882 4094 5882 0 net56
rlabel metal1 3864 6426 3864 6426 0 net57
rlabel metal2 4462 7446 4462 7446 0 net58
rlabel metal1 4968 5882 4968 5882 0 net59
rlabel metal2 36018 4284 36018 4284 0 net6
rlabel metal1 5244 5338 5244 5338 0 net60
rlabel metal1 5520 5882 5520 5882 0 net61
rlabel metal1 6256 5882 6256 5882 0 net62
rlabel metal1 6394 7820 6394 7820 0 net63
rlabel metal1 6210 8500 6210 8500 0 net64
rlabel metal1 6256 5338 6256 5338 0 net65
rlabel metal1 7038 5882 7038 5882 0 net66
rlabel metal1 7590 6426 7590 6426 0 net67
rlabel metal1 8050 6426 8050 6426 0 net68
rlabel metal1 8510 6630 8510 6630 0 net69
rlabel metal1 15134 3400 15134 3400 0 net7
rlabel metal1 10626 6392 10626 6392 0 net70
rlabel metal1 10442 7310 10442 7310 0 net71
rlabel metal2 8418 8840 8418 8840 0 net72
rlabel metal1 9246 7922 9246 7922 0 net73
rlabel metal2 11362 8636 11362 8636 0 net74
rlabel metal1 12006 7888 12006 7888 0 net75
rlabel metal1 12098 8398 12098 8398 0 net76
rlabel metal1 13984 8058 13984 8058 0 net77
rlabel metal1 13018 7820 13018 7820 0 net78
rlabel metal2 19734 8500 19734 8500 0 net79
rlabel metal2 36110 4318 36110 4318 0 net8
rlabel metal2 8694 8704 8694 8704 0 net80
rlabel metal2 11914 7582 11914 7582 0 net81
rlabel metal1 9568 7514 9568 7514 0 net82
rlabel metal1 8326 7990 8326 7990 0 net83
rlabel metal1 9752 7242 9752 7242 0 net84
rlabel metal1 11592 6426 11592 6426 0 net85
rlabel metal1 10764 8466 10764 8466 0 net86
rlabel metal2 10994 6868 10994 6868 0 net87
rlabel metal2 17158 5576 17158 5576 0 net88
rlabel metal2 13202 8143 13202 8143 0 net89
rlabel via2 11454 4539 11454 4539 0 net9
rlabel metal2 19182 7582 19182 7582 0 net90
rlabel metal2 16146 8636 16146 8636 0 net91
rlabel metal2 23138 8228 23138 8228 0 net92
rlabel metal1 17158 8398 17158 8398 0 net93
rlabel metal1 20976 7514 20976 7514 0 net94
rlabel metal2 12190 7072 12190 7072 0 net95
rlabel metal2 13846 7293 13846 7293 0 net96
rlabel metal2 20470 7650 20470 7650 0 net97
rlabel metal1 17066 8296 17066 8296 0 net98
rlabel metal1 14674 7888 14674 7888 0 net99
<< properties >>
string FIXED_BBOX 0 0 41000 11250
<< end >>
