* NGSPICE file created from EF_SRAM.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

.subckt EF_SRAM AD_SRAM0 AD_SRAM1 AD_SRAM2 AD_SRAM3 AD_SRAM4 AD_SRAM5 AD_SRAM6 AD_SRAM7
+ AD_SRAM8 AD_SRAM9 BEN_SRAM0 BEN_SRAM1 BEN_SRAM10 BEN_SRAM11 BEN_SRAM12 BEN_SRAM13
+ BEN_SRAM14 BEN_SRAM15 BEN_SRAM16 BEN_SRAM17 BEN_SRAM18 BEN_SRAM19 BEN_SRAM2 BEN_SRAM20
+ BEN_SRAM21 BEN_SRAM22 BEN_SRAM23 BEN_SRAM24 BEN_SRAM25 BEN_SRAM26 BEN_SRAM27 BEN_SRAM28
+ BEN_SRAM29 BEN_SRAM3 BEN_SRAM30 BEN_SRAM31 BEN_SRAM4 BEN_SRAM5 BEN_SRAM6 BEN_SRAM7
+ BEN_SRAM8 BEN_SRAM9 CLOCK_SRAM DI_SRAM0 DI_SRAM1 DI_SRAM10 DI_SRAM11 DI_SRAM12 DI_SRAM13
+ DI_SRAM14 DI_SRAM15 DI_SRAM16 DI_SRAM17 DI_SRAM18 DI_SRAM19 DI_SRAM2 DI_SRAM20 DI_SRAM21
+ DI_SRAM22 DI_SRAM23 DI_SRAM24 DI_SRAM25 DI_SRAM26 DI_SRAM27 DI_SRAM28 DI_SRAM29
+ DI_SRAM3 DI_SRAM30 DI_SRAM31 DI_SRAM4 DI_SRAM5 DI_SRAM6 DI_SRAM7 DI_SRAM8 DI_SRAM9
+ DO_SRAM0 DO_SRAM1 DO_SRAM10 DO_SRAM11 DO_SRAM12 DO_SRAM13 DO_SRAM14 DO_SRAM15 DO_SRAM16
+ DO_SRAM17 DO_SRAM18 DO_SRAM19 DO_SRAM2 DO_SRAM20 DO_SRAM21 DO_SRAM22 DO_SRAM23 DO_SRAM24
+ DO_SRAM25 DO_SRAM26 DO_SRAM27 DO_SRAM28 DO_SRAM29 DO_SRAM3 DO_SRAM30 DO_SRAM31 DO_SRAM4
+ DO_SRAM5 DO_SRAM6 DO_SRAM7 DO_SRAM8 DO_SRAM9 EN_SRAM R_WB_SRAM Tile_X0Y0_E1END[0]
+ Tile_X0Y0_E1END[1] Tile_X0Y0_E1END[2] Tile_X0Y0_E1END[3] Tile_X0Y0_E2END[0] Tile_X0Y0_E2END[1]
+ Tile_X0Y0_E2END[2] Tile_X0Y0_E2END[3] Tile_X0Y0_E2END[4] Tile_X0Y0_E2END[5] Tile_X0Y0_E2END[6]
+ Tile_X0Y0_E2END[7] Tile_X0Y0_E2MID[0] Tile_X0Y0_E2MID[1] Tile_X0Y0_E2MID[2] Tile_X0Y0_E2MID[3]
+ Tile_X0Y0_E2MID[4] Tile_X0Y0_E2MID[5] Tile_X0Y0_E2MID[6] Tile_X0Y0_E2MID[7] Tile_X0Y0_E6END[0]
+ Tile_X0Y0_E6END[10] Tile_X0Y0_E6END[11] Tile_X0Y0_E6END[1] Tile_X0Y0_E6END[2] Tile_X0Y0_E6END[3]
+ Tile_X0Y0_E6END[4] Tile_X0Y0_E6END[5] Tile_X0Y0_E6END[6] Tile_X0Y0_E6END[7] Tile_X0Y0_E6END[8]
+ Tile_X0Y0_E6END[9] Tile_X0Y0_EE4END[0] Tile_X0Y0_EE4END[10] Tile_X0Y0_EE4END[11]
+ Tile_X0Y0_EE4END[12] Tile_X0Y0_EE4END[13] Tile_X0Y0_EE4END[14] Tile_X0Y0_EE4END[15]
+ Tile_X0Y0_EE4END[1] Tile_X0Y0_EE4END[2] Tile_X0Y0_EE4END[3] Tile_X0Y0_EE4END[4]
+ Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[6] Tile_X0Y0_EE4END[7] Tile_X0Y0_EE4END[8]
+ Tile_X0Y0_EE4END[9] Tile_X0Y0_FrameData[0] Tile_X0Y0_FrameData[10] Tile_X0Y0_FrameData[11]
+ Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData[13] Tile_X0Y0_FrameData[14] Tile_X0Y0_FrameData[15]
+ Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData[17] Tile_X0Y0_FrameData[18] Tile_X0Y0_FrameData[19]
+ Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData[20] Tile_X0Y0_FrameData[21] Tile_X0Y0_FrameData[22]
+ Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData[24] Tile_X0Y0_FrameData[25] Tile_X0Y0_FrameData[26]
+ Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData[28] Tile_X0Y0_FrameData[29] Tile_X0Y0_FrameData[2]
+ Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData[31] Tile_X0Y0_FrameData[3] Tile_X0Y0_FrameData[4]
+ Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData[6] Tile_X0Y0_FrameData[7] Tile_X0Y0_FrameData[8]
+ Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[0] Tile_X0Y0_FrameData_O[10] Tile_X0Y0_FrameData_O[11]
+ Tile_X0Y0_FrameData_O[12] Tile_X0Y0_FrameData_O[13] Tile_X0Y0_FrameData_O[14] Tile_X0Y0_FrameData_O[15]
+ Tile_X0Y0_FrameData_O[16] Tile_X0Y0_FrameData_O[17] Tile_X0Y0_FrameData_O[18] Tile_X0Y0_FrameData_O[19]
+ Tile_X0Y0_FrameData_O[1] Tile_X0Y0_FrameData_O[20] Tile_X0Y0_FrameData_O[21] Tile_X0Y0_FrameData_O[22]
+ Tile_X0Y0_FrameData_O[23] Tile_X0Y0_FrameData_O[24] Tile_X0Y0_FrameData_O[25] Tile_X0Y0_FrameData_O[26]
+ Tile_X0Y0_FrameData_O[27] Tile_X0Y0_FrameData_O[28] Tile_X0Y0_FrameData_O[29] Tile_X0Y0_FrameData_O[2]
+ Tile_X0Y0_FrameData_O[30] Tile_X0Y0_FrameData_O[31] Tile_X0Y0_FrameData_O[3] Tile_X0Y0_FrameData_O[4]
+ Tile_X0Y0_FrameData_O[5] Tile_X0Y0_FrameData_O[6] Tile_X0Y0_FrameData_O[7] Tile_X0Y0_FrameData_O[8]
+ Tile_X0Y0_FrameData_O[9] Tile_X0Y0_FrameStrobe_O[0] Tile_X0Y0_FrameStrobe_O[10]
+ Tile_X0Y0_FrameStrobe_O[11] Tile_X0Y0_FrameStrobe_O[12] Tile_X0Y0_FrameStrobe_O[13]
+ Tile_X0Y0_FrameStrobe_O[14] Tile_X0Y0_FrameStrobe_O[15] Tile_X0Y0_FrameStrobe_O[16]
+ Tile_X0Y0_FrameStrobe_O[17] Tile_X0Y0_FrameStrobe_O[18] Tile_X0Y0_FrameStrobe_O[19]
+ Tile_X0Y0_FrameStrobe_O[1] Tile_X0Y0_FrameStrobe_O[2] Tile_X0Y0_FrameStrobe_O[3]
+ Tile_X0Y0_FrameStrobe_O[4] Tile_X0Y0_FrameStrobe_O[5] Tile_X0Y0_FrameStrobe_O[6]
+ Tile_X0Y0_FrameStrobe_O[7] Tile_X0Y0_FrameStrobe_O[8] Tile_X0Y0_FrameStrobe_O[9]
+ Tile_X0Y0_N1BEG[0] Tile_X0Y0_N1BEG[1] Tile_X0Y0_N1BEG[2] Tile_X0Y0_N1BEG[3] Tile_X0Y0_N2BEG[0]
+ Tile_X0Y0_N2BEG[1] Tile_X0Y0_N2BEG[2] Tile_X0Y0_N2BEG[3] Tile_X0Y0_N2BEG[4] Tile_X0Y0_N2BEG[5]
+ Tile_X0Y0_N2BEG[6] Tile_X0Y0_N2BEG[7] Tile_X0Y0_N2BEGb[0] Tile_X0Y0_N2BEGb[1] Tile_X0Y0_N2BEGb[2]
+ Tile_X0Y0_N2BEGb[3] Tile_X0Y0_N2BEGb[4] Tile_X0Y0_N2BEGb[5] Tile_X0Y0_N2BEGb[6]
+ Tile_X0Y0_N2BEGb[7] Tile_X0Y0_N4BEG[0] Tile_X0Y0_N4BEG[10] Tile_X0Y0_N4BEG[11] Tile_X0Y0_N4BEG[12]
+ Tile_X0Y0_N4BEG[13] Tile_X0Y0_N4BEG[14] Tile_X0Y0_N4BEG[15] Tile_X0Y0_N4BEG[1] Tile_X0Y0_N4BEG[2]
+ Tile_X0Y0_N4BEG[3] Tile_X0Y0_N4BEG[4] Tile_X0Y0_N4BEG[5] Tile_X0Y0_N4BEG[6] Tile_X0Y0_N4BEG[7]
+ Tile_X0Y0_N4BEG[8] Tile_X0Y0_N4BEG[9] Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[1] Tile_X0Y0_S1END[2]
+ Tile_X0Y0_S1END[3] Tile_X0Y0_S2END[0] Tile_X0Y0_S2END[1] Tile_X0Y0_S2END[2] Tile_X0Y0_S2END[3]
+ Tile_X0Y0_S2END[4] Tile_X0Y0_S2END[5] Tile_X0Y0_S2END[6] Tile_X0Y0_S2END[7] Tile_X0Y0_S2MID[0]
+ Tile_X0Y0_S2MID[1] Tile_X0Y0_S2MID[2] Tile_X0Y0_S2MID[3] Tile_X0Y0_S2MID[4] Tile_X0Y0_S2MID[5]
+ Tile_X0Y0_S2MID[6] Tile_X0Y0_S2MID[7] Tile_X0Y0_S4END[0] Tile_X0Y0_S4END[10] Tile_X0Y0_S4END[11]
+ Tile_X0Y0_S4END[12] Tile_X0Y0_S4END[13] Tile_X0Y0_S4END[14] Tile_X0Y0_S4END[15]
+ Tile_X0Y0_S4END[1] Tile_X0Y0_S4END[2] Tile_X0Y0_S4END[3] Tile_X0Y0_S4END[4] Tile_X0Y0_S4END[5]
+ Tile_X0Y0_S4END[6] Tile_X0Y0_S4END[7] Tile_X0Y0_S4END[8] Tile_X0Y0_S4END[9] Tile_X0Y0_UserCLKo
+ Tile_X0Y0_W1BEG[0] Tile_X0Y0_W1BEG[1] Tile_X0Y0_W1BEG[2] Tile_X0Y0_W1BEG[3] Tile_X0Y0_W2BEG[0]
+ Tile_X0Y0_W2BEG[1] Tile_X0Y0_W2BEG[2] Tile_X0Y0_W2BEG[3] Tile_X0Y0_W2BEG[4] Tile_X0Y0_W2BEG[5]
+ Tile_X0Y0_W2BEG[6] Tile_X0Y0_W2BEG[7] Tile_X0Y0_W2BEGb[0] Tile_X0Y0_W2BEGb[1] Tile_X0Y0_W2BEGb[2]
+ Tile_X0Y0_W2BEGb[3] Tile_X0Y0_W2BEGb[4] Tile_X0Y0_W2BEGb[5] Tile_X0Y0_W2BEGb[6]
+ Tile_X0Y0_W2BEGb[7] Tile_X0Y0_W6BEG[0] Tile_X0Y0_W6BEG[10] Tile_X0Y0_W6BEG[11] Tile_X0Y0_W6BEG[1]
+ Tile_X0Y0_W6BEG[2] Tile_X0Y0_W6BEG[3] Tile_X0Y0_W6BEG[4] Tile_X0Y0_W6BEG[5] Tile_X0Y0_W6BEG[6]
+ Tile_X0Y0_W6BEG[7] Tile_X0Y0_W6BEG[8] Tile_X0Y0_W6BEG[9] Tile_X0Y0_WW4BEG[0] Tile_X0Y0_WW4BEG[10]
+ Tile_X0Y0_WW4BEG[11] Tile_X0Y0_WW4BEG[12] Tile_X0Y0_WW4BEG[13] Tile_X0Y0_WW4BEG[14]
+ Tile_X0Y0_WW4BEG[15] Tile_X0Y0_WW4BEG[1] Tile_X0Y0_WW4BEG[2] Tile_X0Y0_WW4BEG[3]
+ Tile_X0Y0_WW4BEG[4] Tile_X0Y0_WW4BEG[5] Tile_X0Y0_WW4BEG[6] Tile_X0Y0_WW4BEG[7]
+ Tile_X0Y0_WW4BEG[8] Tile_X0Y0_WW4BEG[9] Tile_X0Y1_E1END[0] Tile_X0Y1_E1END[1] Tile_X0Y1_E1END[2]
+ Tile_X0Y1_E1END[3] Tile_X0Y1_E2END[0] Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2] Tile_X0Y1_E2END[3]
+ Tile_X0Y1_E2END[4] Tile_X0Y1_E2END[5] Tile_X0Y1_E2END[6] Tile_X0Y1_E2END[7] Tile_X0Y1_E2MID[0]
+ Tile_X0Y1_E2MID[1] Tile_X0Y1_E2MID[2] Tile_X0Y1_E2MID[3] Tile_X0Y1_E2MID[4] Tile_X0Y1_E2MID[5]
+ Tile_X0Y1_E2MID[6] Tile_X0Y1_E2MID[7] Tile_X0Y1_E6END[0] Tile_X0Y1_E6END[10] Tile_X0Y1_E6END[11]
+ Tile_X0Y1_E6END[1] Tile_X0Y1_E6END[2] Tile_X0Y1_E6END[3] Tile_X0Y1_E6END[4] Tile_X0Y1_E6END[5]
+ Tile_X0Y1_E6END[6] Tile_X0Y1_E6END[7] Tile_X0Y1_E6END[8] Tile_X0Y1_E6END[9] Tile_X0Y1_EE4END[0]
+ Tile_X0Y1_EE4END[10] Tile_X0Y1_EE4END[11] Tile_X0Y1_EE4END[12] Tile_X0Y1_EE4END[13]
+ Tile_X0Y1_EE4END[14] Tile_X0Y1_EE4END[15] Tile_X0Y1_EE4END[1] Tile_X0Y1_EE4END[2]
+ Tile_X0Y1_EE4END[3] Tile_X0Y1_EE4END[4] Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[6]
+ Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[8] Tile_X0Y1_EE4END[9] Tile_X0Y1_FrameData[0]
+ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData[13]
+ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData[17]
+ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData[20]
+ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData[24]
+ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData[28]
+ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData[31]
+ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData[6]
+ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[0]
+ Tile_X0Y1_FrameData_O[10] Tile_X0Y1_FrameData_O[11] Tile_X0Y1_FrameData_O[12] Tile_X0Y1_FrameData_O[13]
+ Tile_X0Y1_FrameData_O[14] Tile_X0Y1_FrameData_O[15] Tile_X0Y1_FrameData_O[16] Tile_X0Y1_FrameData_O[17]
+ Tile_X0Y1_FrameData_O[18] Tile_X0Y1_FrameData_O[19] Tile_X0Y1_FrameData_O[1] Tile_X0Y1_FrameData_O[20]
+ Tile_X0Y1_FrameData_O[21] Tile_X0Y1_FrameData_O[22] Tile_X0Y1_FrameData_O[23] Tile_X0Y1_FrameData_O[24]
+ Tile_X0Y1_FrameData_O[25] Tile_X0Y1_FrameData_O[26] Tile_X0Y1_FrameData_O[27] Tile_X0Y1_FrameData_O[28]
+ Tile_X0Y1_FrameData_O[29] Tile_X0Y1_FrameData_O[2] Tile_X0Y1_FrameData_O[30] Tile_X0Y1_FrameData_O[31]
+ Tile_X0Y1_FrameData_O[3] Tile_X0Y1_FrameData_O[4] Tile_X0Y1_FrameData_O[5] Tile_X0Y1_FrameData_O[6]
+ Tile_X0Y1_FrameData_O[7] Tile_X0Y1_FrameData_O[8] Tile_X0Y1_FrameData_O[9] Tile_X0Y1_FrameStrobe[0]
+ Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_FrameStrobe[13]
+ Tile_X0Y1_FrameStrobe[14] Tile_X0Y1_FrameStrobe[15] Tile_X0Y1_FrameStrobe[16] Tile_X0Y1_FrameStrobe[17]
+ Tile_X0Y1_FrameStrobe[18] Tile_X0Y1_FrameStrobe[19] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_FrameStrobe[2]
+ Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_FrameStrobe[6]
+ Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_N1END[0]
+ Tile_X0Y1_N1END[1] Tile_X0Y1_N1END[2] Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[0] Tile_X0Y1_N2END[1]
+ Tile_X0Y1_N2END[2] Tile_X0Y1_N2END[3] Tile_X0Y1_N2END[4] Tile_X0Y1_N2END[5] Tile_X0Y1_N2END[6]
+ Tile_X0Y1_N2END[7] Tile_X0Y1_N2MID[0] Tile_X0Y1_N2MID[1] Tile_X0Y1_N2MID[2] Tile_X0Y1_N2MID[3]
+ Tile_X0Y1_N2MID[4] Tile_X0Y1_N2MID[5] Tile_X0Y1_N2MID[6] Tile_X0Y1_N2MID[7] Tile_X0Y1_N4END[0]
+ Tile_X0Y1_N4END[10] Tile_X0Y1_N4END[11] Tile_X0Y1_N4END[12] Tile_X0Y1_N4END[13]
+ Tile_X0Y1_N4END[14] Tile_X0Y1_N4END[15] Tile_X0Y1_N4END[1] Tile_X0Y1_N4END[2] Tile_X0Y1_N4END[3]
+ Tile_X0Y1_N4END[4] Tile_X0Y1_N4END[5] Tile_X0Y1_N4END[6] Tile_X0Y1_N4END[7] Tile_X0Y1_N4END[8]
+ Tile_X0Y1_N4END[9] Tile_X0Y1_S1BEG[0] Tile_X0Y1_S1BEG[1] Tile_X0Y1_S1BEG[2] Tile_X0Y1_S1BEG[3]
+ Tile_X0Y1_S2BEG[0] Tile_X0Y1_S2BEG[1] Tile_X0Y1_S2BEG[2] Tile_X0Y1_S2BEG[3] Tile_X0Y1_S2BEG[4]
+ Tile_X0Y1_S2BEG[5] Tile_X0Y1_S2BEG[6] Tile_X0Y1_S2BEG[7] Tile_X0Y1_S2BEGb[0] Tile_X0Y1_S2BEGb[1]
+ Tile_X0Y1_S2BEGb[2] Tile_X0Y1_S2BEGb[3] Tile_X0Y1_S2BEGb[4] Tile_X0Y1_S2BEGb[5]
+ Tile_X0Y1_S2BEGb[6] Tile_X0Y1_S2BEGb[7] Tile_X0Y1_S4BEG[0] Tile_X0Y1_S4BEG[10] Tile_X0Y1_S4BEG[11]
+ Tile_X0Y1_S4BEG[12] Tile_X0Y1_S4BEG[13] Tile_X0Y1_S4BEG[14] Tile_X0Y1_S4BEG[15]
+ Tile_X0Y1_S4BEG[1] Tile_X0Y1_S4BEG[2] Tile_X0Y1_S4BEG[3] Tile_X0Y1_S4BEG[4] Tile_X0Y1_S4BEG[5]
+ Tile_X0Y1_S4BEG[6] Tile_X0Y1_S4BEG[7] Tile_X0Y1_S4BEG[8] Tile_X0Y1_S4BEG[9] Tile_X0Y1_UserCLK
+ Tile_X0Y1_W1BEG[0] Tile_X0Y1_W1BEG[1] Tile_X0Y1_W1BEG[2] Tile_X0Y1_W1BEG[3] Tile_X0Y1_W2BEG[0]
+ Tile_X0Y1_W2BEG[1] Tile_X0Y1_W2BEG[2] Tile_X0Y1_W2BEG[3] Tile_X0Y1_W2BEG[4] Tile_X0Y1_W2BEG[5]
+ Tile_X0Y1_W2BEG[6] Tile_X0Y1_W2BEG[7] Tile_X0Y1_W2BEGb[0] Tile_X0Y1_W2BEGb[1] Tile_X0Y1_W2BEGb[2]
+ Tile_X0Y1_W2BEGb[3] Tile_X0Y1_W2BEGb[4] Tile_X0Y1_W2BEGb[5] Tile_X0Y1_W2BEGb[6]
+ Tile_X0Y1_W2BEGb[7] Tile_X0Y1_W6BEG[0] Tile_X0Y1_W6BEG[10] Tile_X0Y1_W6BEG[11] Tile_X0Y1_W6BEG[1]
+ Tile_X0Y1_W6BEG[2] Tile_X0Y1_W6BEG[3] Tile_X0Y1_W6BEG[4] Tile_X0Y1_W6BEG[5] Tile_X0Y1_W6BEG[6]
+ Tile_X0Y1_W6BEG[7] Tile_X0Y1_W6BEG[8] Tile_X0Y1_W6BEG[9] Tile_X0Y1_WW4BEG[0] Tile_X0Y1_WW4BEG[10]
+ Tile_X0Y1_WW4BEG[11] Tile_X0Y1_WW4BEG[12] Tile_X0Y1_WW4BEG[13] Tile_X0Y1_WW4BEG[14]
+ Tile_X0Y1_WW4BEG[15] Tile_X0Y1_WW4BEG[1] Tile_X0Y1_WW4BEG[2] Tile_X0Y1_WW4BEG[3]
+ Tile_X0Y1_WW4BEG[4] Tile_X0Y1_WW4BEG[5] Tile_X0Y1_WW4BEG[6] Tile_X0Y1_WW4BEG[7]
+ Tile_X0Y1_WW4BEG[8] Tile_X0Y1_WW4BEG[9] VGND VPWR
X_0367_ net10 net19 net363 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit24.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit25.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb1
+ sky130_fd_sc_hd__mux4_1
X_0298_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit30.Q _0070_
+ _0002_ _0069_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_65_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1270_ net455 net375 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_95_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0221_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit27.Q VGND
+ VGND VPWR VPWR _0000_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_19_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0985_ net84 net377 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput401 net518 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput412 net529 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput423 net540 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[5] sky130_fd_sc_hd__buf_2
Xoutput434 net551 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[0] sky130_fd_sc_hd__buf_2
Xoutput456 net573 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput445 net562 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[9] sky130_fd_sc_hd__buf_2
Xoutput467 net584 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[14] sky130_fd_sc_hd__buf_2
Xoutput478 net595 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[24] sky130_fd_sc_hd__buf_2
X_1537_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb5 VGND VGND VPWR
+ VPWR net664 sky130_fd_sc_hd__buf_1
Xoutput489 net606 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[5] sky130_fd_sc_hd__buf_2
X_1468_ Tile_X0Y1_FrameData[16] VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1399_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG0 VGND VGND VPWR
+ VPWR net517 sky130_fd_sc_hd__clkbuf_2
X_0419_ net75 net68 net59 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG4
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit6.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit7.Q
+ VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__mux4_1
XFILLER_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0770_ net106 net436 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_154_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1322_ net110 VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__clkbuf_1
X_1253_ net190 net383 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_56_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1184_ net465 net398 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0968_ net469 net377 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0899_ net103 net405 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput253 net253 VGND VGND VPWR VPWR AD_SRAM5 sky130_fd_sc_hd__buf_2
Xoutput286 net286 VGND VGND VPWR VPWR BEN_SRAM6 sky130_fd_sc_hd__buf_2
Xoutput264 net264 VGND VGND VPWR VPWR BEN_SRAM14 sky130_fd_sc_hd__buf_2
Xoutput275 net275 VGND VGND VPWR VPWR BEN_SRAM24 sky130_fd_sc_hd__buf_2
Xoutput297 net297 VGND VGND VPWR VPWR DI_SRAM14 sky130_fd_sc_hd__buf_2
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_122_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_140_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0822_ net87 net420 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0753_ net93 net437 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_115_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0684_ _0052_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG0 _0196_ VGND VGND VPWR
+ VPWR _0197_ sky130_fd_sc_hd__o31a_1
XFILLER_142_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1305_ net458 net370 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_96_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1236_ net453 net382 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1167_ net189 net408 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_143_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1098_ net214 net425 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_306 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1021_ net462 net440 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_75_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0805_ net81 net428 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0736_ net108 net446 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0667_ _0044_ _0182_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q
+ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__a21o_1
XFILLER_103_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0598_ _0026_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q
+ net366 _0152_ VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__a31o_1
X_1219_ net192 net390 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_44_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_5 net272 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0521_ net158 net150 net162 _0078_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_152_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0452_ _0094_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit1.Q
+ _0004_ _0093_ VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__a2bb2o_2
X_0383_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END1 net245 net114
+ net134 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit26.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit27.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG9
+ sky130_fd_sc_hd__mux4_2
XFILLER_26_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1004_ net473 net372 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_34_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0719_ net476 net445 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput120 Tile_X0Y0_S2END[3] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_2
XFILLER_95_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput131 Tile_X0Y0_S2MID[6] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
Xinput142 Tile_X0Y1_E1END[1] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__buf_2
Xinput153 Tile_X0Y1_E2MID[0] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
Xinput186 Tile_X0Y1_EE4END[7] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_2
Xinput175 Tile_X0Y1_EE4END[11] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput164 Tile_X0Y1_E6END[1] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__buf_1
XFILLER_102_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput197 Tile_X0Y1_FrameData[19] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1553_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG1 VGND VGND VPWR
+ VPWR net686 sky130_fd_sc_hd__buf_1
XFILLER_140_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0504_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG7 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit27.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit28.Q
+ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__mux4_1
X_1484_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG0 VGND VGND VPWR
+ VPWR net611 sky130_fd_sc_hd__clkbuf_2
XFILLER_140_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0435_ net75 net68 net59 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG4
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit6.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit7.Q
+ VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__mux4_2
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0366_ net9 net18 net364 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit22.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit23.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb0
+ sky130_fd_sc_hd__mux4_1
XFILLER_39_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0297_ net116 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit31.Q
+ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__nand2_1
XFILLER_22_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0984_ net85 net377 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput402 net519 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[14] sky130_fd_sc_hd__buf_2
XFILLER_8_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput413 net530 VGND VGND VPWR VPWR Tile_X0Y0_UserCLKo sky130_fd_sc_hd__buf_1
Xoutput424 net541 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[6] sky130_fd_sc_hd__buf_2
Xoutput435 net552 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[10] sky130_fd_sc_hd__buf_2
X_1536_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb4 VGND VGND VPWR
+ VPWR net663 sky130_fd_sc_hd__buf_1
Xoutput446 net563 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput457 net574 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput468 net585 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[15] sky130_fd_sc_hd__buf_2
Xoutput479 net596 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[25] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_26_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1467_ net465 VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__buf_4
X_0418_ net74 net67 net58 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG3
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit4.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit5.Q
+ VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__mux4_2
X_1398_ Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_11.A VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__buf_4
XFILLER_86_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0349_ net33 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12 net63
+ _0086_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit27.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit26.Q
+ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__mux4_2
XFILLER_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_146_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1321_ net109 VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__buf_1
XFILLER_68_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1252_ net191 net384 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1183_ net464 net398 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0967_ net468 net379 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0898_ net106 net405 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput254 net254 VGND VGND VPWR VPWR AD_SRAM6 sky130_fd_sc_hd__buf_2
XFILLER_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput265 net265 VGND VGND VPWR VPWR BEN_SRAM15 sky130_fd_sc_hd__buf_2
Xoutput276 net276 VGND VGND VPWR VPWR BEN_SRAM25 sky130_fd_sc_hd__buf_2
X_1519_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG3 VGND VGND VPWR
+ VPWR net637 sky130_fd_sc_hd__buf_1
Xoutput287 net287 VGND VGND VPWR VPWR BEN_SRAM7 sky130_fd_sc_hd__buf_2
Xoutput298 net298 VGND VGND VPWR VPWR DI_SRAM15 sky130_fd_sc_hd__buf_2
XFILLER_99_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout470 net101 VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__clkbuf_4
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0821_ net88 net421 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0752_ net94 net439 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_127_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0683_ net149 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q _0195_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
+ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__o311a_1
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1304_ net457 net370 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_96_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1235_ net452 net383 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_49_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1166_ net198 net409 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_143_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1097_ net215 net425 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1020_ net461 net441 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_75_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0804_ net92 net428 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0735_ net109 net446 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0666_ net142 net177 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q
+ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__mux2_1
XFILLER_69_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0597_ net148 _0026_ _0151_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__o21a_1
XFILLER_69_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1218_ net193 net390 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1149_ net462 net408 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_6 net273 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0520_ net159 net151 net172 _0077_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_152_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0451_ net38 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit0.Q
+ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__nand2_1
X_0382_ net15 net19 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit16.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit17.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG5 sky130_fd_sc_hd__mux4_1
XFILLER_66_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1003_ net472 net372 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_77_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0718_ net475 net445 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0649_ _0035_ _0167_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q
+ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__a21o_1
XFILLER_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput110 Tile_X0Y0_FrameData[7] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_4
Xinput121 Tile_X0Y0_S2END[4] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput132 Tile_X0Y0_S2MID[7] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
Xinput143 Tile_X0Y1_E1END[2] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_2
Xinput154 Tile_X0Y1_E2MID[1] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
Xinput176 Tile_X0Y1_EE4END[12] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_2
Xinput187 Tile_X0Y1_EE4END[8] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_2
Xinput165 Tile_X0Y1_E6END[2] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_1
Xinput198 Tile_X0Y1_FrameData[1] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__buf_4
XFILLER_63_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1552_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG0 VGND VGND VPWR
+ VPWR net679 sky130_fd_sc_hd__clkbuf_2
X_0503_ _0016_ _0131_ _0135_ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG2
+ sky130_fd_sc_hd__o21a_1
X_1483_ net449 VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__buf_2
XFILLER_140_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0434_ net74 net67 net58 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG3
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit4.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit5.Q
+ VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0365_ net17 net26 net364 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit20.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit21.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG7
+ sky130_fd_sc_hd__mux4_1
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0296_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END3 net58 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit30.Q
+ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0983_ net86 net380 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput403 net520 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[15] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_10_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput414 net531 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[0] sky130_fd_sc_hd__buf_2
Xoutput425 net542 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[7] sky130_fd_sc_hd__buf_2
X_1535_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb3 VGND VGND VPWR
+ VPWR net662 sky130_fd_sc_hd__buf_1
Xoutput458 net575 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput447 net564 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput436 net553 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[11] sky130_fd_sc_hd__buf_2
Xoutput469 net586 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[16] sky130_fd_sc_hd__buf_2
X_1466_ net466 VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__buf_4
XFILLER_86_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0417_ net73 net66 net57 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG2
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit2.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit3.Q
+ VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__mux4_2
X_1397_ Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_10.A VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_2_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0348_ _0019_ _0084_ _0085_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_146_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0279_ net34 net64 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13
+ _0057_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit28.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit29.Q
+ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_105_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1320_ net108 VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__clkbuf_2
X_1251_ net192 net383 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1182_ net463 net398 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_91_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0966_ net467 net379 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_133_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0897_ net107 net405 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput255 net255 VGND VGND VPWR VPWR AD_SRAM7 sky130_fd_sc_hd__buf_2
Xoutput266 net266 VGND VGND VPWR VPWR BEN_SRAM16 sky130_fd_sc_hd__buf_2
Xoutput277 net277 VGND VGND VPWR VPWR BEN_SRAM26 sky130_fd_sc_hd__buf_2
XFILLER_99_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1518_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG2 VGND VGND VPWR
+ VPWR net636 sky130_fd_sc_hd__buf_1
Xoutput288 net288 VGND VGND VPWR VPWR BEN_SRAM8 sky130_fd_sc_hd__buf_2
Xoutput299 net299 VGND VGND VPWR VPWR DI_SRAM16 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_98_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1449_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG13 VGND VGND VPWR
+ VPWR net567 sky130_fd_sc_hd__clkbuf_1
XFILLER_114_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout460 net199 VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__clkbuf_4
Xfanout471 net100 VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__buf_4
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0820_ net89 net421 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0751_ net476 net438 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_115_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0682_ net128 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q VGND VGND VPWR
+ VPWR _0195_ sky130_fd_sc_hd__or3b_1
X_1303_ net456 net370 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1234_ net451 net383 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_96_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1165_ net209 net408 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_64_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1096_ net216 net426 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_35_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0949_ net88 net385 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0803_ net103 net428 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_115_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0734_ net110 net446 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0665_ _0043_ _0143_ _0180_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q
+ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__o211a_1
X_0596_ net156 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q VGND VGND VPWR
+ VPWR _0151_ sky130_fd_sc_hd__o21ba_1
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1217_ net466 net390 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1148_ net461 net408 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1079_ net456 net424 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_80_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_119_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_7 net276 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_128_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0450_ net46 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit1.Q
+ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__mux2_1
XFILLER_112_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0381_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END2 net246 net115
+ net135 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit28.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit29.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG10
+ sky130_fd_sc_hd__mux4_2
XFILLER_66_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1002_ net471 net372 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_77_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_137_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0717_ net97 net448 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0648_ net143 net181 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q
+ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__mux2_1
X_0579_ net27 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG11 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG7
+ net369 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG4
+ sky130_fd_sc_hd__mux4_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput100 Tile_X0Y0_FrameData[27] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_2
Xinput111 Tile_X0Y0_FrameData[8] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_4
Xinput133 Tile_X0Y0_S4END[0] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
Xinput122 Tile_X0Y0_S2END[5] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput144 Tile_X0Y1_E1END[3] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_2
Xinput155 Tile_X0Y1_E2MID[2] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput177 Tile_X0Y1_EE4END[13] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput166 Tile_X0Y1_E6END[3] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
Xinput188 Tile_X0Y1_EE4END[9] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__buf_1
Xinput199 Tile_X0Y1_FrameData[20] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__buf_1
XFILLER_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1551_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG11 VGND VGND VPWR
+ VPWR net669 sky130_fd_sc_hd__buf_1
X_0502_ _0132_ _0133_ _0134_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit25.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit26.Q VGND VGND VPWR
+ VPWR _0135_ sky130_fd_sc_hd__a221o_1
X_1482_ net450 VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__buf_2
X_0433_ net73 net66 net57 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG2
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit2.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit3.Q
+ VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__mux4_2
XFILLER_86_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_145_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0364_ net16 net25 net363 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit18.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit19.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG6
+ sky130_fd_sc_hd__mux4_1
X_0295_ net35 net61 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14
+ _0064_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit26.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit27.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG2
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_65_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_154_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0982_ net87 net380 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput404 net521 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_10_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput415 net532 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[1] sky130_fd_sc_hd__buf_2
Xoutput426 net543 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[0] sky130_fd_sc_hd__buf_2
X_1534_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb2 VGND VGND VPWR
+ VPWR net661 sky130_fd_sc_hd__buf_1
Xoutput459 net576 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput448 net565 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput437 net554 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[1] sky130_fd_sc_hd__buf_2
X_1465_ net193 VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__buf_4
X_0416_ net72 net80 net56 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG1
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit0.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit1.Q
+ VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__mux4_2
X_1396_ Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_9.A VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__buf_4
X_0347_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit24.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit25.Q
+ net113 VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__and3b_1
X_0278_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit26.Q _0056_
+ _0000_ _0055_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1250_ net193 net389 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1181_ net462 net400 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_91_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0965_ net81 net387 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0896_ net108 net405 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_133_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput256 net256 VGND VGND VPWR VPWR AD_SRAM8 sky130_fd_sc_hd__buf_2
Xoutput267 net267 VGND VGND VPWR VPWR BEN_SRAM17 sky130_fd_sc_hd__buf_2
Xoutput289 net289 VGND VGND VPWR VPWR BEN_SRAM9 sky130_fd_sc_hd__buf_2
Xoutput278 net278 VGND VGND VPWR VPWR BEN_SRAM27 sky130_fd_sc_hd__buf_2
X_1517_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG1 VGND VGND VPWR
+ VPWR net635 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_98_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1448_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG12 VGND VGND VPWR
+ VPWR net566 sky130_fd_sc_hd__clkbuf_2
XFILLER_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1379_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb0 VGND VGND VPWR
+ VPWR net506 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_81_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout450 net210 VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__buf_4
Xfanout461 net197 VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__clkbuf_4
Xfanout472 net99 VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_100_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0750_ net475 net438 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_127_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0681_ _0191_ _0193_ _0194_ _0051_ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG3
+ sky130_fd_sc_hd__o22a_1
XFILLER_115_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1302_ net455 net370 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_96_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1233_ net450 net381 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1164_ net212 net408 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1095_ net217 net424 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_64_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0948_ net89 net385 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_154_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0879_ net476 net402 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_133_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0802_ net106 net428 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_40_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0733_ net111 net444 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0664_ net168 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q
+ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__or2_1
XFILLER_115_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0595_ _0025_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q
+ net367 _0150_ VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__a31o_1
XFILLER_69_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1216_ net465 net390 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1147_ net460 net407 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1078_ net455 net424 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_115_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_8 net277 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0380_ net14 net18 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG11
+ net361 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit14.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit15.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG4
+ sky130_fd_sc_hd__mux4_1
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1001_ net470 net372 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_34_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0716_ net98 net448 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0647_ _0034_ _0142_ _0165_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q
+ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__o211a_1
XFILLER_103_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0578_ net243 net140 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG8
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG3 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_68_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput101 Tile_X0Y0_FrameData[28] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
Xinput134 Tile_X0Y0_S4END[1] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__buf_2
Xinput123 Tile_X0Y0_S2END[6] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
Xinput112 Tile_X0Y0_FrameData[9] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_4
Xinput145 Tile_X0Y1_E2END[0] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput156 Tile_X0Y1_E2MID[3] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
Xinput178 Tile_X0Y1_EE4END[14] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput167 Tile_X0Y1_E6END[4] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_2
Xinput189 Tile_X0Y1_FrameData[0] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__buf_4
XFILLER_56_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1550_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG10 VGND VGND VPWR
+ VPWR net668 sky130_fd_sc_hd__clkbuf_1
X_0501_ net61 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG2 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit24.Q
+ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__mux2_1
X_1481_ net451 VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__buf_4
X_0432_ net72 net80 net56 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG1
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit0.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit1.Q
+ VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__mux4_2
XFILLER_140_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0363_ net15 net23 net362 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit16.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit17.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG5
+ sky130_fd_sc_hd__mux4_1
XFILLER_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0294_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END2 net246 net115
+ net135 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit4.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit5.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14
+ sky130_fd_sc_hd__mux4_2
XFILLER_47_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0981_ net88 net380 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput405 net522 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_10_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput416 net533 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[2] sky130_fd_sc_hd__buf_2
X_1533_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb1 VGND VGND VPWR
+ VPWR net660 sky130_fd_sc_hd__clkbuf_1
Xoutput427 net544 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput449 net566 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput438 net555 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1464_ net192 VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__buf_4
X_0415_ net65 net79 net53 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG0
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit30.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit31.Q
+ VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__mux4_1
XFILLER_113_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1395_ Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_8.A VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__buf_4
XFILLER_79_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0346_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END0 net53 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit24.Q
+ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__mux2_1
XFILLER_94_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0277_ net114 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit27.Q
+ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__nand2_1
XFILLER_35_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_13_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1180_ net461 net400 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_64_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0964_ net92 net387 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0895_ net109 net405 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1516_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG0 VGND VGND VPWR
+ VPWR net634 sky130_fd_sc_hd__buf_1
Xoutput257 net257 VGND VGND VPWR VPWR AD_SRAM9 sky130_fd_sc_hd__buf_2
Xoutput268 net268 VGND VGND VPWR VPWR BEN_SRAM18 sky130_fd_sc_hd__buf_2
XFILLER_99_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput279 net279 VGND VGND VPWR VPWR BEN_SRAM28 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_98_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1447_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG11 VGND VGND VPWR
+ VPWR net565 sky130_fd_sc_hd__buf_1
X_1378_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG7 VGND VGND VPWR
+ VPWR net505 sky130_fd_sc_hd__buf_4
X_0329_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb4 net129 net236
+ net121 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit17.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit16.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG4
+ sky130_fd_sc_hd__mux4_1
XFILLER_82_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout440 net443 VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__buf_2
Xfanout451 net208 VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__clkbuf_4
Xfanout462 net196 VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__clkbuf_4
Xfanout473 net98 VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__clkbuf_4
XFILLER_104_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0680_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG7
+ _0083_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG11 _0050_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q
+ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__mux4_1
X_1301_ net454 net371 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1232_ net449 net381 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1163_ net213 net409 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_64_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1094_ net218 net424 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_64_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0947_ net90 net388 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_154_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0878_ net475 net402 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0801_ net107 net427 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_40_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0732_ net112 net444 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0663_ _0176_ _0178_ _0179_ _0042_ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG0
+ sky130_fd_sc_hd__o22a_1
X_0594_ net147 _0025_ _0149_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__o21a_1
XFILLER_123_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1215_ net464 net392 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1146_ net459 net408 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_92_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1077_ net454 net426 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 net278 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_5_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1000_ net469 net219 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_34_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0715_ net472 net446 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0646_ net162 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q
+ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__or2_1
X_0577_ net242 net139 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG9
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1129_ net215 net417 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_15_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput102 Tile_X0Y0_FrameData[29] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput124 Tile_X0Y0_S2END[7] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
Xinput113 Tile_X0Y0_S1END[0] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_2
Xinput135 Tile_X0Y0_S4END[2] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput157 Tile_X0Y1_E2MID[4] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
Xinput146 Tile_X0Y1_E2END[1] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_2
Xinput168 Tile_X0Y1_E6END[5] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput179 Tile_X0Y1_EE4END[15] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0500_ net35 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit24.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit25.Q VGND VGND VPWR
+ VPWR _0133_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1480_ net452 VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__buf_4
XFILLER_98_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0431_ net65 net79 net53 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG0
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit30.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit31.Q
+ VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__mux4_1
XFILLER_98_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0362_ net14 net22 net361 net360 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit14.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit15.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG4 sky130_fd_sc_hd__mux4_1
XFILLER_94_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0293_ net143 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14 net169
+ _0068_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit19.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit18.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END2
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_65_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0629_ net182 net175 net163 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG11
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q
+ VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__mux4_2
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_77_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_95_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0980_ net89 net378 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_145_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput406 net523 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_10_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput417 net534 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[3] sky130_fd_sc_hd__buf_2
X_1532_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb0 VGND VGND VPWR
+ VPWR net659 sky130_fd_sc_hd__buf_1
Xoutput428 net545 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput439 net556 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[3] sky130_fd_sc_hd__buf_2
X_1463_ net191 VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__buf_4
XFILLER_79_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0414_ net12 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG0
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit29.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit28.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG11 sky130_fd_sc_hd__mux4_1
X_1394_ Tile_X0Y1_N4END[15] VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__buf_4
X_0345_ net45 net37 net53 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit12.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit13.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG7
+ sky130_fd_sc_hd__mux4_1
X_0276_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END1 net56 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit26.Q
+ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__mux2_1
XFILLER_35_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0963_ net103 net385 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_110_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0894_ net110 net405 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1515_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG3 VGND VGND VPWR
+ VPWR net633 sky130_fd_sc_hd__buf_4
Xoutput258 net258 VGND VGND VPWR VPWR BEN_SRAM0 sky130_fd_sc_hd__buf_2
Xoutput269 net269 VGND VGND VPWR VPWR BEN_SRAM19 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_98_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1446_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG10 VGND VGND VPWR
+ VPWR net564 sky130_fd_sc_hd__clkbuf_1
X_1377_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG6 VGND VGND VPWR
+ VPWR net504 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0328_ net156 net148 net166 _0080_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit30.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit31.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb4 sky130_fd_sc_hd__mux4_1
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0259_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q VGND
+ VGND VPWR VPWR _0038_ sky130_fd_sc_hd__inv_2
XFILLER_82_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout441 net443 VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkbuf_4
Xfanout430 net431 VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__buf_2
Xfanout463 Tile_X0Y1_FrameData[17] VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__buf_4
Xfanout452 net207 VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout474 net97 VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1300_ net453 net371 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1231_ net189 net392 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1162_ net214 net409 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1093_ net190 net426 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_32_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0946_ net91 net388 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_154_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0877_ net474 net404 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_125_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1429_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG5 VGND VGND VPWR
+ VPWR net558 sky130_fd_sc_hd__buf_1
XFILLER_141_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0800_ net108 net427 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_40_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0731_ net82 net444 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_155_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0662_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG4
+ net365 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG8 _0041_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q
+ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__mux4_1
XFILLER_115_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0593_ net155 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q VGND VGND VPWR
+ VPWR _0149_ sky130_fd_sc_hd__o21ba_1
XFILLER_69_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1214_ net463 net392 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1145_ net458 net408 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_92_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1076_ net453 net426 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_40_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0929_ net107 net397 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_114_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0714_ net471 net446 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0645_ _0161_ _0163_ _0164_ _0033_ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_9.A
+ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_115_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0576_ net241 net138 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG10
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1128_ net216 net417 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_124_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1059_ net192 net433 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_133_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput136 Tile_X0Y0_S4END[3] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
Xinput125 Tile_X0Y0_S2MID[0] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
Xinput114 Tile_X0Y0_S1END[1] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__buf_2
Xinput103 Tile_X0Y0_FrameData[2] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput158 Tile_X0Y1_E2MID[5] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput147 Tile_X0Y1_E2END[2] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
Xinput169 Tile_X0Y1_E6END[6] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_2
XFILLER_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0430_ net36 net78 net71 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit28.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit29.Q
+ VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__mux4_2
XFILLER_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0361_ net12 net21 net361 net360 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit12.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit13.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG3 sky130_fd_sc_hd__mux4_1
X_0292_ _0021_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q
+ _0065_ _0067_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__a31o_1
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0628_ net181 net174 net162 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG10
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q
+ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__mux4_2
X_0559_ net223 net243 _0072_ net140 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG7 sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_96_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput407 net524 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_10_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1531_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG7 VGND VGND VPWR
+ VPWR net658 sky130_fd_sc_hd__buf_1
Xoutput418 net535 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput429 net546 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[3] sky130_fd_sc_hd__buf_2
X_1462_ net190 VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__buf_4
X_0413_ net11 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG1
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit27.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit26.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG10 sky130_fd_sc_hd__mux4_1
XFILLER_113_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1393_ Tile_X0Y1_N4END[14] VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__buf_4
X_0344_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb7 net132 net239
+ net124 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit23.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit22.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7
+ sky130_fd_sc_hd__mux4_2
X_0275_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q VGND VGND
+ VPWR VPWR _0054_ sky130_fd_sc_hd__inv_2
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0962_ net106 net385 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_110_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0893_ net111 net404 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_145_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1514_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG2 VGND VGND VPWR
+ VPWR net632 sky130_fd_sc_hd__buf_4
Xoutput248 net248 VGND VGND VPWR VPWR AD_SRAM0 sky130_fd_sc_hd__buf_2
Xoutput259 net259 VGND VGND VPWR VPWR BEN_SRAM1 sky130_fd_sc_hd__buf_2
XFILLER_59_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1445_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG9 VGND VGND VPWR
+ VPWR net578 sky130_fd_sc_hd__buf_1
XFILLER_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1376_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG5 VGND VGND VPWR
+ VPWR net503 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0327_ net236 net228 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG4
+ net129 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q
+ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__mux4_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0258_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q VGND
+ VGND VPWR VPWR _0037_ sky130_fd_sc_hd__inv_1
XFILLER_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout420 net423 VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__buf_2
Xfanout431 Tile_X0Y1_FrameStrobe[2] VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__clkbuf_4
Xfanout475 net96 VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__clkbuf_4
Xfanout464 Tile_X0Y1_FrameData[16] VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__buf_4
XFILLER_48_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout453 net206 VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__clkbuf_4
Xfanout442 net443 VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__buf_2
XFILLER_58_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1230_ net198 net392 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1161_ net215 net407 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1092_ net191 net426 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_52_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0945_ net93 net388 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_154_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0876_ net473 net404 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_125_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1428_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG4 VGND VGND VPWR
+ VPWR net557 sky130_fd_sc_hd__clkbuf_2
X_1359_ Tile_X0Y1_FrameStrobe[12] VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__clkbuf_1
XFILLER_141_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0730_ net83 net444 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_155_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0661_ _0041_ _0177_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q
+ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__a21o_1
X_0592_ _0024_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q
+ net368 _0148_ VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__a31o_1
XFILLER_108_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1213_ net462 net392 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_77_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1144_ net457 net408 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1075_ net452 net431 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_92_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0928_ net108 net397 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0859_ net82 net413 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0713_ net101 net447 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0644_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG5
+ net368 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG9 _0032_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q
+ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__mux4_1
X_0575_ net240 net137 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG11
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1127_ net217 net416 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1058_ net193 net433 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_33_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput126 Tile_X0Y0_S2MID[1] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
Xinput115 Tile_X0Y0_S1END[2] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_2
Xinput104 Tile_X0Y0_FrameData[30] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_2
Xinput137 Tile_X0Y0_S4END[4] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_4
Xinput159 Tile_X0Y1_E2MID[6] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
Xinput148 Tile_X0Y1_E2END[3] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0360_ net11 net20 net362 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit10.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit11.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG2
+ sky130_fd_sc_hd__mux4_1
X_0291_ net165 _0021_ _0066_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__o21a_1
XFILLER_153_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0627_ net180 net188 net172 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG9
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q
+ VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__mux4_2
X_0558_ net30 net4 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG8
+ net369 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG7
+ sky130_fd_sc_hd__mux4_1
X_0489_ net59 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG0 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit18.Q
+ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_22 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput408 net525 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_10_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1530_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG6 VGND VGND VPWR
+ VPWR net657 sky130_fd_sc_hd__buf_1
Xoutput419 net536 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[1] sky130_fd_sc_hd__buf_2
X_1461_ net218 VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__buf_4
X_1392_ Tile_X0Y1_N4END[13] VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__buf_4
XFILLER_79_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0412_ net10 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG6 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG2
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit25.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit24.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG9 sky130_fd_sc_hd__mux4_1
X_0343_ net153 net145 net161 _0083_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb7 sky130_fd_sc_hd__mux4_2
XFILLER_94_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0274_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q VGND VGND
+ VPWR VPWR _0053_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_18_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_151_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0961_ net107 net386 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0892_ net112 net404 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_110_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1513_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG1 VGND VGND VPWR
+ VPWR net646 sky130_fd_sc_hd__buf_4
Xoutput249 net249 VGND VGND VPWR VPWR AD_SRAM1 sky130_fd_sc_hd__buf_2
XFILLER_99_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1444_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG8 VGND VGND VPWR
+ VPWR net577 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1375_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG4 VGND VGND VPWR
+ VPWR net502 sky130_fd_sc_hd__clkbuf_2
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0326_ net33 net40 net48 net360 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit11.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit10.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG4 sky130_fd_sc_hd__mux4_2
X_0257_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q VGND
+ VGND VPWR VPWR _0036_ sky130_fd_sc_hd__inv_1
XFILLER_82_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout421 net423 VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__buf_2
Xfanout432 net433 VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__clkbuf_2
Xfanout410 Tile_X0Y1_FrameStrobe[4] VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__buf_2
Xfanout454 net205 VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__clkbuf_4
Xfanout465 net195 VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__clkbuf_4
Xfanout443 Tile_X0Y1_FrameStrobe[0] VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__clkbuf_2
Xfanout476 net95 VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1160_ net216 net407 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_49_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1091_ net192 net431 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_43_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0944_ net94 net386 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0875_ net472 net402 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_154_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1427_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG3 VGND VGND VPWR
+ VPWR net556 sky130_fd_sc_hd__buf_1
X_1358_ Tile_X0Y1_FrameStrobe[11] VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__clkbuf_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1289_ net215 net375 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0309_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb0 net125 net232
+ net117 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit9.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit8.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG0
+ sky130_fd_sc_hd__mux4_1
XFILLER_70_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0660_ net141 net176 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q
+ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__mux2_1
X_0591_ net146 _0024_ _0147_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__o21a_1
XFILLER_111_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1212_ net461 net392 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1143_ net456 net410 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_77_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1074_ net451 net431 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_52_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0927_ net109 net395 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0858_ net83 net413 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0789_ net88 net428 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_114_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0712_ net102 net447 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0643_ _0032_ _0162_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q
+ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__a21o_1
XFILLER_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0574_ net24 net8 _0144_ net369 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG15 sky130_fd_sc_hd__mux4_1
XFILLER_97_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1126_ net218 net416 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_25_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1057_ net466 net433 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_51_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput127 Tile_X0Y0_S2MID[2] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__buf_2
Xinput116 Tile_X0Y0_S1END[3] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
Xinput105 Tile_X0Y0_FrameData[31] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_2
Xinput138 Tile_X0Y0_S4END[5] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_4
Xinput149 Tile_X0Y1_E2END[4] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__buf_2
XFILLER_71_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0290_ net222 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q VGND VGND VPWR
+ VPWR _0066_ sky130_fd_sc_hd__o21ba_1
XFILLER_94_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0626_ net173 net187 net171 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG8
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q
+ VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__mux4_1
XFILLER_131_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0557_ net220 net240 _0087_ net137 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG8 sky130_fd_sc_hd__mux4_2
XFILLER_85_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0488_ net33 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit18.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit19.Q VGND VGND VPWR
+ VPWR _0123_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_96_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1109_ net454 net419 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_46_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_55_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_64_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput409 net526 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[6] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1460_ net217 VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__buf_4
X_1391_ Tile_X0Y1_N4END[12] VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__buf_4
X_0411_ net9 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG7 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG3
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit23.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit22.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG8 sky130_fd_sc_hd__mux4_1
XFILLER_67_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0342_ net239 net231 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG7
+ net132 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q
+ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__mux4_2
XFILLER_79_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0273_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q VGND VGND
+ VPWR VPWR _0052_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0609_ net186 net179 net170 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG7
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q
+ VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__mux4_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_145_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0960_ net108 net386 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0891_ net82 net404 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_110_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1512_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG0 VGND VGND VPWR
+ VPWR net645 sky130_fd_sc_hd__buf_4
XFILLER_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1443_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG7 VGND VGND VPWR
+ VPWR net576 sky130_fd_sc_hd__buf_1
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1374_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG3 VGND VGND VPWR
+ VPWR net501 sky130_fd_sc_hd__clkbuf_2
X_0325_ net49 net41 net59 net361 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit4.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit5.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG3 sky130_fd_sc_hd__mux4_1
X_0256_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q VGND
+ VGND VPWR VPWR _0035_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_38_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout422 net423 VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__clkbuf_2
Xfanout400 net401 VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__buf_2
XFILLER_48_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout411 net412 VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__clkbuf_2
Xfanout433 net434 VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__clkbuf_2
Xfanout455 net204 VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__buf_4
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout466 net194 VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__buf_4
Xfanout444 net445 VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__clkbuf_2
XFILLER_73_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1090_ net193 net431 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_52_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0943_ net95 net386 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0874_ net471 net402 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_154_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1426_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG2 VGND VGND VPWR
+ VPWR net555 sky130_fd_sc_hd__clkbuf_1
X_1357_ Tile_X0Y1_FrameStrobe[10] VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__clkbuf_1
XFILLER_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0308_ net160 net152 net170 net369 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit22.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit23.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb0 sky130_fd_sc_hd__mux4_1
XFILLER_95_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1288_ net216 net375 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0239_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q VGND
+ VGND VPWR VPWR _0018_ sky130_fd_sc_hd__inv_2
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput570 net687 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f_Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK VGND VGND VPWR VPWR clknet_1_1__leaf_Tile_X0Y1_UserCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_115_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_142_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0590_ net154 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q VGND VGND VPWR
+ VPWR _0147_ sky130_fd_sc_hd__o21ba_1
XFILLER_111_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1211_ net460 net391 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1142_ net455 net410 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1073_ net450 net424 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0926_ net110 net394 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0857_ net84 net414 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_136_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0788_ net89 net428 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1409_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG1 VGND VGND VPWR
+ VPWR net536 sky130_fd_sc_hd__buf_1
XFILLER_28_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0711_ net468 net446 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0642_ net142 net180 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q
+ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__mux2_1
X_0573_ net220 net240 _0087_ net137 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q VGND VGND VPWR
+ VPWR _0144_ sky130_fd_sc_hd__mux4_2
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1125_ net190 net418 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1056_ net465 net433 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_40_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0909_ net474 net396 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput117 Tile_X0Y0_S2END[0] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
Xinput106 Tile_X0Y0_FrameData[3] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput139 Tile_X0Y0_S4END[6] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_4
Xinput128 Tile_X0Y0_S2MID[3] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__buf_2
XFILLER_56_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_90 net596 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0625_ net186 net179 net170 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG7
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q
+ VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__mux4_2
XFILLER_89_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0556_ net29 net3 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG9
+ net368 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG6
+ sky130_fd_sc_hd__mux4_1
X_0487_ net68 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit18.Q
+ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__nand2b_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1108_ net453 net419 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1039_ net189 net441 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_139_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_2_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1390_ Tile_X0Y1_N4END[11] VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__buf_4
X_0410_ net17 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG8
+ net361 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit20.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit21.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG7
+ sky130_fd_sc_hd__mux4_1
X_0341_ net36 net45 net37 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit16.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit17.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG7
+ sky130_fd_sc_hd__mux4_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0272_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q VGND
+ VGND VPWR VPWR _0051_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_18_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0608_ net185 net178 net169 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG6
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q
+ VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__mux4_2
X_0539_ net1 net31 net369 _0083_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb0 sky130_fd_sc_hd__mux4_1
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0890_ net83 net402 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_110_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1511_ Tile_X0Y0_S4END[15] VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__buf_4
X_1442_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG6 VGND VGND VPWR
+ VPWR net575 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1373_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG2 VGND VGND VPWR
+ VPWR net500 sky130_fd_sc_hd__clkbuf_2
XFILLER_67_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0324_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb3 net128 net235
+ net120 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit15.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit14.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG3
+ sky130_fd_sc_hd__mux4_2
X_0255_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q VGND
+ VGND VPWR VPWR _0034_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_38_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout401 net406 VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__clkbuf_2
Xfanout423 Tile_X0Y1_FrameStrobe[3] VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__buf_2
Xfanout412 net413 VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout456 net203 VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__buf_4
Xfanout434 net435 VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__clkbuf_2
Xfanout445 net448 VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_92_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout467 net105 VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__buf_2
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0942_ net96 net385 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_13_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0873_ net470 net402 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_118_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1425_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG1 VGND VGND VPWR
+ VPWR net554 sky130_fd_sc_hd__buf_1
X_1356_ net372 VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__buf_1
XFILLER_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0307_ net232 net224 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG0
+ net125 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q
+ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__mux4_1
XFILLER_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1287_ net217 net375 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0238_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit29.Q VGND
+ VGND VPWR VPWR _0017_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_124_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput560 net677 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[8] sky130_fd_sc_hd__buf_2
Xoutput571 net688 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_132_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_142_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1210_ net459 net391 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_48_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1141_ net454 net410 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_148_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1072_ net449 net424 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0925_ net111 net394 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0856_ net85 net414 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0787_ net90 net429 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1408_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG0 VGND VGND VPWR
+ VPWR net535 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1339_ net474 VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput390 net507 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[1] sky130_fd_sc_hd__buf_2
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0710_ net467 net446 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0641_ _0031_ _0143_ _0160_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q
+ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__o211a_1
X_0572_ net13 net7 _0143_ net368 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG14 sky130_fd_sc_hd__mux4_1
XFILLER_151_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1124_ net191 net418 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1055_ net464 net432 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_121_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0908_ net473 net396 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0839_ net468 net414 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput118 Tile_X0Y0_S2END[1] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
Xinput107 Tile_X0Y0_FrameData[4] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_4
Xinput129 Tile_X0Y0_S2MID[4] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_80 Tile_X0Y1_FrameData[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 net597 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0624_ net185 net178 net169 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG6
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q
+ VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__mux4_2
X_0555_ net221 net241 _0058_ net138 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG9 sky130_fd_sc_hd__mux4_2
XFILLER_85_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0486_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12 net360 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit18.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit19.Q VGND VGND VPWR
+ VPWR _0121_ sky130_fd_sc_hd__mux4_1
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1107_ net452 net419 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1038_ net198 net440 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_112_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0340_ net46 net38 net56 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit10.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit11.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG6
+ sky130_fd_sc_hd__mux4_1
X_0271_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q VGND
+ VGND VPWR VPWR _0050_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_121_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_130_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0607_ net184 net177 net168 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG5
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q
+ VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__mux4_2
X_0538_ net30 net8 net369 _0083_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG7 sky130_fd_sc_hd__mux4_1
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0469_ net72 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit17.Q
+ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_84_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1510_ Tile_X0Y0_S4END[14] VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__buf_4
XFILLER_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1441_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG5 VGND VGND VPWR
+ VPWR net574 sky130_fd_sc_hd__buf_1
XFILLER_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1372_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG1 VGND VGND VPWR
+ VPWR net499 sky130_fd_sc_hd__clkbuf_1
X_0323_ net157 net149 net167 _0079_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit28.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit29.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb3 sky130_fd_sc_hd__mux4_1
XFILLER_67_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0254_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q VGND
+ VGND VPWR VPWR _0033_ sky130_fd_sc_hd__inv_1
XFILLER_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout402 net404 VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__clkbuf_4
Xfanout413 net414 VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout457 net202 VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__clkbuf_4
Xfanout424 net425 VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__clkbuf_2
Xfanout446 net448 VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__buf_2
Xfanout435 Tile_X0Y1_FrameStrobe[1] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__buf_2
Xfanout468 net104 VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__buf_2
XFILLER_120_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0941_ net474 net387 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_13_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0872_ net469 net402 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_118_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1424_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG0 VGND VGND VPWR
+ VPWR net551 sky130_fd_sc_hd__buf_1
X_1355_ net379 VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__buf_1
X_0306_ net52 net44 net63 net364 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit2.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit3.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG0 sky130_fd_sc_hd__mux4_2
X_1286_ net218 net373 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0237_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit26.Q VGND
+ VGND VPWR VPWR _0016_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_124_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput561 net678 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[9] sky130_fd_sc_hd__buf_2
Xoutput550 net667 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[0] sky130_fd_sc_hd__buf_2
Xoutput572 net689 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_75_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1140_ net453 net410 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1071_ net189 net435 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_92_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_170 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0924_ net112 net395 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0855_ net86 net415 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0786_ net91 net428 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_114_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1407_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG3 VGND VGND VPWR
+ VPWR net534 sky130_fd_sc_hd__clkbuf_2
X_1338_ net475 VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__buf_1
XFILLER_45_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1269_ net454 net374 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_24_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput380 net497 VGND VGND VPWR VPWR Tile_X0Y0_N1BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_126_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput391 net508 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[2] sky130_fd_sc_hd__buf_2
XFILLER_142_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0640_ net172 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q
+ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__or2_1
XFILLER_143_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0571_ net221 net241 _0058_ net138 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q VGND VGND VPWR
+ VPWR _0143_ sky130_fd_sc_hd__mux4_2
XFILLER_111_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1123_ net192 net417 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1054_ net463 net432 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_121_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0907_ net472 net396 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0838_ net467 net414 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0769_ net107 net436 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput108 Tile_X0Y0_FrameData[5] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput119 Tile_X0Y0_S2END[2] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_25_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_70 net526 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_92 net598 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_81 Tile_X0Y1_FrameData[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0623_ net184 net177 net168 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG5
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q
+ VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__mux4_2
X_0554_ net28 net32 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG10
+ net367 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG5
+ sky130_fd_sc_hd__mux4_1
X_0485_ _0013_ _0116_ _0120_ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG3
+ sky130_fd_sc_hd__o21a_1
XFILLER_85_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1106_ net451 net417 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_108_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1037_ net209 net441 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput90 Tile_X0Y0_FrameData[18] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_4
XFILLER_115_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0270_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q VGND
+ VGND VPWR VPWR _0049_ sky130_fd_sc_hd__inv_1
XFILLER_67_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0606_ net183 net176 net167 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG4
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q
+ VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__mux4_1
X_0537_ net29 net7 net368 _0082_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG6 sky130_fd_sc_hd__mux4_1
X_0468_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13 net363 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit17.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit18.Q VGND VGND VPWR
+ VPWR _0106_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_84_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0399_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END1 net245 net114
+ net134 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit10.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit11.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG1
+ sky130_fd_sc_hd__mux4_2
XFILLER_26_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1440_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG4 VGND VGND VPWR
+ VPWR net573 sky130_fd_sc_hd__clkbuf_2
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1371_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG0 VGND VGND VPWR
+ VPWR net498 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_98_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0322_ net235 net227 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG3
+ net128 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q
+ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__mux4_1
X_0253_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q VGND
+ VGND VPWR VPWR _0032_ sky130_fd_sc_hd__inv_2
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout414 Tile_X0Y1_FrameStrobe[4] VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__clkbuf_2
Xfanout403 net404 VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout425 net426 VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__buf_2
Xfanout447 net448 VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout436 net437 VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__clkbuf_4
Xfanout458 net201 VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__clkbuf_4
Xfanout469 net102 VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__clkbuf_4
XFILLER_46_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0940_ net473 net387 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0871_ net468 net402 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1423_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb7 VGND VGND VPWR
+ VPWR net550 sky130_fd_sc_hd__clkbuf_2
X_1354_ net387 VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__clkbuf_1
X_0305_ net36 net62 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15
+ _0071_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit28.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit29.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG3
+ sky130_fd_sc_hd__mux4_1
XFILLER_28_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1285_ net190 net373 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0236_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit23.Q VGND
+ VGND VPWR VPWR _0015_ sky130_fd_sc_hd__inv_1
XFILLER_95_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput551 net668 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[10] sky130_fd_sc_hd__buf_2
Xoutput562 net679 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput540 net657 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput573 net690 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_75_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1070_ net198 net435 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_52_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_160 net524 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_171 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0923_ net82 net394 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0854_ net87 net415 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0785_ net93 net427 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1406_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG2 VGND VGND VPWR
+ VPWR net533 sky130_fd_sc_hd__buf_1
XFILLER_68_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1337_ net476 VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__buf_1
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1268_ net453 net374 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1199_ net189 net400 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_54_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_89_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput370 net487 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
XFILLER_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput392 net509 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput381 net498 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_86_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0570_ net2 net6 _0142_ net367 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG13 sky130_fd_sc_hd__mux4_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1122_ net193 net418 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1053_ net462 net434 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_121_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0906_ net471 net396 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0837_ net81 net421 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0768_ net108 net436 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput109 Tile_X0Y0_FrameData[6] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_4
X_0699_ net127 _0054_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__nand2_1
XFILLER_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_60 net525 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 net526 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 net599 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 Tile_X0Y1_FrameData[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0622_ net183 net176 net167 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG4
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q
+ VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__mux4_1
X_0553_ net222 net242 _0065_ net139 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG10 sky130_fd_sc_hd__mux4_2
X_0484_ _0117_ _0118_ _0119_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit24.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit25.Q VGND VGND VPWR
+ VPWR _0120_ sky130_fd_sc_hd__a221o_1
XFILLER_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1105_ net450 net416 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_53_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1036_ net212 net441 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput91 Tile_X0Y0_FrameData[19] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_4
Xinput80 Tile_X0Y0_EE4END[9] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_1
XFILLER_122_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0605_ net182 net175 net166 _0141_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q VGND VGND VPWR
+ VPWR net281 sky130_fd_sc_hd__mux4_1
X_0536_ net28 net6 net367 _0081_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG5 sky130_fd_sc_hd__mux4_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0467_ _0010_ _0101_ _0105_ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG0
+ sky130_fd_sc_hd__o21a_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0398_ net10 net23 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG2
+ net362 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit0.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit1.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG13
+ sky130_fd_sc_hd__mux4_1
XFILLER_81_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1019_ net460 net440 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_92_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1370_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG3 VGND VGND VPWR
+ VPWR net497 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_98_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0321_ net49 net41 net55 net361 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit8.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit9.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG3 sky130_fd_sc_hd__mux4_2
XFILLER_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0252_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q VGND VGND
+ VPWR VPWR _0031_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_81_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout404 net406 VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__buf_2
Xfanout426 net431 VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__buf_2
Xfanout448 Tile_X0Y1_FrameStrobe[0] VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__clkbuf_2
Xfanout415 Tile_X0Y1_FrameStrobe[4] VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__buf_2
Xfanout437 net439 VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__clkbuf_2
Xfanout459 net200 VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__clkbuf_4
X_0519_ net160 net152 net171 _0076_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG0 sky130_fd_sc_hd__mux4_1
X_1499_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG3 VGND VGND VPWR
+ VPWR net626 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_61_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_70_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_109_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0870_ net467 net403 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1422_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb6 VGND VGND VPWR
+ VPWR net549 sky130_fd_sc_hd__clkbuf_1
XFILLER_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1353_ net397 VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_118_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1284_ net191 net376 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0304_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END3 net247 net116
+ net136 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit6.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit7.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15
+ sky130_fd_sc_hd__mux4_2
XFILLER_95_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0235_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit20.Q VGND
+ VGND VPWR VPWR _0014_ sky130_fd_sc_hd__inv_2
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_127_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0999_ net468 net372 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_135_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_136_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput552 net669 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[11] sky130_fd_sc_hd__buf_2
Xoutput563 net680 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput541 net658 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput530 net647 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput574 net691 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_75_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_161 net524 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_150 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_172 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0922_ net83 net394 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0853_ net88 net412 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0784_ net94 net427 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_154_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1405_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG1 VGND VGND VPWR
+ VPWR net532 sky130_fd_sc_hd__buf_1
X_1336_ net94 VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 DO_SRAM0 VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_79_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1267_ net452 net373 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1198_ net198 net400 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_144_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput360 net477 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
Xoutput371 net488 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[4] sky130_fd_sc_hd__buf_2
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput382 net499 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput393 net510 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[4] sky130_fd_sc_hd__buf_2
XFILLER_120_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_153_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1121_ net466 net416 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1052_ net461 net434 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0905_ net470 net396 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0836_ net92 net421 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0767_ net109 net436 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_132_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0698_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q _0209_
+ _0208_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q VGND
+ VGND VPWR VPWR _0210_ sky130_fd_sc_hd__o211a_1
XFILLER_102_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1319_ net107 VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_50 net523 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 net527 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 net525 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_83 Tile_X0Y1_FrameData[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_94 net601 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0621_ net182 net175 net166 _0141_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q VGND VGND VPWR
+ VPWR net314 sky130_fd_sc_hd__mux4_2
XFILLER_109_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0552_ net27 net31 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG11
+ net366 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG4
+ sky130_fd_sc_hd__mux4_1
XFILLER_97_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0483_ net55 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG3 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit23.Q
+ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__mux2_1
X_1104_ net449 net416 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1035_ net213 net441 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput81 Tile_X0Y0_FrameData[0] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_4
Xinput70 Tile_X0Y0_EE4END[14] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dlymetal6s2s_1
X_0819_ net90 net421 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput92 Tile_X0Y0_FrameData[1] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_4
XFILLER_107_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0604_ net181 net174 net165 _0142_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q VGND VGND VPWR
+ VPWR net270 sky130_fd_sc_hd__mux4_2
X_0535_ net27 net5 net366 net365 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG4 sky130_fd_sc_hd__mux4_1
X_0466_ _0102_ _0103_ _0104_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit15.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit16.Q VGND VGND VPWR
+ VPWR _0105_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0397_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END2 net246 net115
+ net135 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit12.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit13.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG2
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_1_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1018_ net459 net440 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_92_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0320_ net50 net42 net60 net362 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit2.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit3.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG2 sky130_fd_sc_hd__mux4_1
X_0251_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q VGND VGND
+ VPWR VPWR _0030_ sky130_fd_sc_hd__inv_1
XFILLER_90_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1567_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG15 VGND VGND VPWR
+ VPWR net685 sky130_fd_sc_hd__buf_1
Xfanout405 net406 VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__buf_2
Xfanout427 net429 VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__clkbuf_4
X_0518_ net144 net163 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15
+ _0075_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG3
+ sky130_fd_sc_hd__mux4_1
XFILLER_58_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout416 net419 VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__clkbuf_2
Xfanout438 Tile_X0Y1_FrameStrobe[1] VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__clkbuf_2
Xfanout449 net211 VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__buf_4
X_1498_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG2 VGND VGND VPWR
+ VPWR net625 sky130_fd_sc_hd__clkbuf_2
X_0449_ _0092_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit31.Q
+ _0003_ _0091_ VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__a2bb2o_1
XFILLER_66_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1421_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb5 VGND VGND VPWR
+ VPWR net548 sky130_fd_sc_hd__buf_1
X_1352_ net406 VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__buf_4
XFILLER_95_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1283_ net192 net376 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0303_ net144 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15 net170
+ _0075_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit21.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit20.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END3
+ sky130_fd_sc_hd__mux4_2
X_0234_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit25.Q VGND
+ VGND VPWR VPWR _0013_ sky130_fd_sc_hd__inv_2
XFILLER_48_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0998_ net467 net372 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_135_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput520 net637 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput553 net670 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[1] sky130_fd_sc_hd__buf_2
Xoutput542 net659 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput531 net648 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[1] sky130_fd_sc_hd__buf_2
Xoutput564 net681 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput575 net692 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_115_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_140 net643 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_151 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_162 net524 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_173 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0921_ net84 net394 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0852_ net89 net412 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0783_ net476 net430 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_154_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1404_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG0 VGND VGND VPWR
+ VPWR net531 sky130_fd_sc_hd__buf_1
X_1335_ net93 VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__buf_1
Xinput2 DO_SRAM1 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1266_ net451 net373 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1197_ net209 net400 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_101_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput361 net478 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[13] sky130_fd_sc_hd__buf_2
XFILLER_126_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput350 net350 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[3] sky130_fd_sc_hd__buf_2
XFILLER_105_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput372 net489 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[5] sky130_fd_sc_hd__buf_2
Xoutput394 net511 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput383 net500 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_126_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1120_ net465 net416 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_65_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1051_ net460 net433 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_76_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0904_ net469 net396 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0835_ net103 net421 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0766_ net110 net436 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_132_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0697_ net149 net128 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
+ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__mux2_1
XFILLER_56_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1318_ net106 VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__clkbuf_2
X_1249_ net194 net389 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_40 net515 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 net527 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 net523 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 net525 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_84 net581 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_95 net606 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0620_ net181 net174 net165 _0142_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q VGND VGND VPWR
+ VPWR net303 sky130_fd_sc_hd__mux4_2
XFILLER_109_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0551_ net223 net243 _0072_ net140 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG11 sky130_fd_sc_hd__mux4_2
XFILLER_97_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0482_ net36 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit23.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit24.Q VGND VGND VPWR
+ VPWR _0118_ sky130_fd_sc_hd__o21ba_1
XFILLER_87_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1103_ net189 net424 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1034_ net214 net441 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput82 Tile_X0Y0_FrameData[10] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_4
Xinput60 Tile_X0Y0_E6END[5] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_2
Xinput71 Tile_X0Y0_EE4END[15] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_2
X_0818_ net91 net423 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput93 Tile_X0Y0_FrameData[20] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_4
X_0749_ net474 net438 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_107_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0603_ net180 net188 net164 _0143_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q VGND VGND VPWR
+ VPWR net259 sky130_fd_sc_hd__mux4_2
X_0534_ net24 net4 net366 net365 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_58_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0465_ net63 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG0 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit14.Q
+ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__mux2_1
X_0396_ net9 net22 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG3
+ net361 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit30.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit31.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG12
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_1_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1017_ net458 net440 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_92_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0250_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q VGND VGND
+ VPWR VPWR _0029_ sky130_fd_sc_hd__inv_2
XFILLER_82_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1566_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG14 VGND VGND VPWR
+ VPWR net684 sky130_fd_sc_hd__clkbuf_1
Xfanout428 net429 VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__buf_2
Xfanout417 net418 VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__clkbuf_2
X_0517_ net143 net162 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14
+ _0068_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit22.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit23.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG2
+ sky130_fd_sc_hd__mux4_1
Xfanout406 Tile_X0Y1_FrameStrobe[5] VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__clkbuf_2
Xfanout439 Tile_X0Y1_FrameStrobe[1] VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1497_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG1 VGND VGND VPWR
+ VPWR net624 sky130_fd_sc_hd__buf_4
X_0448_ net37 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit30.Q
+ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__nand2_1
XFILLER_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0379_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END3 net247 net116
+ net136 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit30.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit31.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG11
+ sky130_fd_sc_hd__mux4_2
XFILLER_64_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1420_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb4 VGND VGND VPWR
+ VPWR net547 sky130_fd_sc_hd__buf_1
XFILLER_141_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1351_ net414 VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__clkbuf_2
X_0302_ _0022_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q
+ _0072_ _0074_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__a31o_1
X_1282_ net193 net376 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0233_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit22.Q VGND
+ VGND VPWR VPWR _0012_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_34_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0997_ net81 net377 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_135_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput510 net627 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput554 net671 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[2] sky130_fd_sc_hd__buf_2
Xoutput543 net660 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput521 net638 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput532 net649 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_120_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput565 net682 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput576 net693 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[8] sky130_fd_sc_hd__buf_2
X_1549_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG9 VGND VGND VPWR
+ VPWR net678 sky130_fd_sc_hd__buf_1
XFILLER_115_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_141 net646 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_130 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_152 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_163 net524 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_174 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0920_ net85 net394 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_81_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0851_ net90 net411 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0782_ net475 net430 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1403_ clknet_1_1__leaf_Tile_X0Y1_UserCLK VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__buf_2
X_1334_ net91 VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__clkbuf_2
XFILLER_28_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1265_ net450 net373 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput3 DO_SRAM10 VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_79_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1196_ net212 net400 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput362 net479 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[14] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput351 net351 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[4] sky130_fd_sc_hd__buf_2
Xoutput340 net340 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[23] sky130_fd_sc_hd__buf_2
XFILLER_105_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput384 net501 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput373 net490 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[6] sky130_fd_sc_hd__buf_2
Xoutput395 net512 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[6] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_58_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1050_ net459 net433 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_85_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0903_ net468 net396 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0834_ net106 net421 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_94_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0765_ net111 net438 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_142_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0696_ _0054_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG0 VGND VGND VPWR VPWR
+ _0208_ sky130_fd_sc_hd__or3_1
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1317_ net103 VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__clkbuf_2
X_1248_ net195 net389 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1179_ net460 net399 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_41 net517 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_30 net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_74 net527 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 net525 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 net523 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_96 Tile_X0Y1_FrameStrobe[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_85 net583 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0550_ net24 net8 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12
+ net365 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG3
+ sky130_fd_sc_hd__mux4_1
XFILLER_124_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0481_ net74 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit23.Q
+ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__nand2b_1
XFILLER_97_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1102_ net198 net424 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1033_ net215 net440 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_53_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0817_ net93 net422 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput61 Tile_X0Y0_E6END[6] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_2
Xinput72 Tile_X0Y0_EE4END[1] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_1
Xinput50 Tile_X0Y0_E2MID[5] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_1
Xinput94 Tile_X0Y0_FrameData[21] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_4
Xinput83 Tile_X0Y0_FrameData[11] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_4
X_0748_ net473 net438 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0679_ _0050_ _0192_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q
+ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__a21o_1
XFILLER_123_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0602_ net173 net187 net161 _0144_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q VGND VGND VPWR
+ VPWR net258 sky130_fd_sc_hd__mux4_1
X_0533_ net13 net3 net367 _0081_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_85_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0464_ net33 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit14.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit15.Q VGND VGND VPWR
+ VPWR _0103_ sky130_fd_sc_hd__o21ba_1
XFILLER_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0395_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END3 net247 net116
+ net136 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit14.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit15.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG3
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_1_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1016_ net457 net440 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_92_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_22_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput240 Tile_X0Y1_N4END[0] VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1565_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG13 VGND VGND VPWR
+ VPWR net683 sky130_fd_sc_hd__buf_1
XFILLER_98_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout407 net408 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__clkbuf_2
Xfanout418 net419 VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__clkbuf_2
X_0516_ net142 net172 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13
+ _0061_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit20.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit21.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG1
+ sky130_fd_sc_hd__mux4_1
Xfanout429 net431 VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__dlymetal6s2s_1
X_1496_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG0 VGND VGND VPWR
+ VPWR net623 sky130_fd_sc_hd__clkbuf_2
X_0447_ net45 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit31.Q
+ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__mux2_1
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0378_ net12 net26 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12
+ net360 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit12.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit13.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG3
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_37_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1350_ net421 VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__clkbuf_2
XFILLER_79_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0301_ net166 _0022_ _0073_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__o21a_1
X_1281_ net466 net376 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0232_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit19.Q VGND
+ VGND VPWR VPWR _0011_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_34_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0996_ net92 net377 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_135_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput511 net628 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput500 net617 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput544 net661 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput522 net639 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput533 net650 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[3] sky130_fd_sc_hd__buf_2
Xoutput555 net672 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[3] sky130_fd_sc_hd__buf_2
Xoutput566 net683 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput577 net694 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[9] sky130_fd_sc_hd__buf_2
X_1548_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG8 VGND VGND VPWR
+ VPWR net677 sky130_fd_sc_hd__clkbuf_2
X_1479_ net453 VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_105_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_114_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_123_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_142 net646 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_131 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_120 Tile_X0Y1_FrameStrobe[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_164 net524 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_153 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0850_ net91 net411 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_139_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0781_ net474 net427 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_154_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1402_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG3 VGND VGND VPWR
+ VPWR net520 sky130_fd_sc_hd__buf_1
XFILLER_114_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1333_ net90 VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1264_ net449 net373 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 DO_SRAM11 VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_79_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1195_ net213 net401 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_36_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0979_ net90 net378 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_145_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput352 net352 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[5] sky130_fd_sc_hd__buf_2
Xoutput330 net330 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[14] sky130_fd_sc_hd__buf_2
Xoutput341 net341 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[24] sky130_fd_sc_hd__buf_2
XFILLER_105_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput374 net491 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[7] sky130_fd_sc_hd__buf_2
Xoutput396 net513 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput385 net502 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput363 net480 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[15] sky130_fd_sc_hd__buf_2
XFILLER_113_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0902_ net467 net397 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0833_ net107 net422 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_132_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0764_ net112 net438 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_142_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0695_ _0203_ _0205_ _0207_ _0201_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q
+ VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__a32o_1
XFILLER_142_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1316_ net92 VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_67_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1247_ net464 net383 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1178_ net459 net399 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_31 net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_20 net350 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 net521 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_75 net527 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 net523 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 net525 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_97 Tile_X0Y1_FrameStrobe[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_86 net588 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0480_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG7 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit23.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit24.Q
+ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__mux4_1
XFILLER_124_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1101_ net209 net425 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1032_ net216 net440 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput40 Tile_X0Y0_E2END[3] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlymetal6s2s_1
X_0816_ net94 net422 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput62 Tile_X0Y0_E6END[7] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_2
Xinput73 Tile_X0Y0_EE4END[2] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_1
Xinput51 Tile_X0Y0_E2MID[6] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_1
Xinput95 Tile_X0Y0_FrameData[22] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_1
Xinput84 Tile_X0Y0_FrameData[12] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_4
X_0747_ net472 net436 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0678_ net144 net179 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q
+ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__mux2_1
XFILLER_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0601_ _0027_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q
+ net365 _0154_ VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__a31o_1
X_0532_ net2 net32 net368 _0082_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_98_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0463_ net65 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit14.Q
+ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__nand2b_1
X_0394_ net17 net21 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG4
+ net360 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit28.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit29.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG11
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_1_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1015_ net203 net441 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_92_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput241 Tile_X0Y1_N4END[1] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_2
Xinput230 Tile_X0Y1_N2END[6] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_2
XFILLER_75_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1564_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG12 VGND VGND VPWR
+ VPWR net682 sky130_fd_sc_hd__buf_1
Xfanout408 net409 VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__buf_2
X_1495_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG7 VGND VGND VPWR
+ VPWR net622 sky130_fd_sc_hd__buf_1
X_0515_ net141 net171 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12
+ _0090_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit18.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit19.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG0
+ sky130_fd_sc_hd__mux4_1
Xfanout419 Tile_X0Y1_FrameStrobe[3] VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_97_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0446_ net36 net78 net71 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit28.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit29.Q
+ VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__mux4_2
X_0377_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END0 net244 net113
+ net133 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit0.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit1.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12
+ sky130_fd_sc_hd__mux4_2
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0300_ net223 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q VGND VGND VPWR
+ VPWR _0073_ sky130_fd_sc_hd__o21ba_1
X_1280_ net465 net375 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_95_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0231_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit16.Q VGND
+ VGND VPWR VPWR _0010_ sky130_fd_sc_hd__inv_2
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0995_ net103 net377 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_135_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput501 net618 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_117_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput545 net662 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput512 net629 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput523 net640 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput534 net651 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput556 net673 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[4] sky130_fd_sc_hd__buf_2
Xoutput567 net684 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[14] sky130_fd_sc_hd__buf_2
XFILLER_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1547_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG7 VGND VGND VPWR
+ VPWR net676 sky130_fd_sc_hd__clkbuf_1
XFILLER_115_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1478_ net454 VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__buf_4
X_0429_ net35 net77 net70 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit26.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit27.Q
+ VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__mux4_2
XFILLER_10_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_110 Tile_X0Y1_FrameStrobe[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_143 net646 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_121 Tile_X0Y1_FrameStrobe[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 net611 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_154 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_176 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0780_ net473 net427 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1401_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG2 VGND VGND VPWR
+ VPWR net519 sky130_fd_sc_hd__buf_1
XFILLER_122_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1332_ net89 VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__clkbuf_2
X_1263_ net189 net381 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput5 DO_SRAM12 VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_79_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1194_ net214 net401 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_36_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0978_ net91 net378 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_126_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput320 net320 VGND VGND VPWR VPWR DI_SRAM7 sky130_fd_sc_hd__buf_2
Xoutput353 net353 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[6] sky130_fd_sc_hd__buf_2
Xoutput331 net331 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[15] sky130_fd_sc_hd__buf_2
Xoutput342 net342 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[25] sky130_fd_sc_hd__buf_2
Xoutput364 net481 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[16] sky130_fd_sc_hd__buf_2
Xoutput375 net492 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[8] sky130_fd_sc_hd__buf_2
Xoutput386 net503 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[5] sky130_fd_sc_hd__buf_2
Xoutput397 net514 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0901_ net81 net405 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0832_ net108 net422 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_132_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0763_ net82 net437 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_142_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0694_ _0052_ _0206_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q
+ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__o21ba_1
XFILLER_142_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1315_ net81 VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__buf_1
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1246_ net463 net383 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_142_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1177_ net458 net398 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_24_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_32 net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 net300 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 net356 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_65 net526 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 net521 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 net523 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 net528 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 Tile_X0Y1_FrameStrobe[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_87 net592 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1100_ net212 net425 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_64_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1031_ net217 net442 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput30 DO_SRAM7 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_2
Xinput63 Tile_X0Y0_E6END[8] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_2
Xinput41 Tile_X0Y0_E2END[4] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_12_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0815_ net476 net420 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput52 Tile_X0Y0_E2MID[7] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_2
Xinput96 Tile_X0Y0_FrameData[23] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput85 Tile_X0Y0_FrameData[13] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_4
Xinput74 Tile_X0Y0_EE4END[3] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
X_0746_ net471 net436 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0677_ _0049_ _0141_ _0190_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q
+ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_4_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_150_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1229_ net209 net392 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_107_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0600_ net149 _0027_ _0153_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__o21a_1
X_0531_ net1 net31 net369 _0083_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0462_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12 net364 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit14.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit15.Q VGND VGND VPWR
+ VPWR _0101_ sky130_fd_sc_hd__mux4_1
XFILLER_112_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0393_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END0 net244 net113
+ net133 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit16.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit17.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG4
+ sky130_fd_sc_hd__mux4_2
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1014_ net204 net441 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_92_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0729_ net84 net444 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_103_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput220 Tile_X0Y1_N1END[0] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__buf_2
Xinput242 Tile_X0Y1_N4END[2] VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_2
Xinput231 Tile_X0Y1_N2END[7] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_126_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1563_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG11 VGND VGND VPWR
+ VPWR net681 sky130_fd_sc_hd__buf_1
Xfanout409 net410 VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__clkbuf_2
X_1494_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG6 VGND VGND VPWR
+ VPWR net621 sky130_fd_sc_hd__clkbuf_2
X_0514_ net33 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12 net59
+ _0086_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit23.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit22.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG0
+ sky130_fd_sc_hd__mux4_1
X_0445_ net35 net77 net70 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit26.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit27.Q
+ VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_97_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0376_ net11 net25 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit10.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit11.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0230_ net127 VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__inv_1
XFILLER_36_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0994_ net106 net377 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput502 net619 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput535 net652 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput513 net630 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput524 net641 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput557 net674 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[5] sky130_fd_sc_hd__buf_2
Xoutput568 net685 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput546 net663 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[4] sky130_fd_sc_hd__buf_2
X_1546_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG6 VGND VGND VPWR
+ VPWR net675 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1477_ net455 VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__buf_4
X_0428_ net34 net76 net69 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit24.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit25.Q
+ VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__mux4_2
XFILLER_39_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0359_ net10 net19 net363 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit8.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit9.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG1
+ sky130_fd_sc_hd__mux4_1
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_19_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_37_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_100 Tile_X0Y1_FrameStrobe[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_111 Tile_X0Y1_FrameStrobe[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_133 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_122 Tile_X0Y1_FrameStrobe[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 net631 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_144 net646 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_155 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_177 net511 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1400_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG1 VGND VGND VPWR
+ VPWR net518 sky130_fd_sc_hd__buf_1
XFILLER_122_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1331_ net88 VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_2
X_1262_ net198 net381 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput6 DO_SRAM13 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_79_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1193_ net215 net399 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_91_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0977_ net93 net378 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput310 net310 VGND VGND VPWR VPWR DI_SRAM26 sky130_fd_sc_hd__buf_2
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput321 net321 VGND VGND VPWR VPWR DI_SRAM8 sky130_fd_sc_hd__buf_2
Xoutput332 net332 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[16] sky130_fd_sc_hd__buf_2
Xoutput343 net343 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[26] sky130_fd_sc_hd__buf_2
Xoutput365 net482 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[17] sky130_fd_sc_hd__buf_2
Xoutput376 net493 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[9] sky130_fd_sc_hd__buf_2
Xoutput387 net504 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[6] sky130_fd_sc_hd__buf_2
Xoutput354 net354 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[7] sky130_fd_sc_hd__buf_2
XFILLER_113_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput398 net515 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[10] sky130_fd_sc_hd__buf_2
X_1529_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG5 VGND VGND VPWR
+ VPWR net656 sky130_fd_sc_hd__buf_1
XFILLER_142_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ net92 net405 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0831_ net109 net420 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0762_ net83 net437 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_132_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0693_ net227 net146 net153 net147 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q VGND VGND VPWR
+ VPWR _0206_ sky130_fd_sc_hd__mux4_1
XFILLER_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1314_ clknet_1_0__leaf_Tile_X0Y1_UserCLK VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_67_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1245_ net462 net384 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1176_ net457 net398 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_112_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_22 net489 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_11 net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_66 net526 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 net521 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 net523 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_99 Tile_X0Y1_FrameStrobe[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 net535 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 net593 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1030_ net218 net442 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_46_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput31 DO_SRAM8 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput20 DO_SRAM26 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_2
X_0814_ net475 net420 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput64 Tile_X0Y0_E6END[9] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput53 Tile_X0Y0_E6END[0] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_2
Xinput42 Tile_X0Y0_E2END[5] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_12_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput97 Tile_X0Y0_FrameData[24] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
Xinput86 Tile_X0Y0_FrameData[14] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_4
Xinput75 Tile_X0Y0_EE4END[4] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_2
X_0745_ net470 net437 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0676_ net170 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q
+ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__or2_1
XFILLER_88_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1228_ net212 net392 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1159_ net217 net407 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_52_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0530_ net223 net2 _0072_ net27 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG3 sky130_fd_sc_hd__mux4_1
X_0461_ net41 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit6.Q
+ _0007_ _0100_ VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__a31o_2
XFILLER_66_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0392_ net16 net20 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG5
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit26.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit27.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG10 sky130_fd_sc_hd__mux4_1
XFILLER_93_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1013_ net205 net442 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_81_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0728_ net85 net444 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0659_ _0040_ _0144_ _0175_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q
+ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__o211a_1
XFILLER_103_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput210 Tile_X0Y1_FrameData[30] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__buf_1
XFILLER_68_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput243 Tile_X0Y1_N4END[3] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_2
Xinput232 Tile_X0Y1_N2MID[0] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__buf_2
Xinput221 Tile_X0Y1_N1END[1] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_2
XFILLER_84_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1562_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG10 VGND VGND VPWR
+ VPWR net680 sky130_fd_sc_hd__clkbuf_1
XFILLER_140_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0513_ net223 net243 _0072_ net140 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15 sky130_fd_sc_hd__mux4_2
X_1493_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG5 VGND VGND VPWR
+ VPWR net620 sky130_fd_sc_hd__clkbuf_2
X_0444_ net34 net76 net69 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit24.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit25.Q
+ VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_97_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0375_ net10 net23 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit8.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit9.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_66_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0993_ net107 net377 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_42_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput536 net653 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput503 net620 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[5] sky130_fd_sc_hd__buf_2
Xoutput514 net631 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput525 net642 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput558 net675 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[6] sky130_fd_sc_hd__buf_2
Xoutput569 net686 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[1] sky130_fd_sc_hd__buf_2
X_1545_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG5 VGND VGND VPWR
+ VPWR net674 sky130_fd_sc_hd__buf_1
Xoutput547 net664 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[5] sky130_fd_sc_hd__buf_2
X_1476_ net456 VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_146_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0427_ net33 net75 net68 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit22.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit23.Q
+ VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__mux4_1
XFILLER_27_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0358_ net9 net18 net364 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit6.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit7.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG0
+ sky130_fd_sc_hd__mux4_1
X_0289_ net35 net54 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14
+ _0064_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit30.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit31.Q
+ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__mux4_2
XFILLER_10_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_112 Tile_X0Y1_FrameStrobe[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_101 Tile_X0Y1_FrameStrobe[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_134 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_123 net615 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_167 net631 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_145 net646 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_156 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1330_ net87 VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__buf_1
XFILLER_122_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1261_ net209 net381 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1192_ net216 net399 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput7 DO_SRAM14 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
X_0976_ net94 net378 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput300 net300 VGND VGND VPWR VPWR DI_SRAM17 sky130_fd_sc_hd__buf_2
Xoutput322 net322 VGND VGND VPWR VPWR DI_SRAM9 sky130_fd_sc_hd__buf_2
Xoutput311 net311 VGND VGND VPWR VPWR DI_SRAM27 sky130_fd_sc_hd__buf_2
Xoutput333 net333 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[17] sky130_fd_sc_hd__buf_2
Xoutput344 net344 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[27] sky130_fd_sc_hd__buf_2
Xoutput366 net483 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[18] sky130_fd_sc_hd__buf_2
Xoutput377 net494 VGND VGND VPWR VPWR Tile_X0Y0_N1BEG[0] sky130_fd_sc_hd__buf_2
Xoutput355 net355 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[8] sky130_fd_sc_hd__buf_2
Xoutput399 net516 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput388 net505 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[7] sky130_fd_sc_hd__buf_2
X_1528_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG4 VGND VGND VPWR
+ VPWR net655 sky130_fd_sc_hd__buf_1
XFILLER_113_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1459_ net216 VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__buf_4
XFILLER_59_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0830_ net110 net420 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0761_ net84 net439 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0692_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ _0204_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__or3_1
X_1313_ net466 net370 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1244_ net461 net384 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1175_ net456 net398 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_75_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_23 net498 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_12 net310 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_45 net521 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 net523 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 net526 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 net539 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_89 net593 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0959_ net109 net386 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_118_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout390 net392 VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0813_ net474 net422 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput10 DO_SRAM17 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_4
Xinput21 DO_SRAM27 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
Xinput54 Tile_X0Y0_E6END[10] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
Xinput43 Tile_X0Y0_E2END[6] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_12_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput32 DO_SRAM9 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_2
Xinput98 Tile_X0Y0_FrameData[25] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_2
Xinput87 Tile_X0Y0_FrameData[15] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_4
Xinput76 Tile_X0Y0_EE4END[5] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_1
Xinput65 Tile_X0Y0_EE4END[0] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_2
X_0744_ net469 net437 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0675_ _0186_ _0188_ _0189_ _0048_ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG2
+ sky130_fd_sc_hd__o22a_1
XFILLER_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1227_ net213 net391 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1158_ net218 net407 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_107_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1089_ net466 net424 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_138_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0460_ _0007_ net360 _0099_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__o21a_1
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0391_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END1 net245 net114
+ net134 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit18.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit19.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG5
+ sky130_fd_sc_hd__mux4_2
XFILLER_78_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1012_ net206 net442 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0727_ net86 net444 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_103_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0658_ net167 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q
+ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__or2_1
XFILLER_103_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_139_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0589_ _0023_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q
+ net369 _0146_ VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__a31o_1
XFILLER_69_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput200 Tile_X0Y1_FrameData[21] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__buf_1
Xinput211 Tile_X0Y1_FrameData[31] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__buf_1
Xinput244 Tile_X0Y1_N4END[4] VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_4
Xinput233 Tile_X0Y1_N2MID[1] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_2
Xinput222 Tile_X0Y1_N1END[2] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__buf_2
XFILLER_63_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1561_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG9 VGND VGND VPWR
+ VPWR net694 sky130_fd_sc_hd__buf_1
XFILLER_140_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0512_ net222 net242 _0065_ net139 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14 sky130_fd_sc_hd__mux4_2
X_1492_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG4 VGND VGND VPWR
+ VPWR net619 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_97_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0443_ net33 net75 net68 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit22.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit23.Q
+ VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__mux4_1
X_0374_ net9 net22 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit6.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit7.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_81_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_147_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_156_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0992_ net108 net377 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_42_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput504 net621 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[6] sky130_fd_sc_hd__buf_2
Xoutput526 net643 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput515 net632 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput559 net676 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[7] sky130_fd_sc_hd__buf_2
X_1544_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG4 VGND VGND VPWR
+ VPWR net673 sky130_fd_sc_hd__clkbuf_2
Xoutput548 net665 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput537 net654 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_140_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1475_ net457 VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_146_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0426_ net74 net67 net55 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit20.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit21.Q
+ VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__mux4_2
XFILLER_27_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0357_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END3 net10 net116 net14
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit5.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit4.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG3
+ sky130_fd_sc_hd__mux4_1
X_0288_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit28.Q _0063_
+ _0001_ _0062_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_102 Tile_X0Y1_FrameStrobe[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_113 Tile_X0Y1_FrameStrobe[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_124 net628 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_135 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_146 net646 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_157 net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_168 net644 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1260_ net212 net382 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1191_ net217 net398 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput8 DO_SRAM15 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0975_ net476 net378 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput301 net301 VGND VGND VPWR VPWR DI_SRAM18 sky130_fd_sc_hd__buf_2
XFILLER_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput312 net312 VGND VGND VPWR VPWR DI_SRAM28 sky130_fd_sc_hd__buf_2
Xoutput323 net323 VGND VGND VPWR VPWR EN_SRAM sky130_fd_sc_hd__buf_2
Xoutput334 net334 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[18] sky130_fd_sc_hd__buf_2
XFILLER_99_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput367 net484 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[19] sky130_fd_sc_hd__buf_2
Xoutput378 net495 VGND VGND VPWR VPWR Tile_X0Y0_N1BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput356 net356 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[9] sky130_fd_sc_hd__buf_2
Xoutput345 net345 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[28] sky130_fd_sc_hd__buf_2
Xoutput389 net506 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[0] sky130_fd_sc_hd__buf_2
X_1527_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG3 VGND VGND VPWR
+ VPWR net654 sky130_fd_sc_hd__buf_1
XFILLER_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1458_ net215 VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__buf_4
XFILLER_74_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0409_ net16 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG9
+ net362 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit18.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit19.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG6
+ sky130_fd_sc_hd__mux4_1
XFILLER_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1389_ Tile_X0Y1_N4END[10] VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_78_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0760_ net85 net439 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0691_ net238 net226 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
+ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__mux2_1
XFILLER_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1312_ net465 net370 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_102_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1243_ net460 net383 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1174_ net455 net398 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_64_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_111_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_13 net323 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 net505 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 net521 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 net523 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_68 net526 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 net547 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0958_ net110 net386 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_137_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0889_ net84 net405 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_118_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_120_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout391 net392 VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout380 Tile_X0Y1_FrameStrobe[8] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__buf_2
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0812_ net473 net422 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput11 DO_SRAM18 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
Xinput22 DO_SRAM28 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
Xinput55 Tile_X0Y0_E6END[11] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
Xinput44 Tile_X0Y0_E2END[7] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_12_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput33 Tile_X0Y0_E1END[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_4
Xinput88 Tile_X0Y0_FrameData[16] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_4
Xinput66 Tile_X0Y0_EE4END[10] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_1
Xinput77 Tile_X0Y0_EE4END[6] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlymetal6s2s_1
X_0743_ net468 net438 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput99 Tile_X0Y0_FrameData[26] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_2
X_0674_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG6
+ _0082_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG10 _0047_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q
+ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__mux4_1
XFILLER_115_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1226_ net214 net391 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1157_ net190 net409 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_107_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1088_ net465 net424 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0390_ net15 net19 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit24.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit25.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG9 sky130_fd_sc_hd__mux4_1
XFILLER_78_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1011_ net207 net442 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0726_ net87 net444 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0657_ _0171_ _0173_ _0174_ _0039_ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_11.A
+ sky130_fd_sc_hd__o22a_1
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0588_ net145 _0023_ _0145_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__o21a_1
XFILLER_69_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1209_ net458 net391 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_72_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput201 Tile_X0Y1_FrameData[22] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput245 Tile_X0Y1_N4END[5] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__buf_2
Xinput234 Tile_X0Y1_N2MID[2] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_2
Xinput223 Tile_X0Y1_N1END[3] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__buf_2
Xinput212 Tile_X0Y1_FrameData[3] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_4
XFILLER_84_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1560_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG8 VGND VGND VPWR
+ VPWR net693 sky130_fd_sc_hd__buf_1
X_0511_ net221 net241 _0058_ net138 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13 sky130_fd_sc_hd__mux4_2
XFILLER_140_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1491_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG3 VGND VGND VPWR
+ VPWR net618 sky130_fd_sc_hd__clkbuf_2
X_0442_ net74 net67 net55 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit20.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit21.Q
+ VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__mux4_2
XFILLER_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0373_ net17 net26 net364 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit4.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit5.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb7
+ sky130_fd_sc_hd__mux4_1
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_144_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0709_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q _0219_
+ _0220_ _0210_ VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__o22a_1
XFILLER_97_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0991_ net109 net380 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_42_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput505 net622 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput527 net644 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput516 net633 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput549 net666 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput538 net655 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[4] sky130_fd_sc_hd__buf_2
X_1543_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG3 VGND VGND VPWR
+ VPWR net672 sky130_fd_sc_hd__buf_1
X_1474_ net458 VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__buf_4
XFILLER_140_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0425_ net73 net66 net54 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit18.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit19.Q
+ VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__mux4_2
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0356_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END2 net9 net115 net15
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit3.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit2.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG2
+ sky130_fd_sc_hd__mux4_1
XFILLER_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0287_ net115 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit29.Q
+ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__nand2_1
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_114 Tile_X0Y1_FrameStrobe[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_103 Tile_X0Y1_FrameStrobe[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_125 net635 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_136 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_147 net646 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_158 net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_169 net692 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1190_ net218 net398 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 DO_SRAM16 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_24_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0974_ net475 net380 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput302 net302 VGND VGND VPWR VPWR DI_SRAM19 sky130_fd_sc_hd__buf_2
Xoutput313 net313 VGND VGND VPWR VPWR DI_SRAM29 sky130_fd_sc_hd__buf_2
Xoutput324 net324 VGND VGND VPWR VPWR R_WB_SRAM sky130_fd_sc_hd__buf_2
Xoutput335 net335 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[19] sky130_fd_sc_hd__buf_2
Xoutput368 net485 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput357 net357 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[0] sky130_fd_sc_hd__buf_2
X_1526_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG2 VGND VGND VPWR
+ VPWR net653 sky130_fd_sc_hd__buf_1
Xoutput346 net346 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[29] sky130_fd_sc_hd__buf_2
Xoutput379 net496 VGND VGND VPWR VPWR Tile_X0Y0_N1BEG[2] sky130_fd_sc_hd__buf_2
X_1457_ net214 VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__buf_4
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1388_ Tile_X0Y1_N4END[9] VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__buf_4
X_0408_ net15 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG10 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG6
+ net363 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit17.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit16.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG5
+ sky130_fd_sc_hd__mux4_1
X_0339_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb6 net131 net238
+ net123 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit21.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit20.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6
+ sky130_fd_sc_hd__mux4_2
XFILLER_27_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0690_ _0202_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q VGND VGND VPWR
+ VPWR _0203_ sky130_fd_sc_hd__or3b_1
X_1311_ net464 net371 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1242_ net459 net383 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1173_ net454 net400 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_75_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_14 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG1 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 net506 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 net521 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_69 net526 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 net523 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0957_ net111 net385 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_133_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0888_ net85 net405 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_133_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1509_ Tile_X0Y0_S4END[13] VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__buf_4
XFILLER_141_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout392 net393 VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__buf_2
Xfanout381 net384 VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__buf_2
Xfanout370 net219 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__buf_2
XFILLER_93_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0811_ net472 net422 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput12 DO_SRAM19 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput23 DO_SRAM29 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_2
Xinput34 Tile_X0Y0_E1END[1] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_2
Xinput45 Tile_X0Y0_E2MID[0] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
X_0742_ net467 net438 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput89 Tile_X0Y0_FrameData[17] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_4
Xinput56 Tile_X0Y0_E6END[1] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_2
Xinput67 Tile_X0Y0_EE4END[11] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
Xinput78 Tile_X0Y0_EE4END[7] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_2
X_0673_ _0047_ _0187_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q
+ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__a21o_1
XFILLER_115_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1225_ net215 net391 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1156_ net191 net409 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1087_ net464 net425 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1010_ net208 net442 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_17_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0725_ net88 net444 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0656_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG7
+ net366 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG11 _0038_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q
+ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__mux4_1
X_0587_ net153 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q VGND VGND VPWR
+ VPWR _0145_ sky130_fd_sc_hd__o21ba_1
XFILLER_57_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1208_ net457 net391 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_0_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1139_ net452 net410 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_91_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput202 Tile_X0Y1_FrameData[23] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput224 Tile_X0Y1_N2END[0] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_2
Xinput235 Tile_X0Y1_N2MID[3] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_2
Xinput213 Tile_X0Y1_FrameData[4] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_4
XFILLER_124_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput246 Tile_X0Y1_N4END[6] VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__buf_2
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0510_ net220 net240 _0087_ net137 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12 sky130_fd_sc_hd__mux4_2
X_1490_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG2 VGND VGND VPWR
+ VPWR net617 sky130_fd_sc_hd__clkbuf_2
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0441_ net73 net66 net54 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit18.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit19.Q
+ VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_97_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0372_ net16 net25 net363 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit2.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit3.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb6
+ sky130_fd_sc_hd__mux4_1
XFILLER_39_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0708_ _0212_ _0213_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q
+ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__o21ai_1
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0639_ _0156_ _0158_ _0159_ _0030_ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_8.A
+ sky130_fd_sc_hd__o22a_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_79_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0990_ net110 net380 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_42_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput506 net623 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput517 net634 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[12] sky130_fd_sc_hd__buf_2
XFILLER_5_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput539 net656 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[5] sky130_fd_sc_hd__buf_2
Xoutput528 net645 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[8] sky130_fd_sc_hd__buf_2
X_1542_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG2 VGND VGND VPWR
+ VPWR net671 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_97_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1473_ net459 VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__buf_4
XFILLER_140_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0424_ net72 net80 net64 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit16.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit17.Q
+ VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__mux4_2
XFILLER_79_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0355_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END1 net12 net114 net16
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit1.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit0.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG1
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0286_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END2 net57 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit28.Q
+ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__mux2_1
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_104 Tile_X0Y1_FrameStrobe[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_115 Tile_X0Y1_FrameStrobe[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_137 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_126 net639 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_148 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_159 net225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0973_ net474 net380 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput303 net303 VGND VGND VPWR VPWR DI_SRAM2 sky130_fd_sc_hd__buf_2
Xoutput314 net314 VGND VGND VPWR VPWR DI_SRAM3 sky130_fd_sc_hd__buf_2
Xoutput325 net325 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[0] sky130_fd_sc_hd__buf_2
Xoutput369 net486 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
Xoutput358 net358 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[10] sky130_fd_sc_hd__buf_2
X_1525_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG1 VGND VGND VPWR
+ VPWR net652 sky130_fd_sc_hd__buf_1
Xoutput336 net336 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[1] sky130_fd_sc_hd__buf_2
Xoutput347 net347 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[2] sky130_fd_sc_hd__buf_2
X_1456_ net213 VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__buf_4
X_1387_ Tile_X0Y1_N4END[8] VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__buf_4
X_0407_ net14 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG11 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG7
+ net364 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit15.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit14.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG4
+ sky130_fd_sc_hd__mux4_1
X_0338_ net154 net146 net164 _0082_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb6 sky130_fd_sc_hd__mux4_1
XFILLER_27_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0269_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q VGND
+ VGND VPWR VPWR _0048_ sky130_fd_sc_hd__inv_1
XFILLER_35_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1310_ net463 net371 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1241_ net458 net383 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1172_ net453 net400 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_64_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_26 net509 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 net515 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 net522 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_15 net326 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_59 net525 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0956_ net112 net385 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0887_ net86 net403 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_133_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1508_ Tile_X0Y0_S4END[12] VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__buf_4
XFILLER_101_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1439_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG3 VGND VGND VPWR
+ VPWR net572 sky130_fd_sc_hd__clkbuf_2
XFILLER_55_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout382 net384 VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkbuf_2
Xfanout371 net219 VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkbuf_2
Xfanout393 Tile_X0Y1_FrameStrobe[6] VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout360 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG4 VGND VGND
+ VPWR VPWR net360 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0810_ net471 net422 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput13 DO_SRAM2 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
Xinput24 DO_SRAM3 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_2
X_0741_ net81 net445 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput35 Tile_X0Y0_E1END[2] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
Xinput46 Tile_X0Y0_E2MID[1] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput57 Tile_X0Y0_E6END[2] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_2
Xinput68 Tile_X0Y0_EE4END[12] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_2
Xinput79 Tile_X0Y0_EE4END[8] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_12_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0672_ net143 net178 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q
+ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__mux2_1
XFILLER_115_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1224_ net216 net391 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1155_ net192 net407 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1086_ net463 net425 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_148_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0939_ net472 net387 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_106_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_60_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0724_ net89 net444 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0655_ _0038_ _0172_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q
+ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__a21o_1
XFILLER_69_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0586_ net24 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG4 _0144_
+ _0083_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG11
+ sky130_fd_sc_hd__mux4_1
XFILLER_57_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1207_ net456 net390 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_72_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1138_ net451 net410 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_92_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1069_ net209 net435 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_91_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_117_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput225 Tile_X0Y1_N2END[1] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_2
Xinput236 Tile_X0Y1_N2MID[4] VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_2
Xinput214 Tile_X0Y1_FrameData[5] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_4
Xinput203 Tile_X0Y1_FrameData[24] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_126_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput247 Tile_X0Y1_N4END[7] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_4
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_135_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0440_ net72 net80 net64 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit16.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit17.Q
+ VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__mux4_2
X_0371_ net15 net23 net362 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit0.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit1.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb5
+ sky130_fd_sc_hd__mux4_1
XFILLER_66_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0707_ _0215_ _0217_ _0218_ _0054_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__o22a_1
X_0638_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG4
+ net369 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG8 _0029_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q
+ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__mux4_1
X_0569_ net222 net242 _0065_ net139 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q VGND VGND VPWR
+ VPWR _0142_ sky130_fd_sc_hd__mux4_2
XFILLER_97_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_143_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput507 net624 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput518 net635 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput529 net646 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_5_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1541_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG1 VGND VGND VPWR
+ VPWR net670 sky130_fd_sc_hd__buf_1
X_1472_ net460 VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__buf_4
XFILLER_113_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0423_ net65 net79 net63 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit14.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit15.Q
+ VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__mux4_1
XFILLER_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0354_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END0 net11 net113 net17
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit31.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit30.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG0
+ sky130_fd_sc_hd__mux4_1
XFILLER_94_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0285_ net34 net60 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13
+ _0057_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit24.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit25.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG1
+ sky130_fd_sc_hd__mux4_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_105 Tile_X0Y1_FrameStrobe[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_116 Tile_X0Y1_FrameStrobe[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_127 net640 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_138 net643 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0972_ net473 net379 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_30_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput304 net304 VGND VGND VPWR VPWR DI_SRAM20 sky130_fd_sc_hd__buf_2
Xoutput315 net315 VGND VGND VPWR VPWR DI_SRAM30 sky130_fd_sc_hd__buf_2
Xoutput326 net326 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[10] sky130_fd_sc_hd__buf_2
Xoutput359 net359 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
X_1524_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG0 VGND VGND VPWR
+ VPWR net651 sky130_fd_sc_hd__clkbuf_2
Xoutput337 net337 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[20] sky130_fd_sc_hd__buf_2
Xoutput348 net348 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[30] sky130_fd_sc_hd__buf_2
X_1455_ net212 VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__buf_4
X_1386_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb7 VGND VGND VPWR
+ VPWR net513 sky130_fd_sc_hd__buf_4
XFILLER_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0406_ net247 net136 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit13.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG3 sky130_fd_sc_hd__mux4_1
X_0337_ net238 net230 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG6
+ net131 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q
+ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_78_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0268_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q VGND
+ VGND VPWR VPWR _0047_ sky130_fd_sc_hd__inv_2
XFILLER_82_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1240_ net457 net383 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1171_ net452 net399 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_27 net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 net515 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_16 net327 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_49 net523 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0955_ net82 net385 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0886_ net87 net403 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_126_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1507_ Tile_X0Y0_S4END[11] VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__buf_4
XFILLER_141_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1438_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG2 VGND VGND VPWR
+ VPWR net571 sky130_fd_sc_hd__clkbuf_1
XFILLER_101_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1369_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG2 VGND VGND VPWR
+ VPWR net496 sky130_fd_sc_hd__buf_1
XFILLER_102_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout361 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG3 VGND VGND
+ VPWR VPWR net361 sky130_fd_sc_hd__buf_2
Xfanout383 net384 VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__clkbuf_2
Xfanout372 net219 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__buf_2
Xfanout394 net395 VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput14 DO_SRAM20 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
Xinput25 DO_SRAM30 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_2
X_0740_ net92 net445 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput36 Tile_X0Y0_E1END[3] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_4
Xinput58 Tile_X0Y0_E6END[3] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_2
Xinput69 Tile_X0Y0_EE4END[13] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_1
Xinput47 Tile_X0Y0_E2MID[2] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_1
X_0671_ _0046_ _0142_ _0185_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q
+ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__o211a_1
XFILLER_115_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1223_ net217 net390 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1154_ net193 net408 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1085_ net196 net426 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_63_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0938_ net471 net388 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0869_ net81 net411 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_87_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0723_ net90 net447 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0654_ net144 net182 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q
+ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__mux2_1
XFILLER_103_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0585_ net13 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG5 _0143_
+ _0082_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG10
+ sky130_fd_sc_hd__mux4_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1206_ net455 net390 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_0_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1137_ net210 net410 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_80_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1068_ net212 net435 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_103_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput226 Tile_X0Y1_N2END[2] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput215 Tile_X0Y1_FrameData[6] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_4
Xinput204 Tile_X0Y1_FrameData[25] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput237 Tile_X0Y1_N2MID[5] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_126_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0370_ net14 net22 net361 net360 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit30.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit31.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb4 sky130_fd_sc_hd__mux4_1
XFILLER_66_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_144_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0706_ net227 net146 net153 net147 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q VGND VGND VPWR
+ VPWR _0218_ sky130_fd_sc_hd__mux4_1
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0637_ _0029_ _0157_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q
+ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__a21o_1
X_0568_ net1 net5 _0141_ net366 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG12 sky130_fd_sc_hd__mux4_1
XFILLER_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0499_ net70 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit24.Q
+ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__nand2b_1
XFILLER_53_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput508 net625 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[2] sky130_fd_sc_hd__buf_2
X_1540_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG0 VGND VGND VPWR
+ VPWR net667 sky130_fd_sc_hd__clkbuf_2
Xoutput519 net636 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[14] sky130_fd_sc_hd__buf_2
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1471_ net461 VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__buf_4
XFILLER_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0422_ net78 net71 net62 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit12.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit13.Q
+ VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__mux4_2
XFILLER_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0353_ net141 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12 net167
+ _0090_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit15.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit14.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END0
+ sky130_fd_sc_hd__mux4_2
XFILLER_39_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0284_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END1 net245 net114
+ net134 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit2.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit3.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_33_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_106 Tile_X0Y1_FrameStrobe[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_128 net640 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_139 net643 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 Tile_X0Y1_FrameStrobe[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0971_ net99 net380 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_145_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput305 net305 VGND VGND VPWR VPWR DI_SRAM21 sky130_fd_sc_hd__buf_2
Xoutput316 net316 VGND VGND VPWR VPWR DI_SRAM31 sky130_fd_sc_hd__buf_2
XFILLER_153_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1523_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG3 VGND VGND VPWR
+ VPWR net650 sky130_fd_sc_hd__clkbuf_2
Xoutput327 net327 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[11] sky130_fd_sc_hd__buf_2
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput338 net338 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[21] sky130_fd_sc_hd__buf_2
Xoutput349 net349 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[31] sky130_fd_sc_hd__buf_2
X_1454_ net209 VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__buf_4
X_0405_ net246 net135 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit10.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit11.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_67_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1385_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb6 VGND VGND VPWR
+ VPWR net512 sky130_fd_sc_hd__clkbuf_2
X_0336_ net35 net46 net38 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit14.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit15.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG6
+ sky130_fd_sc_hd__mux4_1
X_0267_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q VGND
+ VGND VPWR VPWR _0046_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_53_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1170_ net451 net399 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_49_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_28 net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 net515 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 net333 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0954_ net83 net385 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0885_ net88 net404 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_113_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1506_ Tile_X0Y0_S4END[10] VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__buf_4
XFILLER_141_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1437_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG1 VGND VGND VPWR
+ VPWR net570 sky130_fd_sc_hd__clkbuf_1
X_1368_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG1 VGND VGND VPWR
+ VPWR net495 sky130_fd_sc_hd__buf_1
XFILLER_101_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0319_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb2 net127 net234
+ net119 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit13.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit12.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG2
+ sky130_fd_sc_hd__mux4_1
X_1299_ net452 net370 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout373 net374 VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_2
Xfanout384 net389 VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__clkbuf_2
Xfanout362 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG2 VGND VGND
+ VPWR VPWR net362 sky130_fd_sc_hd__clkbuf_4
Xfanout395 net397 VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput15 DO_SRAM21 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
Xinput26 DO_SRAM31 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
Xinput37 Tile_X0Y0_E2END[0] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_2
Xinput59 Tile_X0Y0_E6END[4] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_2
X_0670_ net169 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q
+ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__or2_1
Xinput48 Tile_X0Y0_E2MID[3] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1222_ net218 net390 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1153_ net466 net407 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1084_ net197 net426 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_63_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0937_ net470 net388 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0868_ net92 net411 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0799_ net109 net430 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0722_ net91 net447 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0653_ _0037_ _0141_ _0170_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q
+ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__o211a_1
X_0584_ net2 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG6 _0142_
+ _0081_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG9
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_149_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1205_ net454 net393 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_0_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1136_ net211 net410 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_83_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1067_ net213 net435 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_103_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput227 Tile_X0Y1_N2END[3] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_2
Xinput216 Tile_X0Y1_FrameData[7] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_4
Xinput205 Tile_X0Y1_FrameData[26] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__buf_1
Xinput238 Tile_X0Y1_N2MID[6] VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__buf_2
XFILLER_75_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_144_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0705_ net226 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q _0216_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q
+ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__o311a_1
XFILLER_131_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0636_ net141 net173 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q
+ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0567_ net223 net243 _0072_ net140 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q VGND VGND VPWR
+ VPWR _0141_ sky130_fd_sc_hd__mux4_2
X_0498_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG6 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit24.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit25.Q
+ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__mux4_1
X_1119_ net464 net416 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_13_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput509 net626 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[3] sky130_fd_sc_hd__buf_2
XFILLER_113_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1470_ net462 VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__buf_4
X_0421_ net77 net70 net61 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit10.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit11.Q
+ VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0352_ _0018_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q
+ _0087_ _0089_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_66_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0283_ net142 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13 net168
+ _0061_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit17.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit16.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END1
+ sky130_fd_sc_hd__mux4_2
XFILLER_62_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_75_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0619_ net180 net188 net164 _0143_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q VGND VGND VPWR
+ VPWR net292 sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_84_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_107 Tile_X0Y1_FrameStrobe[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_129 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 Tile_X0Y1_FrameStrobe[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_93_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0970_ net100 net380 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_145_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput317 net317 VGND VGND VPWR VPWR DI_SRAM4 sky130_fd_sc_hd__buf_2
Xoutput306 net306 VGND VGND VPWR VPWR DI_SRAM22 sky130_fd_sc_hd__buf_2
X_1522_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG2 VGND VGND VPWR
+ VPWR net649 sky130_fd_sc_hd__buf_1
Xoutput328 net328 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[12] sky130_fd_sc_hd__buf_2
Xoutput339 net339 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[22] sky130_fd_sc_hd__buf_2
XFILLER_113_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1453_ net198 VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__clkbuf_2
X_0404_ net245 net134 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG1 sky130_fd_sc_hd__mux4_1
X_1384_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb5 VGND VGND VPWR
+ VPWR net511 sky130_fd_sc_hd__clkbuf_2
X_0335_ net47 net39 net57 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit8.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit9.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG5
+ sky130_fd_sc_hd__mux4_1
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0266_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q VGND
+ VGND VPWR VPWR _0045_ sky130_fd_sc_hd__inv_1
XFILLER_82_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_29 net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_18 net335 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0953_ net84 net386 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0884_ net89 net404 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_113_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1505_ Tile_X0Y0_S4END[9] VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__buf_4
XFILLER_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1436_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG0 VGND VGND VPWR
+ VPWR net563 sky130_fd_sc_hd__clkbuf_2
X_1367_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG0 VGND VGND VPWR
+ VPWR net494 sky130_fd_sc_hd__buf_4
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0318_ net158 net150 net168 net367 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit26.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit27.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb2 sky130_fd_sc_hd__mux4_1
X_1298_ net451 net370 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0249_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q VGND VGND
+ VPWR VPWR _0028_ sky130_fd_sc_hd__inv_1
XFILLER_23_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_12_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout374 net376 VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkbuf_2
Xfanout363 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG1 VGND VGND
+ VPWR VPWR net363 sky130_fd_sc_hd__buf_2
Xfanout385 net387 VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_21_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout396 net397 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput27 DO_SRAM4 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
Xinput16 DO_SRAM22 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput49 Tile_X0Y0_E2MID[4] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_2
Xinput38 Tile_X0Y0_E2END[1] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1221_ net190 net393 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1152_ net465 net407 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1083_ net460 net425 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_63_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0936_ net469 net388 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0867_ net103 net411 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0798_ net110 net430 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1419_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb3 VGND VGND VPWR
+ VPWR net546 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_86_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0721_ net93 net447 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0652_ net163 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q
+ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__or2_1
X_0583_ net1 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG7 _0141_
+ net365 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG8
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_149_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1204_ net453 net393 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_0_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1135_ net189 net416 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_83_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1066_ net214 net435 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_33_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0919_ net86 net395 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_108_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput217 Tile_X0Y1_FrameData[8] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__buf_4
Xinput206 Tile_X0Y1_FrameData[27] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__buf_1
XFILLER_102_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput228 Tile_X0Y1_N2END[4] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_2
Xinput239 Tile_X0Y1_N2MID[7] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__buf_2
XFILLER_48_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_113_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_144_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0704_ net159 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q VGND VGND VPWR
+ VPWR _0216_ sky130_fd_sc_hd__or3b_1
X_0635_ _0028_ _0144_ _0155_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q
+ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__o211a_1
XFILLER_131_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0566_ net30 net4 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG4
+ net365 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG11
+ sky130_fd_sc_hd__mux4_1
X_0497_ _0015_ _0126_ _0130_ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG1
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_96_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1118_ net463 net416 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1049_ net458 net432 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_80_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0420_ net76 net69 net60 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG5
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit8.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit9.Q
+ VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__mux4_2
XFILLER_69_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0351_ net161 _0018_ _0088_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__o21a_1
X_0282_ _0020_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q
+ _0058_ _0060_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__a31o_1
XFILLER_85_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0618_ net173 net187 net161 _0144_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR
+ VPWR net291 sky130_fd_sc_hd__mux4_1
X_0549_ net13 net7 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13
+ _0081_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG2
+ sky130_fd_sc_hd__mux4_1
XFILLER_105_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_108 Tile_X0Y1_FrameStrobe[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_119 Tile_X0Y1_FrameStrobe[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput307 net307 VGND VGND VPWR VPWR DI_SRAM23 sky130_fd_sc_hd__buf_2
XFILLER_153_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1521_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG1 VGND VGND VPWR
+ VPWR net648 sky130_fd_sc_hd__clkbuf_1
Xoutput318 net318 VGND VGND VPWR VPWR DI_SRAM5 sky130_fd_sc_hd__buf_2
Xoutput329 net329 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[13] sky130_fd_sc_hd__buf_2
X_1452_ net189 VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0403_ net244 net133 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit6.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit7.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG0 sky130_fd_sc_hd__mux4_1
X_1383_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb4 VGND VGND VPWR
+ VPWR net510 sky130_fd_sc_hd__buf_2
X_0334_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb5 net130 net237
+ net122 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit19.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit18.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5
+ sky130_fd_sc_hd__mux4_2
XFILLER_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0265_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q VGND
+ VGND VPWR VPWR _0044_ sky130_fd_sc_hd__inv_2
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0952_ net85 net386 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_19 net338 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0883_ net90 net402 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_113_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1504_ Tile_X0Y0_S4END[8] VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__buf_4
X_1435_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG11 VGND VGND VPWR
+ VPWR net553 sky130_fd_sc_hd__clkbuf_2
X_1366_ Tile_X0Y1_FrameStrobe[19] VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__clkbuf_1
X_0317_ net234 net226 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG2
+ net127 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q
+ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__mux4_1
X_1297_ net450 net371 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0248_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q VGND
+ VGND VPWR VPWR _0027_ sky130_fd_sc_hd__inv_2
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout375 net376 VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkbuf_2
Xfanout364 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG0 VGND VGND
+ VPWR VPWR net364 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout386 net387 VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__buf_2
Xfanout397 Tile_X0Y1_FrameStrobe[6] VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput28 DO_SRAM5 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_2
Xinput17 DO_SRAM23 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
XFILLER_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput39 Tile_X0Y0_E2END[2] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlymetal6s2s_1
X_1220_ net191 net393 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1151_ net464 net407 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1082_ net459 net425 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_63_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0935_ net104 net388 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0866_ net106 net411 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_11_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0797_ net111 net428 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_114_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1418_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb2 VGND VGND VPWR
+ VPWR net545 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_86_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1349_ net428 VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__clkbuf_2
XFILLER_113_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput490 net607 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[6] sky130_fd_sc_hd__buf_2
XFILLER_154_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0720_ net94 net447 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_155_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0651_ _0166_ _0168_ _0169_ _0036_ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_10.A
+ sky130_fd_sc_hd__o22a_1
X_0582_ net30 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG4 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG8
+ net366 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG7
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_149_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1203_ net452 net390 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_77_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1134_ net198 net416 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_25_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1065_ net215 net435 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_80_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0918_ net87 net395 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0849_ net93 net415 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput218 Tile_X0Y1_FrameData[9] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__buf_4
Xinput207 Tile_X0Y1_FrameData[28] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__buf_1
Xinput229 Tile_X0Y1_N2END[5] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0703_ net238 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q _0214_ _0053_
+ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__o311a_1
X_0634_ net171 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q
+ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__or2_1
XFILLER_99_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0565_ net220 net240 _0087_ net137 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG4 sky130_fd_sc_hd__mux4_2
X_0496_ _0127_ _0128_ _0129_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit22.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit23.Q VGND VGND VPWR
+ VPWR _0130_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_96_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1117_ net462 net418 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_80_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1048_ net457 net432 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_80_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f_Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK VGND VGND VPWR VPWR clknet_1_0__leaf_Tile_X0Y1_UserCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0350_ net220 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q VGND VGND VPWR
+ VPWR _0088_ sky130_fd_sc_hd__o21ba_1
X_0281_ net164 _0020_ _0059_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__o21a_1
XFILLER_94_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0617_ net144 net186 net179 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q
+ VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__mux4_1
X_0548_ net2 net6 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14
+ _0082_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG1
+ sky130_fd_sc_hd__mux4_1
X_0479_ _0012_ _0111_ _0115_ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG2
+ sky130_fd_sc_hd__o21a_1
XANTENNA_109 Tile_X0Y1_FrameStrobe[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_141_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput308 net308 VGND VGND VPWR VPWR DI_SRAM24 sky130_fd_sc_hd__buf_2
XFILLER_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1520_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG0 VGND VGND VPWR
+ VPWR net647 sky130_fd_sc_hd__clkbuf_2
Xoutput319 net319 VGND VGND VPWR VPWR DI_SRAM6 sky130_fd_sc_hd__buf_2
X_1451_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG15 VGND VGND VPWR
+ VPWR net569 sky130_fd_sc_hd__clkbuf_2
X_1382_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb3 VGND VGND VPWR
+ VPWR net509 sky130_fd_sc_hd__buf_4
X_0402_ net12 net26 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG0
+ net364 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit4.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit5.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG15
+ sky130_fd_sc_hd__mux4_1
X_0333_ net155 net147 net165 _0081_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit0.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit1.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb5 sky130_fd_sc_hd__mux4_1
XFILLER_67_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0264_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q VGND
+ VGND VPWR VPWR _0043_ sky130_fd_sc_hd__inv_1
XFILLER_82_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0951_ net86 net386 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0882_ net91 net402 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_118_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1503_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG7 VGND VGND VPWR
+ VPWR net630 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1434_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG10 VGND VGND VPWR
+ VPWR net552 sky130_fd_sc_hd__clkbuf_1
XFILLER_99_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1365_ Tile_X0Y1_FrameStrobe[18] VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__clkbuf_1
X_0316_ net50 net42 net54 net362 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit6.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit7.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG2 sky130_fd_sc_hd__mux4_2
X_1296_ net449 net371 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0247_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q VGND
+ VGND VPWR VPWR _0026_ sky130_fd_sc_hd__inv_2
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout365 _0080_ VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout387 net388 VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__clkbuf_2
Xfanout398 net400 VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__clkbuf_2
Xfanout376 Tile_X0Y1_FrameStrobe[8] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput18 DO_SRAM24 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
XFILLER_52_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 DO_SRAM6 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_2
XFILLER_96_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1150_ net463 net407 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1081_ net458 net426 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_28_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0934_ net105 net388 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0865_ net107 net415 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_11_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0796_ net112 net428 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_114_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1417_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb1 VGND VGND VPWR
+ VPWR net544 sky130_fd_sc_hd__buf_1
XFILLER_114_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1348_ net437 VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__clkbuf_2
XFILLER_113_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1279_ net464 net375 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_94_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput480 net597 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[26] sky130_fd_sc_hd__buf_2
XFILLER_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput491 net608 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[7] sky130_fd_sc_hd__buf_2
XFILLER_27_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0650_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG6
+ net367 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG10 _0035_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q
+ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__mux4_1
XFILLER_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0581_ net29 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG5 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG9
+ net367 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG6
+ sky130_fd_sc_hd__mux4_1
XFILLER_88_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1202_ net451 net390 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1133_ net209 net418 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_92_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1064_ net216 net435 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0917_ net88 net394 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0848_ net94 net415 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0779_ net472 net427 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput208 Tile_X0Y1_FrameData[29] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__buf_1
Xinput219 Tile_X0Y1_FrameStrobe[9] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_4
XFILLER_84_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_18_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0702_ net156 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q VGND VGND VPWR
+ VPWR _0214_ sky130_fd_sc_hd__or3b_1
XFILLER_116_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0633_ net144 net186 net179 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q
+ VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__mux4_2
X_0564_ net29 net3 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG5
+ _0081_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG10
+ sky130_fd_sc_hd__mux4_1
X_0495_ net60 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG1 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit21.Q
+ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__mux2_1
XFILLER_57_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1116_ net461 net418 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_65_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1047_ net456 net432 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0280_ net221 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q VGND VGND VPWR
+ VPWR _0059_ sky130_fd_sc_hd__o21ba_1
XFILLER_94_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_44_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0616_ net143 net185 net178 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q
+ VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__mux4_2
X_0547_ net1 net5 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15
+ _0083_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG0
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0478_ _0112_ _0113_ _0114_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit21.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit22.Q VGND VGND VPWR
+ VPWR _0115_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_53_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput309 net309 VGND VGND VPWR VPWR DI_SRAM25 sky130_fd_sc_hd__buf_2
X_1450_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG14 VGND VGND VPWR
+ VPWR net568 sky130_fd_sc_hd__clkbuf_1
X_1381_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb2 VGND VGND VPWR
+ VPWR net508 sky130_fd_sc_hd__clkbuf_2
X_0401_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END0 net244 net113
+ net133 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit8.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit9.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG0
+ sky130_fd_sc_hd__mux4_2
XFILLER_67_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0332_ net237 net229 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG5
+ net130 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q
+ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__mux4_2
XFILLER_96_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0263_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q VGND
+ VGND VPWR VPWR _0042_ sky130_fd_sc_hd__inv_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_140_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0950_ net87 net385 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0881_ net93 net403 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1502_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG6 VGND VGND VPWR
+ VPWR net629 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1433_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG9 VGND VGND VPWR
+ VPWR net562 sky130_fd_sc_hd__clkbuf_1
X_1364_ Tile_X0Y1_FrameStrobe[17] VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__clkbuf_1
X_1295_ net189 net373 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0315_ net51 net43 net61 net363 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit0.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit1.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG1 sky130_fd_sc_hd__mux4_1
X_0246_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q VGND
+ VGND VPWR VPWR _0025_ sky130_fd_sc_hd__inv_2
XFILLER_70_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout366 _0079_ VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__buf_2
XFILLER_143_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout377 net379 VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__clkbuf_4
Xfanout399 net400 VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__clkbuf_2
Xfanout388 net389 VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__buf_2
XFILLER_100_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput19 DO_SRAM25 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1080_ net457 net426 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0933_ net81 net395 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0864_ net108 net415 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0795_ net82 net427 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_114_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1416_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb0 VGND VGND VPWR
+ VPWR net543 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1347_ net447 VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__buf_4
XFILLER_95_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1278_ net463 net375 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0229_ net150 VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput470 net587 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[17] sky130_fd_sc_hd__buf_2
Xoutput481 net598 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[27] sky130_fd_sc_hd__buf_2
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput492 net609 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[8] sky130_fd_sc_hd__buf_2
XFILLER_47_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0580_ net28 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG10 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG6
+ net368 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG5
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_149_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1201_ net450 net393 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1132_ net212 net418 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1063_ net217 net432 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_0_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0916_ net89 net394 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0847_ net476 net412 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0778_ net471 net429 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput209 Tile_X0Y1_FrameData[2] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__buf_2
XFILLER_75_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0701_ _0008_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q _0211_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q
+ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_155_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0632_ net143 net185 net178 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q
+ VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__mux4_2
XFILLER_143_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0563_ net221 net241 _0058_ net138 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG5 sky130_fd_sc_hd__mux4_2
XFILLER_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0494_ net34 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit21.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit22.Q VGND VGND VPWR
+ VPWR _0128_ sky130_fd_sc_hd__o21ba_1
X_1115_ net199 net417 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1046_ net455 net432 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_143_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0615_ net142 net184 net177 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q
+ VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__mux4_2
XFILLER_124_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0546_ net30 net8 net369 _0083_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb7 sky130_fd_sc_hd__mux4_1
X_0477_ net54 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG2 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit20.Q
+ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_0_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1029_ net190 net442 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_154_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1380_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb1 VGND VGND VPWR
+ VPWR net507 sky130_fd_sc_hd__clkbuf_2
X_0400_ net11 net25 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG1
+ net363 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit2.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit3.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG14
+ sky130_fd_sc_hd__mux4_1
X_0331_ net34 net47 net39 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit12.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit13.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG5
+ sky130_fd_sc_hd__mux4_1
XFILLER_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0262_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q VGND
+ VGND VPWR VPWR _0041_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_78_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0529_ net222 net1 _0065_ net28 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0880_ net94 net403 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_126_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1501_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG5 VGND VGND VPWR
+ VPWR net628 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_81_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1432_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG8 VGND VGND VPWR
+ VPWR net561 sky130_fd_sc_hd__buf_1
X_1363_ Tile_X0Y1_FrameStrobe[16] VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__clkbuf_1
X_1294_ net198 net373 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0314_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb1 net126 net233
+ net118 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit11.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit10.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG1
+ sky130_fd_sc_hd__mux4_1
X_0245_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q VGND
+ VGND VPWR VPWR _0024_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_90_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout378 net379 VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__buf_2
Xfanout367 _0078_ VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__buf_2
Xfanout389 Tile_X0Y1_FrameStrobe[7] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_2
XFILLER_100_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_129_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_138_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0932_ net92 net395 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0863_ net109 net415 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0794_ net83 net429 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1415_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG7 VGND VGND VPWR
+ VPWR net542 sky130_fd_sc_hd__clkbuf_2
X_1346_ net467 VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__buf_1
XFILLER_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1277_ net462 net375 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0228_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit7.Q VGND VGND
+ VPWR VPWR _0007_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput460 net577 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput471 net588 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[18] sky130_fd_sc_hd__buf_2
Xoutput482 net599 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[28] sky130_fd_sc_hd__buf_2
Xoutput493 net610 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[9] sky130_fd_sc_hd__buf_2
XFILLER_120_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_146_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_155_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_149_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1200_ net449 net393 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_77_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1131_ net213 net417 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1062_ net218 net432 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_91_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0915_ net90 net396 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_111_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0846_ net475 net412 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0777_ net470 net430 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1329_ net86 VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkbuf_1
XFILLER_140_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput290 net290 VGND VGND VPWR VPWR CLOCK_SRAM sky130_fd_sc_hd__buf_1
XFILLER_74_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0700_ net148 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q VGND VGND VPWR
+ VPWR _0212_ sky130_fd_sc_hd__nor3_1
XFILLER_128_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0631_ net142 net184 net177 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q
+ VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__mux4_2
XFILLER_99_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0562_ net28 net32 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG6
+ _0082_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG9
+ sky130_fd_sc_hd__mux4_1
XFILLER_151_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0493_ net69 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit21.Q
+ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__nand2b_1
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1114_ net200 net417 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_53_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1045_ net454 net434 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_80_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0829_ net111 net421 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_130_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_143_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0614_ net141 net183 net176 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q
+ VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__mux4_1
XFILLER_116_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0545_ net29 net7 net368 _0082_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb6 sky130_fd_sc_hd__mux4_1
XFILLER_112_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0476_ net35 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit20.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit21.Q VGND VGND VPWR
+ VPWR _0113_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1028_ net191 net442 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_101_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_110_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0330_ net48 net40 net58 net360 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit6.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit7.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG4 sky130_fd_sc_hd__mux4_1
XFILLER_121_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0261_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q VGND
+ VGND VPWR VPWR _0040_ sky130_fd_sc_hd__inv_1
XFILLER_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0528_ net221 net24 _0058_ net29 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_58_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0459_ net49 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit7.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit6.Q VGND VGND VPWR
+ VPWR _0099_ sky130_fd_sc_hd__o21ba_1
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1500_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG4 VGND VGND VPWR
+ VPWR net627 sky130_fd_sc_hd__clkbuf_2
X_1431_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG7 VGND VGND VPWR
+ VPWR net560 sky130_fd_sc_hd__buf_1
XFILLER_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1362_ Tile_X0Y1_FrameStrobe[15] VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__clkbuf_1
XFILLER_95_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1293_ net209 net373 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0313_ net159 net151 net169 net368 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit24.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit25.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb1 sky130_fd_sc_hd__mux4_1
X_0244_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q VGND
+ VGND VPWR VPWR _0023_ sky130_fd_sc_hd__inv_2
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput190 Tile_X0Y1_FrameData[10] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_4
XFILLER_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout379 net380 VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__clkbuf_2
Xfanout368 _0077_ VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkbuf_4
XFILLER_100_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0931_ net103 net397 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0862_ net110 net415 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0793_ net84 net430 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1414_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG6 VGND VGND VPWR
+ VPWR net541 sky130_fd_sc_hd__clkbuf_1
X_1345_ net468 VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__buf_1
X_1276_ net461 net375 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0227_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit4.Q VGND VGND
+ VPWR VPWR _0006_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput461 net578 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput450 net567 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput483 net600 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[29] sky130_fd_sc_hd__buf_2
Xoutput494 net611 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput472 net589 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[19] sky130_fd_sc_hd__buf_2
XFILLER_120_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1130_ net214 net417 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_77_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1061_ net190 net434 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_16_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0914_ net91 net396 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_111_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0845_ net474 net411 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_119_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0776_ net469 net430 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1328_ net85 VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__buf_1
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1259_ net213 net381 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput280 net280 VGND VGND VPWR VPWR BEN_SRAM29 sky130_fd_sc_hd__buf_2
Xoutput291 net291 VGND VGND VPWR VPWR DI_SRAM0 sky130_fd_sc_hd__buf_2
XFILLER_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0630_ net141 net183 net176 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q
+ VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__mux4_1
XFILLER_143_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0561_ net222 net242 _0065_ net139 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG6 sky130_fd_sc_hd__mux4_2
XFILLER_99_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0492_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit21.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit22.Q
+ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__mux4_1
X_1113_ net201 net417 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1044_ net453 net434 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_65_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0828_ net112 net421 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0759_ net86 net437 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_23_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0613_ net182 net175 net163 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG11
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q
+ VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__mux4_1
X_0544_ net28 net6 net367 _0081_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb5 sky130_fd_sc_hd__mux4_1
X_0475_ net73 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit20.Q
+ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__nand2b_1
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1027_ net192 net443 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0260_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q VGND
+ VGND VPWR VPWR _0039_ sky130_fd_sc_hd__inv_1
XFILLER_121_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0527_ net220 net13 _0087_ net30 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_112_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0458_ _0098_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit5.Q
+ _0006_ _0097_ VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__a2bb2o_2
X_0389_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END2 net246 net115
+ net135 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit20.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit21.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG6
+ sky130_fd_sc_hd__mux4_2
XFILLER_14_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1430_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG6 VGND VGND VPWR
+ VPWR net559 sky130_fd_sc_hd__clkbuf_1
X_1361_ Tile_X0Y1_FrameStrobe[14] VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__clkbuf_1
X_0312_ net233 net225 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG1
+ net126 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q
+ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__mux4_1
X_1292_ net212 net373 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput180 Tile_X0Y1_EE4END[1] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__dlymetal6s2s_1
X_0243_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q VGND
+ VGND VPWR VPWR _0022_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput191 Tile_X0Y1_FrameData[11] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_4
XFILLER_16_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1559_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG7 VGND VGND VPWR
+ VPWR net692 sky130_fd_sc_hd__buf_1
Xfanout369 _0076_ VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__clkbuf_4
XFILLER_98_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0930_ net106 net397 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_9_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0861_ net111 net413 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0792_ net85 net430 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1413_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG5 VGND VGND VPWR
+ VPWR net540 sky130_fd_sc_hd__clkbuf_1
X_1344_ net469 VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__buf_1
X_1275_ net460 net374 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_95_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0226_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit2.Q VGND VGND
+ VPWR VPWR _0005_ sky130_fd_sc_hd__inv_2
XFILLER_95_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput451 net568 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput462 net579 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[0] sky130_fd_sc_hd__buf_2
Xoutput440 net557 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[4] sky130_fd_sc_hd__buf_2
Xoutput495 net612 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[1] sky130_fd_sc_hd__buf_2
Xoutput473 net590 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[1] sky130_fd_sc_hd__buf_2
Xoutput484 net601 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[2] sky130_fd_sc_hd__buf_2
XFILLER_86_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_69_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1060_ net191 net434 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_78_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0913_ net93 net395 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_306 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0844_ net473 net411 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_119_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0775_ net468 net427 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1327_ net84 VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_39_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1258_ net214 net381 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1189_ net190 net406 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_82_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_96_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput270 net270 VGND VGND VPWR VPWR BEN_SRAM2 sky130_fd_sc_hd__buf_2
Xoutput281 net281 VGND VGND VPWR VPWR BEN_SRAM3 sky130_fd_sc_hd__buf_2
Xoutput292 net292 VGND VGND VPWR VPWR DI_SRAM1 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0560_ net27 net31 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG7
+ _0083_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG8
+ sky130_fd_sc_hd__mux4_1
X_0491_ _0014_ _0121_ _0125_ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG0
+ sky130_fd_sc_hd__o21a_1
XFILLER_97_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1112_ net202 net417 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1043_ net452 net433 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_125_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0827_ net82 net422 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0758_ net87 net439 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_135_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0689_ net156 net159 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
+ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__mux2_1
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0612_ net181 net174 net162 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG10
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q
+ VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__mux4_2
XFILLER_124_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0543_ net27 net5 net366 net365 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb4 sky130_fd_sc_hd__mux4_1
X_0474_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG6 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14 net362 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit20.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit21.Q VGND VGND VPWR
+ VPWR _0111_ sky130_fd_sc_hd__mux4_1
X_1026_ net193 net443 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_134_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0526_ net144 net145 net153 _0083_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG7 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_69_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0457_ net40 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit4.Q
+ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__nand2_1
XFILLER_112_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0388_ net14 net18 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit22.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit23.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG8 sky130_fd_sc_hd__mux4_1
X_1009_ net450 net440 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_140_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1360_ Tile_X0Y1_FrameStrobe[13] VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_50_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0311_ net51 net43 net64 net363 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit4.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit5.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG1 sky130_fd_sc_hd__mux4_2
X_1291_ net213 net374 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput181 Tile_X0Y1_EE4END[2] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput170 Tile_X0Y1_E6END[7] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__buf_2
X_0242_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q VGND
+ VGND VPWR VPWR _0021_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput192 Tile_X0Y1_FrameData[12] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_4
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1558_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG6 VGND VGND VPWR
+ VPWR net691 sky130_fd_sc_hd__buf_1
XFILLER_143_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0509_ _0017_ _0136_ _0140_ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG3
+ sky130_fd_sc_hd__o21a_1
X_1489_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG1 VGND VGND VPWR
+ VPWR net616 sky130_fd_sc_hd__clkbuf_2
XFILLER_54_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_107_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_116_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0860_ net112 net413 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0791_ net86 net430 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_125_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1412_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG4 VGND VGND VPWR
+ VPWR net539 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1343_ net470 VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__buf_1
XFILLER_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1274_ net459 net374 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_134_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0225_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit0.Q VGND VGND
+ VPWR VPWR _0004_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0989_ net111 net378 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput430 net547 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput452 net569 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[15] sky130_fd_sc_hd__buf_2
XFILLER_105_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput441 net558 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[5] sky130_fd_sc_hd__buf_2
Xoutput485 net602 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[30] sky130_fd_sc_hd__buf_2
Xoutput496 net613 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_59_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput463 net580 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[10] sky130_fd_sc_hd__buf_2
Xoutput474 net591 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[20] sky130_fd_sc_hd__buf_2
XFILLER_113_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0912_ net94 net396 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0843_ net472 net411 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_119_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0774_ net467 net427 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_142_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1326_ net83 VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__buf_2
XFILLER_83_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1257_ net215 net381 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_140_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1188_ net191 net406 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_82_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput260 net260 VGND VGND VPWR VPWR BEN_SRAM10 sky130_fd_sc_hd__buf_2
Xoutput271 net271 VGND VGND VPWR VPWR BEN_SRAM20 sky130_fd_sc_hd__buf_2
XFILLER_59_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput282 net282 VGND VGND VPWR VPWR BEN_SRAM30 sky130_fd_sc_hd__buf_2
Xoutput293 net293 VGND VGND VPWR VPWR DI_SRAM10 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0490_ _0122_ _0123_ _0124_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit19.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit20.Q VGND VGND VPWR
+ VPWR _0125_ sky130_fd_sc_hd__a221o_1
XFILLER_97_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1111_ net456 net419 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1042_ net451 net433 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_125_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0826_ net83 net422 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0757_ net88 net438 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_135_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0688_ _0198_ _0199_ _0200_ _0197_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__a31o_1
XFILLER_29_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1309_ net462 net371 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_56_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0611_ net180 net188 net172 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG9
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q
+ VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__mux4_2
X_0542_ net24 net4 net366 net365 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb3 sky130_fd_sc_hd__mux4_1
X_0473_ _0011_ _0106_ _0110_ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG1
+ sky130_fd_sc_hd__o21a_1
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1025_ net466 net442 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0809_ net470 net423 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_115_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_1 net256 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0525_ net143 net146 net154 _0082_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG6 sky130_fd_sc_hd__mux4_1
X_0456_ net48 net361 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit5.Q
+ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0387_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END3 net247 net116
+ net136 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit22.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit23.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG7
+ sky130_fd_sc_hd__mux4_2
XFILLER_81_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1008_ net449 net440 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0310_ net52 net44 net62 net364 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit30.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit31.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG0 sky130_fd_sc_hd__mux4_1
X_1290_ net214 net374 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput160 Tile_X0Y1_E2MID[7] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_2
Xinput171 Tile_X0Y1_E6END[8] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_2
X_0241_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q VGND
+ VGND VPWR VPWR _0020_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput182 Tile_X0Y1_EE4END[3] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput193 Tile_X0Y1_FrameData[13] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_4
XFILLER_149_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1557_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG5 VGND VGND VPWR
+ VPWR net690 sky130_fd_sc_hd__buf_1
X_0508_ _0137_ _0138_ _0139_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit28.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit29.Q VGND VGND VPWR
+ VPWR _0140_ sky130_fd_sc_hd__a221o_1
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1488_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG0 VGND VGND VPWR
+ VPWR net615 sky130_fd_sc_hd__clkbuf_2
X_0439_ net65 net79 net63 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit14.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit15.Q
+ VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_109_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0790_ net87 net430 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_11_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1411_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG3 VGND VGND VPWR
+ VPWR net538 sky130_fd_sc_hd__buf_1
X_1342_ net471 VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1273_ net458 net376 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0224_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit30.Q VGND
+ VGND VPWR VPWR _0003_ sky130_fd_sc_hd__inv_2
XFILLER_83_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0988_ net112 net378 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput420 net537 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_105_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput431 net548 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput453 net570 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_105_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput442 net559 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[6] sky130_fd_sc_hd__buf_2
Xoutput486 net603 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[31] sky130_fd_sc_hd__buf_2
Xoutput464 net581 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[11] sky130_fd_sc_hd__buf_2
Xoutput475 net592 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[21] sky130_fd_sc_hd__buf_2
Xoutput497 net614 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_59_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0911_ net476 net394 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0842_ net471 net411 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_119_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0773_ net81 net436 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_142_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1325_ net82 VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__clkbuf_2
XFILLER_110_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1256_ net216 net382 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1187_ net192 net399 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_82_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput250 net250 VGND VGND VPWR VPWR AD_SRAM2 sky130_fd_sc_hd__buf_2
Xoutput261 net261 VGND VGND VPWR VPWR BEN_SRAM11 sky130_fd_sc_hd__buf_2
Xoutput272 net272 VGND VGND VPWR VPWR BEN_SRAM21 sky130_fd_sc_hd__buf_2
Xoutput283 net283 VGND VGND VPWR VPWR BEN_SRAM31 sky130_fd_sc_hd__buf_2
Xoutput294 net294 VGND VGND VPWR VPWR DI_SRAM11 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1110_ net455 net419 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_65_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1041_ net450 net432 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_53_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0825_ net84 net420 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0756_ net89 net438 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_142_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0687_ _0009_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q VGND VGND VPWR
+ VPWR _0200_ sky130_fd_sc_hd__a21oi_1
XFILLER_130_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1308_ net461 net371 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1239_ net456 net382 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_44_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_152_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0610_ net173 net187 net171 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG8
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q
+ VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__mux4_1
X_0541_ net13 net3 net367 _0081_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb2 sky130_fd_sc_hd__mux4_1
X_0472_ _0107_ _0108_ _0109_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit18.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit19.Q VGND VGND VPWR
+ VPWR _0110_ sky130_fd_sc_hd__a221o_1
XFILLER_26_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1024_ net465 net442 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0808_ net469 net423 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0739_ net103 net446 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_103_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_2 net267 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0524_ net142 net147 net155 _0081_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG5 sky130_fd_sc_hd__mux4_1
XFILLER_58_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0455_ _0096_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit3.Q
+ _0005_ _0095_ VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_69_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0386_ net17 net21 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG8
+ net364 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit20.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit21.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG7
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_77_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1007_ net476 net372 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_41_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0240_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit25.Q VGND
+ VGND VPWR VPWR _0019_ sky130_fd_sc_hd__inv_1
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput150 Tile_X0Y1_E2END[5] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
Xinput161 Tile_X0Y1_E6END[0] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_2
Xinput172 Tile_X0Y1_E6END[9] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_66_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput183 Tile_X0Y1_EE4END[4] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_2
Xinput194 Tile_X0Y1_FrameData[14] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__buf_1
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1556_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG4 VGND VGND VPWR
+ VPWR net689 sky130_fd_sc_hd__buf_1
XFILLER_140_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0507_ net62 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG3 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit27.Q
+ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__mux2_1
X_1487_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG3 VGND VGND VPWR
+ VPWR net614 sky130_fd_sc_hd__buf_1
XFILLER_98_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0438_ net78 net71 net62 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit12.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit13.Q
+ VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__mux4_2
X_0369_ net12 net21 net361 net360 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit28.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit29.Q VGND VGND VPWR
+ VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb3 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_109_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1410_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG2 VGND VGND VPWR
+ VPWR net537 sky130_fd_sc_hd__clkbuf_1
X_1341_ net472 VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkbuf_2
X_1272_ net457 net376 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_67_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0223_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit31.Q VGND
+ VGND VPWR VPWR _0002_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_106_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0987_ net82 net378 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput410 net527 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput421 net538 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput432 net549 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput443 net560 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_154_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput454 net571 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput487 net604 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[3] sky130_fd_sc_hd__buf_2
Xoutput465 net582 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[12] sky130_fd_sc_hd__buf_2
Xoutput476 net593 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[22] sky130_fd_sc_hd__buf_2
X_1539_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb7 VGND VGND VPWR
+ VPWR net666 sky130_fd_sc_hd__buf_1
Xoutput498 net615 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_59_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0910_ net475 net394 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0841_ net470 net415 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_119_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0772_ net92 net436 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_142_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_47_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1324_ net112 VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1255_ net217 net381 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1186_ net193 net399 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_56_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_65_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput251 net251 VGND VGND VPWR VPWR AD_SRAM3 sky130_fd_sc_hd__buf_2
Xoutput262 net262 VGND VGND VPWR VPWR BEN_SRAM12 sky130_fd_sc_hd__buf_2
XFILLER_59_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput284 net284 VGND VGND VPWR VPWR BEN_SRAM4 sky130_fd_sc_hd__buf_2
Xoutput273 net273 VGND VGND VPWR VPWR BEN_SRAM22 sky130_fd_sc_hd__buf_2
Xoutput295 net295 VGND VGND VPWR VPWR DI_SRAM12 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_74_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1040_ net449 net432 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_73_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0824_ net85 net420 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_127_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0755_ net90 net437 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_142_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0686_ _0008_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q VGND VGND VPWR
+ VPWR _0199_ sky130_fd_sc_hd__o21ai_1
XFILLER_142_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1307_ net460 net370 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1238_ net455 net382 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1169_ net450 net401 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_35_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0540_ net2 net32 net368 _0082_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb1 sky130_fd_sc_hd__mux4_1
XFILLER_124_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0471_ net64 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG1 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit17.Q
+ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__mux2_1
XFILLER_38_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1023_ net464 net443 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_34_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0807_ net468 net420 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0738_ net106 net446 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0669_ _0181_ _0183_ _0184_ _0045_ VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG1
+ sky130_fd_sc_hd__o22a_1
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_3 net268 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0523_ net141 net148 net156 net365 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG4 sky130_fd_sc_hd__mux4_1
X_0454_ net39 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit2.Q
+ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__nand2_1
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0385_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END0 net244 net113
+ net133 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit24.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit25.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG8
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_77_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1006_ net475 net372 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_60_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_151_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput140 Tile_X0Y0_S4END[7] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_4
Xinput151 Tile_X0Y1_E2END[6] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__buf_1
Xinput162 Tile_X0Y1_E6END[10] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_2
Xinput173 Tile_X0Y1_EE4END[0] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_2
Xinput184 Tile_X0Y1_EE4END[5] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__buf_1
XFILLER_48_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput195 Tile_X0Y1_FrameData[15] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_74_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1555_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG3 VGND VGND VPWR
+ VPWR net688 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0506_ net36 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit27.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit28.Q VGND VGND VPWR
+ VPWR _0138_ sky130_fd_sc_hd__o21ba_1
X_1486_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG2 VGND VGND VPWR
+ VPWR net613 sky130_fd_sc_hd__buf_1
X_0437_ net77 net70 net61 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit10.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit11.Q
+ VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__mux4_2
X_0368_ net11 net20 net362 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit26.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit27.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb2
+ sky130_fd_sc_hd__mux4_1
XFILLER_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0299_ net36 net55 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15
+ _0071_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit0.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit1.Q
+ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__mux4_2
XFILLER_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1340_ net473 VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__clkbuf_2
XFILLER_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1271_ net456 net375 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_95_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0222_ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit29.Q VGND
+ VGND VPWR VPWR _0001_ sky130_fd_sc_hd__inv_1
XFILLER_51_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_103_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_Tile_X0Y1_UserCLK Tile_X0Y1_UserCLK VGND VGND VPWR VPWR clknet_0_Tile_X0Y1_UserCLK
+ sky130_fd_sc_hd__clkbuf_16
X_0986_ net83 net378 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput400 net517 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput411 net528 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput422 net539 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput433 net550 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput444 net561 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[8] sky130_fd_sc_hd__buf_2
Xoutput455 net572 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput466 net583 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[13] sky130_fd_sc_hd__buf_2
Xoutput477 net594 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput499 net616 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[1] sky130_fd_sc_hd__buf_2
X_1538_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb6 VGND VGND VPWR
+ VPWR net665 sky130_fd_sc_hd__buf_1
Xoutput488 net605 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[4] sky130_fd_sc_hd__buf_2
X_1469_ Tile_X0Y1_FrameData[17] VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_2_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0840_ net469 net415 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0771_ net103 net436 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1323_ net111 VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__clkbuf_2
X_1254_ net218 net381 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1185_ net466 net398 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0969_ net470 net377 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput252 net252 VGND VGND VPWR VPWR AD_SRAM4 sky130_fd_sc_hd__buf_2
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput285 net285 VGND VGND VPWR VPWR BEN_SRAM5 sky130_fd_sc_hd__buf_2
Xoutput263 net263 VGND VGND VPWR VPWR BEN_SRAM13 sky130_fd_sc_hd__buf_2
Xoutput274 net274 VGND VGND VPWR VPWR BEN_SRAM23 sky130_fd_sc_hd__buf_2
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput296 net296 VGND VGND VPWR VPWR DI_SRAM13 sky130_fd_sc_hd__buf_2
XFILLER_74_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0823_ net86 net420 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_136_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0754_ net91 net437 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0685_ net148 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q VGND VGND VPWR
+ VPWR _0198_ sky130_fd_sc_hd__or3_1
XFILLER_142_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1306_ net459 net370 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_96_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1237_ net454 net382 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1168_ net449 net401 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_35_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1099_ net213 net425 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_12_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0470_ net34 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit17.Q
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit18.Q VGND VGND VPWR
+ VPWR _0108_ sky130_fd_sc_hd__o21ba_1
X_1022_ net463 net443 VGND VGND VPWR VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_34_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0806_ net467 net420 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0737_ net107 net446 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_115_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0668_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG5
+ _0081_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG9 _0044_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q
+ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__mux4_1
X_0599_ net157 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q VGND VGND VPWR
+ VPWR _0153_ sky130_fd_sc_hd__o21ba_1
XFILLER_69_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_4 net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0522_ net157 net149 net163 net366 Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q
+ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q VGND VGND VPWR
+ VPWR Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0453_ net47 net362 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit3.Q
+ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__mux2_1
XFILLER_112_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0384_ net16 net20 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG9
+ net363 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit18.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit19.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG6
+ sky130_fd_sc_hd__mux4_1
XFILLER_66_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1005_ net474 net372 VGND VGND VPWR VPWR Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_149_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput130 Tile_X0Y0_S2MID[5] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
Xinput141 Tile_X0Y1_E1END[0] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__buf_2
Xinput152 Tile_X0Y1_E2END[7] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
Xinput163 Tile_X0Y1_E6END[11] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
Xinput185 Tile_X0Y1_EE4END[6] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__buf_1
Xinput174 Tile_X0Y1_EE4END[10] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__buf_1
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput196 Tile_X0Y1_FrameData[18] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1554_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG2 VGND VGND VPWR
+ VPWR net687 sky130_fd_sc_hd__buf_1
XFILLER_140_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0505_ net71 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit27.Q
+ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__nand2b_1
XFILLER_125_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1485_ Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG1 VGND VGND VPWR
+ VPWR net612 sky130_fd_sc_hd__clkbuf_2
X_0436_ net76 net69 net60 Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG5
+ Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit8.Q Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit9.Q
+ VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__mux4_2
.ends

