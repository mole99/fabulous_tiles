module N_term_DSP (UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1END,
    N2END,
    N2MID,
    N4END,
    NN4END,
    S1BEG,
    S2BEG,
    S2BEGb,
    S4BEG,
    SS4BEG);
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] N1END;
 input [7:0] N2END;
 input [7:0] N2MID;
 input [15:0] N4END;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 output [15:0] S4BEG;
 output [15:0] SS4BEG;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;

 sky130_fd_sc_hd__buf_1 _000_ (.A(FrameData[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 _001_ (.A(FrameData[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 _002_ (.A(FrameData[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 _003_ (.A(FrameData[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 _004_ (.A(FrameData[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 _005_ (.A(FrameData[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 _006_ (.A(FrameData[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 _007_ (.A(FrameData[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 _008_ (.A(FrameData[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 _009_ (.A(FrameData[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 _010_ (.A(FrameData[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 _011_ (.A(FrameData[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 _012_ (.A(FrameData[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 _013_ (.A(FrameData[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 _014_ (.A(FrameData[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 _015_ (.A(FrameData[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 _016_ (.A(FrameData[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 _017_ (.A(FrameData[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 _018_ (.A(FrameData[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 _019_ (.A(FrameData[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 _020_ (.A(FrameData[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 _021_ (.A(FrameData[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 _022_ (.A(FrameData[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 _023_ (.A(FrameData[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 _024_ (.A(FrameData[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 _025_ (.A(FrameData[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 _026_ (.A(FrameData[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 _027_ (.A(FrameData[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 _028_ (.A(FrameData[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 _029_ (.A(FrameData[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 _030_ (.A(FrameData[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 _031_ (.A(FrameData[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 _032_ (.A(FrameStrobe[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 _033_ (.A(FrameStrobe[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 _034_ (.A(FrameStrobe[2]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 _035_ (.A(FrameStrobe[3]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 _036_ (.A(FrameStrobe[4]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 _037_ (.A(FrameStrobe[5]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 _038_ (.A(FrameStrobe[6]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 _039_ (.A(FrameStrobe[7]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 _040_ (.A(FrameStrobe[8]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 _041_ (.A(FrameStrobe[9]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 _042_ (.A(FrameStrobe[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 _043_ (.A(FrameStrobe[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 _044_ (.A(FrameStrobe[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 _045_ (.A(FrameStrobe[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 _046_ (.A(FrameStrobe[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 _047_ (.A(FrameStrobe[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 _048_ (.A(FrameStrobe[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 _049_ (.A(FrameStrobe[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 _050_ (.A(FrameStrobe[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 _051_ (.A(FrameStrobe[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 _052_ (.A(N1END[3]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 _053_ (.A(N1END[2]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 _054_ (.A(N1END[1]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 _055_ (.A(N1END[0]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 _056_ (.A(N2MID[7]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 _057_ (.A(N2MID[6]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 _058_ (.A(N2MID[5]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 _059_ (.A(N2MID[4]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 _060_ (.A(N2MID[3]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 _061_ (.A(N2MID[2]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 _062_ (.A(N2MID[1]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 _063_ (.A(N2MID[0]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 _064_ (.A(N2END[7]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 _065_ (.A(N2END[6]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 _066_ (.A(N2END[5]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _067_ (.A(N2END[4]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _068_ (.A(N2END[3]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _069_ (.A(N2END[2]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _070_ (.A(N2END[1]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 _071_ (.A(N2END[0]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _072_ (.A(N4END[15]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 _073_ (.A(N4END[14]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _074_ (.A(N4END[13]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 _075_ (.A(N4END[12]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _076_ (.A(N4END[11]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 _077_ (.A(N4END[10]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 _078_ (.A(N4END[9]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _079_ (.A(N4END[8]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 _080_ (.A(N4END[7]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 _081_ (.A(N4END[6]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 _082_ (.A(N4END[5]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 _083_ (.A(N4END[4]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _084_ (.A(N4END[3]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _085_ (.A(N4END[2]),
    .X(net77));
 sky130_fd_sc_hd__buf_1 _086_ (.A(N4END[1]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 _087_ (.A(N4END[0]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _088_ (.A(NN4END[15]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 _089_ (.A(NN4END[14]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _090_ (.A(NN4END[13]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _091_ (.A(NN4END[12]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 _092_ (.A(NN4END[11]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 _093_ (.A(NN4END[10]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 _094_ (.A(NN4END[9]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 _095_ (.A(NN4END[8]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 _096_ (.A(NN4END[7]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 _097_ (.A(NN4END[6]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 _098_ (.A(NN4END[5]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 _099_ (.A(NN4END[4]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 _100_ (.A(NN4END[3]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 _101_ (.A(NN4END[2]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 _102_ (.A(NN4END[1]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 _103_ (.A(NN4END[0]),
    .X(net95));
 sky130_fd_sc_hd__buf_2 _104_ (.A(UserCLK),
    .X(net105));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_135 ();
 sky130_fd_sc_hd__buf_2 output1 (.A(net1),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output2 (.A(net2),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(S1BEG[0]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(S1BEG[1]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(S1BEG[2]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(S1BEG[3]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(S2BEG[0]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(S2BEG[1]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(S2BEG[2]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(S2BEG[3]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(S2BEG[4]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(S2BEG[5]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(S2BEG[6]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(S2BEG[7]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(S2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(S2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(S2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(S2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(S2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(S2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(S2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(S4BEG[0]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(S4BEG[10]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(S4BEG[11]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(S4BEG[12]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(S4BEG[13]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(S4BEG[14]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(S4BEG[15]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(S4BEG[1]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(S4BEG[2]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(S4BEG[3]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(S4BEG[4]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(S4BEG[5]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(S4BEG[6]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(S4BEG[7]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(S4BEG[8]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(S4BEG[9]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(SS4BEG[0]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(SS4BEG[10]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(SS4BEG[11]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(SS4BEG[12]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(SS4BEG[13]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(SS4BEG[14]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(SS4BEG[15]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(SS4BEG[1]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(SS4BEG[2]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(SS4BEG[3]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(SS4BEG[4]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(SS4BEG[5]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(SS4BEG[6]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(SS4BEG[7]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(SS4BEG[8]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(SS4BEG[9]));
 sky130_fd_sc_hd__buf_1 output105 (.A(net105),
    .X(UserCLKo));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(FrameData[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(FrameData[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(FrameData[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(FrameData[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(FrameData[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(FrameData[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(FrameData[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(FrameData[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(FrameData[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(FrameData[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(FrameData[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(FrameData[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(FrameData[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(FrameData[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(FrameData[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(FrameData[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(FrameData[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(FrameData[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(FrameData[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(FrameData[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(FrameData[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(FrameData[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(FrameData[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(FrameData[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(FrameData[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(FrameData[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(FrameData[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(FrameStrobe[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(FrameStrobe[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(FrameStrobe[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(NN4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(NN4END[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(NN4END[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(NN4END[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(NN4END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(NN4END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(NN4END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(NN4END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(NN4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(NN4END[9]));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_449 ();
endmodule
