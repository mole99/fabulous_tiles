magic
tech sky130A
magscale 1 2
timestamp 1740383373
<< viali >>
rect 1409 8585 1443 8619
rect 3249 8585 3283 8619
rect 5181 8585 5215 8619
rect 7113 8585 7147 8619
rect 9045 8585 9079 8619
rect 10977 8585 11011 8619
rect 12909 8585 12943 8619
rect 14841 8585 14875 8619
rect 16773 8585 16807 8619
rect 18705 8585 18739 8619
rect 20637 8585 20671 8619
rect 22569 8585 22603 8619
rect 24501 8585 24535 8619
rect 26525 8585 26559 8619
rect 28457 8585 28491 8619
rect 30389 8585 30423 8619
rect 32321 8585 32355 8619
rect 34253 8585 34287 8619
rect 36185 8585 36219 8619
rect 37013 8585 37047 8619
rect 37749 8585 37783 8619
rect 38117 8585 38151 8619
rect 38669 8585 38703 8619
rect 1593 8449 1627 8483
rect 3433 8449 3467 8483
rect 5365 8449 5399 8483
rect 7297 8449 7331 8483
rect 9229 8449 9263 8483
rect 11161 8449 11195 8483
rect 13093 8449 13127 8483
rect 15025 8449 15059 8483
rect 16957 8449 16991 8483
rect 18889 8449 18923 8483
rect 20821 8449 20855 8483
rect 22753 8449 22787 8483
rect 24685 8449 24719 8483
rect 26341 8449 26375 8483
rect 28273 8449 28307 8483
rect 30205 8449 30239 8483
rect 32137 8449 32171 8483
rect 34069 8449 34103 8483
rect 36001 8449 36035 8483
rect 36829 8449 36863 8483
rect 37565 8449 37599 8483
rect 37933 8449 37967 8483
rect 38485 8449 38519 8483
rect 38853 8449 38887 8483
rect 39221 8449 39255 8483
rect 39037 8313 39071 8347
rect 39405 8313 39439 8347
rect 38301 8041 38335 8075
rect 38669 8041 38703 8075
rect 37749 7837 37783 7871
rect 38117 7837 38151 7871
rect 38485 7837 38519 7871
rect 38853 7837 38887 7871
rect 39221 7837 39255 7871
rect 37933 7701 37967 7735
rect 39037 7701 39071 7735
rect 39405 7701 39439 7735
rect 16221 7497 16255 7531
rect 17417 7497 17451 7531
rect 17969 7497 18003 7531
rect 18153 7497 18187 7531
rect 18705 7497 18739 7531
rect 18889 7497 18923 7531
rect 19257 7497 19291 7531
rect 19349 7497 19383 7531
rect 20177 7497 20211 7531
rect 20453 7497 20487 7531
rect 20729 7497 20763 7531
rect 20821 7497 20855 7531
rect 21097 7497 21131 7531
rect 22109 7497 22143 7531
rect 22569 7497 22603 7531
rect 22937 7497 22971 7531
rect 39037 7497 39071 7531
rect 16129 7429 16163 7463
rect 16313 7429 16347 7463
rect 16405 7361 16439 7395
rect 16681 7361 16715 7395
rect 16957 7361 16991 7395
rect 17233 7361 17267 7395
rect 17785 7361 17819 7395
rect 18337 7361 18371 7395
rect 18981 7361 19015 7395
rect 19073 7361 19107 7395
rect 19533 7361 19567 7395
rect 19625 7361 19659 7395
rect 19993 7361 20027 7395
rect 20453 7361 20487 7395
rect 20545 7361 20579 7395
rect 21005 7361 21039 7395
rect 21281 7361 21315 7395
rect 22109 7361 22143 7395
rect 22201 7361 22235 7395
rect 22661 7361 22695 7395
rect 22753 7361 22787 7395
rect 23029 7361 23063 7395
rect 26157 7361 26191 7395
rect 27353 7361 27387 7395
rect 27721 7361 27755 7395
rect 27997 7361 28031 7395
rect 28273 7361 28307 7395
rect 28549 7361 28583 7395
rect 28825 7361 28859 7395
rect 38853 7361 38887 7395
rect 39221 7361 39255 7395
rect 17509 7293 17543 7327
rect 21465 7293 21499 7327
rect 16865 7225 16899 7259
rect 23213 7225 23247 7259
rect 17141 7157 17175 7191
rect 18429 7157 18463 7191
rect 18797 7157 18831 7191
rect 19809 7157 19843 7191
rect 21373 7157 21407 7191
rect 22385 7157 22419 7191
rect 25973 7157 26007 7191
rect 27169 7157 27203 7191
rect 27537 7157 27571 7191
rect 27813 7157 27847 7191
rect 28089 7157 28123 7191
rect 28365 7157 28399 7191
rect 28641 7157 28675 7191
rect 39405 7157 39439 7191
rect 10609 6885 10643 6919
rect 17877 6885 17911 6919
rect 17509 6817 17543 6851
rect 9045 6749 9079 6783
rect 9321 6749 9355 6783
rect 9597 6749 9631 6783
rect 9965 6749 9999 6783
rect 10425 6749 10459 6783
rect 10701 6749 10735 6783
rect 11069 6749 11103 6783
rect 11437 6749 11471 6783
rect 11713 6749 11747 6783
rect 17601 6749 17635 6783
rect 17693 6749 17727 6783
rect 22109 6749 22143 6783
rect 22385 6749 22419 6783
rect 38853 6749 38887 6783
rect 39221 6749 39255 6783
rect 9229 6613 9263 6647
rect 9505 6613 9539 6647
rect 9781 6613 9815 6647
rect 10149 6613 10183 6647
rect 10885 6613 10919 6647
rect 11253 6613 11287 6647
rect 11621 6613 11655 6647
rect 11897 6613 11931 6647
rect 21925 6613 21959 6647
rect 22201 6613 22235 6647
rect 39037 6613 39071 6647
rect 39405 6613 39439 6647
rect 27445 6409 27479 6443
rect 39405 6409 39439 6443
rect 8861 6273 8895 6307
rect 13645 6273 13679 6307
rect 13921 6273 13955 6307
rect 14197 6273 14231 6307
rect 27629 6273 27663 6307
rect 38853 6273 38887 6307
rect 39221 6273 39255 6307
rect 9045 6137 9079 6171
rect 13829 6137 13863 6171
rect 14105 6069 14139 6103
rect 14381 6069 14415 6103
rect 39037 6069 39071 6103
rect 9229 5865 9263 5899
rect 15117 5865 15151 5899
rect 19533 5865 19567 5899
rect 26341 5865 26375 5899
rect 7757 5797 7791 5831
rect 14473 5797 14507 5831
rect 19901 5797 19935 5831
rect 39405 5797 39439 5831
rect 7573 5661 7607 5695
rect 9045 5661 9079 5695
rect 13461 5661 13495 5695
rect 13737 5661 13771 5695
rect 14289 5661 14323 5695
rect 14565 5661 14599 5695
rect 14933 5661 14967 5695
rect 19625 5661 19659 5695
rect 19717 5661 19751 5695
rect 26157 5661 26191 5695
rect 38853 5661 38887 5695
rect 39221 5661 39255 5695
rect 13645 5525 13679 5559
rect 13921 5525 13955 5559
rect 14749 5525 14783 5559
rect 39037 5525 39071 5559
rect 3157 5321 3191 5355
rect 6193 5321 6227 5355
rect 16129 5321 16163 5355
rect 17969 5321 18003 5355
rect 36921 5321 36955 5355
rect 39405 5321 39439 5355
rect 2697 5185 2731 5219
rect 2973 5185 3007 5219
rect 3249 5185 3283 5219
rect 6009 5185 6043 5219
rect 15393 5185 15427 5219
rect 15669 5185 15703 5219
rect 15945 5185 15979 5219
rect 17601 5185 17635 5219
rect 17785 5185 17819 5219
rect 22385 5185 22419 5219
rect 37105 5185 37139 5219
rect 38853 5185 38887 5219
rect 39221 5185 39255 5219
rect 15853 5049 15887 5083
rect 2881 4981 2915 5015
rect 3433 4981 3467 5015
rect 15577 4981 15611 5015
rect 22569 4981 22603 5015
rect 39037 4981 39071 5015
rect 16773 4777 16807 4811
rect 23213 4777 23247 4811
rect 23489 4777 23523 4811
rect 27629 4777 27663 4811
rect 29377 4777 29411 4811
rect 31401 4777 31435 4811
rect 33333 4777 33367 4811
rect 4905 4709 4939 4743
rect 23857 4709 23891 4743
rect 27261 4709 27295 4743
rect 29837 4709 29871 4743
rect 39405 4709 39439 4743
rect 20085 4641 20119 4675
rect 22845 4641 22879 4675
rect 31585 4641 31619 4675
rect 2973 4573 3007 4607
rect 4261 4573 4295 4607
rect 4721 4573 4755 4607
rect 16589 4573 16623 4607
rect 20177 4573 20211 4607
rect 20269 4573 20303 4607
rect 22937 4573 22971 4607
rect 23029 4573 23063 4607
rect 23581 4573 23615 4607
rect 23673 4573 23707 4607
rect 24041 4573 24075 4607
rect 24409 4573 24443 4607
rect 25421 4573 25455 4607
rect 26525 4573 26559 4607
rect 27353 4573 27387 4607
rect 27445 4573 27479 4607
rect 28733 4573 28767 4607
rect 29101 4573 29135 4607
rect 29193 4573 29227 4607
rect 29653 4573 29687 4607
rect 29929 4573 29963 4607
rect 30205 4573 30239 4607
rect 30297 4573 30331 4607
rect 30849 4573 30883 4607
rect 31953 4573 31987 4607
rect 32229 4573 32263 4607
rect 32505 4573 32539 4607
rect 33149 4573 33183 4607
rect 35725 4573 35759 4607
rect 38853 4573 38887 4607
rect 39221 4573 39255 4607
rect 30113 4505 30147 4539
rect 3157 4437 3191 4471
rect 4445 4437 4479 4471
rect 20453 4437 20487 4471
rect 24225 4437 24259 4471
rect 25605 4437 25639 4471
rect 26709 4437 26743 4471
rect 28917 4437 28951 4471
rect 29009 4437 29043 4471
rect 30481 4437 30515 4471
rect 31033 4437 31067 4471
rect 31769 4437 31803 4471
rect 32045 4437 32079 4471
rect 32321 4437 32355 4471
rect 35909 4437 35943 4471
rect 39037 4437 39071 4471
rect 4721 4097 4755 4131
rect 17049 4097 17083 4131
rect 17509 4097 17543 4131
rect 19441 4097 19475 4131
rect 21557 4097 21591 4131
rect 21833 4097 21867 4131
rect 22201 4097 22235 4131
rect 22477 4097 22511 4131
rect 24317 4097 24351 4131
rect 24409 4097 24443 4131
rect 27261 4097 27295 4131
rect 27353 4097 27387 4131
rect 28181 4097 28215 4131
rect 29101 4097 29135 4131
rect 29377 4097 29411 4131
rect 29929 4097 29963 4131
rect 30205 4097 30239 4131
rect 30849 4097 30883 4131
rect 31033 4097 31067 4131
rect 31309 4097 31343 4131
rect 31585 4097 31619 4131
rect 38853 4097 38887 4131
rect 39221 4097 39255 4131
rect 17693 3961 17727 3995
rect 22017 3961 22051 3995
rect 22385 3961 22419 3995
rect 24593 3961 24627 3995
rect 30665 3961 30699 3995
rect 31401 3961 31435 3995
rect 39405 3961 39439 3995
rect 4905 3893 4939 3927
rect 17233 3893 17267 3927
rect 19625 3893 19659 3927
rect 24225 3893 24259 3927
rect 27169 3893 27203 3927
rect 27537 3893 27571 3927
rect 28365 3893 28399 3927
rect 29009 3893 29043 3927
rect 29193 3893 29227 3927
rect 29837 3893 29871 3927
rect 30021 3893 30055 3927
rect 31033 3893 31067 3927
rect 31125 3893 31159 3927
rect 39037 3893 39071 3927
rect 19533 3689 19567 3723
rect 22201 3689 22235 3723
rect 25421 3689 25455 3723
rect 25789 3689 25823 3723
rect 23673 3621 23707 3655
rect 24593 3621 24627 3655
rect 25145 3621 25179 3655
rect 39405 3621 39439 3655
rect 24225 3553 24259 3587
rect 18337 3485 18371 3519
rect 18429 3485 18463 3519
rect 18705 3485 18739 3519
rect 19257 3485 19291 3519
rect 21741 3485 21775 3519
rect 22293 3485 22327 3519
rect 22385 3485 22419 3519
rect 22753 3485 22787 3519
rect 22845 3485 22879 3519
rect 23121 3485 23155 3519
rect 23397 3485 23431 3519
rect 23857 3485 23891 3519
rect 24409 3485 24443 3519
rect 24685 3485 24719 3519
rect 24961 3485 24995 3519
rect 25237 3485 25271 3519
rect 25605 3485 25639 3519
rect 26525 3485 26559 3519
rect 38853 3485 38887 3519
rect 39221 3485 39255 3519
rect 18245 3349 18279 3383
rect 18613 3349 18647 3383
rect 18889 3349 18923 3383
rect 19441 3349 19475 3383
rect 21925 3349 21959 3383
rect 22569 3349 22603 3383
rect 22661 3349 22695 3383
rect 23029 3349 23063 3383
rect 23305 3349 23339 3383
rect 23581 3349 23615 3383
rect 24133 3349 24167 3383
rect 24869 3349 24903 3383
rect 26709 3349 26743 3383
rect 39037 3349 39071 3383
rect 23765 3145 23799 3179
rect 39405 3145 39439 3179
rect 18245 3009 18279 3043
rect 19073 3009 19107 3043
rect 19625 3009 19659 3043
rect 23213 3009 23247 3043
rect 23581 3009 23615 3043
rect 24593 3009 24627 3043
rect 25697 3009 25731 3043
rect 26065 3009 26099 3043
rect 26985 3009 27019 3043
rect 27905 3009 27939 3043
rect 28733 3009 28767 3043
rect 29285 3009 29319 3043
rect 30389 3009 30423 3043
rect 30941 3009 30975 3043
rect 31309 3009 31343 3043
rect 38485 3009 38519 3043
rect 38853 3009 38887 3043
rect 39221 3009 39255 3043
rect 38669 2873 38703 2907
rect 18429 2805 18463 2839
rect 19257 2805 19291 2839
rect 19809 2805 19843 2839
rect 23397 2805 23431 2839
rect 24777 2805 24811 2839
rect 25881 2805 25915 2839
rect 26249 2805 26283 2839
rect 27169 2805 27203 2839
rect 28089 2805 28123 2839
rect 28549 2805 28583 2839
rect 29101 2805 29135 2839
rect 30205 2805 30239 2839
rect 31125 2805 31159 2839
rect 31493 2805 31527 2839
rect 39037 2805 39071 2839
rect 23489 2601 23523 2635
rect 25329 2601 25363 2635
rect 28273 2601 28307 2635
rect 30757 2601 30791 2635
rect 22385 2533 22419 2567
rect 23121 2533 23155 2567
rect 24593 2533 24627 2567
rect 25697 2533 25731 2567
rect 27169 2533 27203 2567
rect 29009 2533 29043 2567
rect 30021 2533 30055 2567
rect 31125 2533 31159 2567
rect 32321 2533 32355 2567
rect 39405 2533 39439 2567
rect 17693 2397 17727 2431
rect 18061 2397 18095 2431
rect 18429 2397 18463 2431
rect 18797 2397 18831 2431
rect 19441 2397 19475 2431
rect 19809 2397 19843 2431
rect 20177 2397 20211 2431
rect 20545 2397 20579 2431
rect 20913 2397 20947 2431
rect 21281 2397 21315 2431
rect 21833 2397 21867 2431
rect 22201 2397 22235 2431
rect 22569 2397 22603 2431
rect 22937 2397 22971 2431
rect 23305 2397 23339 2431
rect 23673 2397 23707 2431
rect 24409 2397 24443 2431
rect 24777 2397 24811 2431
rect 25145 2397 25179 2431
rect 25513 2397 25547 2431
rect 25881 2397 25915 2431
rect 26249 2397 26283 2431
rect 26985 2397 27019 2431
rect 27359 2397 27393 2431
rect 27721 2397 27755 2431
rect 28089 2397 28123 2431
rect 28457 2397 28491 2431
rect 28825 2397 28859 2431
rect 29837 2397 29871 2431
rect 30205 2397 30239 2431
rect 30573 2397 30607 2431
rect 30941 2397 30975 2431
rect 31309 2397 31343 2431
rect 31401 2397 31435 2431
rect 32137 2397 32171 2431
rect 32505 2397 32539 2431
rect 32873 2397 32907 2431
rect 37749 2397 37783 2431
rect 38117 2397 38151 2431
rect 38485 2397 38519 2431
rect 39129 2397 39163 2431
rect 39221 2397 39255 2431
rect 17877 2261 17911 2295
rect 18245 2261 18279 2295
rect 18613 2261 18647 2295
rect 18981 2261 19015 2295
rect 19625 2261 19659 2295
rect 19993 2261 20027 2295
rect 20361 2261 20395 2295
rect 20729 2261 20763 2295
rect 21097 2261 21131 2295
rect 21465 2261 21499 2295
rect 22017 2261 22051 2295
rect 22753 2261 22787 2295
rect 23857 2261 23891 2295
rect 24961 2261 24995 2295
rect 26065 2261 26099 2295
rect 26433 2261 26467 2295
rect 27537 2261 27571 2295
rect 27905 2261 27939 2295
rect 28641 2261 28675 2295
rect 29653 2261 29687 2295
rect 30389 2261 30423 2295
rect 31585 2261 31619 2295
rect 32689 2261 32723 2295
rect 33057 2261 33091 2295
rect 37933 2261 37967 2295
rect 38301 2261 38335 2295
rect 38669 2261 38703 2295
rect 39037 2261 39071 2295
<< metal1 >>
rect 1302 9324 1308 9376
rect 1360 9364 1366 9376
rect 23014 9364 23020 9376
rect 1360 9336 23020 9364
rect 1360 9324 1366 9336
rect 23014 9324 23020 9336
rect 23072 9324 23078 9376
rect 20714 9256 20720 9308
rect 20772 9296 20778 9308
rect 20772 9268 39896 9296
rect 20772 9256 20778 9268
rect 20806 9228 20812 9240
rect 3436 9200 20812 9228
rect 3436 8832 3464 9200
rect 20806 9188 20812 9200
rect 20864 9188 20870 9240
rect 25774 9188 25780 9240
rect 25832 9228 25838 9240
rect 30190 9228 30196 9240
rect 25832 9200 30196 9228
rect 25832 9188 25838 9200
rect 30190 9188 30196 9200
rect 30248 9188 30254 9240
rect 18874 9120 18880 9172
rect 18932 9160 18938 9172
rect 27430 9160 27436 9172
rect 18932 9132 27436 9160
rect 18932 9120 18938 9132
rect 27430 9120 27436 9132
rect 27488 9120 27494 9172
rect 16850 9052 16856 9104
rect 16908 9092 16914 9104
rect 27798 9092 27804 9104
rect 16908 9064 27804 9092
rect 16908 9052 16914 9064
rect 27798 9052 27804 9064
rect 27856 9052 27862 9104
rect 13078 8984 13084 9036
rect 13136 9024 13142 9036
rect 27522 9024 27528 9036
rect 13136 8996 27528 9024
rect 13136 8984 13142 8996
rect 27522 8984 27528 8996
rect 27580 8984 27586 9036
rect 16942 8916 16948 8968
rect 17000 8956 17006 8968
rect 28074 8956 28080 8968
rect 17000 8928 28080 8956
rect 17000 8916 17006 8928
rect 28074 8916 28080 8928
rect 28132 8916 28138 8968
rect 36998 8916 37004 8968
rect 37056 8956 37062 8968
rect 39758 8956 39764 8968
rect 37056 8928 39764 8956
rect 37056 8916 37062 8928
rect 39758 8916 39764 8928
rect 39816 8916 39822 8968
rect 17954 8848 17960 8900
rect 18012 8888 18018 8900
rect 37550 8888 37556 8900
rect 18012 8860 37556 8888
rect 18012 8848 18018 8860
rect 37550 8848 37556 8860
rect 37608 8848 37614 8900
rect 3418 8780 3424 8832
rect 3476 8780 3482 8832
rect 5350 8780 5356 8832
rect 5408 8820 5414 8832
rect 18138 8820 18144 8832
rect 5408 8792 18144 8820
rect 5408 8780 5414 8792
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 20346 8780 20352 8832
rect 20404 8820 20410 8832
rect 33778 8820 33784 8832
rect 20404 8792 33784 8820
rect 20404 8780 20410 8792
rect 33778 8780 33784 8792
rect 33836 8780 33842 8832
rect 1104 8730 39836 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 39010 8730
rect 39062 8678 39074 8730
rect 39126 8678 39138 8730
rect 39190 8678 39202 8730
rect 39254 8678 39266 8730
rect 39318 8678 39836 8730
rect 1104 8656 39836 8678
rect 1118 8576 1124 8628
rect 1176 8616 1182 8628
rect 1397 8619 1455 8625
rect 1397 8616 1409 8619
rect 1176 8588 1409 8616
rect 1176 8576 1182 8588
rect 1397 8585 1409 8588
rect 1443 8585 1455 8619
rect 1397 8579 1455 8585
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 3237 8619 3295 8625
rect 3237 8616 3249 8619
rect 2924 8588 3249 8616
rect 2924 8576 2930 8588
rect 3237 8585 3249 8588
rect 3283 8585 3295 8619
rect 3237 8579 3295 8585
rect 3418 8576 3424 8628
rect 3476 8576 3482 8628
rect 4982 8576 4988 8628
rect 5040 8616 5046 8628
rect 5169 8619 5227 8625
rect 5169 8616 5181 8619
rect 5040 8588 5181 8616
rect 5040 8576 5046 8588
rect 5169 8585 5181 8588
rect 5215 8585 5227 8619
rect 5169 8579 5227 8585
rect 6914 8576 6920 8628
rect 6972 8616 6978 8628
rect 7101 8619 7159 8625
rect 7101 8616 7113 8619
rect 6972 8588 7113 8616
rect 6972 8576 6978 8588
rect 7101 8585 7113 8588
rect 7147 8585 7159 8619
rect 7101 8579 7159 8585
rect 8846 8576 8852 8628
rect 8904 8616 8910 8628
rect 9033 8619 9091 8625
rect 9033 8616 9045 8619
rect 8904 8588 9045 8616
rect 8904 8576 8910 8588
rect 9033 8585 9045 8588
rect 9079 8585 9091 8619
rect 9033 8579 9091 8585
rect 10778 8576 10784 8628
rect 10836 8616 10842 8628
rect 10965 8619 11023 8625
rect 10965 8616 10977 8619
rect 10836 8588 10977 8616
rect 10836 8576 10842 8588
rect 10965 8585 10977 8588
rect 11011 8585 11023 8619
rect 10965 8579 11023 8585
rect 12710 8576 12716 8628
rect 12768 8616 12774 8628
rect 12897 8619 12955 8625
rect 12897 8616 12909 8619
rect 12768 8588 12909 8616
rect 12768 8576 12774 8588
rect 12897 8585 12909 8588
rect 12943 8585 12955 8619
rect 12897 8579 12955 8585
rect 14642 8576 14648 8628
rect 14700 8616 14706 8628
rect 14829 8619 14887 8625
rect 14829 8616 14841 8619
rect 14700 8588 14841 8616
rect 14700 8576 14706 8588
rect 14829 8585 14841 8588
rect 14875 8585 14887 8619
rect 14829 8579 14887 8585
rect 16574 8576 16580 8628
rect 16632 8616 16638 8628
rect 16761 8619 16819 8625
rect 16761 8616 16773 8619
rect 16632 8588 16773 8616
rect 16632 8576 16638 8588
rect 16761 8585 16773 8588
rect 16807 8585 16819 8619
rect 16761 8579 16819 8585
rect 18506 8576 18512 8628
rect 18564 8616 18570 8628
rect 18693 8619 18751 8625
rect 18693 8616 18705 8619
rect 18564 8588 18705 8616
rect 18564 8576 18570 8588
rect 18693 8585 18705 8588
rect 18739 8585 18751 8619
rect 18693 8579 18751 8585
rect 20438 8576 20444 8628
rect 20496 8616 20502 8628
rect 20625 8619 20683 8625
rect 20625 8616 20637 8619
rect 20496 8588 20637 8616
rect 20496 8576 20502 8588
rect 20625 8585 20637 8588
rect 20671 8585 20683 8619
rect 20625 8579 20683 8585
rect 22370 8576 22376 8628
rect 22428 8616 22434 8628
rect 22557 8619 22615 8625
rect 22557 8616 22569 8619
rect 22428 8588 22569 8616
rect 22428 8576 22434 8588
rect 22557 8585 22569 8588
rect 22603 8585 22615 8619
rect 22557 8579 22615 8585
rect 24302 8576 24308 8628
rect 24360 8616 24366 8628
rect 24489 8619 24547 8625
rect 24489 8616 24501 8619
rect 24360 8588 24501 8616
rect 24360 8576 24366 8588
rect 24489 8585 24501 8588
rect 24535 8585 24547 8619
rect 24489 8579 24547 8585
rect 26234 8576 26240 8628
rect 26292 8616 26298 8628
rect 26513 8619 26571 8625
rect 26513 8616 26525 8619
rect 26292 8588 26525 8616
rect 26292 8576 26298 8588
rect 26513 8585 26525 8588
rect 26559 8585 26571 8619
rect 26513 8579 26571 8585
rect 28166 8576 28172 8628
rect 28224 8616 28230 8628
rect 28445 8619 28503 8625
rect 28445 8616 28457 8619
rect 28224 8588 28457 8616
rect 28224 8576 28230 8588
rect 28445 8585 28457 8588
rect 28491 8585 28503 8619
rect 28445 8579 28503 8585
rect 30098 8576 30104 8628
rect 30156 8616 30162 8628
rect 30377 8619 30435 8625
rect 30377 8616 30389 8619
rect 30156 8588 30389 8616
rect 30156 8576 30162 8588
rect 30377 8585 30389 8588
rect 30423 8585 30435 8619
rect 30377 8579 30435 8585
rect 32030 8576 32036 8628
rect 32088 8616 32094 8628
rect 32309 8619 32367 8625
rect 32309 8616 32321 8619
rect 32088 8588 32321 8616
rect 32088 8576 32094 8588
rect 32309 8585 32321 8588
rect 32355 8585 32367 8619
rect 32309 8579 32367 8585
rect 33962 8576 33968 8628
rect 34020 8616 34026 8628
rect 34241 8619 34299 8625
rect 34241 8616 34253 8619
rect 34020 8588 34253 8616
rect 34020 8576 34026 8588
rect 34241 8585 34253 8588
rect 34287 8585 34299 8619
rect 34241 8579 34299 8585
rect 35894 8576 35900 8628
rect 35952 8616 35958 8628
rect 36173 8619 36231 8625
rect 36173 8616 36185 8619
rect 35952 8588 36185 8616
rect 35952 8576 35958 8588
rect 36173 8585 36185 8588
rect 36219 8585 36231 8619
rect 36173 8579 36231 8585
rect 36998 8576 37004 8628
rect 37056 8576 37062 8628
rect 37734 8576 37740 8628
rect 37792 8576 37798 8628
rect 37826 8576 37832 8628
rect 37884 8616 37890 8628
rect 38105 8619 38163 8625
rect 38105 8616 38117 8619
rect 37884 8588 38117 8616
rect 37884 8576 37890 8588
rect 38105 8585 38117 8588
rect 38151 8585 38163 8619
rect 38105 8579 38163 8585
rect 38654 8576 38660 8628
rect 38712 8576 38718 8628
rect 1578 8440 1584 8492
rect 1636 8440 1642 8492
rect 3436 8489 3464 8576
rect 25866 8548 25872 8560
rect 12406 8520 25872 8548
rect 3421 8483 3479 8489
rect 3421 8449 3433 8483
rect 3467 8449 3479 8483
rect 3421 8443 3479 8449
rect 5350 8440 5356 8492
rect 5408 8440 5414 8492
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 11149 8483 11207 8489
rect 11149 8449 11161 8483
rect 11195 8480 11207 8483
rect 12406 8480 12434 8520
rect 25866 8508 25872 8520
rect 25924 8508 25930 8560
rect 25976 8520 28994 8548
rect 11195 8452 12434 8480
rect 11195 8449 11207 8452
rect 11149 8443 11207 8449
rect 7300 8344 7328 8443
rect 9232 8412 9260 8443
rect 13078 8440 13084 8492
rect 13136 8440 13142 8492
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8480 15071 8483
rect 16850 8480 16856 8492
rect 15059 8452 16856 8480
rect 15059 8449 15071 8452
rect 15013 8443 15071 8449
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 16942 8440 16948 8492
rect 17000 8440 17006 8492
rect 18874 8440 18880 8492
rect 18932 8440 18938 8492
rect 20809 8483 20867 8489
rect 20809 8449 20821 8483
rect 20855 8480 20867 8483
rect 20855 8452 22094 8480
rect 20855 8449 20867 8452
rect 20809 8443 20867 8449
rect 16574 8412 16580 8424
rect 9232 8384 16580 8412
rect 16574 8372 16580 8384
rect 16632 8372 16638 8424
rect 22066 8412 22094 8452
rect 22738 8440 22744 8492
rect 22796 8440 22802 8492
rect 24670 8440 24676 8492
rect 24728 8440 24734 8492
rect 24762 8440 24768 8492
rect 24820 8480 24826 8492
rect 25976 8480 26004 8520
rect 24820 8452 26004 8480
rect 24820 8440 24826 8452
rect 26326 8440 26332 8492
rect 26384 8440 26390 8492
rect 28261 8483 28319 8489
rect 28261 8449 28273 8483
rect 28307 8449 28319 8483
rect 28966 8480 28994 8520
rect 29564 8520 34192 8548
rect 29564 8480 29592 8520
rect 28966 8452 29592 8480
rect 28261 8443 28319 8449
rect 25406 8412 25412 8424
rect 22066 8384 25412 8412
rect 25406 8372 25412 8384
rect 25464 8372 25470 8424
rect 25590 8372 25596 8424
rect 25648 8412 25654 8424
rect 28276 8412 28304 8443
rect 30190 8440 30196 8492
rect 30248 8440 30254 8492
rect 32125 8483 32183 8489
rect 32125 8449 32137 8483
rect 32171 8480 32183 8483
rect 32582 8480 32588 8492
rect 32171 8452 32588 8480
rect 32171 8449 32183 8452
rect 32125 8443 32183 8449
rect 32582 8440 32588 8452
rect 32640 8440 32646 8492
rect 34057 8483 34115 8489
rect 34057 8449 34069 8483
rect 34103 8449 34115 8483
rect 34057 8443 34115 8449
rect 25648 8384 28304 8412
rect 25648 8372 25654 8384
rect 31018 8372 31024 8424
rect 31076 8412 31082 8424
rect 34072 8412 34100 8443
rect 31076 8384 34100 8412
rect 34164 8412 34192 8520
rect 35986 8440 35992 8492
rect 36044 8440 36050 8492
rect 36814 8440 36820 8492
rect 36872 8440 36878 8492
rect 37550 8440 37556 8492
rect 37608 8440 37614 8492
rect 37642 8440 37648 8492
rect 37700 8480 37706 8492
rect 37921 8483 37979 8489
rect 37921 8480 37933 8483
rect 37700 8452 37933 8480
rect 37700 8440 37706 8452
rect 37921 8449 37933 8452
rect 37967 8449 37979 8483
rect 37921 8443 37979 8449
rect 38473 8483 38531 8489
rect 38473 8449 38485 8483
rect 38519 8449 38531 8483
rect 38473 8443 38531 8449
rect 38841 8483 38899 8489
rect 38841 8449 38853 8483
rect 38887 8449 38899 8483
rect 38841 8443 38899 8449
rect 39209 8483 39267 8489
rect 39209 8449 39221 8483
rect 39255 8480 39267 8483
rect 39868 8480 39896 9268
rect 39255 8452 39896 8480
rect 39255 8449 39267 8452
rect 39209 8443 39267 8449
rect 38488 8412 38516 8443
rect 34164 8384 38516 8412
rect 31076 8372 31082 8384
rect 22186 8344 22192 8356
rect 7300 8316 22192 8344
rect 22186 8304 22192 8316
rect 22244 8304 22250 8356
rect 22738 8304 22744 8356
rect 22796 8344 22802 8356
rect 26878 8344 26884 8356
rect 22796 8316 26884 8344
rect 22796 8304 22802 8316
rect 26878 8304 26884 8316
rect 26936 8304 26942 8356
rect 33778 8304 33784 8356
rect 33836 8344 33842 8356
rect 38856 8344 38884 8443
rect 33836 8316 38884 8344
rect 33836 8304 33842 8316
rect 39022 8304 39028 8356
rect 39080 8304 39086 8356
rect 39390 8304 39396 8356
rect 39448 8304 39454 8356
rect 1104 8186 39836 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 37950 8186
rect 38002 8134 38014 8186
rect 38066 8134 38078 8186
rect 38130 8134 38142 8186
rect 38194 8134 38206 8186
rect 38258 8134 39836 8186
rect 1104 8112 39836 8134
rect 16482 8032 16488 8084
rect 16540 8072 16546 8084
rect 18874 8072 18880 8084
rect 16540 8044 18880 8072
rect 16540 8032 16546 8044
rect 18874 8032 18880 8044
rect 18932 8032 18938 8084
rect 19242 8032 19248 8084
rect 19300 8072 19306 8084
rect 19300 8044 22968 8072
rect 19300 8032 19306 8044
rect 17126 7964 17132 8016
rect 17184 8004 17190 8016
rect 17184 7976 22876 8004
rect 17184 7964 17190 7976
rect 16114 7896 16120 7948
rect 16172 7936 16178 7948
rect 18322 7936 18328 7948
rect 16172 7908 18328 7936
rect 16172 7896 16178 7908
rect 18322 7896 18328 7908
rect 18380 7936 18386 7948
rect 22462 7936 22468 7948
rect 18380 7908 22468 7936
rect 18380 7896 18386 7908
rect 22462 7896 22468 7908
rect 22520 7896 22526 7948
rect 16390 7828 16396 7880
rect 16448 7868 16454 7880
rect 19978 7868 19984 7880
rect 16448 7840 19984 7868
rect 16448 7828 16454 7840
rect 19978 7828 19984 7840
rect 20036 7868 20042 7880
rect 20898 7868 20904 7880
rect 20036 7840 20904 7868
rect 20036 7828 20042 7840
rect 20898 7828 20904 7840
rect 20956 7828 20962 7880
rect 22848 7868 22876 7976
rect 22940 7936 22968 8044
rect 38286 8032 38292 8084
rect 38344 8032 38350 8084
rect 38657 8075 38715 8081
rect 38657 8041 38669 8075
rect 38703 8072 38715 8075
rect 39482 8072 39488 8084
rect 38703 8044 39488 8072
rect 38703 8041 38715 8044
rect 38657 8035 38715 8041
rect 39482 8032 39488 8044
rect 39540 8032 39546 8084
rect 23198 7964 23204 8016
rect 23256 8004 23262 8016
rect 23256 7976 38884 8004
rect 23256 7964 23262 7976
rect 22940 7908 38516 7936
rect 22848 7840 31754 7868
rect 16574 7760 16580 7812
rect 16632 7800 16638 7812
rect 19334 7800 19340 7812
rect 16632 7772 19340 7800
rect 16632 7760 16638 7772
rect 19334 7760 19340 7772
rect 19392 7760 19398 7812
rect 31726 7800 31754 7840
rect 37734 7828 37740 7880
rect 37792 7828 37798 7880
rect 38102 7828 38108 7880
rect 38160 7828 38166 7880
rect 38488 7877 38516 7908
rect 38856 7877 38884 7976
rect 38473 7871 38531 7877
rect 38473 7837 38485 7871
rect 38519 7837 38531 7871
rect 38473 7831 38531 7837
rect 38841 7871 38899 7877
rect 38841 7837 38853 7871
rect 38887 7837 38899 7871
rect 38841 7831 38899 7837
rect 39209 7871 39267 7877
rect 39209 7837 39221 7871
rect 39255 7837 39267 7871
rect 39209 7831 39267 7837
rect 37826 7800 37832 7812
rect 31726 7772 37832 7800
rect 37826 7760 37832 7772
rect 37884 7760 37890 7812
rect 38010 7760 38016 7812
rect 38068 7800 38074 7812
rect 39224 7800 39252 7831
rect 38068 7772 39252 7800
rect 38068 7760 38074 7772
rect 14826 7692 14832 7744
rect 14884 7732 14890 7744
rect 17770 7732 17776 7744
rect 14884 7704 17776 7732
rect 14884 7692 14890 7704
rect 17770 7692 17776 7704
rect 17828 7692 17834 7744
rect 19058 7692 19064 7744
rect 19116 7732 19122 7744
rect 20438 7732 20444 7744
rect 19116 7704 20444 7732
rect 19116 7692 19122 7704
rect 20438 7692 20444 7704
rect 20496 7692 20502 7744
rect 25406 7692 25412 7744
rect 25464 7732 25470 7744
rect 26142 7732 26148 7744
rect 25464 7704 26148 7732
rect 25464 7692 25470 7704
rect 26142 7692 26148 7704
rect 26200 7692 26206 7744
rect 27430 7692 27436 7744
rect 27488 7732 27494 7744
rect 28350 7732 28356 7744
rect 27488 7704 28356 7732
rect 27488 7692 27494 7704
rect 28350 7692 28356 7704
rect 28408 7692 28414 7744
rect 37921 7735 37979 7741
rect 37921 7701 37933 7735
rect 37967 7732 37979 7735
rect 38378 7732 38384 7744
rect 37967 7704 38384 7732
rect 37967 7701 37979 7704
rect 37921 7695 37979 7701
rect 38378 7692 38384 7704
rect 38436 7692 38442 7744
rect 38930 7692 38936 7744
rect 38988 7732 38994 7744
rect 39025 7735 39083 7741
rect 39025 7732 39037 7735
rect 38988 7704 39037 7732
rect 38988 7692 38994 7704
rect 39025 7701 39037 7704
rect 39071 7701 39083 7735
rect 39025 7695 39083 7701
rect 39390 7692 39396 7744
rect 39448 7692 39454 7744
rect 1104 7642 39836 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 39010 7642
rect 39062 7590 39074 7642
rect 39126 7590 39138 7642
rect 39190 7590 39202 7642
rect 39254 7590 39266 7642
rect 39318 7590 39836 7642
rect 1104 7568 39836 7590
rect 14918 7488 14924 7540
rect 14976 7528 14982 7540
rect 16209 7531 16267 7537
rect 16209 7528 16221 7531
rect 14976 7500 16221 7528
rect 14976 7488 14982 7500
rect 16209 7497 16221 7500
rect 16255 7497 16267 7531
rect 16209 7491 16267 7497
rect 17405 7531 17463 7537
rect 17405 7497 17417 7531
rect 17451 7528 17463 7531
rect 17451 7500 17908 7528
rect 17451 7497 17463 7500
rect 17405 7491 17463 7497
rect 16114 7420 16120 7472
rect 16172 7420 16178 7472
rect 16301 7463 16359 7469
rect 16301 7429 16313 7463
rect 16347 7460 16359 7463
rect 16347 7432 17264 7460
rect 16347 7429 16359 7432
rect 16301 7423 16359 7429
rect 15102 7352 15108 7404
rect 15160 7392 15166 7404
rect 17236 7401 17264 7432
rect 16393 7395 16451 7401
rect 16393 7392 16405 7395
rect 15160 7364 16405 7392
rect 15160 7352 15166 7364
rect 16393 7361 16405 7364
rect 16439 7392 16451 7395
rect 16669 7395 16727 7401
rect 16669 7392 16681 7395
rect 16439 7364 16681 7392
rect 16439 7361 16451 7364
rect 16393 7355 16451 7361
rect 16669 7361 16681 7364
rect 16715 7361 16727 7395
rect 16669 7355 16727 7361
rect 16945 7395 17003 7401
rect 16945 7361 16957 7395
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 17221 7395 17279 7401
rect 17221 7361 17233 7395
rect 17267 7361 17279 7395
rect 17221 7355 17279 7361
rect 16482 7284 16488 7336
rect 16540 7324 16546 7336
rect 16960 7324 16988 7355
rect 17770 7352 17776 7404
rect 17828 7352 17834 7404
rect 17880 7392 17908 7500
rect 17954 7488 17960 7540
rect 18012 7488 18018 7540
rect 18138 7488 18144 7540
rect 18196 7488 18202 7540
rect 18690 7488 18696 7540
rect 18748 7488 18754 7540
rect 18874 7488 18880 7540
rect 18932 7488 18938 7540
rect 19242 7488 19248 7540
rect 19300 7488 19306 7540
rect 19334 7488 19340 7540
rect 19392 7488 19398 7540
rect 20165 7531 20223 7537
rect 20165 7497 20177 7531
rect 20211 7528 20223 7531
rect 20346 7528 20352 7540
rect 20211 7500 20352 7528
rect 20211 7497 20223 7500
rect 20165 7491 20223 7497
rect 20346 7488 20352 7500
rect 20404 7488 20410 7540
rect 20438 7488 20444 7540
rect 20496 7488 20502 7540
rect 20714 7488 20720 7540
rect 20772 7488 20778 7540
rect 20806 7488 20812 7540
rect 20864 7488 20870 7540
rect 20898 7488 20904 7540
rect 20956 7528 20962 7540
rect 21085 7531 21143 7537
rect 21085 7528 21097 7531
rect 20956 7500 21097 7528
rect 20956 7488 20962 7500
rect 21085 7497 21097 7500
rect 21131 7497 21143 7531
rect 21085 7491 21143 7497
rect 22094 7488 22100 7540
rect 22152 7488 22158 7540
rect 22554 7488 22560 7540
rect 22612 7488 22618 7540
rect 22925 7531 22983 7537
rect 22925 7497 22937 7531
rect 22971 7528 22983 7531
rect 39025 7531 39083 7537
rect 22971 7500 31754 7528
rect 22971 7497 22983 7500
rect 22925 7491 22983 7497
rect 18248 7432 26556 7460
rect 18248 7392 18276 7432
rect 17880 7364 18276 7392
rect 18322 7352 18328 7404
rect 18380 7352 18386 7404
rect 18969 7395 19027 7401
rect 18969 7361 18981 7395
rect 19015 7392 19027 7395
rect 19061 7395 19119 7401
rect 19061 7392 19073 7395
rect 19015 7364 19073 7392
rect 19015 7361 19027 7364
rect 18969 7355 19027 7361
rect 19061 7361 19073 7364
rect 19107 7361 19119 7395
rect 19061 7355 19119 7361
rect 19521 7395 19579 7401
rect 19521 7361 19533 7395
rect 19567 7361 19579 7395
rect 19521 7355 19579 7361
rect 17497 7327 17555 7333
rect 17497 7324 17509 7327
rect 16540 7296 17509 7324
rect 16540 7284 16546 7296
rect 17497 7293 17509 7296
rect 17543 7293 17555 7327
rect 19536 7324 19564 7355
rect 19610 7352 19616 7404
rect 19668 7352 19674 7404
rect 19978 7352 19984 7404
rect 20036 7352 20042 7404
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7392 20499 7395
rect 20533 7395 20591 7401
rect 20533 7392 20545 7395
rect 20487 7364 20545 7392
rect 20487 7361 20499 7364
rect 20441 7355 20499 7361
rect 20533 7361 20545 7364
rect 20579 7361 20591 7395
rect 20533 7355 20591 7361
rect 20993 7395 21051 7401
rect 20993 7361 21005 7395
rect 21039 7392 21051 7395
rect 21269 7395 21327 7401
rect 21269 7392 21281 7395
rect 21039 7364 21281 7392
rect 21039 7361 21051 7364
rect 20993 7355 21051 7361
rect 21269 7361 21281 7364
rect 21315 7361 21327 7395
rect 21269 7355 21327 7361
rect 22097 7395 22155 7401
rect 22097 7361 22109 7395
rect 22143 7392 22155 7395
rect 22189 7395 22247 7401
rect 22189 7392 22201 7395
rect 22143 7364 22201 7392
rect 22143 7361 22155 7364
rect 22097 7355 22155 7361
rect 22189 7361 22201 7364
rect 22235 7361 22247 7395
rect 22189 7355 22247 7361
rect 22649 7395 22707 7401
rect 22649 7361 22661 7395
rect 22695 7392 22707 7395
rect 22741 7395 22799 7401
rect 22741 7392 22753 7395
rect 22695 7364 22753 7392
rect 22695 7361 22707 7364
rect 22649 7355 22707 7361
rect 22741 7361 22753 7364
rect 22787 7361 22799 7395
rect 22741 7355 22799 7361
rect 23014 7352 23020 7404
rect 23072 7352 23078 7404
rect 23198 7352 23204 7404
rect 23256 7352 23262 7404
rect 25222 7352 25228 7404
rect 25280 7392 25286 7404
rect 26145 7395 26203 7401
rect 26145 7392 26157 7395
rect 25280 7364 26157 7392
rect 25280 7352 25286 7364
rect 26145 7361 26157 7364
rect 26191 7361 26203 7395
rect 26145 7355 26203 7361
rect 21453 7327 21511 7333
rect 21453 7324 21465 7327
rect 17497 7287 17555 7293
rect 17880 7296 19334 7324
rect 19536 7296 21465 7324
rect 16853 7259 16911 7265
rect 16853 7225 16865 7259
rect 16899 7256 16911 7259
rect 17880 7256 17908 7296
rect 16899 7228 17908 7256
rect 19306 7256 19334 7296
rect 21453 7293 21465 7296
rect 21499 7324 21511 7327
rect 22922 7324 22928 7336
rect 21499 7296 22928 7324
rect 21499 7293 21511 7296
rect 21453 7287 21511 7293
rect 22922 7284 22928 7296
rect 22980 7284 22986 7336
rect 23106 7256 23112 7268
rect 19306 7228 23112 7256
rect 16899 7225 16911 7228
rect 16853 7219 16911 7225
rect 23106 7216 23112 7228
rect 23164 7216 23170 7268
rect 23216 7265 23244 7352
rect 26528 7324 26556 7432
rect 26878 7420 26884 7472
rect 26936 7460 26942 7472
rect 28442 7460 28448 7472
rect 26936 7432 28448 7460
rect 26936 7420 26942 7432
rect 28442 7420 28448 7432
rect 28500 7420 28506 7472
rect 31726 7460 31754 7500
rect 39025 7497 39037 7531
rect 39071 7528 39083 7531
rect 39574 7528 39580 7540
rect 39071 7500 39580 7528
rect 39071 7497 39083 7500
rect 39025 7491 39083 7497
rect 39574 7488 39580 7500
rect 39632 7488 39638 7540
rect 37734 7460 37740 7472
rect 28552 7432 30144 7460
rect 31726 7432 37740 7460
rect 27338 7352 27344 7404
rect 27396 7352 27402 7404
rect 27706 7352 27712 7404
rect 27764 7352 27770 7404
rect 27982 7352 27988 7404
rect 28040 7352 28046 7404
rect 28258 7352 28264 7404
rect 28316 7352 28322 7404
rect 28552 7401 28580 7432
rect 28537 7395 28595 7401
rect 28537 7361 28549 7395
rect 28583 7361 28595 7395
rect 28537 7355 28595 7361
rect 28810 7352 28816 7404
rect 28868 7352 28874 7404
rect 30116 7392 30144 7432
rect 37734 7420 37740 7432
rect 37792 7420 37798 7472
rect 37826 7420 37832 7472
rect 37884 7460 37890 7472
rect 37884 7432 39252 7460
rect 37884 7420 37890 7432
rect 34698 7392 34704 7404
rect 30116 7364 34704 7392
rect 34698 7352 34704 7364
rect 34756 7352 34762 7404
rect 38838 7352 38844 7404
rect 38896 7352 38902 7404
rect 39224 7401 39252 7432
rect 39209 7395 39267 7401
rect 39209 7361 39221 7395
rect 39255 7361 39267 7395
rect 39209 7355 39267 7361
rect 38102 7324 38108 7336
rect 26528 7296 38108 7324
rect 38102 7284 38108 7296
rect 38160 7284 38166 7336
rect 23201 7259 23259 7265
rect 23201 7225 23213 7259
rect 23247 7225 23259 7259
rect 23201 7219 23259 7225
rect 23290 7216 23296 7268
rect 23348 7256 23354 7268
rect 38010 7256 38016 7268
rect 23348 7228 38016 7256
rect 23348 7216 23354 7228
rect 38010 7216 38016 7228
rect 38068 7216 38074 7268
rect 17126 7148 17132 7200
rect 17184 7148 17190 7200
rect 17770 7148 17776 7200
rect 17828 7188 17834 7200
rect 18417 7191 18475 7197
rect 18417 7188 18429 7191
rect 17828 7160 18429 7188
rect 17828 7148 17834 7160
rect 18417 7157 18429 7160
rect 18463 7157 18475 7191
rect 18417 7151 18475 7157
rect 18785 7191 18843 7197
rect 18785 7157 18797 7191
rect 18831 7188 18843 7191
rect 19610 7188 19616 7200
rect 18831 7160 19616 7188
rect 18831 7157 18843 7160
rect 18785 7151 18843 7157
rect 19610 7148 19616 7160
rect 19668 7148 19674 7200
rect 19794 7148 19800 7200
rect 19852 7148 19858 7200
rect 21358 7148 21364 7200
rect 21416 7148 21422 7200
rect 22373 7191 22431 7197
rect 22373 7157 22385 7191
rect 22419 7188 22431 7191
rect 24762 7188 24768 7200
rect 22419 7160 24768 7188
rect 22419 7157 22431 7160
rect 22373 7151 22431 7157
rect 24762 7148 24768 7160
rect 24820 7148 24826 7200
rect 25866 7148 25872 7200
rect 25924 7188 25930 7200
rect 25961 7191 26019 7197
rect 25961 7188 25973 7191
rect 25924 7160 25973 7188
rect 25924 7148 25930 7160
rect 25961 7157 25973 7160
rect 26007 7157 26019 7191
rect 25961 7151 26019 7157
rect 26142 7148 26148 7200
rect 26200 7188 26206 7200
rect 27157 7191 27215 7197
rect 27157 7188 27169 7191
rect 26200 7160 27169 7188
rect 26200 7148 26206 7160
rect 27157 7157 27169 7160
rect 27203 7157 27215 7191
rect 27157 7151 27215 7157
rect 27522 7148 27528 7200
rect 27580 7148 27586 7200
rect 27798 7148 27804 7200
rect 27856 7148 27862 7200
rect 28074 7148 28080 7200
rect 28132 7148 28138 7200
rect 28350 7148 28356 7200
rect 28408 7148 28414 7200
rect 28442 7148 28448 7200
rect 28500 7188 28506 7200
rect 28629 7191 28687 7197
rect 28629 7188 28641 7191
rect 28500 7160 28641 7188
rect 28500 7148 28506 7160
rect 28629 7157 28641 7160
rect 28675 7157 28687 7191
rect 28629 7151 28687 7157
rect 39390 7148 39396 7200
rect 39448 7148 39454 7200
rect 1104 7098 39836 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 37950 7098
rect 38002 7046 38014 7098
rect 38066 7046 38078 7098
rect 38130 7046 38142 7098
rect 38194 7046 38206 7098
rect 38258 7046 39836 7098
rect 1104 7024 39836 7046
rect 19794 6944 19800 6996
rect 19852 6984 19858 6996
rect 38838 6984 38844 6996
rect 19852 6956 38844 6984
rect 19852 6944 19858 6956
rect 38838 6944 38844 6956
rect 38896 6944 38902 6996
rect 9122 6876 9128 6928
rect 9180 6916 9186 6928
rect 10597 6919 10655 6925
rect 9180 6888 9444 6916
rect 9180 6876 9186 6888
rect 7742 6808 7748 6860
rect 7800 6848 7806 6860
rect 9416 6848 9444 6888
rect 10597 6885 10609 6919
rect 10643 6916 10655 6919
rect 10643 6888 11560 6916
rect 10643 6885 10655 6888
rect 10597 6879 10655 6885
rect 7800 6820 9352 6848
rect 9416 6820 10456 6848
rect 7800 6808 7806 6820
rect 7834 6740 7840 6792
rect 7892 6780 7898 6792
rect 9324 6789 9352 6820
rect 9033 6783 9091 6789
rect 9033 6780 9045 6783
rect 7892 6752 9045 6780
rect 7892 6740 7898 6752
rect 9033 6749 9045 6752
rect 9079 6749 9091 6783
rect 9033 6743 9091 6749
rect 9309 6783 9367 6789
rect 9309 6749 9321 6783
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 9582 6740 9588 6792
rect 9640 6740 9646 6792
rect 9950 6740 9956 6792
rect 10008 6740 10014 6792
rect 10428 6789 10456 6820
rect 10778 6808 10784 6860
rect 10836 6848 10842 6860
rect 11532 6848 11560 6888
rect 17420 6888 17632 6916
rect 17420 6848 17448 6888
rect 10836 6820 11468 6848
rect 11532 6820 17448 6848
rect 10836 6808 10842 6820
rect 10413 6783 10471 6789
rect 10413 6749 10425 6783
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 10502 6740 10508 6792
rect 10560 6780 10566 6792
rect 10689 6783 10747 6789
rect 10689 6780 10701 6783
rect 10560 6752 10701 6780
rect 10560 6740 10566 6752
rect 10689 6749 10701 6752
rect 10735 6749 10747 6783
rect 10689 6743 10747 6749
rect 10870 6740 10876 6792
rect 10928 6780 10934 6792
rect 11440 6789 11468 6820
rect 17494 6808 17500 6860
rect 17552 6808 17558 6860
rect 17604 6848 17632 6888
rect 17862 6876 17868 6928
rect 17920 6876 17926 6928
rect 21358 6876 21364 6928
rect 21416 6916 21422 6928
rect 26878 6916 26884 6928
rect 21416 6888 26884 6916
rect 21416 6876 21422 6888
rect 26878 6876 26884 6888
rect 26936 6876 26942 6928
rect 27706 6876 27712 6928
rect 27764 6916 27770 6928
rect 33870 6916 33876 6928
rect 27764 6888 33876 6916
rect 27764 6876 27770 6888
rect 33870 6876 33876 6888
rect 33928 6876 33934 6928
rect 18414 6848 18420 6860
rect 17604 6820 18420 6848
rect 18414 6808 18420 6820
rect 18472 6808 18478 6860
rect 32306 6848 32312 6860
rect 22112 6820 32312 6848
rect 11057 6783 11115 6789
rect 11057 6780 11069 6783
rect 10928 6752 11069 6780
rect 10928 6740 10934 6752
rect 11057 6749 11069 6752
rect 11103 6749 11115 6783
rect 11057 6743 11115 6749
rect 11425 6783 11483 6789
rect 11425 6749 11437 6783
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 11698 6740 11704 6792
rect 11756 6740 11762 6792
rect 22112 6789 22140 6820
rect 32306 6808 32312 6820
rect 32364 6808 32370 6860
rect 17589 6783 17647 6789
rect 17589 6749 17601 6783
rect 17635 6780 17647 6783
rect 17681 6783 17739 6789
rect 17681 6780 17693 6783
rect 17635 6752 17693 6780
rect 17635 6749 17647 6752
rect 17589 6743 17647 6749
rect 17681 6749 17693 6752
rect 17727 6749 17739 6783
rect 17681 6743 17739 6749
rect 22097 6783 22155 6789
rect 22097 6749 22109 6783
rect 22143 6749 22155 6783
rect 22097 6743 22155 6749
rect 22373 6783 22431 6789
rect 22373 6749 22385 6783
rect 22419 6780 22431 6783
rect 32766 6780 32772 6792
rect 22419 6752 32772 6780
rect 22419 6749 22431 6752
rect 22373 6743 22431 6749
rect 32766 6740 32772 6752
rect 32824 6740 32830 6792
rect 38841 6783 38899 6789
rect 38841 6780 38853 6783
rect 38626 6752 38853 6780
rect 1578 6672 1584 6724
rect 1636 6712 1642 6724
rect 1636 6684 21956 6712
rect 1636 6672 1642 6684
rect 4614 6604 4620 6656
rect 4672 6644 4678 6656
rect 9122 6644 9128 6656
rect 4672 6616 9128 6644
rect 4672 6604 4678 6616
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 9217 6647 9275 6653
rect 9217 6613 9229 6647
rect 9263 6644 9275 6647
rect 9398 6644 9404 6656
rect 9263 6616 9404 6644
rect 9263 6613 9275 6616
rect 9217 6607 9275 6613
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 9490 6604 9496 6656
rect 9548 6604 9554 6656
rect 9766 6604 9772 6656
rect 9824 6604 9830 6656
rect 10137 6647 10195 6653
rect 10137 6613 10149 6647
rect 10183 6644 10195 6647
rect 10226 6644 10232 6656
rect 10183 6616 10232 6644
rect 10183 6613 10195 6616
rect 10137 6607 10195 6613
rect 10226 6604 10232 6616
rect 10284 6604 10290 6656
rect 10686 6604 10692 6656
rect 10744 6644 10750 6656
rect 10873 6647 10931 6653
rect 10873 6644 10885 6647
rect 10744 6616 10885 6644
rect 10744 6604 10750 6616
rect 10873 6613 10885 6616
rect 10919 6613 10931 6647
rect 10873 6607 10931 6613
rect 11238 6604 11244 6656
rect 11296 6604 11302 6656
rect 11422 6604 11428 6656
rect 11480 6644 11486 6656
rect 11609 6647 11667 6653
rect 11609 6644 11621 6647
rect 11480 6616 11621 6644
rect 11480 6604 11486 6616
rect 11609 6613 11621 6616
rect 11655 6613 11667 6647
rect 11609 6607 11667 6613
rect 11882 6604 11888 6656
rect 11940 6604 11946 6656
rect 11974 6604 11980 6656
rect 12032 6644 12038 6656
rect 18690 6644 18696 6656
rect 12032 6616 18696 6644
rect 12032 6604 12038 6616
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 21928 6653 21956 6684
rect 31570 6672 31576 6724
rect 31628 6712 31634 6724
rect 38626 6712 38654 6752
rect 38841 6749 38853 6752
rect 38887 6749 38899 6783
rect 38841 6743 38899 6749
rect 39206 6740 39212 6792
rect 39264 6740 39270 6792
rect 39942 6712 39948 6724
rect 31628 6684 38654 6712
rect 39040 6684 39948 6712
rect 31628 6672 31634 6684
rect 21913 6647 21971 6653
rect 21913 6613 21925 6647
rect 21959 6613 21971 6647
rect 21913 6607 21971 6613
rect 22186 6604 22192 6656
rect 22244 6604 22250 6656
rect 39040 6653 39068 6684
rect 39942 6672 39948 6684
rect 40000 6672 40006 6724
rect 39025 6647 39083 6653
rect 39025 6613 39037 6647
rect 39071 6613 39083 6647
rect 39025 6607 39083 6613
rect 39390 6604 39396 6656
rect 39448 6604 39454 6656
rect 1104 6554 39836 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 39010 6554
rect 39062 6502 39074 6554
rect 39126 6502 39138 6554
rect 39190 6502 39202 6554
rect 39254 6502 39266 6554
rect 39318 6502 39836 6554
rect 1104 6480 39836 6502
rect 6546 6400 6552 6452
rect 6604 6440 6610 6452
rect 6604 6412 8984 6440
rect 6604 6400 6610 6412
rect 8478 6264 8484 6316
rect 8536 6304 8542 6316
rect 8849 6307 8907 6313
rect 8849 6304 8861 6307
rect 8536 6276 8861 6304
rect 8536 6264 8542 6276
rect 8849 6273 8861 6276
rect 8895 6273 8907 6307
rect 8956 6304 8984 6412
rect 9398 6400 9404 6452
rect 9456 6440 9462 6452
rect 22278 6440 22284 6452
rect 9456 6412 22284 6440
rect 9456 6400 9462 6412
rect 22278 6400 22284 6412
rect 22336 6400 22342 6452
rect 24670 6400 24676 6452
rect 24728 6440 24734 6452
rect 27433 6443 27491 6449
rect 27433 6440 27445 6443
rect 24728 6412 27445 6440
rect 24728 6400 24734 6412
rect 27433 6409 27445 6412
rect 27479 6409 27491 6443
rect 27433 6403 27491 6409
rect 39390 6400 39396 6452
rect 39448 6400 39454 6452
rect 9122 6332 9128 6384
rect 9180 6372 9186 6384
rect 9582 6372 9588 6384
rect 9180 6344 9588 6372
rect 9180 6332 9186 6344
rect 9582 6332 9588 6344
rect 9640 6332 9646 6384
rect 11514 6332 11520 6384
rect 11572 6372 11578 6384
rect 11572 6344 14228 6372
rect 11572 6332 11578 6344
rect 11698 6304 11704 6316
rect 8956 6276 11704 6304
rect 8849 6267 8907 6273
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 11790 6264 11796 6316
rect 11848 6304 11854 6316
rect 14200 6313 14228 6344
rect 17954 6332 17960 6384
rect 18012 6372 18018 6384
rect 18012 6344 22094 6372
rect 18012 6332 18018 6344
rect 13633 6307 13691 6313
rect 13633 6304 13645 6307
rect 11848 6276 13645 6304
rect 11848 6264 11854 6276
rect 13633 6273 13645 6276
rect 13679 6273 13691 6307
rect 13633 6267 13691 6273
rect 13909 6307 13967 6313
rect 13909 6273 13921 6307
rect 13955 6273 13967 6307
rect 13909 6267 13967 6273
rect 14185 6307 14243 6313
rect 14185 6273 14197 6307
rect 14231 6273 14243 6307
rect 14185 6267 14243 6273
rect 7374 6196 7380 6248
rect 7432 6236 7438 6248
rect 9950 6236 9956 6248
rect 7432 6208 9956 6236
rect 7432 6196 7438 6208
rect 9950 6196 9956 6208
rect 10008 6196 10014 6248
rect 12066 6196 12072 6248
rect 12124 6236 12130 6248
rect 13924 6236 13952 6267
rect 12124 6208 13952 6236
rect 12124 6196 12130 6208
rect 13998 6196 14004 6248
rect 14056 6236 14062 6248
rect 21358 6236 21364 6248
rect 14056 6208 21364 6236
rect 14056 6196 14062 6208
rect 21358 6196 21364 6208
rect 21416 6196 21422 6248
rect 22066 6236 22094 6344
rect 27617 6307 27675 6313
rect 27617 6273 27629 6307
rect 27663 6304 27675 6307
rect 35526 6304 35532 6316
rect 27663 6276 35532 6304
rect 27663 6273 27675 6276
rect 27617 6267 27675 6273
rect 35526 6264 35532 6276
rect 35584 6264 35590 6316
rect 38654 6264 38660 6316
rect 38712 6304 38718 6316
rect 38841 6307 38899 6313
rect 38841 6304 38853 6307
rect 38712 6276 38853 6304
rect 38712 6264 38718 6276
rect 38841 6273 38853 6276
rect 38887 6273 38899 6307
rect 38841 6267 38899 6273
rect 39209 6307 39267 6313
rect 39209 6273 39221 6307
rect 39255 6273 39267 6307
rect 39209 6267 39267 6273
rect 39224 6236 39252 6267
rect 22066 6208 39252 6236
rect 9033 6171 9091 6177
rect 9033 6137 9045 6171
rect 9079 6168 9091 6171
rect 13817 6171 13875 6177
rect 9079 6140 13768 6168
rect 9079 6137 9091 6140
rect 9033 6131 9091 6137
rect 7650 6060 7656 6112
rect 7708 6100 7714 6112
rect 9122 6100 9128 6112
rect 7708 6072 9128 6100
rect 7708 6060 7714 6072
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 13630 6100 13636 6112
rect 9548 6072 13636 6100
rect 9548 6060 9554 6072
rect 13630 6060 13636 6072
rect 13688 6060 13694 6112
rect 13740 6100 13768 6140
rect 13817 6137 13829 6171
rect 13863 6168 13875 6171
rect 20714 6168 20720 6180
rect 13863 6140 20720 6168
rect 13863 6137 13875 6140
rect 13817 6131 13875 6137
rect 20714 6128 20720 6140
rect 20772 6128 20778 6180
rect 22922 6128 22928 6180
rect 22980 6168 22986 6180
rect 33502 6168 33508 6180
rect 22980 6140 33508 6168
rect 22980 6128 22986 6140
rect 33502 6128 33508 6140
rect 33560 6128 33566 6180
rect 13998 6100 14004 6112
rect 13740 6072 14004 6100
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 14093 6103 14151 6109
rect 14093 6069 14105 6103
rect 14139 6100 14151 6103
rect 14274 6100 14280 6112
rect 14139 6072 14280 6100
rect 14139 6069 14151 6072
rect 14093 6063 14151 6069
rect 14274 6060 14280 6072
rect 14332 6060 14338 6112
rect 14369 6103 14427 6109
rect 14369 6069 14381 6103
rect 14415 6100 14427 6103
rect 14918 6100 14924 6112
rect 14415 6072 14924 6100
rect 14415 6069 14427 6072
rect 14369 6063 14427 6069
rect 14918 6060 14924 6072
rect 14976 6060 14982 6112
rect 15010 6060 15016 6112
rect 15068 6100 15074 6112
rect 21818 6100 21824 6112
rect 15068 6072 21824 6100
rect 15068 6060 15074 6072
rect 21818 6060 21824 6072
rect 21876 6060 21882 6112
rect 39022 6060 39028 6112
rect 39080 6060 39086 6112
rect 1104 6010 39836 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 37950 6010
rect 38002 5958 38014 6010
rect 38066 5958 38078 6010
rect 38130 5958 38142 6010
rect 38194 5958 38206 6010
rect 38258 5958 39836 6010
rect 1104 5936 39836 5958
rect 9217 5899 9275 5905
rect 9217 5865 9229 5899
rect 9263 5896 9275 5899
rect 11974 5896 11980 5908
rect 9263 5868 11980 5896
rect 9263 5865 9275 5868
rect 9217 5859 9275 5865
rect 11974 5856 11980 5868
rect 12032 5856 12038 5908
rect 13630 5856 13636 5908
rect 13688 5896 13694 5908
rect 15010 5896 15016 5908
rect 13688 5868 15016 5896
rect 13688 5856 13694 5868
rect 15010 5856 15016 5868
rect 15068 5856 15074 5908
rect 15105 5899 15163 5905
rect 15105 5865 15117 5899
rect 15151 5896 15163 5899
rect 15151 5868 17356 5896
rect 15151 5865 15163 5868
rect 15105 5859 15163 5865
rect 7745 5831 7803 5837
rect 7745 5797 7757 5831
rect 7791 5828 7803 5831
rect 14461 5831 14519 5837
rect 7791 5800 14412 5828
rect 7791 5797 7803 5800
rect 7745 5791 7803 5797
rect 7098 5720 7104 5772
rect 7156 5760 7162 5772
rect 10502 5760 10508 5772
rect 7156 5732 10508 5760
rect 7156 5720 7162 5732
rect 10502 5720 10508 5732
rect 10560 5720 10566 5772
rect 12526 5720 12532 5772
rect 12584 5760 12590 5772
rect 14384 5760 14412 5800
rect 14461 5797 14473 5831
rect 14507 5828 14519 5831
rect 16114 5828 16120 5840
rect 14507 5800 16120 5828
rect 14507 5797 14519 5800
rect 14461 5791 14519 5797
rect 16114 5788 16120 5800
rect 16172 5788 16178 5840
rect 17328 5760 17356 5868
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 19521 5899 19579 5905
rect 19521 5896 19533 5899
rect 17460 5868 19533 5896
rect 17460 5856 17466 5868
rect 19521 5865 19533 5868
rect 19567 5865 19579 5899
rect 19521 5859 19579 5865
rect 22066 5868 26280 5896
rect 19889 5831 19947 5837
rect 19889 5797 19901 5831
rect 19935 5828 19947 5831
rect 22066 5828 22094 5868
rect 19935 5800 22094 5828
rect 19935 5797 19947 5800
rect 19889 5791 19947 5797
rect 20806 5760 20812 5772
rect 12584 5732 14320 5760
rect 14384 5732 16068 5760
rect 17328 5732 20812 5760
rect 12584 5720 12590 5732
rect 5166 5652 5172 5704
rect 5224 5692 5230 5704
rect 7561 5695 7619 5701
rect 7561 5692 7573 5695
rect 5224 5664 7573 5692
rect 5224 5652 5230 5664
rect 7561 5661 7573 5664
rect 7607 5661 7619 5695
rect 7561 5655 7619 5661
rect 9033 5695 9091 5701
rect 9033 5661 9045 5695
rect 9079 5661 9091 5695
rect 9033 5655 9091 5661
rect 4982 5584 4988 5636
rect 5040 5624 5046 5636
rect 9048 5624 9076 5655
rect 11238 5652 11244 5704
rect 11296 5692 11302 5704
rect 13449 5695 13507 5701
rect 13449 5692 13461 5695
rect 11296 5664 13461 5692
rect 11296 5652 11302 5664
rect 13449 5661 13461 5664
rect 13495 5661 13507 5695
rect 13449 5655 13507 5661
rect 13722 5652 13728 5704
rect 13780 5652 13786 5704
rect 14292 5701 14320 5732
rect 14277 5695 14335 5701
rect 14277 5661 14289 5695
rect 14323 5661 14335 5695
rect 14277 5655 14335 5661
rect 14550 5652 14556 5704
rect 14608 5652 14614 5704
rect 14921 5695 14979 5701
rect 14921 5692 14933 5695
rect 14660 5664 14933 5692
rect 5040 5596 9076 5624
rect 5040 5584 5046 5596
rect 12618 5584 12624 5636
rect 12676 5624 12682 5636
rect 14660 5624 14688 5664
rect 14921 5661 14933 5664
rect 14967 5661 14979 5695
rect 16040 5692 16068 5732
rect 20806 5720 20812 5732
rect 20864 5720 20870 5772
rect 26252 5760 26280 5868
rect 26326 5856 26332 5908
rect 26384 5856 26390 5908
rect 39390 5788 39396 5840
rect 39448 5788 39454 5840
rect 31570 5760 31576 5772
rect 26252 5732 31576 5760
rect 31570 5720 31576 5732
rect 31628 5720 31634 5772
rect 19518 5692 19524 5704
rect 16040 5664 19524 5692
rect 14921 5655 14979 5661
rect 19518 5652 19524 5664
rect 19576 5652 19582 5704
rect 19613 5695 19671 5701
rect 19613 5661 19625 5695
rect 19659 5692 19671 5695
rect 19705 5695 19763 5701
rect 19705 5692 19717 5695
rect 19659 5664 19717 5692
rect 19659 5661 19671 5664
rect 19613 5655 19671 5661
rect 19705 5661 19717 5664
rect 19751 5661 19763 5695
rect 19705 5655 19763 5661
rect 26145 5695 26203 5701
rect 26145 5661 26157 5695
rect 26191 5692 26203 5695
rect 35802 5692 35808 5704
rect 26191 5664 35808 5692
rect 26191 5661 26203 5664
rect 26145 5655 26203 5661
rect 35802 5652 35808 5664
rect 35860 5652 35866 5704
rect 38838 5652 38844 5704
rect 38896 5652 38902 5704
rect 39209 5695 39267 5701
rect 39209 5661 39221 5695
rect 39255 5661 39267 5695
rect 39209 5655 39267 5661
rect 12676 5596 14688 5624
rect 14752 5596 20024 5624
rect 12676 5584 12682 5596
rect 6822 5516 6828 5568
rect 6880 5556 6886 5568
rect 10870 5556 10876 5568
rect 6880 5528 10876 5556
rect 6880 5516 6886 5528
rect 10870 5516 10876 5528
rect 10928 5516 10934 5568
rect 13630 5516 13636 5568
rect 13688 5516 13694 5568
rect 13909 5559 13967 5565
rect 13909 5525 13921 5559
rect 13955 5556 13967 5559
rect 14366 5556 14372 5568
rect 13955 5528 14372 5556
rect 13955 5525 13967 5528
rect 13909 5519 13967 5525
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 14752 5565 14780 5596
rect 14737 5559 14795 5565
rect 14737 5525 14749 5559
rect 14783 5525 14795 5559
rect 19996 5556 20024 5596
rect 20438 5584 20444 5636
rect 20496 5624 20502 5636
rect 39224 5624 39252 5655
rect 20496 5596 39252 5624
rect 20496 5584 20502 5596
rect 24854 5556 24860 5568
rect 19996 5528 24860 5556
rect 14737 5519 14795 5525
rect 24854 5516 24860 5528
rect 24912 5516 24918 5568
rect 39025 5559 39083 5565
rect 39025 5525 39037 5559
rect 39071 5556 39083 5559
rect 39942 5556 39948 5568
rect 39071 5528 39948 5556
rect 39071 5525 39083 5528
rect 39025 5519 39083 5525
rect 39942 5516 39948 5528
rect 40000 5516 40006 5568
rect 1104 5466 39836 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 39010 5466
rect 39062 5414 39074 5466
rect 39126 5414 39138 5466
rect 39190 5414 39202 5466
rect 39254 5414 39266 5466
rect 39318 5414 39836 5466
rect 1104 5392 39836 5414
rect 3145 5355 3203 5361
rect 3145 5321 3157 5355
rect 3191 5352 3203 5355
rect 6086 5352 6092 5364
rect 3191 5324 6092 5352
rect 3191 5321 3203 5324
rect 3145 5315 3203 5321
rect 6086 5312 6092 5324
rect 6144 5312 6150 5364
rect 6181 5355 6239 5361
rect 6181 5321 6193 5355
rect 6227 5352 6239 5355
rect 9582 5352 9588 5364
rect 6227 5324 9588 5352
rect 6227 5321 6239 5324
rect 6181 5315 6239 5321
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 11054 5312 11060 5364
rect 11112 5352 11118 5364
rect 16117 5355 16175 5361
rect 11112 5324 16068 5352
rect 11112 5312 11118 5324
rect 10134 5244 10140 5296
rect 10192 5284 10198 5296
rect 10192 5256 15976 5284
rect 10192 5244 10198 5256
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5185 2743 5219
rect 2685 5179 2743 5185
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5185 3019 5219
rect 2961 5179 3019 5185
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5216 3295 5219
rect 3510 5216 3516 5228
rect 3283 5188 3516 5216
rect 3283 5185 3295 5188
rect 3237 5179 3295 5185
rect 2700 5080 2728 5179
rect 2976 5148 3004 5179
rect 3510 5176 3516 5188
rect 3568 5176 3574 5228
rect 5442 5176 5448 5228
rect 5500 5216 5506 5228
rect 5997 5219 6055 5225
rect 5997 5216 6009 5219
rect 5500 5188 6009 5216
rect 5500 5176 5506 5188
rect 5997 5185 6009 5188
rect 6043 5185 6055 5219
rect 5997 5179 6055 5185
rect 10410 5176 10416 5228
rect 10468 5216 10474 5228
rect 15948 5225 15976 5256
rect 15381 5219 15439 5225
rect 15381 5216 15393 5219
rect 10468 5188 15393 5216
rect 10468 5176 10474 5188
rect 15381 5185 15393 5188
rect 15427 5185 15439 5219
rect 15381 5179 15439 5185
rect 15657 5219 15715 5225
rect 15657 5185 15669 5219
rect 15703 5185 15715 5219
rect 15657 5179 15715 5185
rect 15933 5219 15991 5225
rect 15933 5185 15945 5219
rect 15979 5185 15991 5219
rect 16040 5216 16068 5324
rect 16117 5321 16129 5355
rect 16163 5321 16175 5355
rect 16117 5315 16175 5321
rect 16132 5284 16160 5315
rect 17954 5312 17960 5364
rect 18012 5312 18018 5364
rect 22002 5312 22008 5364
rect 22060 5352 22066 5364
rect 22060 5324 31754 5352
rect 22060 5312 22066 5324
rect 24118 5284 24124 5296
rect 16132 5256 24124 5284
rect 24118 5244 24124 5256
rect 24176 5244 24182 5296
rect 31726 5284 31754 5324
rect 36814 5312 36820 5364
rect 36872 5352 36878 5364
rect 36909 5355 36967 5361
rect 36909 5352 36921 5355
rect 36872 5324 36921 5352
rect 36872 5312 36878 5324
rect 36909 5321 36921 5324
rect 36955 5321 36967 5355
rect 36909 5315 36967 5321
rect 39390 5312 39396 5364
rect 39448 5312 39454 5364
rect 31726 5256 38884 5284
rect 17589 5219 17647 5225
rect 17589 5216 17601 5219
rect 16040 5188 17601 5216
rect 15933 5179 15991 5185
rect 17589 5185 17601 5188
rect 17635 5216 17647 5219
rect 17773 5219 17831 5225
rect 17773 5216 17785 5219
rect 17635 5188 17785 5216
rect 17635 5185 17647 5188
rect 17589 5179 17647 5185
rect 17773 5185 17785 5188
rect 17819 5185 17831 5219
rect 17773 5179 17831 5185
rect 4062 5148 4068 5160
rect 2976 5120 4068 5148
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 12894 5108 12900 5160
rect 12952 5148 12958 5160
rect 15672 5148 15700 5179
rect 22370 5176 22376 5228
rect 22428 5176 22434 5228
rect 28074 5176 28080 5228
rect 28132 5216 28138 5228
rect 31386 5216 31392 5228
rect 28132 5188 31392 5216
rect 28132 5176 28138 5188
rect 31386 5176 31392 5188
rect 31444 5176 31450 5228
rect 37093 5219 37151 5225
rect 37093 5185 37105 5219
rect 37139 5216 37151 5219
rect 37734 5216 37740 5228
rect 37139 5188 37740 5216
rect 37139 5185 37151 5188
rect 37093 5179 37151 5185
rect 37734 5176 37740 5188
rect 37792 5176 37798 5228
rect 38856 5225 38884 5256
rect 38841 5219 38899 5225
rect 38841 5185 38853 5219
rect 38887 5185 38899 5219
rect 38841 5179 38899 5185
rect 39206 5176 39212 5228
rect 39264 5176 39270 5228
rect 27430 5148 27436 5160
rect 12952 5120 15700 5148
rect 22066 5120 27436 5148
rect 12952 5108 12958 5120
rect 3786 5080 3792 5092
rect 2700 5052 3792 5080
rect 3786 5040 3792 5052
rect 3844 5040 3850 5092
rect 15841 5083 15899 5089
rect 15841 5049 15853 5083
rect 15887 5080 15899 5083
rect 15887 5052 21680 5080
rect 15887 5049 15899 5052
rect 15841 5043 15899 5049
rect 2869 5015 2927 5021
rect 2869 4981 2881 5015
rect 2915 5012 2927 5015
rect 3050 5012 3056 5024
rect 2915 4984 3056 5012
rect 2915 4981 2927 4984
rect 2869 4975 2927 4981
rect 3050 4972 3056 4984
rect 3108 4972 3114 5024
rect 3421 5015 3479 5021
rect 3421 4981 3433 5015
rect 3467 5012 3479 5015
rect 5350 5012 5356 5024
rect 3467 4984 5356 5012
rect 3467 4981 3479 4984
rect 3421 4975 3479 4981
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 5534 4972 5540 5024
rect 5592 5012 5598 5024
rect 11146 5012 11152 5024
rect 5592 4984 11152 5012
rect 5592 4972 5598 4984
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 15562 4972 15568 5024
rect 15620 4972 15626 5024
rect 21652 5012 21680 5052
rect 21726 5040 21732 5092
rect 21784 5080 21790 5092
rect 22066 5080 22094 5120
rect 27430 5108 27436 5120
rect 27488 5108 27494 5160
rect 27614 5108 27620 5160
rect 27672 5148 27678 5160
rect 32490 5148 32496 5160
rect 27672 5120 32496 5148
rect 27672 5108 27678 5120
rect 32490 5108 32496 5120
rect 32548 5108 32554 5160
rect 21784 5052 22094 5080
rect 21784 5040 21790 5052
rect 23198 5040 23204 5092
rect 23256 5080 23262 5092
rect 33778 5080 33784 5092
rect 23256 5052 33784 5080
rect 23256 5040 23262 5052
rect 33778 5040 33784 5052
rect 33836 5040 33842 5092
rect 22462 5012 22468 5024
rect 21652 4984 22468 5012
rect 22462 4972 22468 4984
rect 22520 4972 22526 5024
rect 22557 5015 22615 5021
rect 22557 4981 22569 5015
rect 22603 5012 22615 5015
rect 38654 5012 38660 5024
rect 22603 4984 38660 5012
rect 22603 4981 22615 4984
rect 22557 4975 22615 4981
rect 38654 4972 38660 4984
rect 38712 4972 38718 5024
rect 39022 4972 39028 5024
rect 39080 4972 39086 5024
rect 1104 4922 39836 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 37950 4922
rect 38002 4870 38014 4922
rect 38066 4870 38078 4922
rect 38130 4870 38142 4922
rect 38194 4870 38206 4922
rect 38258 4870 39836 4922
rect 1104 4848 39836 4870
rect 6086 4768 6092 4820
rect 6144 4808 6150 4820
rect 16666 4808 16672 4820
rect 6144 4780 16672 4808
rect 6144 4768 6150 4780
rect 16666 4768 16672 4780
rect 16724 4768 16730 4820
rect 16761 4811 16819 4817
rect 16761 4777 16773 4811
rect 16807 4808 16819 4811
rect 21726 4808 21732 4820
rect 16807 4780 21732 4808
rect 16807 4777 16819 4780
rect 16761 4771 16819 4777
rect 21726 4768 21732 4780
rect 21784 4768 21790 4820
rect 23198 4768 23204 4820
rect 23256 4768 23262 4820
rect 23474 4768 23480 4820
rect 23532 4768 23538 4820
rect 23750 4768 23756 4820
rect 23808 4808 23814 4820
rect 23808 4780 27568 4808
rect 23808 4768 23814 4780
rect 4890 4700 4896 4752
rect 4948 4700 4954 4752
rect 15562 4700 15568 4752
rect 15620 4740 15626 4752
rect 23845 4743 23903 4749
rect 15620 4712 22094 4740
rect 15620 4700 15626 4712
rect 5350 4632 5356 4684
rect 5408 4672 5414 4684
rect 17770 4672 17776 4684
rect 5408 4644 17776 4672
rect 5408 4632 5414 4644
rect 17770 4632 17776 4644
rect 17828 4632 17834 4684
rect 19794 4632 19800 4684
rect 19852 4672 19858 4684
rect 20073 4675 20131 4681
rect 20073 4672 20085 4675
rect 19852 4644 20085 4672
rect 19852 4632 19858 4644
rect 20073 4641 20085 4644
rect 20119 4641 20131 4675
rect 20073 4635 20131 4641
rect 2866 4564 2872 4616
rect 2924 4604 2930 4616
rect 2961 4607 3019 4613
rect 2961 4604 2973 4607
rect 2924 4576 2973 4604
rect 2924 4564 2930 4576
rect 2961 4573 2973 4576
rect 3007 4573 3019 4607
rect 2961 4567 3019 4573
rect 4246 4564 4252 4616
rect 4304 4564 4310 4616
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4604 4767 4607
rect 5718 4604 5724 4616
rect 4755 4576 5724 4604
rect 4755 4573 4767 4576
rect 4709 4567 4767 4573
rect 5718 4564 5724 4576
rect 5776 4564 5782 4616
rect 8662 4564 8668 4616
rect 8720 4604 8726 4616
rect 9858 4604 9864 4616
rect 8720 4576 9864 4604
rect 8720 4564 8726 4576
rect 9858 4564 9864 4576
rect 9916 4564 9922 4616
rect 16574 4564 16580 4616
rect 16632 4564 16638 4616
rect 20165 4607 20223 4613
rect 20165 4573 20177 4607
rect 20211 4604 20223 4607
rect 20257 4607 20315 4613
rect 20257 4604 20269 4607
rect 20211 4576 20269 4604
rect 20211 4573 20223 4576
rect 20165 4567 20223 4573
rect 20257 4573 20269 4576
rect 20303 4573 20315 4607
rect 20257 4567 20315 4573
rect 3050 4496 3056 4548
rect 3108 4536 3114 4548
rect 17954 4536 17960 4548
rect 3108 4508 17960 4536
rect 3108 4496 3114 4508
rect 17954 4496 17960 4508
rect 18012 4496 18018 4548
rect 22066 4536 22094 4712
rect 23845 4709 23857 4743
rect 23891 4709 23903 4743
rect 23845 4703 23903 4709
rect 22830 4632 22836 4684
rect 22888 4632 22894 4684
rect 23860 4672 23888 4703
rect 25038 4700 25044 4752
rect 25096 4740 25102 4752
rect 27249 4743 27307 4749
rect 27249 4740 27261 4743
rect 25096 4712 27261 4740
rect 25096 4700 25102 4712
rect 27249 4709 27261 4712
rect 27295 4709 27307 4743
rect 27540 4740 27568 4780
rect 27614 4768 27620 4820
rect 27672 4768 27678 4820
rect 29365 4811 29423 4817
rect 29365 4777 29377 4811
rect 29411 4808 29423 4811
rect 31294 4808 31300 4820
rect 29411 4780 31300 4808
rect 29411 4777 29423 4780
rect 29365 4771 29423 4777
rect 31294 4768 31300 4780
rect 31352 4768 31358 4820
rect 31386 4768 31392 4820
rect 31444 4808 31450 4820
rect 33321 4811 33379 4817
rect 31444 4780 32168 4808
rect 31444 4768 31450 4780
rect 29825 4743 29883 4749
rect 27540 4712 29684 4740
rect 27249 4703 27307 4709
rect 23860 4644 29500 4672
rect 22925 4607 22983 4613
rect 22925 4573 22937 4607
rect 22971 4604 22983 4607
rect 23017 4607 23075 4613
rect 23017 4604 23029 4607
rect 22971 4576 23029 4604
rect 22971 4573 22983 4576
rect 22925 4567 22983 4573
rect 23017 4573 23029 4576
rect 23063 4573 23075 4607
rect 23017 4567 23075 4573
rect 23569 4607 23627 4613
rect 23569 4573 23581 4607
rect 23615 4604 23627 4607
rect 23661 4607 23719 4613
rect 23661 4604 23673 4607
rect 23615 4576 23673 4604
rect 23615 4573 23627 4576
rect 23569 4567 23627 4573
rect 23661 4573 23673 4576
rect 23707 4573 23719 4607
rect 23661 4567 23719 4573
rect 24026 4564 24032 4616
rect 24084 4604 24090 4616
rect 24397 4607 24455 4613
rect 24397 4604 24409 4607
rect 24084 4576 24409 4604
rect 24084 4564 24090 4576
rect 24397 4573 24409 4576
rect 24443 4573 24455 4607
rect 24397 4567 24455 4573
rect 25409 4607 25467 4613
rect 25409 4573 25421 4607
rect 25455 4604 25467 4607
rect 25682 4604 25688 4616
rect 25455 4576 25688 4604
rect 25455 4573 25467 4576
rect 25409 4567 25467 4573
rect 25682 4564 25688 4576
rect 25740 4564 25746 4616
rect 26513 4607 26571 4613
rect 26513 4573 26525 4607
rect 26559 4604 26571 4607
rect 26602 4604 26608 4616
rect 26559 4576 26608 4604
rect 26559 4573 26571 4576
rect 26513 4567 26571 4573
rect 26602 4564 26608 4576
rect 26660 4564 26666 4616
rect 27341 4607 27399 4613
rect 27341 4573 27353 4607
rect 27387 4604 27399 4607
rect 27433 4607 27491 4613
rect 27433 4604 27445 4607
rect 27387 4576 27445 4604
rect 27387 4573 27399 4576
rect 27341 4567 27399 4573
rect 27433 4573 27445 4576
rect 27479 4573 27491 4607
rect 27433 4567 27491 4573
rect 28721 4607 28779 4613
rect 28721 4573 28733 4607
rect 28767 4573 28779 4607
rect 28721 4567 28779 4573
rect 29089 4607 29147 4613
rect 29089 4573 29101 4607
rect 29135 4604 29147 4607
rect 29181 4607 29239 4613
rect 29181 4604 29193 4607
rect 29135 4576 29193 4604
rect 29135 4573 29147 4576
rect 29089 4567 29147 4573
rect 29181 4573 29193 4576
rect 29227 4573 29239 4607
rect 29181 4567 29239 4573
rect 25866 4536 25872 4548
rect 22066 4508 25872 4536
rect 25866 4496 25872 4508
rect 25924 4496 25930 4548
rect 26786 4496 26792 4548
rect 26844 4536 26850 4548
rect 28736 4536 28764 4567
rect 26844 4508 28764 4536
rect 26844 4496 26850 4508
rect 3145 4471 3203 4477
rect 3145 4437 3157 4471
rect 3191 4468 3203 4471
rect 4338 4468 4344 4480
rect 3191 4440 4344 4468
rect 3191 4437 3203 4440
rect 3145 4431 3203 4437
rect 4338 4428 4344 4440
rect 4396 4428 4402 4480
rect 4433 4471 4491 4477
rect 4433 4437 4445 4471
rect 4479 4468 4491 4471
rect 11054 4468 11060 4480
rect 4479 4440 11060 4468
rect 4479 4437 4491 4440
rect 4433 4431 4491 4437
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 20438 4428 20444 4480
rect 20496 4428 20502 4480
rect 24210 4428 24216 4480
rect 24268 4428 24274 4480
rect 25590 4428 25596 4480
rect 25648 4428 25654 4480
rect 26418 4428 26424 4480
rect 26476 4468 26482 4480
rect 26697 4471 26755 4477
rect 26697 4468 26709 4471
rect 26476 4440 26709 4468
rect 26476 4428 26482 4440
rect 26697 4437 26709 4440
rect 26743 4437 26755 4471
rect 26697 4431 26755 4437
rect 28534 4428 28540 4480
rect 28592 4468 28598 4480
rect 28905 4471 28963 4477
rect 28905 4468 28917 4471
rect 28592 4440 28917 4468
rect 28592 4428 28598 4440
rect 28905 4437 28917 4440
rect 28951 4437 28963 4471
rect 28905 4431 28963 4437
rect 28994 4428 29000 4480
rect 29052 4428 29058 4480
rect 29472 4468 29500 4644
rect 29656 4613 29684 4712
rect 29825 4709 29837 4743
rect 29871 4740 29883 4743
rect 30834 4740 30840 4752
rect 29871 4712 30840 4740
rect 29871 4709 29883 4712
rect 29825 4703 29883 4709
rect 30834 4700 30840 4712
rect 30892 4700 30898 4752
rect 31570 4632 31576 4684
rect 31628 4632 31634 4684
rect 31754 4632 31760 4684
rect 31812 4672 31818 4684
rect 31812 4644 31984 4672
rect 31812 4632 31818 4644
rect 29641 4607 29699 4613
rect 29641 4573 29653 4607
rect 29687 4604 29699 4607
rect 29917 4607 29975 4613
rect 29917 4604 29929 4607
rect 29687 4576 29929 4604
rect 29687 4573 29699 4576
rect 29641 4567 29699 4573
rect 29917 4573 29929 4576
rect 29963 4573 29975 4607
rect 29917 4567 29975 4573
rect 30193 4607 30251 4613
rect 30193 4573 30205 4607
rect 30239 4604 30251 4607
rect 30285 4607 30343 4613
rect 30285 4604 30297 4607
rect 30239 4576 30297 4604
rect 30239 4573 30251 4576
rect 30193 4567 30251 4573
rect 30285 4573 30297 4576
rect 30331 4573 30343 4607
rect 30285 4567 30343 4573
rect 30837 4607 30895 4613
rect 30837 4573 30849 4607
rect 30883 4604 30895 4607
rect 31846 4604 31852 4616
rect 30883 4576 31852 4604
rect 30883 4573 30895 4576
rect 30837 4567 30895 4573
rect 31846 4564 31852 4576
rect 31904 4564 31910 4616
rect 31956 4613 31984 4644
rect 31941 4607 31999 4613
rect 31941 4573 31953 4607
rect 31987 4573 31999 4607
rect 32140 4604 32168 4780
rect 33321 4777 33333 4811
rect 33367 4808 33379 4811
rect 35986 4808 35992 4820
rect 33367 4780 35992 4808
rect 33367 4777 33379 4780
rect 33321 4771 33379 4777
rect 35986 4768 35992 4780
rect 36044 4768 36050 4820
rect 33778 4700 33784 4752
rect 33836 4740 33842 4752
rect 33836 4712 39252 4740
rect 33836 4700 33842 4712
rect 37090 4672 37096 4684
rect 33152 4644 37096 4672
rect 32217 4607 32275 4613
rect 32217 4604 32229 4607
rect 32140 4576 32229 4604
rect 31941 4567 31999 4573
rect 32217 4573 32229 4576
rect 32263 4573 32275 4607
rect 32217 4567 32275 4573
rect 32493 4607 32551 4613
rect 32493 4573 32505 4607
rect 32539 4604 32551 4607
rect 32674 4604 32680 4616
rect 32539 4576 32680 4604
rect 32539 4573 32551 4576
rect 32493 4567 32551 4573
rect 32674 4564 32680 4576
rect 32732 4564 32738 4616
rect 33152 4613 33180 4644
rect 37090 4632 37096 4644
rect 37148 4632 37154 4684
rect 33137 4607 33195 4613
rect 33137 4573 33149 4607
rect 33183 4573 33195 4607
rect 33137 4567 33195 4573
rect 35713 4607 35771 4613
rect 35713 4573 35725 4607
rect 35759 4604 35771 4607
rect 37458 4604 37464 4616
rect 35759 4576 37464 4604
rect 35759 4573 35771 4576
rect 35713 4567 35771 4573
rect 37458 4564 37464 4576
rect 37516 4564 37522 4616
rect 39224 4613 39252 4712
rect 39390 4700 39396 4752
rect 39448 4700 39454 4752
rect 38841 4607 38899 4613
rect 38841 4573 38853 4607
rect 38887 4573 38899 4607
rect 38841 4567 38899 4573
rect 39209 4607 39267 4613
rect 39209 4573 39221 4607
rect 39255 4573 39267 4607
rect 39209 4567 39267 4573
rect 29546 4496 29552 4548
rect 29604 4536 29610 4548
rect 30101 4539 30159 4545
rect 30101 4536 30113 4539
rect 29604 4508 30113 4536
rect 29604 4496 29610 4508
rect 30101 4505 30113 4508
rect 30147 4505 30159 4539
rect 38856 4536 38884 4567
rect 30101 4499 30159 4505
rect 30208 4508 38884 4536
rect 30208 4468 30236 4508
rect 29472 4440 30236 4468
rect 30469 4471 30527 4477
rect 30469 4437 30481 4471
rect 30515 4468 30527 4471
rect 30926 4468 30932 4480
rect 30515 4440 30932 4468
rect 30515 4437 30527 4440
rect 30469 4431 30527 4437
rect 30926 4428 30932 4440
rect 30984 4428 30990 4480
rect 31018 4428 31024 4480
rect 31076 4428 31082 4480
rect 31754 4428 31760 4480
rect 31812 4428 31818 4480
rect 31846 4428 31852 4480
rect 31904 4468 31910 4480
rect 32033 4471 32091 4477
rect 32033 4468 32045 4471
rect 31904 4440 32045 4468
rect 31904 4428 31910 4440
rect 32033 4437 32045 4440
rect 32079 4437 32091 4471
rect 32033 4431 32091 4437
rect 32309 4471 32367 4477
rect 32309 4437 32321 4471
rect 32355 4468 32367 4471
rect 32398 4468 32404 4480
rect 32355 4440 32404 4468
rect 32355 4437 32367 4440
rect 32309 4431 32367 4437
rect 32398 4428 32404 4440
rect 32456 4428 32462 4480
rect 35897 4471 35955 4477
rect 35897 4437 35909 4471
rect 35943 4468 35955 4471
rect 37182 4468 37188 4480
rect 35943 4440 37188 4468
rect 35943 4437 35955 4440
rect 35897 4431 35955 4437
rect 37182 4428 37188 4440
rect 37240 4428 37246 4480
rect 39025 4471 39083 4477
rect 39025 4437 39037 4471
rect 39071 4468 39083 4471
rect 39942 4468 39948 4480
rect 39071 4440 39948 4468
rect 39071 4437 39083 4440
rect 39025 4431 39083 4437
rect 39942 4428 39948 4440
rect 40000 4428 40006 4480
rect 1104 4378 39836 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 39010 4378
rect 39062 4326 39074 4378
rect 39126 4326 39138 4378
rect 39190 4326 39202 4378
rect 39254 4326 39266 4378
rect 39318 4326 39836 4378
rect 1104 4304 39836 4326
rect 4890 4224 4896 4276
rect 4948 4264 4954 4276
rect 9674 4264 9680 4276
rect 4948 4236 9680 4264
rect 4948 4224 4954 4236
rect 9674 4224 9680 4236
rect 9732 4224 9738 4276
rect 9858 4224 9864 4276
rect 9916 4264 9922 4276
rect 21910 4264 21916 4276
rect 9916 4236 21916 4264
rect 9916 4224 9922 4236
rect 21910 4224 21916 4236
rect 21968 4224 21974 4276
rect 24210 4224 24216 4276
rect 24268 4264 24274 4276
rect 35894 4264 35900 4276
rect 24268 4236 35900 4264
rect 24268 4224 24274 4236
rect 35894 4224 35900 4236
rect 35952 4224 35958 4276
rect 4338 4156 4344 4208
rect 4396 4196 4402 4208
rect 10870 4196 10876 4208
rect 4396 4168 10876 4196
rect 4396 4156 4402 4168
rect 10870 4156 10876 4168
rect 10928 4156 10934 4208
rect 11146 4156 11152 4208
rect 11204 4196 11210 4208
rect 21726 4196 21732 4208
rect 11204 4168 21732 4196
rect 11204 4156 11210 4168
rect 21726 4156 21732 4168
rect 21784 4156 21790 4208
rect 23658 4156 23664 4208
rect 23716 4196 23722 4208
rect 28994 4196 29000 4208
rect 23716 4168 29000 4196
rect 23716 4156 23722 4168
rect 28994 4156 29000 4168
rect 29052 4156 29058 4208
rect 29840 4168 31708 4196
rect 4709 4131 4767 4137
rect 4709 4097 4721 4131
rect 4755 4128 4767 4131
rect 6270 4128 6276 4140
rect 4755 4100 6276 4128
rect 4755 4097 4767 4100
rect 4709 4091 4767 4097
rect 6270 4088 6276 4100
rect 6328 4088 6334 4140
rect 9490 4088 9496 4140
rect 9548 4128 9554 4140
rect 17037 4131 17095 4137
rect 17037 4128 17049 4131
rect 9548 4100 17049 4128
rect 9548 4088 9554 4100
rect 17037 4097 17049 4100
rect 17083 4097 17095 4131
rect 17037 4091 17095 4097
rect 17497 4131 17555 4137
rect 17497 4097 17509 4131
rect 17543 4097 17555 4131
rect 17497 4091 17555 4097
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 17512 4060 17540 4091
rect 19426 4088 19432 4140
rect 19484 4088 19490 4140
rect 21542 4088 21548 4140
rect 21600 4128 21606 4140
rect 21821 4131 21879 4137
rect 21821 4128 21833 4131
rect 21600 4100 21833 4128
rect 21600 4088 21606 4100
rect 21821 4097 21833 4100
rect 21867 4097 21879 4131
rect 21821 4091 21879 4097
rect 22094 4088 22100 4140
rect 22152 4128 22158 4140
rect 22189 4131 22247 4137
rect 22189 4128 22201 4131
rect 22152 4100 22201 4128
rect 22152 4088 22158 4100
rect 22189 4097 22201 4100
rect 22235 4128 22247 4131
rect 22465 4131 22523 4137
rect 22465 4128 22477 4131
rect 22235 4100 22477 4128
rect 22235 4097 22247 4100
rect 22189 4091 22247 4097
rect 22465 4097 22477 4100
rect 22511 4097 22523 4131
rect 22465 4091 22523 4097
rect 24305 4131 24363 4137
rect 24305 4097 24317 4131
rect 24351 4128 24363 4131
rect 24397 4131 24455 4137
rect 24397 4128 24409 4131
rect 24351 4100 24409 4128
rect 24351 4097 24363 4100
rect 24305 4091 24363 4097
rect 24397 4097 24409 4100
rect 24443 4097 24455 4131
rect 25406 4128 25412 4140
rect 24397 4091 24455 4097
rect 24504 4100 25412 4128
rect 24504 4060 24532 4100
rect 25406 4088 25412 4100
rect 25464 4088 25470 4140
rect 27249 4131 27307 4137
rect 27249 4097 27261 4131
rect 27295 4128 27307 4131
rect 27341 4131 27399 4137
rect 27341 4128 27353 4131
rect 27295 4100 27353 4128
rect 27295 4097 27307 4100
rect 27249 4091 27307 4097
rect 27341 4097 27353 4100
rect 27387 4097 27399 4131
rect 27341 4091 27399 4097
rect 28166 4088 28172 4140
rect 28224 4088 28230 4140
rect 29089 4131 29147 4137
rect 29089 4097 29101 4131
rect 29135 4128 29147 4131
rect 29365 4131 29423 4137
rect 29365 4128 29377 4131
rect 29135 4100 29377 4128
rect 29135 4097 29147 4100
rect 29089 4091 29147 4097
rect 29365 4097 29377 4100
rect 29411 4097 29423 4131
rect 29365 4091 29423 4097
rect 29454 4088 29460 4140
rect 29512 4128 29518 4140
rect 29840 4128 29868 4168
rect 29512 4100 29868 4128
rect 29917 4131 29975 4137
rect 29512 4088 29518 4100
rect 29917 4097 29929 4131
rect 29963 4128 29975 4131
rect 30193 4131 30251 4137
rect 30193 4128 30205 4131
rect 29963 4100 30205 4128
rect 29963 4097 29975 4100
rect 29917 4091 29975 4097
rect 30193 4097 30205 4100
rect 30239 4097 30251 4131
rect 30193 4091 30251 4097
rect 30374 4088 30380 4140
rect 30432 4128 30438 4140
rect 30837 4131 30895 4137
rect 30837 4128 30849 4131
rect 30432 4100 30849 4128
rect 30432 4088 30438 4100
rect 30837 4097 30849 4100
rect 30883 4097 30895 4131
rect 30837 4091 30895 4097
rect 31021 4131 31079 4137
rect 31021 4097 31033 4131
rect 31067 4128 31079 4131
rect 31297 4131 31355 4137
rect 31297 4128 31309 4131
rect 31067 4100 31309 4128
rect 31067 4097 31079 4100
rect 31021 4091 31079 4097
rect 31297 4097 31309 4100
rect 31343 4097 31355 4131
rect 31297 4091 31355 4097
rect 31570 4088 31576 4140
rect 31628 4088 31634 4140
rect 31680 4128 31708 4168
rect 31938 4156 31944 4208
rect 31996 4196 32002 4208
rect 36906 4196 36912 4208
rect 31996 4168 36912 4196
rect 31996 4156 32002 4168
rect 36906 4156 36912 4168
rect 36964 4156 36970 4208
rect 38841 4131 38899 4137
rect 38841 4128 38853 4131
rect 31680 4100 38853 4128
rect 38841 4097 38853 4100
rect 38887 4097 38899 4131
rect 38841 4091 38899 4097
rect 39209 4131 39267 4137
rect 39209 4097 39221 4131
rect 39255 4097 39267 4131
rect 39209 4091 39267 4097
rect 9456 4032 17540 4060
rect 19306 4032 24532 4060
rect 24596 4032 29408 4060
rect 9456 4020 9462 4032
rect 10686 3952 10692 4004
rect 10744 3992 10750 4004
rect 10962 3992 10968 4004
rect 10744 3964 10968 3992
rect 10744 3952 10750 3964
rect 10962 3952 10968 3964
rect 11020 3952 11026 4004
rect 17681 3995 17739 4001
rect 17681 3961 17693 3995
rect 17727 3992 17739 3995
rect 19306 3992 19334 4032
rect 17727 3964 19334 3992
rect 17727 3961 17739 3964
rect 17681 3955 17739 3961
rect 22002 3952 22008 4004
rect 22060 3952 22066 4004
rect 24596 4001 24624 4032
rect 22373 3995 22431 4001
rect 22373 3961 22385 3995
rect 22419 3992 22431 3995
rect 24581 3995 24639 4001
rect 22419 3964 24532 3992
rect 22419 3961 22431 3964
rect 22373 3955 22431 3961
rect 4890 3884 4896 3936
rect 4948 3884 4954 3936
rect 11882 3884 11888 3936
rect 11940 3924 11946 3936
rect 17126 3924 17132 3936
rect 11940 3896 17132 3924
rect 11940 3884 11946 3896
rect 17126 3884 17132 3896
rect 17184 3884 17190 3936
rect 17221 3927 17279 3933
rect 17221 3893 17233 3927
rect 17267 3924 17279 3927
rect 19518 3924 19524 3936
rect 17267 3896 19524 3924
rect 17267 3893 17279 3896
rect 17221 3887 17279 3893
rect 19518 3884 19524 3896
rect 19576 3884 19582 3936
rect 19610 3884 19616 3936
rect 19668 3884 19674 3936
rect 24210 3884 24216 3936
rect 24268 3884 24274 3936
rect 24504 3924 24532 3964
rect 24581 3961 24593 3995
rect 24627 3961 24639 3995
rect 29270 3992 29276 4004
rect 24581 3955 24639 3961
rect 26252 3964 29276 3992
rect 26252 3924 26280 3964
rect 29270 3952 29276 3964
rect 29328 3952 29334 4004
rect 24504 3896 26280 3924
rect 26326 3884 26332 3936
rect 26384 3924 26390 3936
rect 27157 3927 27215 3933
rect 27157 3924 27169 3927
rect 26384 3896 27169 3924
rect 26384 3884 26390 3896
rect 27157 3893 27169 3896
rect 27203 3893 27215 3927
rect 27157 3887 27215 3893
rect 27525 3927 27583 3933
rect 27525 3893 27537 3927
rect 27571 3924 27583 3927
rect 27890 3924 27896 3936
rect 27571 3896 27896 3924
rect 27571 3893 27583 3896
rect 27525 3887 27583 3893
rect 27890 3884 27896 3896
rect 27948 3884 27954 3936
rect 28353 3927 28411 3933
rect 28353 3893 28365 3927
rect 28399 3924 28411 3927
rect 28626 3924 28632 3936
rect 28399 3896 28632 3924
rect 28399 3893 28411 3896
rect 28353 3887 28411 3893
rect 28626 3884 28632 3896
rect 28684 3884 28690 3936
rect 28994 3884 29000 3936
rect 29052 3884 29058 3936
rect 29178 3884 29184 3936
rect 29236 3884 29242 3936
rect 29380 3924 29408 4032
rect 30024 4032 31754 4060
rect 30024 3992 30052 4032
rect 29564 3964 30052 3992
rect 29564 3924 29592 3964
rect 30098 3952 30104 4004
rect 30156 3992 30162 4004
rect 30653 3995 30711 4001
rect 30653 3992 30665 3995
rect 30156 3964 30665 3992
rect 30156 3952 30162 3964
rect 30653 3961 30665 3964
rect 30699 3961 30711 3995
rect 30653 3955 30711 3961
rect 30742 3952 30748 4004
rect 30800 3992 30806 4004
rect 31389 3995 31447 4001
rect 31389 3992 31401 3995
rect 30800 3964 31401 3992
rect 30800 3952 30806 3964
rect 31389 3961 31401 3964
rect 31435 3961 31447 3995
rect 31726 3992 31754 4032
rect 35894 4020 35900 4072
rect 35952 4060 35958 4072
rect 39224 4060 39252 4091
rect 35952 4032 39252 4060
rect 35952 4020 35958 4032
rect 39206 3992 39212 4004
rect 31726 3964 39212 3992
rect 31389 3955 31447 3961
rect 39206 3952 39212 3964
rect 39264 3952 39270 4004
rect 39390 3952 39396 4004
rect 39448 3952 39454 4004
rect 29380 3896 29592 3924
rect 29822 3884 29828 3936
rect 29880 3884 29886 3936
rect 30006 3884 30012 3936
rect 30064 3884 30070 3936
rect 31018 3884 31024 3936
rect 31076 3884 31082 3936
rect 31110 3884 31116 3936
rect 31168 3884 31174 3936
rect 39022 3884 39028 3936
rect 39080 3884 39086 3936
rect 1104 3834 39836 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 37950 3834
rect 38002 3782 38014 3834
rect 38066 3782 38078 3834
rect 38130 3782 38142 3834
rect 38194 3782 38206 3834
rect 38258 3782 39836 3834
rect 1104 3760 39836 3782
rect 19150 3680 19156 3732
rect 19208 3720 19214 3732
rect 19521 3723 19579 3729
rect 19521 3720 19533 3723
rect 19208 3692 19533 3720
rect 19208 3680 19214 3692
rect 19521 3689 19533 3692
rect 19567 3689 19579 3723
rect 19521 3683 19579 3689
rect 21910 3680 21916 3732
rect 21968 3720 21974 3732
rect 22189 3723 22247 3729
rect 22189 3720 22201 3723
rect 21968 3692 22201 3720
rect 21968 3680 21974 3692
rect 22189 3689 22201 3692
rect 22235 3689 22247 3723
rect 22189 3683 22247 3689
rect 22738 3680 22744 3732
rect 22796 3720 22802 3732
rect 24302 3720 24308 3732
rect 22796 3692 24308 3720
rect 22796 3680 22802 3692
rect 24302 3680 24308 3692
rect 24360 3680 24366 3732
rect 24394 3680 24400 3732
rect 24452 3720 24458 3732
rect 25409 3723 25467 3729
rect 25409 3720 25421 3723
rect 24452 3692 25421 3720
rect 24452 3680 24458 3692
rect 25409 3689 25421 3692
rect 25455 3689 25467 3723
rect 25409 3683 25467 3689
rect 25774 3680 25780 3732
rect 25832 3680 25838 3732
rect 30190 3680 30196 3732
rect 30248 3720 30254 3732
rect 31110 3720 31116 3732
rect 30248 3692 31116 3720
rect 30248 3680 30254 3692
rect 31110 3680 31116 3692
rect 31168 3680 31174 3732
rect 566 3612 572 3664
rect 624 3652 630 3664
rect 19426 3652 19432 3664
rect 624 3624 19432 3652
rect 624 3612 630 3624
rect 19426 3612 19432 3624
rect 19484 3612 19490 3664
rect 20714 3612 20720 3664
rect 20772 3652 20778 3664
rect 22830 3652 22836 3664
rect 20772 3624 22836 3652
rect 20772 3612 20778 3624
rect 22830 3612 22836 3624
rect 22888 3612 22894 3664
rect 23106 3612 23112 3664
rect 23164 3652 23170 3664
rect 23661 3655 23719 3661
rect 23661 3652 23673 3655
rect 23164 3624 23673 3652
rect 23164 3612 23170 3624
rect 23661 3621 23673 3624
rect 23707 3621 23719 3655
rect 23661 3615 23719 3621
rect 24581 3655 24639 3661
rect 24581 3621 24593 3655
rect 24627 3621 24639 3655
rect 24581 3615 24639 3621
rect 25133 3655 25191 3661
rect 25133 3621 25145 3655
rect 25179 3652 25191 3655
rect 38838 3652 38844 3664
rect 25179 3624 38844 3652
rect 25179 3621 25191 3624
rect 25133 3615 25191 3621
rect 17126 3544 17132 3596
rect 17184 3584 17190 3596
rect 24213 3587 24271 3593
rect 17184 3556 23428 3584
rect 17184 3544 17190 3556
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 18230 3516 18236 3528
rect 11112 3488 18236 3516
rect 11112 3476 11118 3488
rect 18230 3476 18236 3488
rect 18288 3476 18294 3528
rect 18325 3519 18383 3525
rect 18325 3485 18337 3519
rect 18371 3516 18383 3519
rect 18417 3519 18475 3525
rect 18417 3516 18429 3519
rect 18371 3488 18429 3516
rect 18371 3485 18383 3488
rect 18325 3479 18383 3485
rect 18417 3485 18429 3488
rect 18463 3485 18475 3519
rect 18417 3479 18475 3485
rect 18506 3476 18512 3528
rect 18564 3516 18570 3528
rect 18693 3519 18751 3525
rect 18693 3516 18705 3519
rect 18564 3488 18705 3516
rect 18564 3476 18570 3488
rect 18693 3485 18705 3488
rect 18739 3485 18751 3519
rect 18693 3479 18751 3485
rect 19150 3476 19156 3528
rect 19208 3516 19214 3528
rect 19245 3519 19303 3525
rect 19245 3516 19257 3519
rect 19208 3488 19257 3516
rect 19208 3476 19214 3488
rect 19245 3485 19257 3488
rect 19291 3485 19303 3519
rect 19245 3479 19303 3485
rect 19518 3476 19524 3528
rect 19576 3516 19582 3528
rect 19576 3488 19748 3516
rect 19576 3476 19582 3488
rect 9674 3408 9680 3460
rect 9732 3448 9738 3460
rect 19610 3448 19616 3460
rect 9732 3420 19616 3448
rect 9732 3408 9738 3420
rect 19610 3408 19616 3420
rect 19668 3408 19674 3460
rect 19720 3448 19748 3488
rect 21726 3476 21732 3528
rect 21784 3476 21790 3528
rect 22281 3519 22339 3525
rect 22281 3485 22293 3519
rect 22327 3516 22339 3519
rect 22373 3519 22431 3525
rect 22373 3516 22385 3519
rect 22327 3488 22385 3516
rect 22327 3485 22339 3488
rect 22281 3479 22339 3485
rect 22373 3485 22385 3488
rect 22419 3485 22431 3519
rect 22373 3479 22431 3485
rect 22741 3519 22799 3525
rect 22741 3485 22753 3519
rect 22787 3516 22799 3519
rect 22833 3519 22891 3525
rect 22833 3516 22845 3519
rect 22787 3488 22845 3516
rect 22787 3485 22799 3488
rect 22741 3479 22799 3485
rect 22833 3485 22845 3488
rect 22879 3485 22891 3519
rect 22833 3479 22891 3485
rect 23106 3476 23112 3528
rect 23164 3476 23170 3528
rect 23400 3525 23428 3556
rect 24213 3553 24225 3587
rect 24259 3584 24271 3587
rect 24596 3584 24624 3615
rect 38838 3612 38844 3624
rect 38896 3612 38902 3664
rect 39390 3612 39396 3664
rect 39448 3612 39454 3664
rect 24259 3556 24532 3584
rect 24596 3556 31754 3584
rect 24259 3553 24271 3556
rect 24213 3547 24271 3553
rect 23385 3519 23443 3525
rect 23385 3485 23397 3519
rect 23431 3516 23443 3519
rect 23845 3519 23903 3525
rect 23845 3516 23857 3519
rect 23431 3488 23857 3516
rect 23431 3485 23443 3488
rect 23385 3479 23443 3485
rect 23845 3485 23857 3488
rect 23891 3485 23903 3519
rect 23845 3479 23903 3485
rect 24394 3476 24400 3528
rect 24452 3476 24458 3528
rect 24504 3516 24532 3556
rect 24673 3519 24731 3525
rect 24673 3516 24685 3519
rect 24504 3488 24685 3516
rect 24673 3485 24685 3488
rect 24719 3485 24731 3519
rect 24673 3479 24731 3485
rect 24946 3476 24952 3528
rect 25004 3516 25010 3528
rect 25225 3519 25283 3525
rect 25225 3516 25237 3519
rect 25004 3488 25237 3516
rect 25004 3476 25010 3488
rect 25225 3485 25237 3488
rect 25271 3485 25283 3519
rect 25225 3479 25283 3485
rect 25593 3519 25651 3525
rect 25593 3485 25605 3519
rect 25639 3516 25651 3519
rect 26142 3516 26148 3528
rect 25639 3488 26148 3516
rect 25639 3485 25651 3488
rect 25593 3479 25651 3485
rect 26142 3476 26148 3488
rect 26200 3476 26206 3528
rect 26510 3476 26516 3528
rect 26568 3476 26574 3528
rect 29914 3476 29920 3528
rect 29972 3516 29978 3528
rect 31018 3516 31024 3528
rect 29972 3488 31024 3516
rect 29972 3476 29978 3488
rect 31018 3476 31024 3488
rect 31076 3476 31082 3528
rect 31726 3516 31754 3556
rect 38841 3519 38899 3525
rect 38841 3516 38853 3519
rect 31726 3488 38853 3516
rect 38841 3485 38853 3488
rect 38887 3485 38899 3519
rect 38841 3479 38899 3485
rect 39206 3476 39212 3528
rect 39264 3476 39270 3528
rect 23474 3448 23480 3460
rect 19720 3420 23480 3448
rect 23474 3408 23480 3420
rect 23532 3408 23538 3460
rect 24762 3448 24768 3460
rect 23584 3420 24768 3448
rect 18230 3340 18236 3392
rect 18288 3340 18294 3392
rect 18598 3340 18604 3392
rect 18656 3340 18662 3392
rect 18877 3383 18935 3389
rect 18877 3349 18889 3383
rect 18923 3380 18935 3383
rect 19334 3380 19340 3392
rect 18923 3352 19340 3380
rect 18923 3349 18935 3352
rect 18877 3343 18935 3349
rect 19334 3340 19340 3352
rect 19392 3340 19398 3392
rect 19426 3340 19432 3392
rect 19484 3340 19490 3392
rect 21910 3340 21916 3392
rect 21968 3340 21974 3392
rect 22554 3340 22560 3392
rect 22612 3340 22618 3392
rect 22646 3340 22652 3392
rect 22704 3340 22710 3392
rect 23014 3340 23020 3392
rect 23072 3340 23078 3392
rect 23198 3340 23204 3392
rect 23256 3380 23262 3392
rect 23584 3389 23612 3420
rect 24762 3408 24768 3420
rect 24820 3408 24826 3460
rect 38930 3448 38936 3460
rect 24872 3420 38936 3448
rect 23293 3383 23351 3389
rect 23293 3380 23305 3383
rect 23256 3352 23305 3380
rect 23256 3340 23262 3352
rect 23293 3349 23305 3352
rect 23339 3349 23351 3383
rect 23293 3343 23351 3349
rect 23569 3383 23627 3389
rect 23569 3349 23581 3383
rect 23615 3349 23627 3383
rect 23569 3343 23627 3349
rect 24118 3340 24124 3392
rect 24176 3340 24182 3392
rect 24872 3389 24900 3420
rect 38930 3408 38936 3420
rect 38988 3408 38994 3460
rect 24857 3383 24915 3389
rect 24857 3349 24869 3383
rect 24903 3349 24915 3383
rect 24857 3343 24915 3349
rect 26697 3383 26755 3389
rect 26697 3349 26709 3383
rect 26743 3380 26755 3383
rect 32582 3380 32588 3392
rect 26743 3352 32588 3380
rect 26743 3349 26755 3352
rect 26697 3343 26755 3349
rect 32582 3340 32588 3352
rect 32640 3340 32646 3392
rect 39025 3383 39083 3389
rect 39025 3349 39037 3383
rect 39071 3380 39083 3383
rect 39942 3380 39948 3392
rect 39071 3352 39948 3380
rect 39071 3349 39083 3352
rect 39025 3343 39083 3349
rect 39942 3340 39948 3352
rect 40000 3340 40006 3392
rect 1104 3290 39836 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 39010 3290
rect 39062 3238 39074 3290
rect 39126 3238 39138 3290
rect 39190 3238 39202 3290
rect 39254 3238 39266 3290
rect 39318 3238 39836 3290
rect 1104 3216 39836 3238
rect 8846 3136 8852 3188
rect 8904 3176 8910 3188
rect 18230 3176 18236 3188
rect 8904 3148 18236 3176
rect 8904 3136 8910 3148
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 18598 3136 18604 3188
rect 18656 3176 18662 3188
rect 23290 3176 23296 3188
rect 18656 3148 23296 3176
rect 18656 3136 18662 3148
rect 23290 3136 23296 3148
rect 23348 3136 23354 3188
rect 23382 3136 23388 3188
rect 23440 3176 23446 3188
rect 23753 3179 23811 3185
rect 23753 3176 23765 3179
rect 23440 3148 23765 3176
rect 23440 3136 23446 3148
rect 23753 3145 23765 3148
rect 23799 3145 23811 3179
rect 23753 3139 23811 3145
rect 24302 3136 24308 3188
rect 24360 3176 24366 3188
rect 24360 3148 24716 3176
rect 24360 3136 24366 3148
rect 4890 3068 4896 3120
rect 4948 3108 4954 3120
rect 4948 3080 19104 3108
rect 4948 3068 4954 3080
rect 17954 3000 17960 3052
rect 18012 3040 18018 3052
rect 18233 3043 18291 3049
rect 18233 3040 18245 3043
rect 18012 3012 18245 3040
rect 18012 3000 18018 3012
rect 18233 3009 18245 3012
rect 18279 3009 18291 3043
rect 18233 3003 18291 3009
rect 18322 3000 18328 3052
rect 18380 3040 18386 3052
rect 18782 3040 18788 3052
rect 18380 3012 18788 3040
rect 18380 3000 18386 3012
rect 18782 3000 18788 3012
rect 18840 3000 18846 3052
rect 19076 3049 19104 3080
rect 19334 3068 19340 3120
rect 19392 3108 19398 3120
rect 22738 3108 22744 3120
rect 19392 3080 22744 3108
rect 19392 3068 19398 3080
rect 22738 3068 22744 3080
rect 22796 3068 22802 3120
rect 22830 3068 22836 3120
rect 22888 3108 22894 3120
rect 24688 3108 24716 3148
rect 24762 3136 24768 3188
rect 24820 3176 24826 3188
rect 24820 3148 38516 3176
rect 24820 3136 24826 3148
rect 28442 3108 28448 3120
rect 22888 3080 24624 3108
rect 24688 3080 28448 3108
rect 22888 3068 22894 3080
rect 19061 3043 19119 3049
rect 19061 3009 19073 3043
rect 19107 3009 19119 3043
rect 19061 3003 19119 3009
rect 19610 3000 19616 3052
rect 19668 3000 19674 3052
rect 24596 3049 24624 3080
rect 28442 3068 28448 3080
rect 28500 3068 28506 3120
rect 32398 3108 32404 3120
rect 30392 3080 32404 3108
rect 23201 3043 23259 3049
rect 23201 3040 23213 3043
rect 22066 3012 23213 3040
rect 11974 2932 11980 2984
rect 12032 2972 12038 2984
rect 22066 2972 22094 3012
rect 23201 3009 23213 3012
rect 23247 3009 23259 3043
rect 23569 3043 23627 3049
rect 23569 3040 23581 3043
rect 23201 3003 23259 3009
rect 23308 3012 23581 3040
rect 12032 2944 22094 2972
rect 12032 2932 12038 2944
rect 22462 2932 22468 2984
rect 22520 2972 22526 2984
rect 23308 2972 23336 3012
rect 23569 3009 23581 3012
rect 23615 3009 23627 3043
rect 23569 3003 23627 3009
rect 24581 3043 24639 3049
rect 24581 3009 24593 3043
rect 24627 3009 24639 3043
rect 24581 3003 24639 3009
rect 24854 3000 24860 3052
rect 24912 3040 24918 3052
rect 25685 3043 25743 3049
rect 25685 3040 25697 3043
rect 24912 3012 25697 3040
rect 24912 3000 24918 3012
rect 25685 3009 25697 3012
rect 25731 3009 25743 3043
rect 25685 3003 25743 3009
rect 25866 3000 25872 3052
rect 25924 3040 25930 3052
rect 26053 3043 26111 3049
rect 26053 3040 26065 3043
rect 25924 3012 26065 3040
rect 25924 3000 25930 3012
rect 26053 3009 26065 3012
rect 26099 3009 26111 3043
rect 26053 3003 26111 3009
rect 26973 3043 27031 3049
rect 26973 3009 26985 3043
rect 27019 3009 27031 3043
rect 26973 3003 27031 3009
rect 22520 2944 23336 2972
rect 22520 2932 22526 2944
rect 23474 2932 23480 2984
rect 23532 2972 23538 2984
rect 26988 2972 27016 3003
rect 27890 3000 27896 3052
rect 27948 3000 27954 3052
rect 28721 3043 28779 3049
rect 28721 3009 28733 3043
rect 28767 3040 28779 3043
rect 29178 3040 29184 3052
rect 28767 3012 29184 3040
rect 28767 3009 28779 3012
rect 28721 3003 28779 3009
rect 29178 3000 29184 3012
rect 29236 3000 29242 3052
rect 29273 3043 29331 3049
rect 29273 3009 29285 3043
rect 29319 3040 29331 3043
rect 30098 3040 30104 3052
rect 29319 3012 30104 3040
rect 29319 3009 29331 3012
rect 29273 3003 29331 3009
rect 30098 3000 30104 3012
rect 30156 3000 30162 3052
rect 30392 3049 30420 3080
rect 32398 3068 32404 3080
rect 32456 3068 32462 3120
rect 30377 3043 30435 3049
rect 30377 3009 30389 3043
rect 30423 3009 30435 3043
rect 30377 3003 30435 3009
rect 30834 3000 30840 3052
rect 30892 3040 30898 3052
rect 30929 3043 30987 3049
rect 30929 3040 30941 3043
rect 30892 3012 30941 3040
rect 30892 3000 30898 3012
rect 30929 3009 30941 3012
rect 30975 3009 30987 3043
rect 30929 3003 30987 3009
rect 31294 3000 31300 3052
rect 31352 3000 31358 3052
rect 38488 3049 38516 3148
rect 39390 3136 39396 3188
rect 39448 3136 39454 3188
rect 38473 3043 38531 3049
rect 38473 3009 38485 3043
rect 38519 3009 38531 3043
rect 38473 3003 38531 3009
rect 38838 3000 38844 3052
rect 38896 3000 38902 3052
rect 38930 3000 38936 3052
rect 38988 3040 38994 3052
rect 39209 3043 39267 3049
rect 39209 3040 39221 3043
rect 38988 3012 39221 3040
rect 38988 3000 38994 3012
rect 39209 3009 39221 3012
rect 39255 3009 39267 3043
rect 39209 3003 39267 3009
rect 23532 2944 27016 2972
rect 23532 2932 23538 2944
rect 9582 2864 9588 2916
rect 9640 2904 9646 2916
rect 22646 2904 22652 2916
rect 9640 2876 22652 2904
rect 9640 2864 9646 2876
rect 22646 2864 22652 2876
rect 22704 2864 22710 2916
rect 23290 2864 23296 2916
rect 23348 2904 23354 2916
rect 25498 2904 25504 2916
rect 23348 2876 25504 2904
rect 23348 2864 23354 2876
rect 25498 2864 25504 2876
rect 25556 2864 25562 2916
rect 26142 2864 26148 2916
rect 26200 2904 26206 2916
rect 27706 2904 27712 2916
rect 26200 2876 27712 2904
rect 26200 2864 26206 2876
rect 27706 2864 27712 2876
rect 27764 2864 27770 2916
rect 38657 2907 38715 2913
rect 38657 2873 38669 2907
rect 38703 2904 38715 2907
rect 40402 2904 40408 2916
rect 38703 2876 40408 2904
rect 38703 2873 38715 2876
rect 38657 2867 38715 2873
rect 40402 2864 40408 2876
rect 40460 2864 40466 2916
rect 18138 2796 18144 2848
rect 18196 2836 18202 2848
rect 18417 2839 18475 2845
rect 18417 2836 18429 2839
rect 18196 2808 18429 2836
rect 18196 2796 18202 2808
rect 18417 2805 18429 2808
rect 18463 2805 18475 2839
rect 18417 2799 18475 2805
rect 18966 2796 18972 2848
rect 19024 2836 19030 2848
rect 19245 2839 19303 2845
rect 19245 2836 19257 2839
rect 19024 2808 19257 2836
rect 19024 2796 19030 2808
rect 19245 2805 19257 2808
rect 19291 2805 19303 2839
rect 19245 2799 19303 2805
rect 19518 2796 19524 2848
rect 19576 2836 19582 2848
rect 19797 2839 19855 2845
rect 19797 2836 19809 2839
rect 19576 2808 19809 2836
rect 19576 2796 19582 2808
rect 19797 2805 19809 2808
rect 19843 2805 19855 2839
rect 19797 2799 19855 2805
rect 23106 2796 23112 2848
rect 23164 2836 23170 2848
rect 23385 2839 23443 2845
rect 23385 2836 23397 2839
rect 23164 2808 23397 2836
rect 23164 2796 23170 2808
rect 23385 2805 23397 2808
rect 23431 2805 23443 2839
rect 23385 2799 23443 2805
rect 23474 2796 23480 2848
rect 23532 2836 23538 2848
rect 23658 2836 23664 2848
rect 23532 2808 23664 2836
rect 23532 2796 23538 2808
rect 23658 2796 23664 2808
rect 23716 2796 23722 2848
rect 24486 2796 24492 2848
rect 24544 2836 24550 2848
rect 24765 2839 24823 2845
rect 24765 2836 24777 2839
rect 24544 2808 24777 2836
rect 24544 2796 24550 2808
rect 24765 2805 24777 2808
rect 24811 2805 24823 2839
rect 24765 2799 24823 2805
rect 25590 2796 25596 2848
rect 25648 2836 25654 2848
rect 25869 2839 25927 2845
rect 25869 2836 25881 2839
rect 25648 2808 25881 2836
rect 25648 2796 25654 2808
rect 25869 2805 25881 2808
rect 25915 2805 25927 2839
rect 25869 2799 25927 2805
rect 26237 2839 26295 2845
rect 26237 2805 26249 2839
rect 26283 2836 26295 2839
rect 26326 2836 26332 2848
rect 26283 2808 26332 2836
rect 26283 2805 26295 2808
rect 26237 2799 26295 2805
rect 26326 2796 26332 2808
rect 26384 2796 26390 2848
rect 26694 2796 26700 2848
rect 26752 2836 26758 2848
rect 27157 2839 27215 2845
rect 27157 2836 27169 2839
rect 26752 2808 27169 2836
rect 26752 2796 26758 2808
rect 27157 2805 27169 2808
rect 27203 2805 27215 2839
rect 27157 2799 27215 2805
rect 27798 2796 27804 2848
rect 27856 2836 27862 2848
rect 28077 2839 28135 2845
rect 28077 2836 28089 2839
rect 27856 2808 28089 2836
rect 27856 2796 27862 2808
rect 28077 2805 28089 2808
rect 28123 2805 28135 2839
rect 28077 2799 28135 2805
rect 28350 2796 28356 2848
rect 28408 2836 28414 2848
rect 28537 2839 28595 2845
rect 28537 2836 28549 2839
rect 28408 2808 28549 2836
rect 28408 2796 28414 2808
rect 28537 2805 28549 2808
rect 28583 2805 28595 2839
rect 28537 2799 28595 2805
rect 28902 2796 28908 2848
rect 28960 2836 28966 2848
rect 29089 2839 29147 2845
rect 29089 2836 29101 2839
rect 28960 2808 29101 2836
rect 28960 2796 28966 2808
rect 29089 2805 29101 2808
rect 29135 2805 29147 2839
rect 29089 2799 29147 2805
rect 30098 2796 30104 2848
rect 30156 2836 30162 2848
rect 30193 2839 30251 2845
rect 30193 2836 30205 2839
rect 30156 2808 30205 2836
rect 30156 2796 30162 2808
rect 30193 2805 30205 2808
rect 30239 2805 30251 2839
rect 30193 2799 30251 2805
rect 30834 2796 30840 2848
rect 30892 2836 30898 2848
rect 31113 2839 31171 2845
rect 31113 2836 31125 2839
rect 30892 2808 31125 2836
rect 30892 2796 30898 2808
rect 31113 2805 31125 2808
rect 31159 2805 31171 2839
rect 31113 2799 31171 2805
rect 31202 2796 31208 2848
rect 31260 2836 31266 2848
rect 31481 2839 31539 2845
rect 31481 2836 31493 2839
rect 31260 2808 31493 2836
rect 31260 2796 31266 2808
rect 31481 2805 31493 2808
rect 31527 2805 31539 2839
rect 31481 2799 31539 2805
rect 39022 2796 39028 2848
rect 39080 2796 39086 2848
rect 1104 2746 39836 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 37950 2746
rect 38002 2694 38014 2746
rect 38066 2694 38078 2746
rect 38130 2694 38142 2746
rect 38194 2694 38206 2746
rect 38258 2694 39836 2746
rect 1104 2672 39836 2694
rect 7742 2592 7748 2644
rect 7800 2632 7806 2644
rect 8202 2632 8208 2644
rect 7800 2604 8208 2632
rect 7800 2592 7806 2604
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 10962 2592 10968 2644
rect 11020 2632 11026 2644
rect 13722 2632 13728 2644
rect 11020 2604 13728 2632
rect 11020 2592 11026 2604
rect 13722 2592 13728 2604
rect 13780 2592 13786 2644
rect 21174 2632 21180 2644
rect 17236 2604 21180 2632
rect 10594 2524 10600 2576
rect 10652 2564 10658 2576
rect 17236 2564 17264 2604
rect 21174 2592 21180 2604
rect 21232 2592 21238 2644
rect 22002 2592 22008 2644
rect 22060 2632 22066 2644
rect 22186 2632 22192 2644
rect 22060 2604 22192 2632
rect 22060 2592 22066 2604
rect 22186 2592 22192 2604
rect 22244 2592 22250 2644
rect 22554 2592 22560 2644
rect 22612 2632 22618 2644
rect 23477 2635 23535 2641
rect 23477 2632 23489 2635
rect 22612 2604 23489 2632
rect 22612 2592 22618 2604
rect 23477 2601 23489 2604
rect 23523 2601 23535 2635
rect 23477 2595 23535 2601
rect 24210 2592 24216 2644
rect 24268 2632 24274 2644
rect 25317 2635 25375 2641
rect 25317 2632 25329 2635
rect 24268 2604 25329 2632
rect 24268 2592 24274 2604
rect 25317 2601 25329 2604
rect 25363 2601 25375 2635
rect 25317 2595 25375 2601
rect 25406 2592 25412 2644
rect 25464 2632 25470 2644
rect 25464 2604 27292 2632
rect 25464 2592 25470 2604
rect 10652 2536 17264 2564
rect 10652 2524 10658 2536
rect 18322 2524 18328 2576
rect 18380 2564 18386 2576
rect 20070 2564 20076 2576
rect 18380 2536 20076 2564
rect 18380 2524 18386 2536
rect 20070 2524 20076 2536
rect 20128 2524 20134 2576
rect 21100 2536 21312 2564
rect 10226 2456 10232 2508
rect 10284 2496 10290 2508
rect 21100 2496 21128 2536
rect 10284 2468 21128 2496
rect 21284 2496 21312 2536
rect 21726 2524 21732 2576
rect 21784 2564 21790 2576
rect 22373 2567 22431 2573
rect 22373 2564 22385 2567
rect 21784 2536 22385 2564
rect 21784 2524 21790 2536
rect 22373 2533 22385 2536
rect 22419 2533 22431 2567
rect 22373 2527 22431 2533
rect 22462 2524 22468 2576
rect 22520 2564 22526 2576
rect 23109 2567 23167 2573
rect 23109 2564 23121 2567
rect 22520 2536 23121 2564
rect 22520 2524 22526 2536
rect 23109 2533 23121 2536
rect 23155 2533 23167 2567
rect 23109 2527 23167 2533
rect 23658 2524 23664 2576
rect 23716 2564 23722 2576
rect 24581 2567 24639 2573
rect 24581 2564 24593 2567
rect 23716 2536 24593 2564
rect 23716 2524 23722 2536
rect 24581 2533 24593 2536
rect 24627 2533 24639 2567
rect 24581 2527 24639 2533
rect 24762 2524 24768 2576
rect 24820 2564 24826 2576
rect 25685 2567 25743 2573
rect 25685 2564 25697 2567
rect 24820 2536 25697 2564
rect 24820 2524 24826 2536
rect 25685 2533 25697 2536
rect 25731 2533 25743 2567
rect 27157 2567 27215 2573
rect 27157 2564 27169 2567
rect 25685 2527 25743 2533
rect 26436 2536 27169 2564
rect 21284 2468 22968 2496
rect 10284 2456 10290 2468
rect 16666 2388 16672 2440
rect 16724 2428 16730 2440
rect 17681 2431 17739 2437
rect 17681 2428 17693 2431
rect 16724 2400 17693 2428
rect 16724 2388 16730 2400
rect 17681 2397 17693 2400
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 17770 2388 17776 2440
rect 17828 2428 17834 2440
rect 18049 2431 18107 2437
rect 18049 2428 18061 2431
rect 17828 2400 18061 2428
rect 17828 2388 17834 2400
rect 18049 2397 18061 2400
rect 18095 2397 18107 2431
rect 18049 2391 18107 2397
rect 18417 2431 18475 2437
rect 18417 2397 18429 2431
rect 18463 2397 18475 2431
rect 18417 2391 18475 2397
rect 10870 2320 10876 2372
rect 10928 2360 10934 2372
rect 18432 2360 18460 2391
rect 18690 2388 18696 2440
rect 18748 2388 18754 2440
rect 18782 2388 18788 2440
rect 18840 2388 18846 2440
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 19702 2388 19708 2440
rect 19760 2428 19766 2440
rect 19797 2431 19855 2437
rect 19797 2428 19809 2431
rect 19760 2400 19809 2428
rect 19760 2388 19766 2400
rect 19797 2397 19809 2400
rect 19843 2397 19855 2431
rect 19797 2391 19855 2397
rect 20165 2431 20223 2437
rect 20165 2397 20177 2431
rect 20211 2397 20223 2431
rect 20165 2391 20223 2397
rect 10928 2332 18460 2360
rect 18708 2360 18736 2388
rect 20180 2360 20208 2391
rect 20254 2388 20260 2440
rect 20312 2428 20318 2440
rect 20533 2431 20591 2437
rect 20533 2428 20545 2431
rect 20312 2400 20545 2428
rect 20312 2388 20318 2400
rect 20533 2397 20545 2400
rect 20579 2397 20591 2431
rect 20533 2391 20591 2397
rect 20714 2388 20720 2440
rect 20772 2428 20778 2440
rect 20901 2431 20959 2437
rect 20901 2428 20913 2431
rect 20772 2400 20913 2428
rect 20772 2388 20778 2400
rect 20901 2397 20913 2400
rect 20947 2397 20959 2431
rect 20901 2391 20959 2397
rect 21269 2431 21327 2437
rect 21269 2397 21281 2431
rect 21315 2428 21327 2431
rect 21358 2428 21364 2440
rect 21315 2400 21364 2428
rect 21315 2397 21327 2400
rect 21269 2391 21327 2397
rect 21358 2388 21364 2400
rect 21416 2388 21422 2440
rect 21818 2388 21824 2440
rect 21876 2388 21882 2440
rect 22189 2431 22247 2437
rect 22189 2397 22201 2431
rect 22235 2428 22247 2431
rect 22278 2428 22284 2440
rect 22235 2400 22284 2428
rect 22235 2397 22247 2400
rect 22189 2391 22247 2397
rect 22278 2388 22284 2400
rect 22336 2388 22342 2440
rect 22370 2388 22376 2440
rect 22428 2428 22434 2440
rect 22940 2437 22968 2468
rect 24854 2456 24860 2508
rect 24912 2496 24918 2508
rect 24912 2468 25636 2496
rect 24912 2456 24918 2468
rect 22557 2431 22615 2437
rect 22557 2428 22569 2431
rect 22428 2400 22569 2428
rect 22428 2388 22434 2400
rect 22557 2397 22569 2400
rect 22603 2397 22615 2431
rect 22557 2391 22615 2397
rect 22925 2431 22983 2437
rect 22925 2397 22937 2431
rect 22971 2397 22983 2431
rect 22925 2391 22983 2397
rect 23293 2431 23351 2437
rect 23293 2397 23305 2431
rect 23339 2397 23351 2431
rect 23293 2391 23351 2397
rect 18708 2332 20208 2360
rect 10928 2320 10934 2332
rect 21174 2320 21180 2372
rect 21232 2360 21238 2372
rect 23308 2360 23336 2391
rect 23566 2388 23572 2440
rect 23624 2428 23630 2440
rect 23661 2431 23719 2437
rect 23661 2428 23673 2431
rect 23624 2400 23673 2428
rect 23624 2388 23630 2400
rect 23661 2397 23673 2400
rect 23707 2397 23719 2431
rect 23661 2391 23719 2397
rect 24394 2388 24400 2440
rect 24452 2388 24458 2440
rect 24578 2388 24584 2440
rect 24636 2428 24642 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 24636 2400 24777 2428
rect 24636 2388 24642 2400
rect 24765 2397 24777 2400
rect 24811 2397 24823 2431
rect 24765 2391 24823 2397
rect 25130 2388 25136 2440
rect 25188 2388 25194 2440
rect 25222 2388 25228 2440
rect 25280 2428 25286 2440
rect 25501 2431 25559 2437
rect 25501 2428 25513 2431
rect 25280 2400 25513 2428
rect 25280 2388 25286 2400
rect 25501 2397 25513 2400
rect 25547 2397 25559 2431
rect 25608 2428 25636 2468
rect 26142 2456 26148 2508
rect 26200 2496 26206 2508
rect 26436 2496 26464 2536
rect 27157 2533 27169 2536
rect 27203 2533 27215 2567
rect 27264 2564 27292 2604
rect 27614 2592 27620 2644
rect 27672 2632 27678 2644
rect 28261 2635 28319 2641
rect 28261 2632 28273 2635
rect 27672 2604 28273 2632
rect 27672 2592 27678 2604
rect 28261 2601 28273 2604
rect 28307 2601 28319 2635
rect 28261 2595 28319 2601
rect 29730 2592 29736 2644
rect 29788 2632 29794 2644
rect 30745 2635 30803 2641
rect 30745 2632 30757 2635
rect 29788 2604 30757 2632
rect 29788 2592 29794 2604
rect 30745 2601 30757 2604
rect 30791 2601 30803 2635
rect 30745 2595 30803 2601
rect 31018 2592 31024 2644
rect 31076 2632 31082 2644
rect 31386 2632 31392 2644
rect 31076 2604 31392 2632
rect 31076 2592 31082 2604
rect 31386 2592 31392 2604
rect 31444 2592 31450 2644
rect 27264 2536 27752 2564
rect 27157 2527 27215 2533
rect 27430 2496 27436 2508
rect 26200 2468 26464 2496
rect 27356 2468 27436 2496
rect 26200 2456 26206 2468
rect 25869 2431 25927 2437
rect 25869 2428 25881 2431
rect 25608 2400 25881 2428
rect 25501 2391 25559 2397
rect 25869 2397 25881 2400
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 26050 2388 26056 2440
rect 26108 2428 26114 2440
rect 27356 2437 27384 2468
rect 27430 2456 27436 2468
rect 27488 2456 27494 2508
rect 27724 2437 27752 2536
rect 28074 2524 28080 2576
rect 28132 2564 28138 2576
rect 28997 2567 29055 2573
rect 28997 2564 29009 2567
rect 28132 2536 29009 2564
rect 28132 2524 28138 2536
rect 28997 2533 29009 2536
rect 29043 2533 29055 2567
rect 28997 2527 29055 2533
rect 29178 2524 29184 2576
rect 29236 2564 29242 2576
rect 30009 2567 30067 2573
rect 30009 2564 30021 2567
rect 29236 2536 30021 2564
rect 29236 2524 29242 2536
rect 30009 2533 30021 2536
rect 30055 2533 30067 2567
rect 30009 2527 30067 2533
rect 30282 2524 30288 2576
rect 30340 2564 30346 2576
rect 31113 2567 31171 2573
rect 31113 2564 31125 2567
rect 30340 2536 31125 2564
rect 30340 2524 30346 2536
rect 31113 2533 31125 2536
rect 31159 2533 31171 2567
rect 31113 2527 31171 2533
rect 31478 2524 31484 2576
rect 31536 2564 31542 2576
rect 32309 2567 32367 2573
rect 32309 2564 32321 2567
rect 31536 2536 32321 2564
rect 31536 2524 31542 2536
rect 32309 2533 32321 2536
rect 32355 2533 32367 2567
rect 32309 2527 32367 2533
rect 39390 2524 39396 2576
rect 39448 2524 39454 2576
rect 31754 2496 31760 2508
rect 31312 2468 31760 2496
rect 26237 2431 26295 2437
rect 26237 2428 26249 2431
rect 26108 2400 26249 2428
rect 26108 2388 26114 2400
rect 26237 2397 26249 2400
rect 26283 2397 26295 2431
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26237 2391 26295 2397
rect 26344 2400 26985 2428
rect 21232 2332 23336 2360
rect 21232 2320 21238 2332
rect 24302 2320 24308 2372
rect 24360 2360 24366 2372
rect 26344 2360 26372 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 27347 2431 27405 2437
rect 27347 2397 27359 2431
rect 27393 2397 27405 2431
rect 27347 2391 27405 2397
rect 27709 2431 27767 2437
rect 27709 2397 27721 2431
rect 27755 2397 27767 2431
rect 27709 2391 27767 2397
rect 27890 2388 27896 2440
rect 27948 2428 27954 2440
rect 28077 2431 28135 2437
rect 27948 2400 28028 2428
rect 27948 2388 27954 2400
rect 24360 2332 25084 2360
rect 24360 2320 24366 2332
rect 17862 2252 17868 2304
rect 17920 2252 17926 2304
rect 18233 2295 18291 2301
rect 18233 2261 18245 2295
rect 18279 2292 18291 2295
rect 18414 2292 18420 2304
rect 18279 2264 18420 2292
rect 18279 2261 18291 2264
rect 18233 2255 18291 2261
rect 18414 2252 18420 2264
rect 18472 2252 18478 2304
rect 18601 2295 18659 2301
rect 18601 2261 18613 2295
rect 18647 2292 18659 2295
rect 18690 2292 18696 2304
rect 18647 2264 18696 2292
rect 18647 2261 18659 2264
rect 18601 2255 18659 2261
rect 18690 2252 18696 2264
rect 18748 2252 18754 2304
rect 18969 2295 19027 2301
rect 18969 2261 18981 2295
rect 19015 2292 19027 2295
rect 19242 2292 19248 2304
rect 19015 2264 19248 2292
rect 19015 2261 19027 2264
rect 18969 2255 19027 2261
rect 19242 2252 19248 2264
rect 19300 2252 19306 2304
rect 19613 2295 19671 2301
rect 19613 2261 19625 2295
rect 19659 2292 19671 2295
rect 19794 2292 19800 2304
rect 19659 2264 19800 2292
rect 19659 2261 19671 2264
rect 19613 2255 19671 2261
rect 19794 2252 19800 2264
rect 19852 2252 19858 2304
rect 19981 2295 20039 2301
rect 19981 2261 19993 2295
rect 20027 2292 20039 2295
rect 20070 2292 20076 2304
rect 20027 2264 20076 2292
rect 20027 2261 20039 2264
rect 19981 2255 20039 2261
rect 20070 2252 20076 2264
rect 20128 2252 20134 2304
rect 20346 2252 20352 2304
rect 20404 2252 20410 2304
rect 20622 2252 20628 2304
rect 20680 2292 20686 2304
rect 20717 2295 20775 2301
rect 20717 2292 20729 2295
rect 20680 2264 20729 2292
rect 20680 2252 20686 2264
rect 20717 2261 20729 2264
rect 20763 2261 20775 2295
rect 20717 2255 20775 2261
rect 20898 2252 20904 2304
rect 20956 2292 20962 2304
rect 21085 2295 21143 2301
rect 21085 2292 21097 2295
rect 20956 2264 21097 2292
rect 20956 2252 20962 2264
rect 21085 2261 21097 2264
rect 21131 2261 21143 2295
rect 21085 2255 21143 2261
rect 21358 2252 21364 2304
rect 21416 2292 21422 2304
rect 21453 2295 21511 2301
rect 21453 2292 21465 2295
rect 21416 2264 21465 2292
rect 21416 2252 21422 2264
rect 21453 2261 21465 2264
rect 21499 2261 21511 2295
rect 21453 2255 21511 2261
rect 21542 2252 21548 2304
rect 21600 2292 21606 2304
rect 22005 2295 22063 2301
rect 22005 2292 22017 2295
rect 21600 2264 22017 2292
rect 21600 2252 21606 2264
rect 22005 2261 22017 2264
rect 22051 2261 22063 2295
rect 22005 2255 22063 2261
rect 22186 2252 22192 2304
rect 22244 2292 22250 2304
rect 22741 2295 22799 2301
rect 22741 2292 22753 2295
rect 22244 2264 22753 2292
rect 22244 2252 22250 2264
rect 22741 2261 22753 2264
rect 22787 2261 22799 2295
rect 22741 2255 22799 2261
rect 22830 2252 22836 2304
rect 22888 2292 22894 2304
rect 23845 2295 23903 2301
rect 23845 2292 23857 2295
rect 22888 2264 23857 2292
rect 22888 2252 22894 2264
rect 23845 2261 23857 2264
rect 23891 2261 23903 2295
rect 23845 2255 23903 2261
rect 23934 2252 23940 2304
rect 23992 2292 23998 2304
rect 24949 2295 25007 2301
rect 24949 2292 24961 2295
rect 23992 2264 24961 2292
rect 23992 2252 23998 2264
rect 24949 2261 24961 2264
rect 24995 2261 25007 2295
rect 25056 2292 25084 2332
rect 25976 2332 26372 2360
rect 25976 2292 26004 2332
rect 26878 2320 26884 2372
rect 26936 2360 26942 2372
rect 26936 2332 27936 2360
rect 26936 2320 26942 2332
rect 25056 2264 26004 2292
rect 24949 2255 25007 2261
rect 26050 2252 26056 2304
rect 26108 2252 26114 2304
rect 26234 2252 26240 2304
rect 26292 2292 26298 2304
rect 26421 2295 26479 2301
rect 26421 2292 26433 2295
rect 26292 2264 26433 2292
rect 26292 2252 26298 2264
rect 26421 2261 26433 2264
rect 26467 2261 26479 2295
rect 26421 2255 26479 2261
rect 26510 2252 26516 2304
rect 26568 2292 26574 2304
rect 27908 2301 27936 2332
rect 27525 2295 27583 2301
rect 27525 2292 27537 2295
rect 26568 2264 27537 2292
rect 26568 2252 26574 2264
rect 27525 2261 27537 2264
rect 27571 2261 27583 2295
rect 27525 2255 27583 2261
rect 27893 2295 27951 2301
rect 27893 2261 27905 2295
rect 27939 2261 27951 2295
rect 28000 2292 28028 2400
rect 28077 2397 28089 2431
rect 28123 2428 28135 2431
rect 28166 2428 28172 2440
rect 28123 2400 28172 2428
rect 28123 2397 28135 2400
rect 28077 2391 28135 2397
rect 28166 2388 28172 2400
rect 28224 2388 28230 2440
rect 28442 2388 28448 2440
rect 28500 2388 28506 2440
rect 28626 2388 28632 2440
rect 28684 2428 28690 2440
rect 28813 2431 28871 2437
rect 28813 2428 28825 2431
rect 28684 2400 28825 2428
rect 28684 2388 28690 2400
rect 28813 2397 28825 2400
rect 28859 2397 28871 2431
rect 28813 2391 28871 2397
rect 29825 2431 29883 2437
rect 29825 2397 29837 2431
rect 29871 2428 29883 2431
rect 30006 2428 30012 2440
rect 29871 2400 30012 2428
rect 29871 2397 29883 2400
rect 29825 2391 29883 2397
rect 30006 2388 30012 2400
rect 30064 2388 30070 2440
rect 30190 2388 30196 2440
rect 30248 2388 30254 2440
rect 30561 2431 30619 2437
rect 30561 2397 30573 2431
rect 30607 2428 30619 2431
rect 30650 2428 30656 2440
rect 30607 2400 30656 2428
rect 30607 2397 30619 2400
rect 30561 2391 30619 2397
rect 30650 2388 30656 2400
rect 30708 2388 30714 2440
rect 31312 2437 31340 2468
rect 31754 2456 31760 2468
rect 31812 2456 31818 2508
rect 32030 2456 32036 2508
rect 32088 2496 32094 2508
rect 32088 2468 38148 2496
rect 32088 2456 32094 2468
rect 30929 2431 30987 2437
rect 30929 2397 30941 2431
rect 30975 2397 30987 2431
rect 30929 2391 30987 2397
rect 31297 2431 31355 2437
rect 31297 2397 31309 2431
rect 31343 2397 31355 2431
rect 31297 2391 31355 2397
rect 29454 2320 29460 2372
rect 29512 2360 29518 2372
rect 30944 2360 30972 2391
rect 31386 2388 31392 2440
rect 31444 2388 31450 2440
rect 32122 2388 32128 2440
rect 32180 2388 32186 2440
rect 32490 2388 32496 2440
rect 32548 2388 32554 2440
rect 32858 2388 32864 2440
rect 32916 2388 32922 2440
rect 33410 2388 33416 2440
rect 33468 2428 33474 2440
rect 38120 2437 38148 2468
rect 37737 2431 37795 2437
rect 37737 2428 37749 2431
rect 33468 2400 37749 2428
rect 33468 2388 33474 2400
rect 37737 2397 37749 2400
rect 37783 2397 37795 2431
rect 37737 2391 37795 2397
rect 38105 2431 38163 2437
rect 38105 2397 38117 2431
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 38470 2388 38476 2440
rect 38528 2388 38534 2440
rect 39117 2431 39175 2437
rect 39117 2397 39129 2431
rect 39163 2428 39175 2431
rect 39209 2431 39267 2437
rect 39209 2428 39221 2431
rect 39163 2400 39221 2428
rect 39163 2397 39175 2400
rect 39117 2391 39175 2397
rect 39209 2397 39221 2400
rect 39255 2397 39267 2431
rect 39209 2391 39267 2397
rect 31846 2360 31852 2372
rect 29512 2332 30420 2360
rect 29512 2320 29518 2332
rect 28629 2295 28687 2301
rect 28629 2292 28641 2295
rect 28000 2264 28641 2292
rect 27893 2255 27951 2261
rect 28629 2261 28641 2264
rect 28675 2261 28687 2295
rect 28629 2255 28687 2261
rect 28718 2252 28724 2304
rect 28776 2292 28782 2304
rect 30392 2301 30420 2332
rect 30576 2332 30880 2360
rect 30944 2332 31852 2360
rect 30576 2304 30604 2332
rect 29641 2295 29699 2301
rect 29641 2292 29653 2295
rect 28776 2264 29653 2292
rect 28776 2252 28782 2264
rect 29641 2261 29653 2264
rect 29687 2261 29699 2295
rect 29641 2255 29699 2261
rect 30377 2295 30435 2301
rect 30377 2261 30389 2295
rect 30423 2261 30435 2295
rect 30377 2255 30435 2261
rect 30558 2252 30564 2304
rect 30616 2252 30622 2304
rect 30852 2292 30880 2332
rect 31846 2320 31852 2332
rect 31904 2320 31910 2372
rect 31938 2320 31944 2372
rect 31996 2360 32002 2372
rect 31996 2332 33088 2360
rect 31996 2320 32002 2332
rect 31573 2295 31631 2301
rect 31573 2292 31585 2295
rect 30852 2264 31585 2292
rect 31573 2261 31585 2264
rect 31619 2261 31631 2295
rect 31573 2255 31631 2261
rect 31662 2252 31668 2304
rect 31720 2292 31726 2304
rect 33060 2301 33088 2332
rect 32677 2295 32735 2301
rect 32677 2292 32689 2295
rect 31720 2264 32689 2292
rect 31720 2252 31726 2264
rect 32677 2261 32689 2264
rect 32723 2261 32735 2295
rect 32677 2255 32735 2261
rect 33045 2295 33103 2301
rect 33045 2261 33057 2295
rect 33091 2261 33103 2295
rect 33045 2255 33103 2261
rect 37918 2252 37924 2304
rect 37976 2252 37982 2304
rect 38286 2252 38292 2304
rect 38344 2252 38350 2304
rect 38654 2252 38660 2304
rect 38712 2252 38718 2304
rect 38930 2252 38936 2304
rect 38988 2292 38994 2304
rect 39025 2295 39083 2301
rect 39025 2292 39037 2295
rect 38988 2264 39037 2292
rect 38988 2252 38994 2264
rect 39025 2261 39037 2264
rect 39071 2261 39083 2295
rect 39025 2255 39083 2261
rect 1104 2202 39836 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 39010 2202
rect 39062 2150 39074 2202
rect 39126 2150 39138 2202
rect 39190 2150 39202 2202
rect 39254 2150 39266 2202
rect 39318 2150 39836 2202
rect 1104 2128 39836 2150
rect 14274 2048 14280 2100
rect 14332 2088 14338 2100
rect 25130 2088 25136 2100
rect 14332 2060 25136 2088
rect 14332 2048 14338 2060
rect 25130 2048 25136 2060
rect 25188 2048 25194 2100
rect 25498 2048 25504 2100
rect 25556 2088 25562 2100
rect 28166 2088 28172 2100
rect 25556 2060 28172 2088
rect 25556 2048 25562 2060
rect 28166 2048 28172 2060
rect 28224 2048 28230 2100
rect 33410 2088 33416 2100
rect 28276 2060 33416 2088
rect 9766 1980 9772 2032
rect 9824 2020 9830 2032
rect 9824 1992 17264 2020
rect 9824 1980 9830 1992
rect 11422 1912 11428 1964
rect 11480 1952 11486 1964
rect 11480 1924 12434 1952
rect 11480 1912 11486 1924
rect 12406 1816 12434 1924
rect 17236 1884 17264 1992
rect 23198 1980 23204 2032
rect 23256 2020 23262 2032
rect 28276 2020 28304 2060
rect 33410 2048 33416 2060
rect 33468 2048 33474 2100
rect 38470 2088 38476 2100
rect 35866 2060 38476 2088
rect 23256 1992 28304 2020
rect 23256 1980 23262 1992
rect 28442 1980 28448 2032
rect 28500 2020 28506 2032
rect 32030 2020 32036 2032
rect 28500 1992 32036 2020
rect 28500 1980 28506 1992
rect 32030 1980 32036 1992
rect 32088 1980 32094 2032
rect 35866 2020 35894 2060
rect 38470 2048 38476 2060
rect 38528 2048 38534 2100
rect 32232 1992 35894 2020
rect 21910 1912 21916 1964
rect 21968 1952 21974 1964
rect 21968 1924 28580 1952
rect 21968 1912 21974 1924
rect 22370 1884 22376 1896
rect 17236 1856 22376 1884
rect 22370 1844 22376 1856
rect 22428 1844 22434 1896
rect 25314 1844 25320 1896
rect 25372 1884 25378 1896
rect 26234 1884 26240 1896
rect 25372 1856 26240 1884
rect 25372 1844 25378 1856
rect 26234 1844 26240 1856
rect 26292 1844 26298 1896
rect 27246 1844 27252 1896
rect 27304 1884 27310 1896
rect 27614 1884 27620 1896
rect 27304 1856 27620 1884
rect 27304 1844 27310 1856
rect 27614 1844 27620 1856
rect 27672 1844 27678 1896
rect 20714 1816 20720 1828
rect 12406 1788 20720 1816
rect 20714 1776 20720 1788
rect 20772 1776 20778 1828
rect 23014 1776 23020 1828
rect 23072 1816 23078 1828
rect 28442 1816 28448 1828
rect 23072 1788 28448 1816
rect 23072 1776 23078 1788
rect 28442 1776 28448 1788
rect 28500 1776 28506 1828
rect 28552 1816 28580 1924
rect 28626 1912 28632 1964
rect 28684 1952 28690 1964
rect 32122 1952 32128 1964
rect 28684 1924 32128 1952
rect 28684 1912 28690 1924
rect 32122 1912 32128 1924
rect 32180 1912 32186 1964
rect 32232 1816 32260 1992
rect 32766 1912 32772 1964
rect 32824 1952 32830 1964
rect 33042 1952 33048 1964
rect 32824 1924 33048 1952
rect 32824 1912 32830 1924
rect 33042 1912 33048 1924
rect 33100 1912 33106 1964
rect 38930 1952 38936 1964
rect 35866 1924 38936 1952
rect 28552 1788 32260 1816
rect 16114 1708 16120 1760
rect 16172 1748 16178 1760
rect 24578 1748 24584 1760
rect 16172 1720 24584 1748
rect 16172 1708 16178 1720
rect 24578 1708 24584 1720
rect 24636 1708 24642 1760
rect 27982 1748 27988 1760
rect 25056 1720 27988 1748
rect 15378 1640 15384 1692
rect 15436 1680 15442 1692
rect 25056 1680 25084 1720
rect 27982 1708 27988 1720
rect 28040 1708 28046 1760
rect 35866 1748 35894 1924
rect 38930 1912 38936 1924
rect 38988 1912 38994 1964
rect 28184 1720 35894 1748
rect 15436 1652 25084 1680
rect 15436 1640 15442 1652
rect 27522 1640 27528 1692
rect 27580 1680 27586 1692
rect 27890 1680 27896 1692
rect 27580 1652 27896 1680
rect 27580 1640 27586 1652
rect 27890 1640 27896 1652
rect 27948 1640 27954 1692
rect 14918 1572 14924 1624
rect 14976 1612 14982 1624
rect 25222 1612 25228 1624
rect 14976 1584 25228 1612
rect 14976 1572 14982 1584
rect 25222 1572 25228 1584
rect 25280 1572 25286 1624
rect 20806 1504 20812 1556
rect 20864 1544 20870 1556
rect 24394 1544 24400 1556
rect 20864 1516 24400 1544
rect 20864 1504 20870 1516
rect 24394 1504 24400 1516
rect 24452 1504 24458 1556
rect 25038 1504 25044 1556
rect 25096 1544 25102 1556
rect 26050 1544 26056 1556
rect 25096 1516 26056 1544
rect 25096 1504 25102 1516
rect 26050 1504 26056 1516
rect 26108 1504 26114 1556
rect 22646 1436 22652 1488
rect 22704 1476 22710 1488
rect 28184 1476 28212 1720
rect 32858 1680 32864 1692
rect 22704 1448 28212 1476
rect 31726 1652 32864 1680
rect 22704 1436 22710 1448
rect 26418 1368 26424 1420
rect 26476 1408 26482 1420
rect 31726 1408 31754 1652
rect 32858 1640 32864 1652
rect 32916 1640 32922 1692
rect 26476 1380 31754 1408
rect 26476 1368 26482 1380
rect 15102 1300 15108 1352
rect 15160 1340 15166 1352
rect 22922 1340 22928 1352
rect 15160 1312 22928 1340
rect 15160 1300 15166 1312
rect 22922 1300 22928 1312
rect 22980 1300 22986 1352
rect 28810 1300 28816 1352
rect 28868 1340 28874 1352
rect 35250 1340 35256 1352
rect 28868 1312 35256 1340
rect 28868 1300 28874 1312
rect 35250 1300 35256 1312
rect 35308 1300 35314 1352
rect 4246 1232 4252 1284
rect 4304 1272 4310 1284
rect 5994 1272 6000 1284
rect 4304 1244 6000 1272
rect 4304 1232 4310 1244
rect 5994 1232 6000 1244
rect 6052 1232 6058 1284
rect 26786 1232 26792 1284
rect 26844 1272 26850 1284
rect 32490 1272 32496 1284
rect 26844 1244 32496 1272
rect 26844 1232 26850 1244
rect 32490 1232 32496 1244
rect 32548 1232 32554 1284
rect 13998 484 14004 536
rect 14056 524 14062 536
rect 23474 524 23480 536
rect 14056 496 23480 524
rect 14056 484 14062 496
rect 23474 484 23480 496
rect 23532 484 23538 536
rect 25406 484 25412 536
rect 25464 524 25470 536
rect 33594 524 33600 536
rect 25464 496 33600 524
rect 25464 484 25470 496
rect 33594 484 33600 496
rect 33652 484 33658 536
rect 14274 416 14280 468
rect 14332 456 14338 468
rect 23750 456 23756 468
rect 14332 428 23756 456
rect 14332 416 14338 428
rect 23750 416 23756 428
rect 23808 416 23814 468
rect 25682 416 25688 468
rect 25740 456 25746 468
rect 36078 456 36084 468
rect 25740 428 36084 456
rect 25740 416 25746 428
rect 36078 416 36084 428
rect 36136 416 36142 468
rect 13446 348 13452 400
rect 13504 388 13510 400
rect 24946 388 24952 400
rect 13504 360 24952 388
rect 13504 348 13510 360
rect 24946 348 24952 360
rect 25004 348 25010 400
rect 27706 348 27712 400
rect 27764 388 27770 400
rect 36354 388 36360 400
rect 27764 360 36360 388
rect 27764 348 27770 360
rect 36354 348 36360 360
rect 36412 348 36418 400
rect 15930 280 15936 332
rect 15988 320 15994 332
rect 29914 320 29920 332
rect 15988 292 29920 320
rect 15988 280 15994 292
rect 29914 280 29920 292
rect 29972 280 29978 332
rect 16482 212 16488 264
rect 16540 252 16546 264
rect 29822 252 29828 264
rect 16540 224 29828 252
rect 16540 212 16546 224
rect 29822 212 29828 224
rect 29880 212 29886 264
rect 15102 144 15108 196
rect 15160 144 15166 196
rect 15654 144 15660 196
rect 15712 184 15718 196
rect 31570 184 31576 196
rect 15712 156 31576 184
rect 15712 144 15718 156
rect 31570 144 31576 156
rect 31628 144 31634 196
rect 4430 8 4436 60
rect 4488 48 4494 60
rect 10778 48 10784 60
rect 4488 20 10784 48
rect 4488 8 4494 20
rect 10778 8 10784 20
rect 10836 8 10842 60
rect 15120 48 15148 144
rect 16298 76 16304 128
rect 16356 116 16362 128
rect 30374 116 30380 128
rect 16356 88 30380 116
rect 16356 76 16362 88
rect 30374 76 30380 88
rect 30432 76 30438 128
rect 32674 48 32680 60
rect 15120 20 32680 48
rect 32674 8 32680 20
rect 32732 8 32738 60
<< via1 >>
rect 1308 9324 1360 9376
rect 23020 9324 23072 9376
rect 20720 9256 20772 9308
rect 20812 9188 20864 9240
rect 25780 9188 25832 9240
rect 30196 9188 30248 9240
rect 18880 9120 18932 9172
rect 27436 9120 27488 9172
rect 16856 9052 16908 9104
rect 27804 9052 27856 9104
rect 13084 8984 13136 9036
rect 27528 8984 27580 9036
rect 16948 8916 17000 8968
rect 28080 8916 28132 8968
rect 37004 8916 37056 8968
rect 39764 8916 39816 8968
rect 17960 8848 18012 8900
rect 37556 8848 37608 8900
rect 3424 8780 3476 8832
rect 5356 8780 5408 8832
rect 18144 8780 18196 8832
rect 20352 8780 20404 8832
rect 33784 8780 33836 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 39010 8678 39062 8730
rect 39074 8678 39126 8730
rect 39138 8678 39190 8730
rect 39202 8678 39254 8730
rect 39266 8678 39318 8730
rect 1124 8576 1176 8628
rect 2872 8576 2924 8628
rect 3424 8576 3476 8628
rect 4988 8576 5040 8628
rect 6920 8576 6972 8628
rect 8852 8576 8904 8628
rect 10784 8576 10836 8628
rect 12716 8576 12768 8628
rect 14648 8576 14700 8628
rect 16580 8576 16632 8628
rect 18512 8576 18564 8628
rect 20444 8576 20496 8628
rect 22376 8576 22428 8628
rect 24308 8576 24360 8628
rect 26240 8576 26292 8628
rect 28172 8576 28224 8628
rect 30104 8576 30156 8628
rect 32036 8576 32088 8628
rect 33968 8576 34020 8628
rect 35900 8576 35952 8628
rect 37004 8619 37056 8628
rect 37004 8585 37013 8619
rect 37013 8585 37047 8619
rect 37047 8585 37056 8619
rect 37004 8576 37056 8585
rect 37740 8619 37792 8628
rect 37740 8585 37749 8619
rect 37749 8585 37783 8619
rect 37783 8585 37792 8619
rect 37740 8576 37792 8585
rect 37832 8576 37884 8628
rect 38660 8619 38712 8628
rect 38660 8585 38669 8619
rect 38669 8585 38703 8619
rect 38703 8585 38712 8619
rect 38660 8576 38712 8585
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 25872 8508 25924 8560
rect 13084 8483 13136 8492
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 16856 8440 16908 8492
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 18880 8483 18932 8492
rect 18880 8449 18889 8483
rect 18889 8449 18923 8483
rect 18923 8449 18932 8483
rect 18880 8440 18932 8449
rect 16580 8372 16632 8424
rect 22744 8483 22796 8492
rect 22744 8449 22753 8483
rect 22753 8449 22787 8483
rect 22787 8449 22796 8483
rect 22744 8440 22796 8449
rect 24676 8483 24728 8492
rect 24676 8449 24685 8483
rect 24685 8449 24719 8483
rect 24719 8449 24728 8483
rect 24676 8440 24728 8449
rect 24768 8440 24820 8492
rect 26332 8483 26384 8492
rect 26332 8449 26341 8483
rect 26341 8449 26375 8483
rect 26375 8449 26384 8483
rect 26332 8440 26384 8449
rect 25412 8372 25464 8424
rect 25596 8372 25648 8424
rect 30196 8483 30248 8492
rect 30196 8449 30205 8483
rect 30205 8449 30239 8483
rect 30239 8449 30248 8483
rect 30196 8440 30248 8449
rect 32588 8440 32640 8492
rect 31024 8372 31076 8424
rect 35992 8483 36044 8492
rect 35992 8449 36001 8483
rect 36001 8449 36035 8483
rect 36035 8449 36044 8483
rect 35992 8440 36044 8449
rect 36820 8483 36872 8492
rect 36820 8449 36829 8483
rect 36829 8449 36863 8483
rect 36863 8449 36872 8483
rect 36820 8440 36872 8449
rect 37556 8483 37608 8492
rect 37556 8449 37565 8483
rect 37565 8449 37599 8483
rect 37599 8449 37608 8483
rect 37556 8440 37608 8449
rect 37648 8440 37700 8492
rect 22192 8304 22244 8356
rect 22744 8304 22796 8356
rect 26884 8304 26936 8356
rect 33784 8304 33836 8356
rect 39028 8347 39080 8356
rect 39028 8313 39037 8347
rect 39037 8313 39071 8347
rect 39071 8313 39080 8347
rect 39028 8304 39080 8313
rect 39396 8347 39448 8356
rect 39396 8313 39405 8347
rect 39405 8313 39439 8347
rect 39439 8313 39448 8347
rect 39396 8304 39448 8313
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 37950 8134 38002 8186
rect 38014 8134 38066 8186
rect 38078 8134 38130 8186
rect 38142 8134 38194 8186
rect 38206 8134 38258 8186
rect 16488 8032 16540 8084
rect 18880 8032 18932 8084
rect 19248 8032 19300 8084
rect 17132 7964 17184 8016
rect 16120 7896 16172 7948
rect 18328 7896 18380 7948
rect 22468 7896 22520 7948
rect 16396 7828 16448 7880
rect 19984 7828 20036 7880
rect 20904 7828 20956 7880
rect 38292 8075 38344 8084
rect 38292 8041 38301 8075
rect 38301 8041 38335 8075
rect 38335 8041 38344 8075
rect 38292 8032 38344 8041
rect 39488 8032 39540 8084
rect 23204 7964 23256 8016
rect 16580 7760 16632 7812
rect 19340 7760 19392 7812
rect 37740 7871 37792 7880
rect 37740 7837 37749 7871
rect 37749 7837 37783 7871
rect 37783 7837 37792 7871
rect 37740 7828 37792 7837
rect 38108 7871 38160 7880
rect 38108 7837 38117 7871
rect 38117 7837 38151 7871
rect 38151 7837 38160 7871
rect 38108 7828 38160 7837
rect 37832 7760 37884 7812
rect 38016 7760 38068 7812
rect 14832 7692 14884 7744
rect 17776 7692 17828 7744
rect 19064 7692 19116 7744
rect 20444 7692 20496 7744
rect 25412 7692 25464 7744
rect 26148 7692 26200 7744
rect 27436 7692 27488 7744
rect 28356 7692 28408 7744
rect 38384 7692 38436 7744
rect 38936 7692 38988 7744
rect 39396 7735 39448 7744
rect 39396 7701 39405 7735
rect 39405 7701 39439 7735
rect 39439 7701 39448 7735
rect 39396 7692 39448 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 39010 7590 39062 7642
rect 39074 7590 39126 7642
rect 39138 7590 39190 7642
rect 39202 7590 39254 7642
rect 39266 7590 39318 7642
rect 14924 7488 14976 7540
rect 16120 7463 16172 7472
rect 16120 7429 16129 7463
rect 16129 7429 16163 7463
rect 16163 7429 16172 7463
rect 16120 7420 16172 7429
rect 15108 7352 15160 7404
rect 16488 7284 16540 7336
rect 17776 7395 17828 7404
rect 17776 7361 17785 7395
rect 17785 7361 17819 7395
rect 17819 7361 17828 7395
rect 17776 7352 17828 7361
rect 17960 7531 18012 7540
rect 17960 7497 17969 7531
rect 17969 7497 18003 7531
rect 18003 7497 18012 7531
rect 17960 7488 18012 7497
rect 18144 7531 18196 7540
rect 18144 7497 18153 7531
rect 18153 7497 18187 7531
rect 18187 7497 18196 7531
rect 18144 7488 18196 7497
rect 18696 7531 18748 7540
rect 18696 7497 18705 7531
rect 18705 7497 18739 7531
rect 18739 7497 18748 7531
rect 18696 7488 18748 7497
rect 18880 7531 18932 7540
rect 18880 7497 18889 7531
rect 18889 7497 18923 7531
rect 18923 7497 18932 7531
rect 18880 7488 18932 7497
rect 19248 7531 19300 7540
rect 19248 7497 19257 7531
rect 19257 7497 19291 7531
rect 19291 7497 19300 7531
rect 19248 7488 19300 7497
rect 19340 7531 19392 7540
rect 19340 7497 19349 7531
rect 19349 7497 19383 7531
rect 19383 7497 19392 7531
rect 19340 7488 19392 7497
rect 20352 7488 20404 7540
rect 20444 7531 20496 7540
rect 20444 7497 20453 7531
rect 20453 7497 20487 7531
rect 20487 7497 20496 7531
rect 20444 7488 20496 7497
rect 20720 7531 20772 7540
rect 20720 7497 20729 7531
rect 20729 7497 20763 7531
rect 20763 7497 20772 7531
rect 20720 7488 20772 7497
rect 20812 7531 20864 7540
rect 20812 7497 20821 7531
rect 20821 7497 20855 7531
rect 20855 7497 20864 7531
rect 20812 7488 20864 7497
rect 20904 7488 20956 7540
rect 22100 7531 22152 7540
rect 22100 7497 22109 7531
rect 22109 7497 22143 7531
rect 22143 7497 22152 7531
rect 22100 7488 22152 7497
rect 22560 7531 22612 7540
rect 22560 7497 22569 7531
rect 22569 7497 22603 7531
rect 22603 7497 22612 7531
rect 22560 7488 22612 7497
rect 18328 7395 18380 7404
rect 18328 7361 18337 7395
rect 18337 7361 18371 7395
rect 18371 7361 18380 7395
rect 18328 7352 18380 7361
rect 19616 7395 19668 7404
rect 19616 7361 19625 7395
rect 19625 7361 19659 7395
rect 19659 7361 19668 7395
rect 19616 7352 19668 7361
rect 19984 7395 20036 7404
rect 19984 7361 19993 7395
rect 19993 7361 20027 7395
rect 20027 7361 20036 7395
rect 19984 7352 20036 7361
rect 23020 7395 23072 7404
rect 23020 7361 23029 7395
rect 23029 7361 23063 7395
rect 23063 7361 23072 7395
rect 23020 7352 23072 7361
rect 23204 7352 23256 7404
rect 25228 7352 25280 7404
rect 22928 7284 22980 7336
rect 23112 7216 23164 7268
rect 26884 7420 26936 7472
rect 28448 7420 28500 7472
rect 39580 7488 39632 7540
rect 27344 7395 27396 7404
rect 27344 7361 27353 7395
rect 27353 7361 27387 7395
rect 27387 7361 27396 7395
rect 27344 7352 27396 7361
rect 27712 7395 27764 7404
rect 27712 7361 27721 7395
rect 27721 7361 27755 7395
rect 27755 7361 27764 7395
rect 27712 7352 27764 7361
rect 27988 7395 28040 7404
rect 27988 7361 27997 7395
rect 27997 7361 28031 7395
rect 28031 7361 28040 7395
rect 27988 7352 28040 7361
rect 28264 7395 28316 7404
rect 28264 7361 28273 7395
rect 28273 7361 28307 7395
rect 28307 7361 28316 7395
rect 28264 7352 28316 7361
rect 28816 7395 28868 7404
rect 28816 7361 28825 7395
rect 28825 7361 28859 7395
rect 28859 7361 28868 7395
rect 28816 7352 28868 7361
rect 37740 7420 37792 7472
rect 37832 7420 37884 7472
rect 34704 7352 34756 7404
rect 38844 7395 38896 7404
rect 38844 7361 38853 7395
rect 38853 7361 38887 7395
rect 38887 7361 38896 7395
rect 38844 7352 38896 7361
rect 38108 7284 38160 7336
rect 23296 7216 23348 7268
rect 38016 7216 38068 7268
rect 17132 7191 17184 7200
rect 17132 7157 17141 7191
rect 17141 7157 17175 7191
rect 17175 7157 17184 7191
rect 17132 7148 17184 7157
rect 17776 7148 17828 7200
rect 19616 7148 19668 7200
rect 19800 7191 19852 7200
rect 19800 7157 19809 7191
rect 19809 7157 19843 7191
rect 19843 7157 19852 7191
rect 19800 7148 19852 7157
rect 21364 7191 21416 7200
rect 21364 7157 21373 7191
rect 21373 7157 21407 7191
rect 21407 7157 21416 7191
rect 21364 7148 21416 7157
rect 24768 7148 24820 7200
rect 25872 7148 25924 7200
rect 26148 7148 26200 7200
rect 27528 7191 27580 7200
rect 27528 7157 27537 7191
rect 27537 7157 27571 7191
rect 27571 7157 27580 7191
rect 27528 7148 27580 7157
rect 27804 7191 27856 7200
rect 27804 7157 27813 7191
rect 27813 7157 27847 7191
rect 27847 7157 27856 7191
rect 27804 7148 27856 7157
rect 28080 7191 28132 7200
rect 28080 7157 28089 7191
rect 28089 7157 28123 7191
rect 28123 7157 28132 7191
rect 28080 7148 28132 7157
rect 28356 7191 28408 7200
rect 28356 7157 28365 7191
rect 28365 7157 28399 7191
rect 28399 7157 28408 7191
rect 28356 7148 28408 7157
rect 28448 7148 28500 7200
rect 39396 7191 39448 7200
rect 39396 7157 39405 7191
rect 39405 7157 39439 7191
rect 39439 7157 39448 7191
rect 39396 7148 39448 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 37950 7046 38002 7098
rect 38014 7046 38066 7098
rect 38078 7046 38130 7098
rect 38142 7046 38194 7098
rect 38206 7046 38258 7098
rect 19800 6944 19852 6996
rect 38844 6944 38896 6996
rect 9128 6876 9180 6928
rect 7748 6808 7800 6860
rect 7840 6740 7892 6792
rect 9588 6783 9640 6792
rect 9588 6749 9597 6783
rect 9597 6749 9631 6783
rect 9631 6749 9640 6783
rect 9588 6740 9640 6749
rect 9956 6783 10008 6792
rect 9956 6749 9965 6783
rect 9965 6749 9999 6783
rect 9999 6749 10008 6783
rect 9956 6740 10008 6749
rect 10784 6808 10836 6860
rect 10508 6740 10560 6792
rect 10876 6740 10928 6792
rect 17500 6851 17552 6860
rect 17500 6817 17509 6851
rect 17509 6817 17543 6851
rect 17543 6817 17552 6851
rect 17500 6808 17552 6817
rect 17868 6919 17920 6928
rect 17868 6885 17877 6919
rect 17877 6885 17911 6919
rect 17911 6885 17920 6919
rect 17868 6876 17920 6885
rect 21364 6876 21416 6928
rect 26884 6876 26936 6928
rect 27712 6876 27764 6928
rect 33876 6876 33928 6928
rect 18420 6808 18472 6860
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 32312 6808 32364 6860
rect 32772 6740 32824 6792
rect 1584 6672 1636 6724
rect 4620 6604 4672 6656
rect 9128 6604 9180 6656
rect 9404 6604 9456 6656
rect 9496 6647 9548 6656
rect 9496 6613 9505 6647
rect 9505 6613 9539 6647
rect 9539 6613 9548 6647
rect 9496 6604 9548 6613
rect 9772 6647 9824 6656
rect 9772 6613 9781 6647
rect 9781 6613 9815 6647
rect 9815 6613 9824 6647
rect 9772 6604 9824 6613
rect 10232 6604 10284 6656
rect 10692 6604 10744 6656
rect 11244 6647 11296 6656
rect 11244 6613 11253 6647
rect 11253 6613 11287 6647
rect 11287 6613 11296 6647
rect 11244 6604 11296 6613
rect 11428 6604 11480 6656
rect 11888 6647 11940 6656
rect 11888 6613 11897 6647
rect 11897 6613 11931 6647
rect 11931 6613 11940 6647
rect 11888 6604 11940 6613
rect 11980 6604 12032 6656
rect 18696 6604 18748 6656
rect 31576 6672 31628 6724
rect 39212 6783 39264 6792
rect 39212 6749 39221 6783
rect 39221 6749 39255 6783
rect 39255 6749 39264 6783
rect 39212 6740 39264 6749
rect 22192 6647 22244 6656
rect 22192 6613 22201 6647
rect 22201 6613 22235 6647
rect 22235 6613 22244 6647
rect 22192 6604 22244 6613
rect 39948 6672 40000 6724
rect 39396 6647 39448 6656
rect 39396 6613 39405 6647
rect 39405 6613 39439 6647
rect 39439 6613 39448 6647
rect 39396 6604 39448 6613
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 39010 6502 39062 6554
rect 39074 6502 39126 6554
rect 39138 6502 39190 6554
rect 39202 6502 39254 6554
rect 39266 6502 39318 6554
rect 6552 6400 6604 6452
rect 8484 6264 8536 6316
rect 9404 6400 9456 6452
rect 22284 6400 22336 6452
rect 24676 6400 24728 6452
rect 39396 6443 39448 6452
rect 39396 6409 39405 6443
rect 39405 6409 39439 6443
rect 39439 6409 39448 6443
rect 39396 6400 39448 6409
rect 9128 6332 9180 6384
rect 9588 6332 9640 6384
rect 11520 6332 11572 6384
rect 11704 6264 11756 6316
rect 11796 6264 11848 6316
rect 17960 6332 18012 6384
rect 7380 6196 7432 6248
rect 9956 6196 10008 6248
rect 12072 6196 12124 6248
rect 14004 6196 14056 6248
rect 21364 6196 21416 6248
rect 35532 6264 35584 6316
rect 38660 6264 38712 6316
rect 7656 6060 7708 6112
rect 9128 6060 9180 6112
rect 9496 6060 9548 6112
rect 13636 6060 13688 6112
rect 20720 6128 20772 6180
rect 22928 6128 22980 6180
rect 33508 6128 33560 6180
rect 14004 6060 14056 6112
rect 14280 6060 14332 6112
rect 14924 6060 14976 6112
rect 15016 6060 15068 6112
rect 21824 6060 21876 6112
rect 39028 6103 39080 6112
rect 39028 6069 39037 6103
rect 39037 6069 39071 6103
rect 39071 6069 39080 6103
rect 39028 6060 39080 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 37950 5958 38002 6010
rect 38014 5958 38066 6010
rect 38078 5958 38130 6010
rect 38142 5958 38194 6010
rect 38206 5958 38258 6010
rect 11980 5856 12032 5908
rect 13636 5856 13688 5908
rect 15016 5856 15068 5908
rect 7104 5720 7156 5772
rect 10508 5720 10560 5772
rect 12532 5720 12584 5772
rect 16120 5788 16172 5840
rect 17408 5856 17460 5908
rect 5172 5652 5224 5704
rect 4988 5584 5040 5636
rect 11244 5652 11296 5704
rect 13728 5695 13780 5704
rect 13728 5661 13737 5695
rect 13737 5661 13771 5695
rect 13771 5661 13780 5695
rect 13728 5652 13780 5661
rect 14556 5695 14608 5704
rect 14556 5661 14565 5695
rect 14565 5661 14599 5695
rect 14599 5661 14608 5695
rect 14556 5652 14608 5661
rect 12624 5584 12676 5636
rect 20812 5720 20864 5772
rect 26332 5899 26384 5908
rect 26332 5865 26341 5899
rect 26341 5865 26375 5899
rect 26375 5865 26384 5899
rect 26332 5856 26384 5865
rect 39396 5831 39448 5840
rect 39396 5797 39405 5831
rect 39405 5797 39439 5831
rect 39439 5797 39448 5831
rect 39396 5788 39448 5797
rect 31576 5720 31628 5772
rect 19524 5652 19576 5704
rect 35808 5652 35860 5704
rect 38844 5695 38896 5704
rect 38844 5661 38853 5695
rect 38853 5661 38887 5695
rect 38887 5661 38896 5695
rect 38844 5652 38896 5661
rect 6828 5516 6880 5568
rect 10876 5516 10928 5568
rect 13636 5559 13688 5568
rect 13636 5525 13645 5559
rect 13645 5525 13679 5559
rect 13679 5525 13688 5559
rect 13636 5516 13688 5525
rect 14372 5516 14424 5568
rect 20444 5584 20496 5636
rect 24860 5516 24912 5568
rect 39948 5516 40000 5568
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 39010 5414 39062 5466
rect 39074 5414 39126 5466
rect 39138 5414 39190 5466
rect 39202 5414 39254 5466
rect 39266 5414 39318 5466
rect 6092 5312 6144 5364
rect 9588 5312 9640 5364
rect 11060 5312 11112 5364
rect 10140 5244 10192 5296
rect 3516 5176 3568 5228
rect 5448 5176 5500 5228
rect 10416 5176 10468 5228
rect 17960 5355 18012 5364
rect 17960 5321 17969 5355
rect 17969 5321 18003 5355
rect 18003 5321 18012 5355
rect 17960 5312 18012 5321
rect 22008 5312 22060 5364
rect 24124 5244 24176 5296
rect 36820 5312 36872 5364
rect 39396 5355 39448 5364
rect 39396 5321 39405 5355
rect 39405 5321 39439 5355
rect 39439 5321 39448 5355
rect 39396 5312 39448 5321
rect 4068 5108 4120 5160
rect 12900 5108 12952 5160
rect 22376 5219 22428 5228
rect 22376 5185 22385 5219
rect 22385 5185 22419 5219
rect 22419 5185 22428 5219
rect 22376 5176 22428 5185
rect 28080 5176 28132 5228
rect 31392 5176 31444 5228
rect 37740 5176 37792 5228
rect 39212 5219 39264 5228
rect 39212 5185 39221 5219
rect 39221 5185 39255 5219
rect 39255 5185 39264 5219
rect 39212 5176 39264 5185
rect 3792 5040 3844 5092
rect 3056 4972 3108 5024
rect 5356 4972 5408 5024
rect 5540 4972 5592 5024
rect 11152 4972 11204 5024
rect 15568 5015 15620 5024
rect 15568 4981 15577 5015
rect 15577 4981 15611 5015
rect 15611 4981 15620 5015
rect 15568 4972 15620 4981
rect 21732 5040 21784 5092
rect 27436 5108 27488 5160
rect 27620 5108 27672 5160
rect 32496 5108 32548 5160
rect 23204 5040 23256 5092
rect 33784 5040 33836 5092
rect 22468 4972 22520 5024
rect 38660 4972 38712 5024
rect 39028 5015 39080 5024
rect 39028 4981 39037 5015
rect 39037 4981 39071 5015
rect 39071 4981 39080 5015
rect 39028 4972 39080 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 37950 4870 38002 4922
rect 38014 4870 38066 4922
rect 38078 4870 38130 4922
rect 38142 4870 38194 4922
rect 38206 4870 38258 4922
rect 6092 4768 6144 4820
rect 16672 4768 16724 4820
rect 21732 4768 21784 4820
rect 23204 4811 23256 4820
rect 23204 4777 23213 4811
rect 23213 4777 23247 4811
rect 23247 4777 23256 4811
rect 23204 4768 23256 4777
rect 23480 4811 23532 4820
rect 23480 4777 23489 4811
rect 23489 4777 23523 4811
rect 23523 4777 23532 4811
rect 23480 4768 23532 4777
rect 23756 4768 23808 4820
rect 4896 4743 4948 4752
rect 4896 4709 4905 4743
rect 4905 4709 4939 4743
rect 4939 4709 4948 4743
rect 4896 4700 4948 4709
rect 15568 4700 15620 4752
rect 5356 4632 5408 4684
rect 17776 4632 17828 4684
rect 19800 4632 19852 4684
rect 2872 4564 2924 4616
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 5724 4564 5776 4616
rect 8668 4564 8720 4616
rect 9864 4564 9916 4616
rect 16580 4607 16632 4616
rect 16580 4573 16589 4607
rect 16589 4573 16623 4607
rect 16623 4573 16632 4607
rect 16580 4564 16632 4573
rect 3056 4496 3108 4548
rect 17960 4496 18012 4548
rect 22836 4675 22888 4684
rect 22836 4641 22845 4675
rect 22845 4641 22879 4675
rect 22879 4641 22888 4675
rect 22836 4632 22888 4641
rect 25044 4700 25096 4752
rect 27620 4811 27672 4820
rect 27620 4777 27629 4811
rect 27629 4777 27663 4811
rect 27663 4777 27672 4811
rect 27620 4768 27672 4777
rect 31300 4768 31352 4820
rect 31392 4811 31444 4820
rect 31392 4777 31401 4811
rect 31401 4777 31435 4811
rect 31435 4777 31444 4811
rect 31392 4768 31444 4777
rect 24032 4607 24084 4616
rect 24032 4573 24041 4607
rect 24041 4573 24075 4607
rect 24075 4573 24084 4607
rect 24032 4564 24084 4573
rect 25688 4564 25740 4616
rect 26608 4564 26660 4616
rect 25872 4496 25924 4548
rect 26792 4496 26844 4548
rect 4344 4428 4396 4480
rect 11060 4428 11112 4480
rect 20444 4471 20496 4480
rect 20444 4437 20453 4471
rect 20453 4437 20487 4471
rect 20487 4437 20496 4471
rect 20444 4428 20496 4437
rect 24216 4471 24268 4480
rect 24216 4437 24225 4471
rect 24225 4437 24259 4471
rect 24259 4437 24268 4471
rect 24216 4428 24268 4437
rect 25596 4471 25648 4480
rect 25596 4437 25605 4471
rect 25605 4437 25639 4471
rect 25639 4437 25648 4471
rect 25596 4428 25648 4437
rect 26424 4428 26476 4480
rect 28540 4428 28592 4480
rect 29000 4471 29052 4480
rect 29000 4437 29009 4471
rect 29009 4437 29043 4471
rect 29043 4437 29052 4471
rect 29000 4428 29052 4437
rect 30840 4700 30892 4752
rect 31576 4675 31628 4684
rect 31576 4641 31585 4675
rect 31585 4641 31619 4675
rect 31619 4641 31628 4675
rect 31576 4632 31628 4641
rect 31760 4632 31812 4684
rect 31852 4564 31904 4616
rect 35992 4768 36044 4820
rect 33784 4700 33836 4752
rect 32680 4564 32732 4616
rect 37096 4632 37148 4684
rect 37464 4564 37516 4616
rect 39396 4743 39448 4752
rect 39396 4709 39405 4743
rect 39405 4709 39439 4743
rect 39439 4709 39448 4743
rect 39396 4700 39448 4709
rect 29552 4496 29604 4548
rect 30932 4428 30984 4480
rect 31024 4471 31076 4480
rect 31024 4437 31033 4471
rect 31033 4437 31067 4471
rect 31067 4437 31076 4471
rect 31024 4428 31076 4437
rect 31760 4471 31812 4480
rect 31760 4437 31769 4471
rect 31769 4437 31803 4471
rect 31803 4437 31812 4471
rect 31760 4428 31812 4437
rect 31852 4428 31904 4480
rect 32404 4428 32456 4480
rect 37188 4428 37240 4480
rect 39948 4428 40000 4480
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 39010 4326 39062 4378
rect 39074 4326 39126 4378
rect 39138 4326 39190 4378
rect 39202 4326 39254 4378
rect 39266 4326 39318 4378
rect 4896 4224 4948 4276
rect 9680 4224 9732 4276
rect 9864 4224 9916 4276
rect 21916 4224 21968 4276
rect 24216 4224 24268 4276
rect 35900 4224 35952 4276
rect 4344 4156 4396 4208
rect 10876 4156 10928 4208
rect 11152 4156 11204 4208
rect 21732 4156 21784 4208
rect 23664 4156 23716 4208
rect 29000 4156 29052 4208
rect 6276 4088 6328 4140
rect 9496 4088 9548 4140
rect 9404 4020 9456 4072
rect 19432 4131 19484 4140
rect 19432 4097 19441 4131
rect 19441 4097 19475 4131
rect 19475 4097 19484 4131
rect 19432 4088 19484 4097
rect 21548 4131 21600 4140
rect 21548 4097 21557 4131
rect 21557 4097 21591 4131
rect 21591 4097 21600 4131
rect 21548 4088 21600 4097
rect 22100 4088 22152 4140
rect 25412 4088 25464 4140
rect 28172 4131 28224 4140
rect 28172 4097 28181 4131
rect 28181 4097 28215 4131
rect 28215 4097 28224 4131
rect 28172 4088 28224 4097
rect 29460 4088 29512 4140
rect 30380 4088 30432 4140
rect 31576 4131 31628 4140
rect 31576 4097 31585 4131
rect 31585 4097 31619 4131
rect 31619 4097 31628 4131
rect 31576 4088 31628 4097
rect 31944 4156 31996 4208
rect 36912 4156 36964 4208
rect 10692 3952 10744 4004
rect 10968 3952 11020 4004
rect 22008 3995 22060 4004
rect 22008 3961 22017 3995
rect 22017 3961 22051 3995
rect 22051 3961 22060 3995
rect 22008 3952 22060 3961
rect 4896 3927 4948 3936
rect 4896 3893 4905 3927
rect 4905 3893 4939 3927
rect 4939 3893 4948 3927
rect 4896 3884 4948 3893
rect 11888 3884 11940 3936
rect 17132 3884 17184 3936
rect 19524 3884 19576 3936
rect 19616 3927 19668 3936
rect 19616 3893 19625 3927
rect 19625 3893 19659 3927
rect 19659 3893 19668 3927
rect 19616 3884 19668 3893
rect 24216 3927 24268 3936
rect 24216 3893 24225 3927
rect 24225 3893 24259 3927
rect 24259 3893 24268 3927
rect 24216 3884 24268 3893
rect 29276 3952 29328 4004
rect 26332 3884 26384 3936
rect 27896 3884 27948 3936
rect 28632 3884 28684 3936
rect 29000 3927 29052 3936
rect 29000 3893 29009 3927
rect 29009 3893 29043 3927
rect 29043 3893 29052 3927
rect 29000 3884 29052 3893
rect 29184 3927 29236 3936
rect 29184 3893 29193 3927
rect 29193 3893 29227 3927
rect 29227 3893 29236 3927
rect 29184 3884 29236 3893
rect 30104 3952 30156 4004
rect 30748 3952 30800 4004
rect 35900 4020 35952 4072
rect 39212 3952 39264 4004
rect 39396 3995 39448 4004
rect 39396 3961 39405 3995
rect 39405 3961 39439 3995
rect 39439 3961 39448 3995
rect 39396 3952 39448 3961
rect 29828 3927 29880 3936
rect 29828 3893 29837 3927
rect 29837 3893 29871 3927
rect 29871 3893 29880 3927
rect 29828 3884 29880 3893
rect 30012 3927 30064 3936
rect 30012 3893 30021 3927
rect 30021 3893 30055 3927
rect 30055 3893 30064 3927
rect 30012 3884 30064 3893
rect 31024 3927 31076 3936
rect 31024 3893 31033 3927
rect 31033 3893 31067 3927
rect 31067 3893 31076 3927
rect 31024 3884 31076 3893
rect 31116 3927 31168 3936
rect 31116 3893 31125 3927
rect 31125 3893 31159 3927
rect 31159 3893 31168 3927
rect 31116 3884 31168 3893
rect 39028 3927 39080 3936
rect 39028 3893 39037 3927
rect 39037 3893 39071 3927
rect 39071 3893 39080 3927
rect 39028 3884 39080 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 37950 3782 38002 3834
rect 38014 3782 38066 3834
rect 38078 3782 38130 3834
rect 38142 3782 38194 3834
rect 38206 3782 38258 3834
rect 19156 3680 19208 3732
rect 21916 3680 21968 3732
rect 22744 3680 22796 3732
rect 24308 3680 24360 3732
rect 24400 3680 24452 3732
rect 25780 3723 25832 3732
rect 25780 3689 25789 3723
rect 25789 3689 25823 3723
rect 25823 3689 25832 3723
rect 25780 3680 25832 3689
rect 30196 3680 30248 3732
rect 31116 3680 31168 3732
rect 572 3612 624 3664
rect 19432 3612 19484 3664
rect 20720 3612 20772 3664
rect 22836 3612 22888 3664
rect 23112 3612 23164 3664
rect 17132 3544 17184 3596
rect 11060 3476 11112 3528
rect 18236 3476 18288 3528
rect 18512 3476 18564 3528
rect 19156 3476 19208 3528
rect 19524 3476 19576 3528
rect 9680 3408 9732 3460
rect 19616 3408 19668 3460
rect 21732 3519 21784 3528
rect 21732 3485 21741 3519
rect 21741 3485 21775 3519
rect 21775 3485 21784 3519
rect 21732 3476 21784 3485
rect 23112 3519 23164 3528
rect 23112 3485 23121 3519
rect 23121 3485 23155 3519
rect 23155 3485 23164 3519
rect 23112 3476 23164 3485
rect 38844 3612 38896 3664
rect 39396 3655 39448 3664
rect 39396 3621 39405 3655
rect 39405 3621 39439 3655
rect 39439 3621 39448 3655
rect 39396 3612 39448 3621
rect 24400 3519 24452 3528
rect 24400 3485 24409 3519
rect 24409 3485 24443 3519
rect 24443 3485 24452 3519
rect 24400 3476 24452 3485
rect 24952 3519 25004 3528
rect 24952 3485 24961 3519
rect 24961 3485 24995 3519
rect 24995 3485 25004 3519
rect 24952 3476 25004 3485
rect 26148 3476 26200 3528
rect 26516 3519 26568 3528
rect 26516 3485 26525 3519
rect 26525 3485 26559 3519
rect 26559 3485 26568 3519
rect 26516 3476 26568 3485
rect 29920 3476 29972 3528
rect 31024 3476 31076 3528
rect 39212 3519 39264 3528
rect 39212 3485 39221 3519
rect 39221 3485 39255 3519
rect 39255 3485 39264 3519
rect 39212 3476 39264 3485
rect 23480 3408 23532 3460
rect 18236 3383 18288 3392
rect 18236 3349 18245 3383
rect 18245 3349 18279 3383
rect 18279 3349 18288 3383
rect 18236 3340 18288 3349
rect 18604 3383 18656 3392
rect 18604 3349 18613 3383
rect 18613 3349 18647 3383
rect 18647 3349 18656 3383
rect 18604 3340 18656 3349
rect 19340 3340 19392 3392
rect 19432 3383 19484 3392
rect 19432 3349 19441 3383
rect 19441 3349 19475 3383
rect 19475 3349 19484 3383
rect 19432 3340 19484 3349
rect 21916 3383 21968 3392
rect 21916 3349 21925 3383
rect 21925 3349 21959 3383
rect 21959 3349 21968 3383
rect 21916 3340 21968 3349
rect 22560 3383 22612 3392
rect 22560 3349 22569 3383
rect 22569 3349 22603 3383
rect 22603 3349 22612 3383
rect 22560 3340 22612 3349
rect 22652 3383 22704 3392
rect 22652 3349 22661 3383
rect 22661 3349 22695 3383
rect 22695 3349 22704 3383
rect 22652 3340 22704 3349
rect 23020 3383 23072 3392
rect 23020 3349 23029 3383
rect 23029 3349 23063 3383
rect 23063 3349 23072 3383
rect 23020 3340 23072 3349
rect 23204 3340 23256 3392
rect 24768 3408 24820 3460
rect 24124 3383 24176 3392
rect 24124 3349 24133 3383
rect 24133 3349 24167 3383
rect 24167 3349 24176 3383
rect 24124 3340 24176 3349
rect 38936 3408 38988 3460
rect 32588 3340 32640 3392
rect 39948 3340 40000 3392
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 39010 3238 39062 3290
rect 39074 3238 39126 3290
rect 39138 3238 39190 3290
rect 39202 3238 39254 3290
rect 39266 3238 39318 3290
rect 8852 3136 8904 3188
rect 18236 3136 18288 3188
rect 18604 3136 18656 3188
rect 23296 3136 23348 3188
rect 23388 3136 23440 3188
rect 24308 3136 24360 3188
rect 4896 3068 4948 3120
rect 17960 3000 18012 3052
rect 18328 3000 18380 3052
rect 18788 3000 18840 3052
rect 19340 3068 19392 3120
rect 22744 3068 22796 3120
rect 22836 3068 22888 3120
rect 24768 3136 24820 3188
rect 19616 3043 19668 3052
rect 19616 3009 19625 3043
rect 19625 3009 19659 3043
rect 19659 3009 19668 3043
rect 19616 3000 19668 3009
rect 28448 3068 28500 3120
rect 11980 2932 12032 2984
rect 22468 2932 22520 2984
rect 24860 3000 24912 3052
rect 25872 3000 25924 3052
rect 23480 2932 23532 2984
rect 27896 3043 27948 3052
rect 27896 3009 27905 3043
rect 27905 3009 27939 3043
rect 27939 3009 27948 3043
rect 27896 3000 27948 3009
rect 29184 3000 29236 3052
rect 30104 3000 30156 3052
rect 32404 3068 32456 3120
rect 30840 3000 30892 3052
rect 31300 3043 31352 3052
rect 31300 3009 31309 3043
rect 31309 3009 31343 3043
rect 31343 3009 31352 3043
rect 31300 3000 31352 3009
rect 39396 3179 39448 3188
rect 39396 3145 39405 3179
rect 39405 3145 39439 3179
rect 39439 3145 39448 3179
rect 39396 3136 39448 3145
rect 38844 3043 38896 3052
rect 38844 3009 38853 3043
rect 38853 3009 38887 3043
rect 38887 3009 38896 3043
rect 38844 3000 38896 3009
rect 38936 3000 38988 3052
rect 9588 2864 9640 2916
rect 22652 2864 22704 2916
rect 23296 2864 23348 2916
rect 25504 2864 25556 2916
rect 26148 2864 26200 2916
rect 27712 2864 27764 2916
rect 40408 2864 40460 2916
rect 18144 2796 18196 2848
rect 18972 2796 19024 2848
rect 19524 2796 19576 2848
rect 23112 2796 23164 2848
rect 23480 2796 23532 2848
rect 23664 2796 23716 2848
rect 24492 2796 24544 2848
rect 25596 2796 25648 2848
rect 26332 2796 26384 2848
rect 26700 2796 26752 2848
rect 27804 2796 27856 2848
rect 28356 2796 28408 2848
rect 28908 2796 28960 2848
rect 30104 2796 30156 2848
rect 30840 2796 30892 2848
rect 31208 2796 31260 2848
rect 39028 2839 39080 2848
rect 39028 2805 39037 2839
rect 39037 2805 39071 2839
rect 39071 2805 39080 2839
rect 39028 2796 39080 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 37950 2694 38002 2746
rect 38014 2694 38066 2746
rect 38078 2694 38130 2746
rect 38142 2694 38194 2746
rect 38206 2694 38258 2746
rect 7748 2592 7800 2644
rect 8208 2592 8260 2644
rect 10968 2592 11020 2644
rect 13728 2592 13780 2644
rect 10600 2524 10652 2576
rect 21180 2592 21232 2644
rect 22008 2592 22060 2644
rect 22192 2592 22244 2644
rect 22560 2592 22612 2644
rect 24216 2592 24268 2644
rect 25412 2592 25464 2644
rect 18328 2524 18380 2576
rect 20076 2524 20128 2576
rect 10232 2456 10284 2508
rect 21732 2524 21784 2576
rect 22468 2524 22520 2576
rect 23664 2524 23716 2576
rect 24768 2524 24820 2576
rect 16672 2388 16724 2440
rect 17776 2388 17828 2440
rect 10876 2320 10928 2372
rect 18696 2388 18748 2440
rect 18788 2431 18840 2440
rect 18788 2397 18797 2431
rect 18797 2397 18831 2431
rect 18831 2397 18840 2431
rect 18788 2388 18840 2397
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 19708 2388 19760 2440
rect 20260 2388 20312 2440
rect 20720 2388 20772 2440
rect 21364 2388 21416 2440
rect 21824 2431 21876 2440
rect 21824 2397 21833 2431
rect 21833 2397 21867 2431
rect 21867 2397 21876 2431
rect 21824 2388 21876 2397
rect 22284 2388 22336 2440
rect 22376 2388 22428 2440
rect 24860 2456 24912 2508
rect 21180 2320 21232 2372
rect 23572 2388 23624 2440
rect 24400 2431 24452 2440
rect 24400 2397 24409 2431
rect 24409 2397 24443 2431
rect 24443 2397 24452 2431
rect 24400 2388 24452 2397
rect 24584 2388 24636 2440
rect 25136 2431 25188 2440
rect 25136 2397 25145 2431
rect 25145 2397 25179 2431
rect 25179 2397 25188 2431
rect 25136 2388 25188 2397
rect 25228 2388 25280 2440
rect 26148 2456 26200 2508
rect 27620 2592 27672 2644
rect 29736 2592 29788 2644
rect 31024 2592 31076 2644
rect 31392 2592 31444 2644
rect 26056 2388 26108 2440
rect 27436 2456 27488 2508
rect 28080 2524 28132 2576
rect 29184 2524 29236 2576
rect 30288 2524 30340 2576
rect 31484 2524 31536 2576
rect 39396 2567 39448 2576
rect 39396 2533 39405 2567
rect 39405 2533 39439 2567
rect 39439 2533 39448 2567
rect 39396 2524 39448 2533
rect 24308 2320 24360 2372
rect 27896 2388 27948 2440
rect 17868 2295 17920 2304
rect 17868 2261 17877 2295
rect 17877 2261 17911 2295
rect 17911 2261 17920 2295
rect 17868 2252 17920 2261
rect 18420 2252 18472 2304
rect 18696 2252 18748 2304
rect 19248 2252 19300 2304
rect 19800 2252 19852 2304
rect 20076 2252 20128 2304
rect 20352 2295 20404 2304
rect 20352 2261 20361 2295
rect 20361 2261 20395 2295
rect 20395 2261 20404 2295
rect 20352 2252 20404 2261
rect 20628 2252 20680 2304
rect 20904 2252 20956 2304
rect 21364 2252 21416 2304
rect 21548 2252 21600 2304
rect 22192 2252 22244 2304
rect 22836 2252 22888 2304
rect 23940 2252 23992 2304
rect 26884 2320 26936 2372
rect 26056 2295 26108 2304
rect 26056 2261 26065 2295
rect 26065 2261 26099 2295
rect 26099 2261 26108 2295
rect 26056 2252 26108 2261
rect 26240 2252 26292 2304
rect 26516 2252 26568 2304
rect 28172 2388 28224 2440
rect 28448 2431 28500 2440
rect 28448 2397 28457 2431
rect 28457 2397 28491 2431
rect 28491 2397 28500 2431
rect 28448 2388 28500 2397
rect 28632 2388 28684 2440
rect 30012 2388 30064 2440
rect 30196 2431 30248 2440
rect 30196 2397 30205 2431
rect 30205 2397 30239 2431
rect 30239 2397 30248 2431
rect 30196 2388 30248 2397
rect 30656 2388 30708 2440
rect 31760 2456 31812 2508
rect 32036 2456 32088 2508
rect 29460 2320 29512 2372
rect 31392 2431 31444 2440
rect 31392 2397 31401 2431
rect 31401 2397 31435 2431
rect 31435 2397 31444 2431
rect 31392 2388 31444 2397
rect 32128 2431 32180 2440
rect 32128 2397 32137 2431
rect 32137 2397 32171 2431
rect 32171 2397 32180 2431
rect 32128 2388 32180 2397
rect 32496 2431 32548 2440
rect 32496 2397 32505 2431
rect 32505 2397 32539 2431
rect 32539 2397 32548 2431
rect 32496 2388 32548 2397
rect 32864 2431 32916 2440
rect 32864 2397 32873 2431
rect 32873 2397 32907 2431
rect 32907 2397 32916 2431
rect 32864 2388 32916 2397
rect 33416 2388 33468 2440
rect 38476 2431 38528 2440
rect 38476 2397 38485 2431
rect 38485 2397 38519 2431
rect 38519 2397 38528 2431
rect 38476 2388 38528 2397
rect 28724 2252 28776 2304
rect 30564 2252 30616 2304
rect 31852 2320 31904 2372
rect 31944 2320 31996 2372
rect 31668 2252 31720 2304
rect 37924 2295 37976 2304
rect 37924 2261 37933 2295
rect 37933 2261 37967 2295
rect 37967 2261 37976 2295
rect 37924 2252 37976 2261
rect 38292 2295 38344 2304
rect 38292 2261 38301 2295
rect 38301 2261 38335 2295
rect 38335 2261 38344 2295
rect 38292 2252 38344 2261
rect 38660 2295 38712 2304
rect 38660 2261 38669 2295
rect 38669 2261 38703 2295
rect 38703 2261 38712 2295
rect 38660 2252 38712 2261
rect 38936 2252 38988 2304
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 39010 2150 39062 2202
rect 39074 2150 39126 2202
rect 39138 2150 39190 2202
rect 39202 2150 39254 2202
rect 39266 2150 39318 2202
rect 14280 2048 14332 2100
rect 25136 2048 25188 2100
rect 25504 2048 25556 2100
rect 28172 2048 28224 2100
rect 9772 1980 9824 2032
rect 11428 1912 11480 1964
rect 23204 1980 23256 2032
rect 33416 2048 33468 2100
rect 28448 1980 28500 2032
rect 32036 1980 32088 2032
rect 38476 2048 38528 2100
rect 21916 1912 21968 1964
rect 22376 1844 22428 1896
rect 25320 1844 25372 1896
rect 26240 1844 26292 1896
rect 27252 1844 27304 1896
rect 27620 1844 27672 1896
rect 20720 1776 20772 1828
rect 23020 1776 23072 1828
rect 28448 1776 28500 1828
rect 28632 1912 28684 1964
rect 32128 1912 32180 1964
rect 32772 1912 32824 1964
rect 33048 1912 33100 1964
rect 16120 1708 16172 1760
rect 24584 1708 24636 1760
rect 15384 1640 15436 1692
rect 27988 1708 28040 1760
rect 38936 1912 38988 1964
rect 27528 1640 27580 1692
rect 27896 1640 27948 1692
rect 14924 1572 14976 1624
rect 25228 1572 25280 1624
rect 20812 1504 20864 1556
rect 24400 1504 24452 1556
rect 25044 1504 25096 1556
rect 26056 1504 26108 1556
rect 22652 1436 22704 1488
rect 26424 1368 26476 1420
rect 32864 1640 32916 1692
rect 15108 1300 15160 1352
rect 22928 1300 22980 1352
rect 28816 1300 28868 1352
rect 35256 1300 35308 1352
rect 4252 1232 4304 1284
rect 6000 1232 6052 1284
rect 26792 1232 26844 1284
rect 32496 1232 32548 1284
rect 14004 484 14056 536
rect 23480 484 23532 536
rect 25412 484 25464 536
rect 33600 484 33652 536
rect 14280 416 14332 468
rect 23756 416 23808 468
rect 25688 416 25740 468
rect 36084 416 36136 468
rect 13452 348 13504 400
rect 24952 348 25004 400
rect 27712 348 27764 400
rect 36360 348 36412 400
rect 15936 280 15988 332
rect 29920 280 29972 332
rect 16488 212 16540 264
rect 29828 212 29880 264
rect 15108 144 15160 196
rect 15660 144 15712 196
rect 31576 144 31628 196
rect 4436 8 4488 60
rect 10784 8 10836 60
rect 16304 76 16356 128
rect 30380 76 30432 128
rect 32680 8 32732 60
<< metal2 >>
rect 1122 11194 1178 11250
rect 3054 11194 3110 11250
rect 4986 11194 5042 11250
rect 6918 11194 6974 11250
rect 8850 11194 8906 11250
rect 10782 11194 10838 11250
rect 12714 11194 12770 11250
rect 14646 11194 14702 11250
rect 16578 11194 16634 11250
rect 18510 11194 18566 11250
rect 20442 11194 20498 11250
rect 22374 11194 22430 11250
rect 24306 11194 24362 11250
rect 26238 11194 26294 11250
rect 28170 11194 28226 11250
rect 30102 11194 30158 11250
rect 32034 11194 32090 11250
rect 33966 11194 34022 11250
rect 35898 11194 35954 11250
rect 37830 11194 37886 11250
rect 39762 11194 39818 11250
rect 1136 8634 1164 11194
rect 1308 9376 1360 9382
rect 1308 9318 1360 9324
rect 1124 8628 1176 8634
rect 1124 8570 1176 8576
rect 1320 7449 1348 9318
rect 3068 8922 3096 11194
rect 2884 8894 3096 8922
rect 2778 8800 2834 8809
rect 2778 8735 2834 8744
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1306 7440 1362 7449
rect 1306 7375 1362 7384
rect 1596 6730 1624 8434
rect 2792 8401 2820 8735
rect 2884 8634 2912 8894
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 3436 8634 3464 8774
rect 5000 8634 5028 11194
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5368 8498 5396 8774
rect 6932 8634 6960 11194
rect 8864 8634 8892 11194
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 10796 8634 10824 11194
rect 12728 8634 12756 11194
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 13096 8498 13124 8978
rect 14660 8634 14688 11194
rect 14830 9616 14886 9625
rect 14830 9551 14886 9560
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 2778 8392 2834 8401
rect 2778 8327 2834 8336
rect 1766 8256 1822 8265
rect 1766 8191 1822 8200
rect 1780 7857 1808 8191
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 1766 7848 1822 7857
rect 1766 7783 1822 7792
rect 14844 7750 14872 9551
rect 14922 9344 14978 9353
rect 14922 9279 14978 9288
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 14936 7546 14964 9279
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 16592 8634 16620 11194
rect 16856 9104 16908 9110
rect 16856 9046 16908 9052
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16868 8498 16896 9046
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 16960 8498 16988 8910
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16580 8424 16632 8430
rect 16486 8392 16542 8401
rect 16580 8366 16632 8372
rect 16486 8327 16542 8336
rect 16500 8090 16528 8327
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16120 7948 16172 7954
rect 16120 7890 16172 7896
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 16132 7478 16160 7890
rect 16396 7880 16448 7886
rect 16394 7848 16396 7857
rect 16448 7848 16450 7857
rect 16592 7818 16620 8366
rect 17132 8016 17184 8022
rect 17132 7958 17184 7964
rect 16394 7783 16450 7792
rect 16580 7812 16632 7818
rect 16580 7754 16632 7760
rect 16120 7472 16172 7478
rect 15106 7440 15162 7449
rect 16120 7414 16172 7420
rect 15106 7375 15108 7384
rect 15160 7375 15162 7384
rect 15108 7346 15160 7352
rect 16488 7336 16540 7342
rect 16486 7304 16488 7313
rect 16540 7304 16542 7313
rect 16486 7239 16542 7248
rect 17144 7206 17172 7958
rect 17776 7744 17828 7750
rect 17776 7686 17828 7692
rect 17788 7410 17816 7686
rect 17972 7546 18000 8842
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18156 7546 18184 8774
rect 18524 8634 18552 11194
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 18694 9072 18750 9081
rect 18694 9007 18750 9016
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18328 7948 18380 7954
rect 18328 7890 18380 7896
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 18144 7540 18196 7546
rect 18144 7482 18196 7488
rect 18340 7410 18368 7890
rect 18708 7546 18736 9007
rect 18892 8498 18920 9114
rect 20352 8832 20404 8838
rect 20352 8774 20404 8780
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 19950 8188 20258 8197
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 18892 7546 18920 8026
rect 19062 7984 19118 7993
rect 19062 7919 19118 7928
rect 19076 7750 19104 7919
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 19260 7546 19288 8026
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19340 7812 19392 7818
rect 19340 7754 19392 7760
rect 19352 7546 19380 7754
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19996 7410 20024 7822
rect 20364 7546 20392 8774
rect 20456 8634 20484 11194
rect 20720 9308 20772 9314
rect 20720 9250 20772 9256
rect 20444 8628 20496 8634
rect 20444 8570 20496 8576
rect 20444 7744 20496 7750
rect 20444 7686 20496 7692
rect 20456 7546 20484 7686
rect 20732 7546 20760 9250
rect 20812 9240 20864 9246
rect 20812 9182 20864 9188
rect 20824 7546 20852 9182
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 22388 8634 22416 11194
rect 22558 9888 22614 9897
rect 22558 9823 22614 9832
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 22098 8528 22154 8537
rect 22098 8463 22154 8472
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 20916 7546 20944 7822
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 22112 7546 22140 8463
rect 22192 8356 22244 8362
rect 22192 8298 22244 8304
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 22100 7540 22152 7546
rect 22100 7482 22152 7488
rect 17776 7404 17828 7410
rect 17776 7346 17828 7352
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 19616 7404 19668 7410
rect 19616 7346 19668 7352
rect 19984 7404 20036 7410
rect 19984 7346 20036 7352
rect 17788 7206 17816 7346
rect 19628 7206 19656 7346
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 19616 7200 19668 7206
rect 19616 7142 19668 7148
rect 19800 7200 19852 7206
rect 19800 7142 19852 7148
rect 21364 7200 21416 7206
rect 21364 7142 21416 7148
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 19812 7002 19840 7142
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 19800 6996 19852 7002
rect 19800 6938 19852 6944
rect 21376 6934 21404 7142
rect 9128 6928 9180 6934
rect 17868 6928 17920 6934
rect 9128 6870 9180 6876
rect 17498 6896 17554 6905
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 1584 6724 1636 6730
rect 1584 6666 1636 6672
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 570 5536 626 5545
rect 570 5471 626 5480
rect 584 3670 612 5471
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 2778 5128 2834 5137
rect 2778 5063 2834 5072
rect 1766 4992 1822 5001
rect 1766 4927 1822 4936
rect 1780 4593 1808 4927
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 1766 4584 1822 4593
rect 1766 4519 1822 4528
rect 2792 4457 2820 5063
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2778 4448 2834 4457
rect 2778 4383 2834 4392
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 572 3664 624 3670
rect 572 3606 624 3612
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2884 42 2912 4558
rect 3068 4554 3096 4966
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 3160 56 3280 82
rect 3528 56 3556 5170
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 3792 5092 3844 5098
rect 3792 5034 3844 5040
rect 3804 56 3832 5034
rect 4080 56 4108 5102
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4264 1290 4292 4558
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4356 4214 4384 4422
rect 4344 4208 4396 4214
rect 4344 4150 4396 4156
rect 4252 1284 4304 1290
rect 4252 1226 4304 1232
rect 4356 66 4476 82
rect 4356 60 4488 66
rect 4356 56 4436 60
rect 3160 54 3294 56
rect 3160 42 3188 54
rect 2884 14 3188 42
rect 3238 0 3294 54
rect 3514 0 3570 56
rect 3790 0 3846 56
rect 4066 0 4122 56
rect 4342 54 4436 56
rect 4342 0 4398 54
rect 4632 56 4660 6598
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 4988 5636 5040 5642
rect 4988 5578 5040 5584
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 4908 4282 4936 4694
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 3126 4936 3878
rect 4896 3120 4948 3126
rect 4896 3062 4948 3068
rect 5000 2774 5028 5578
rect 4908 2746 5028 2774
rect 4908 56 4936 2746
rect 5184 56 5212 5646
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5368 4690 5396 4966
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5460 56 5488 5170
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5552 1465 5580 4966
rect 6104 4826 6132 5306
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5538 1456 5594 1465
rect 5538 1391 5594 1400
rect 5736 56 5764 4558
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6000 1284 6052 1290
rect 6000 1226 6052 1232
rect 6012 56 6040 1226
rect 6288 56 6316 4082
rect 6564 56 6592 6394
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6840 56 6868 5510
rect 7116 56 7144 5714
rect 7392 56 7420 6190
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7668 56 7696 6054
rect 7760 2650 7788 6802
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 7852 2530 7880 6734
rect 9140 6662 9168 6870
rect 10784 6860 10836 6866
rect 17868 6870 17920 6876
rect 21364 6928 21416 6934
rect 21364 6870 21416 6876
rect 17498 6831 17500 6840
rect 10784 6802 10836 6808
rect 17552 6831 17554 6840
rect 17500 6802 17552 6808
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 9416 6458 9444 6598
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9128 6384 9180 6390
rect 9128 6326 9180 6332
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 7852 2502 7972 2530
rect 7944 56 7972 2502
rect 8220 56 8248 2586
rect 8496 56 8524 6258
rect 9140 6118 9168 6326
rect 9508 6118 9536 6598
rect 9600 6390 9628 6734
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9678 6488 9734 6497
rect 9678 6423 9734 6432
rect 9588 6384 9640 6390
rect 9588 6326 9640 6332
rect 9692 6202 9720 6423
rect 9600 6174 9720 6202
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 9600 5370 9628 6174
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8680 2553 8708 4558
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8666 2544 8722 2553
rect 8666 2479 8722 2488
rect 8758 1592 8814 1601
rect 8758 1527 8814 1536
rect 8772 56 8800 1527
rect 4436 2 4488 8
rect 4618 0 4674 56
rect 4894 0 4950 56
rect 5170 0 5226 56
rect 5446 0 5502 56
rect 5722 0 5778 56
rect 5998 0 6054 56
rect 6274 0 6330 56
rect 6550 0 6606 56
rect 6826 0 6882 56
rect 7102 0 7158 56
rect 7378 0 7434 56
rect 7654 0 7710 56
rect 7930 0 7986 56
rect 8206 0 8262 56
rect 8482 0 8538 56
rect 8758 0 8814 56
rect 8864 42 8892 3130
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 9416 1986 9444 4014
rect 9324 1958 9444 1986
rect 8956 56 9076 82
rect 9324 56 9352 1958
rect 9508 1578 9536 4082
rect 9692 3466 9720 4218
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9588 2916 9640 2922
rect 9588 2858 9640 2864
rect 9600 1737 9628 2858
rect 9784 2038 9812 6598
rect 9968 6254 9996 6734
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9876 4282 9904 4558
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9862 2272 9918 2281
rect 9862 2207 9918 2216
rect 9772 2032 9824 2038
rect 9772 1974 9824 1980
rect 9586 1728 9642 1737
rect 9586 1663 9642 1672
rect 9508 1550 9628 1578
rect 9600 56 9628 1550
rect 9876 56 9904 2207
rect 10152 56 10180 5238
rect 10244 2514 10272 6598
rect 10520 5778 10548 6734
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 10428 56 10456 5170
rect 10704 4706 10732 6598
rect 10612 4678 10732 4706
rect 10612 2582 10640 4678
rect 10692 4004 10744 4010
rect 10692 3946 10744 3952
rect 10600 2576 10652 2582
rect 10600 2518 10652 2524
rect 10704 56 10732 3946
rect 10796 66 10824 6802
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 11704 6792 11756 6798
rect 17880 6769 17908 6870
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 11704 6734 11756 6740
rect 17406 6760 17462 6769
rect 10888 5574 10916 6734
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 11256 6361 11284 6598
rect 11058 6352 11114 6361
rect 11058 6287 11114 6296
rect 11242 6352 11298 6361
rect 11242 6287 11298 6296
rect 10966 5672 11022 5681
rect 10966 5607 11022 5616
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10888 2378 10916 4150
rect 10980 4010 11008 5607
rect 11072 5370 11100 6287
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 11072 3534 11100 4422
rect 11164 4214 11192 4966
rect 11152 4208 11204 4214
rect 11152 4150 11204 4156
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 10876 2372 10928 2378
rect 10876 2314 10928 2320
rect 10784 60 10836 66
rect 8956 54 9090 56
rect 8956 42 8984 54
rect 8864 14 8984 42
rect 9034 0 9090 54
rect 9310 0 9366 56
rect 9586 0 9642 56
rect 9862 0 9918 56
rect 10138 0 10194 56
rect 10414 0 10470 56
rect 10690 0 10746 56
rect 10980 56 11008 2586
rect 11256 56 11284 5646
rect 11440 1970 11468 6598
rect 11520 6384 11572 6390
rect 11520 6326 11572 6332
rect 11428 1964 11480 1970
rect 11428 1906 11480 1912
rect 11532 56 11560 6326
rect 11716 6322 11744 6734
rect 17406 6695 17462 6704
rect 17866 6760 17922 6769
rect 17866 6695 17922 6704
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11808 56 11836 6258
rect 11900 4026 11928 6598
rect 11992 5914 12020 6598
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 14830 6488 14886 6497
rect 15010 6491 15318 6500
rect 14830 6423 14886 6432
rect 12072 6248 12124 6254
rect 12072 6190 12124 6196
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11900 3998 12020 4026
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11900 2417 11928 3878
rect 11992 2990 12020 3998
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 11886 2408 11942 2417
rect 11886 2343 11942 2352
rect 12084 56 12112 6190
rect 14016 6118 14044 6190
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14280 6112 14332 6118
rect 14844 6089 14872 6423
rect 14924 6112 14976 6118
rect 14280 6054 14332 6060
rect 14830 6080 14886 6089
rect 13648 5914 13676 6054
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12544 4162 12572 5714
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 12624 5636 12676 5642
rect 12624 5578 12676 5584
rect 12360 4134 12572 4162
rect 12360 56 12388 4134
rect 12636 56 12664 5578
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 12912 56 12940 5102
rect 13174 1864 13230 1873
rect 13174 1799 13230 1808
rect 13188 56 13216 1799
rect 13648 1737 13676 5510
rect 13740 2650 13768 5646
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 14292 2106 14320 6054
rect 14924 6054 14976 6060
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 14830 6015 14886 6024
rect 14556 5704 14608 5710
rect 14554 5672 14556 5681
rect 14608 5672 14610 5681
rect 14554 5607 14610 5616
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14384 2553 14412 5510
rect 14370 2544 14426 2553
rect 14370 2479 14426 2488
rect 14280 2100 14332 2106
rect 14280 2042 14332 2048
rect 13634 1728 13690 1737
rect 13634 1663 13690 1672
rect 14936 1630 14964 6054
rect 15028 5914 15056 6054
rect 17420 5914 17448 6695
rect 17960 6384 18012 6390
rect 17960 6326 18012 6332
rect 15016 5908 15068 5914
rect 15016 5850 15068 5856
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 16120 5840 16172 5846
rect 16120 5782 16172 5788
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 15580 4758 15608 4966
rect 15568 4752 15620 4758
rect 15568 4694 15620 4700
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 15010 3227 15318 3236
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 15106 2000 15162 2009
rect 15106 1935 15162 1944
rect 15290 2000 15346 2009
rect 15290 1935 15346 1944
rect 14924 1624 14976 1630
rect 14924 1566 14976 1572
rect 15120 1358 15148 1935
rect 15304 1737 15332 1935
rect 16132 1766 16160 5782
rect 17972 5370 18000 6326
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16592 2417 16620 4558
rect 16684 2446 16712 4762
rect 17776 4684 17828 4690
rect 17776 4626 17828 4632
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 17144 3602 17172 3878
rect 17132 3596 17184 3602
rect 17132 3538 17184 3544
rect 17314 3360 17370 3369
rect 17314 3295 17370 3304
rect 17038 3224 17094 3233
rect 17038 3159 17094 3168
rect 16672 2440 16724 2446
rect 16578 2408 16634 2417
rect 16672 2382 16724 2388
rect 16762 2408 16818 2417
rect 16578 2343 16634 2352
rect 16762 2343 16818 2352
rect 16120 1760 16172 1766
rect 15290 1728 15346 1737
rect 16120 1702 16172 1708
rect 15290 1663 15346 1672
rect 15384 1692 15436 1698
rect 15384 1634 15436 1640
rect 15108 1352 15160 1358
rect 15108 1294 15160 1300
rect 14004 536 14056 542
rect 14004 478 14056 484
rect 13452 400 13504 406
rect 13452 342 13504 348
rect 13726 368 13782 377
rect 13464 56 13492 342
rect 13726 303 13782 312
rect 13740 56 13768 303
rect 14016 56 14044 478
rect 14280 468 14332 474
rect 14280 410 14332 416
rect 14292 56 14320 410
rect 14554 232 14610 241
rect 14554 167 14610 176
rect 15108 196 15160 202
rect 14568 56 14596 167
rect 15108 138 15160 144
rect 14830 96 14886 105
rect 10784 2 10836 8
rect 10966 0 11022 56
rect 11242 0 11298 56
rect 11518 0 11574 56
rect 11794 0 11850 56
rect 12070 0 12126 56
rect 12346 0 12402 56
rect 12622 0 12678 56
rect 12898 0 12954 56
rect 13174 0 13230 56
rect 13450 0 13506 56
rect 13726 0 13782 56
rect 14002 0 14058 56
rect 14278 0 14334 56
rect 14554 0 14610 56
rect 15120 56 15148 138
rect 15396 56 15424 1634
rect 15936 332 15988 338
rect 15936 274 15988 280
rect 15660 196 15712 202
rect 15660 138 15712 144
rect 15672 56 15700 138
rect 15948 56 15976 274
rect 16488 264 16540 270
rect 16488 206 16540 212
rect 16304 128 16356 134
rect 16224 76 16304 82
rect 16224 70 16356 76
rect 16224 56 16344 70
rect 16500 56 16528 206
rect 16776 56 16804 2343
rect 17052 56 17080 3159
rect 17328 56 17356 3295
rect 17788 2446 17816 4626
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 17972 3058 18000 4490
rect 18236 3528 18288 3534
rect 18288 3476 18368 3482
rect 18236 3470 18368 3476
rect 18248 3454 18368 3470
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 18248 3194 18276 3334
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18340 3058 18368 3454
rect 17960 3052 18012 3058
rect 17960 2994 18012 3000
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 17880 56 17908 2246
rect 18156 56 18184 2790
rect 18432 2774 18460 6802
rect 22204 6662 22232 8298
rect 22468 7948 22520 7954
rect 22468 7890 22520 7896
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18340 2746 18460 2774
rect 18340 2582 18368 2746
rect 18328 2576 18380 2582
rect 18328 2518 18380 2524
rect 18420 2304 18472 2310
rect 18420 2246 18472 2252
rect 18432 56 18460 2246
rect 18524 1601 18552 3470
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18616 3194 18644 3334
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18708 2446 18736 6598
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 22284 6452 22336 6458
rect 22284 6394 22336 6400
rect 21364 6248 21416 6254
rect 21364 6190 21416 6196
rect 20720 6180 20772 6186
rect 20720 6122 20772 6128
rect 19338 6080 19394 6089
rect 19338 6015 19394 6024
rect 19352 5386 19380 6015
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 19798 5808 19854 5817
rect 19536 5766 19748 5794
rect 19536 5710 19564 5766
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19614 5672 19670 5681
rect 19614 5607 19670 5616
rect 19260 5358 19380 5386
rect 19154 5264 19210 5273
rect 19154 5199 19210 5208
rect 19168 3738 19196 5199
rect 19156 3732 19208 3738
rect 19156 3674 19208 3680
rect 19168 3534 19196 3674
rect 19156 3528 19208 3534
rect 19156 3470 19208 3476
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 18800 2446 18828 2994
rect 19260 2972 19288 5358
rect 19338 5264 19394 5273
rect 19338 5199 19394 5208
rect 19352 3482 19380 5199
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19444 3670 19472 4082
rect 19628 3942 19656 5607
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19616 3936 19668 3942
rect 19616 3878 19668 3884
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 19536 3534 19564 3878
rect 19524 3528 19576 3534
rect 19352 3454 19472 3482
rect 19524 3470 19576 3476
rect 19444 3398 19472 3454
rect 19616 3460 19668 3466
rect 19616 3402 19668 3408
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19352 3126 19380 3334
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 19628 3058 19656 3402
rect 19616 3052 19668 3058
rect 19616 2994 19668 3000
rect 19260 2944 19472 2972
rect 18972 2848 19024 2854
rect 18972 2790 19024 2796
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 18510 1592 18566 1601
rect 18510 1527 18566 1536
rect 18708 56 18736 2246
rect 18984 56 19012 2790
rect 19444 2446 19472 2944
rect 19524 2848 19576 2854
rect 19524 2790 19576 2796
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19248 2304 19300 2310
rect 19248 2246 19300 2252
rect 19260 56 19288 2246
rect 19536 56 19564 2790
rect 19720 2446 19748 5766
rect 19798 5743 19854 5752
rect 19812 4690 19840 5743
rect 20444 5636 20496 5642
rect 20444 5578 20496 5584
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 19800 4684 19852 4690
rect 19800 4626 19852 4632
rect 20456 4486 20484 5578
rect 20444 4480 20496 4486
rect 20444 4422 20496 4428
rect 20626 4040 20682 4049
rect 20626 3975 20682 3984
rect 20442 3904 20498 3913
rect 19950 3836 20258 3845
rect 20442 3839 20498 3848
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 20350 3768 20406 3777
rect 20350 3703 20406 3712
rect 20364 3369 20392 3703
rect 20350 3360 20406 3369
rect 20350 3295 20406 3304
rect 20456 3233 20484 3839
rect 20442 3224 20498 3233
rect 20442 3159 20498 3168
rect 20640 2961 20668 3975
rect 20732 3670 20760 6122
rect 20812 5772 20864 5778
rect 20812 5714 20864 5720
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 20626 2952 20682 2961
rect 20626 2887 20682 2896
rect 19950 2748 20258 2757
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 20076 2576 20128 2582
rect 20076 2518 20128 2524
rect 19708 2440 19760 2446
rect 20088 2428 20116 2518
rect 20260 2440 20312 2446
rect 20088 2400 20260 2428
rect 19708 2382 19760 2388
rect 20260 2382 20312 2388
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 19800 2304 19852 2310
rect 19800 2246 19852 2252
rect 20076 2304 20128 2310
rect 20076 2246 20128 2252
rect 20352 2304 20404 2310
rect 20352 2246 20404 2252
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 19812 56 19840 2246
rect 20088 56 20116 2246
rect 20364 56 20392 2246
rect 20640 56 20668 2246
rect 20732 1834 20760 2382
rect 20720 1828 20772 1834
rect 20720 1770 20772 1776
rect 20824 1562 20852 5714
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 21180 2644 21232 2650
rect 21180 2586 21232 2592
rect 21192 2378 21220 2586
rect 21376 2446 21404 6190
rect 21824 6112 21876 6118
rect 21824 6054 21876 6060
rect 21732 5092 21784 5098
rect 21732 5034 21784 5040
rect 21744 4826 21772 5034
rect 21732 4820 21784 4826
rect 21732 4762 21784 4768
rect 21546 4584 21602 4593
rect 21546 4519 21602 4528
rect 21560 4146 21588 4519
rect 21732 4208 21784 4214
rect 21732 4150 21784 4156
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 21744 3534 21772 4150
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 21732 2576 21784 2582
rect 21732 2518 21784 2524
rect 21364 2440 21416 2446
rect 21364 2382 21416 2388
rect 21180 2372 21232 2378
rect 21180 2314 21232 2320
rect 20904 2304 20956 2310
rect 20904 2246 20956 2252
rect 21364 2304 21416 2310
rect 21548 2304 21600 2310
rect 21364 2246 21416 2252
rect 21468 2264 21548 2292
rect 20812 1556 20864 1562
rect 20812 1498 20864 1504
rect 20916 56 20944 2246
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 21192 56 21312 82
rect 14830 0 14886 40
rect 15106 0 15162 56
rect 15382 0 15438 56
rect 15658 0 15714 56
rect 15934 0 15990 56
rect 16210 54 16344 56
rect 16210 0 16266 54
rect 16486 0 16542 56
rect 16762 0 16818 56
rect 17038 0 17094 56
rect 17314 0 17370 56
rect 17590 0 17646 56
rect 17866 0 17922 56
rect 18142 0 18198 56
rect 18418 0 18474 56
rect 18694 0 18750 56
rect 18970 0 19026 56
rect 19246 0 19302 56
rect 19522 0 19578 56
rect 19798 0 19854 56
rect 20074 0 20130 56
rect 20350 0 20406 56
rect 20626 0 20682 56
rect 20902 0 20958 56
rect 21178 54 21312 56
rect 21178 0 21234 54
rect 21284 42 21312 54
rect 21376 42 21404 2246
rect 21468 56 21496 2264
rect 21548 2246 21600 2252
rect 21744 56 21772 2518
rect 21836 2446 21864 6054
rect 22008 5364 22060 5370
rect 22008 5306 22060 5312
rect 21916 4276 21968 4282
rect 21916 4218 21968 4224
rect 21928 3738 21956 4218
rect 22020 4010 22048 5306
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22008 4004 22060 4010
rect 22008 3946 22060 3952
rect 21916 3732 21968 3738
rect 21916 3674 21968 3680
rect 21916 3392 21968 3398
rect 21916 3334 21968 3340
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 21928 1970 21956 3334
rect 22112 2961 22140 4082
rect 22098 2952 22154 2961
rect 22098 2887 22154 2896
rect 22008 2644 22060 2650
rect 22008 2586 22060 2592
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 21916 1964 21968 1970
rect 21916 1906 21968 1912
rect 22020 56 22048 2586
rect 22204 2310 22232 2586
rect 22296 2446 22324 6394
rect 22374 6216 22430 6225
rect 22374 6151 22430 6160
rect 22388 5234 22416 6151
rect 22376 5228 22428 5234
rect 22376 5170 22428 5176
rect 22480 5114 22508 7890
rect 22572 7546 22600 9823
rect 23020 9376 23072 9382
rect 23020 9318 23072 9324
rect 22744 8492 22796 8498
rect 22744 8434 22796 8440
rect 22756 8362 22784 8434
rect 22744 8356 22796 8362
rect 22744 8298 22796 8304
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 23032 7410 23060 9318
rect 24320 8634 24348 11194
rect 25780 9240 25832 9246
rect 25780 9182 25832 9188
rect 24308 8628 24360 8634
rect 24308 8570 24360 8576
rect 24676 8492 24728 8498
rect 24676 8434 24728 8440
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 23204 8016 23256 8022
rect 23204 7958 23256 7964
rect 23216 7410 23244 7958
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 23204 7404 23256 7410
rect 23204 7346 23256 7352
rect 22928 7336 22980 7342
rect 22928 7278 22980 7284
rect 22940 6186 22968 7278
rect 23124 7274 23336 7290
rect 23112 7268 23348 7274
rect 23164 7262 23296 7268
rect 23112 7210 23164 7216
rect 23296 7210 23348 7216
rect 24688 6458 24716 8434
rect 24780 7206 24808 8434
rect 25412 8424 25464 8430
rect 25412 8366 25464 8372
rect 25596 8424 25648 8430
rect 25596 8366 25648 8372
rect 25424 7750 25452 8366
rect 25412 7744 25464 7750
rect 25412 7686 25464 7692
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 24768 7200 24820 7206
rect 24768 7142 24820 7148
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 23570 6352 23626 6361
rect 23570 6287 23626 6296
rect 22928 6180 22980 6186
rect 22928 6122 22980 6128
rect 22388 5086 22508 5114
rect 23478 5128 23534 5137
rect 23204 5092 23256 5098
rect 22388 2774 22416 5086
rect 23478 5063 23534 5072
rect 23204 5034 23256 5040
rect 22468 5024 22520 5030
rect 22468 4966 22520 4972
rect 22480 2990 22508 4966
rect 23216 4826 23244 5034
rect 23492 4826 23520 5063
rect 23204 4820 23256 4826
rect 23204 4762 23256 4768
rect 23480 4820 23532 4826
rect 23480 4762 23532 4768
rect 22834 4720 22890 4729
rect 22834 4655 22836 4664
rect 22888 4655 22890 4664
rect 22836 4626 22888 4632
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 22560 3392 22612 3398
rect 22560 3334 22612 3340
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 22468 2984 22520 2990
rect 22468 2926 22520 2932
rect 22572 2774 22600 3334
rect 22664 2922 22692 3334
rect 22756 3126 22784 3674
rect 22836 3664 22888 3670
rect 22836 3606 22888 3612
rect 23112 3664 23164 3670
rect 23112 3606 23164 3612
rect 22848 3126 22876 3606
rect 23124 3534 23152 3606
rect 23112 3528 23164 3534
rect 22940 3488 23112 3516
rect 22744 3120 22796 3126
rect 22744 3062 22796 3068
rect 22836 3120 22888 3126
rect 22836 3062 22888 3068
rect 22652 2916 22704 2922
rect 22652 2858 22704 2864
rect 22388 2746 22508 2774
rect 22572 2746 22692 2774
rect 22480 2689 22508 2746
rect 22466 2680 22522 2689
rect 22466 2615 22522 2624
rect 22560 2644 22612 2650
rect 22560 2586 22612 2592
rect 22468 2576 22520 2582
rect 22468 2518 22520 2524
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 22376 2440 22428 2446
rect 22376 2382 22428 2388
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 22388 1902 22416 2382
rect 22376 1896 22428 1902
rect 22376 1838 22428 1844
rect 22296 56 22416 82
rect 21284 14 21404 42
rect 21454 0 21510 56
rect 21730 0 21786 56
rect 22006 0 22062 56
rect 22282 54 22416 56
rect 22282 0 22338 54
rect 22388 42 22416 54
rect 22480 42 22508 2518
rect 22572 56 22600 2586
rect 22664 1494 22692 2746
rect 22742 2680 22798 2689
rect 22742 2615 22798 2624
rect 22756 1737 22784 2615
rect 22836 2304 22888 2310
rect 22836 2246 22888 2252
rect 22742 1728 22798 1737
rect 22742 1663 22798 1672
rect 22652 1488 22704 1494
rect 22652 1430 22704 1436
rect 22848 56 22876 2246
rect 22940 1358 22968 3488
rect 23112 3470 23164 3476
rect 23480 3460 23532 3466
rect 23480 3402 23532 3408
rect 23020 3392 23072 3398
rect 23020 3334 23072 3340
rect 23204 3392 23256 3398
rect 23204 3334 23256 3340
rect 23032 1834 23060 3334
rect 23112 2848 23164 2854
rect 23112 2790 23164 2796
rect 23020 1828 23072 1834
rect 23020 1770 23072 1776
rect 22928 1352 22980 1358
rect 22928 1294 22980 1300
rect 23124 56 23152 2790
rect 23216 2038 23244 3334
rect 23296 3188 23348 3194
rect 23296 3130 23348 3136
rect 23388 3188 23440 3194
rect 23388 3130 23440 3136
rect 23308 2922 23336 3130
rect 23296 2916 23348 2922
rect 23296 2858 23348 2864
rect 23204 2032 23256 2038
rect 23204 1974 23256 1980
rect 23400 56 23428 3130
rect 23492 2990 23520 3402
rect 23480 2984 23532 2990
rect 23480 2926 23532 2932
rect 23480 2848 23532 2854
rect 23480 2790 23532 2796
rect 23492 542 23520 2790
rect 23584 2446 23612 6287
rect 24860 5568 24912 5574
rect 24860 5510 24912 5516
rect 24124 5296 24176 5302
rect 24124 5238 24176 5244
rect 23756 4820 23808 4826
rect 23756 4762 23808 4768
rect 23664 4208 23716 4214
rect 23664 4150 23716 4156
rect 23676 2854 23704 4150
rect 23664 2848 23716 2854
rect 23664 2790 23716 2796
rect 23664 2576 23716 2582
rect 23664 2518 23716 2524
rect 23572 2440 23624 2446
rect 23572 2382 23624 2388
rect 23480 536 23532 542
rect 23480 478 23532 484
rect 23676 56 23704 2518
rect 23768 474 23796 4762
rect 24032 4616 24084 4622
rect 24032 4558 24084 4564
rect 24044 4185 24072 4558
rect 24030 4176 24086 4185
rect 24030 4111 24086 4120
rect 24136 3516 24164 5238
rect 24216 4480 24268 4486
rect 24216 4422 24268 4428
rect 24228 4282 24256 4422
rect 24216 4276 24268 4282
rect 24216 4218 24268 4224
rect 24216 3936 24268 3942
rect 24216 3878 24268 3884
rect 24228 3641 24256 3878
rect 24308 3732 24360 3738
rect 24308 3674 24360 3680
rect 24400 3732 24452 3738
rect 24400 3674 24452 3680
rect 24214 3632 24270 3641
rect 24214 3567 24270 3576
rect 24136 3488 24256 3516
rect 24124 3392 24176 3398
rect 24124 3334 24176 3340
rect 24136 3097 24164 3334
rect 24122 3088 24178 3097
rect 24122 3023 24178 3032
rect 24228 2774 24256 3488
rect 24320 3194 24348 3674
rect 24412 3534 24440 3674
rect 24400 3528 24452 3534
rect 24398 3496 24400 3505
rect 24452 3496 24454 3505
rect 24398 3431 24454 3440
rect 24768 3460 24820 3466
rect 24768 3402 24820 3408
rect 24780 3194 24808 3402
rect 24308 3188 24360 3194
rect 24308 3130 24360 3136
rect 24768 3188 24820 3194
rect 24768 3130 24820 3136
rect 24872 3058 24900 5510
rect 25044 4752 25096 4758
rect 25044 4694 25096 4700
rect 24952 3528 25004 3534
rect 24952 3470 25004 3476
rect 24860 3052 24912 3058
rect 24860 2994 24912 3000
rect 24492 2848 24544 2854
rect 24964 2825 24992 3470
rect 24492 2790 24544 2796
rect 24950 2816 25006 2825
rect 24228 2746 24348 2774
rect 24216 2644 24268 2650
rect 24216 2586 24268 2592
rect 23940 2304 23992 2310
rect 23940 2246 23992 2252
rect 23756 468 23808 474
rect 23756 410 23808 416
rect 23952 56 23980 2246
rect 24228 56 24256 2586
rect 24320 2378 24348 2746
rect 24400 2440 24452 2446
rect 24400 2382 24452 2388
rect 24308 2372 24360 2378
rect 24308 2314 24360 2320
rect 24412 1562 24440 2382
rect 24400 1556 24452 1562
rect 24400 1498 24452 1504
rect 24504 56 24532 2790
rect 24950 2751 25006 2760
rect 24768 2576 24820 2582
rect 24768 2518 24820 2524
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24596 1766 24624 2382
rect 24584 1760 24636 1766
rect 24584 1702 24636 1708
rect 24780 56 24808 2518
rect 24860 2508 24912 2514
rect 25056 2496 25084 4694
rect 25240 2530 25268 7346
rect 25608 4486 25636 8366
rect 25688 4616 25740 4622
rect 25688 4558 25740 4564
rect 25596 4480 25648 4486
rect 25596 4422 25648 4428
rect 25412 4140 25464 4146
rect 25412 4082 25464 4088
rect 25424 2650 25452 4082
rect 25504 2916 25556 2922
rect 25504 2858 25556 2864
rect 25412 2644 25464 2650
rect 25412 2586 25464 2592
rect 25240 2502 25452 2530
rect 24860 2450 24912 2456
rect 24964 2468 25084 2496
rect 24872 2009 24900 2450
rect 24858 2000 24914 2009
rect 24858 1935 24914 1944
rect 24964 406 24992 2468
rect 25136 2440 25188 2446
rect 25136 2382 25188 2388
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 25148 2106 25176 2382
rect 25136 2100 25188 2106
rect 25136 2042 25188 2048
rect 25240 1630 25268 2382
rect 25320 1896 25372 1902
rect 25320 1838 25372 1844
rect 25228 1624 25280 1630
rect 25228 1566 25280 1572
rect 25044 1556 25096 1562
rect 25044 1498 25096 1504
rect 24952 400 25004 406
rect 24952 342 25004 348
rect 25056 56 25084 1498
rect 25332 56 25360 1838
rect 25424 542 25452 2502
rect 25516 2106 25544 2858
rect 25596 2848 25648 2854
rect 25596 2790 25648 2796
rect 25504 2100 25556 2106
rect 25504 2042 25556 2048
rect 25412 536 25464 542
rect 25412 478 25464 484
rect 25608 56 25636 2790
rect 25700 474 25728 4558
rect 25792 3738 25820 9182
rect 26252 8634 26280 11194
rect 27436 9172 27488 9178
rect 27436 9114 27488 9120
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 26240 8628 26292 8634
rect 26240 8570 26292 8576
rect 25872 8560 25924 8566
rect 25872 8502 25924 8508
rect 25884 7206 25912 8502
rect 26332 8492 26384 8498
rect 26332 8434 26384 8440
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 26148 7744 26200 7750
rect 26148 7686 26200 7692
rect 26160 7206 26188 7686
rect 25872 7200 25924 7206
rect 25872 7142 25924 7148
rect 26148 7200 26200 7206
rect 26148 7142 26200 7148
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 26344 5914 26372 8434
rect 26884 8356 26936 8362
rect 26884 8298 26936 8304
rect 26896 7478 26924 8298
rect 27448 7750 27476 9114
rect 27804 9104 27856 9110
rect 27804 9046 27856 9052
rect 27528 9036 27580 9042
rect 27528 8978 27580 8984
rect 27436 7744 27488 7750
rect 27436 7686 27488 7692
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 26884 7472 26936 7478
rect 26884 7414 26936 7420
rect 27344 7404 27396 7410
rect 27344 7346 27396 7352
rect 26884 6928 26936 6934
rect 26884 6870 26936 6876
rect 26332 5908 26384 5914
rect 26332 5850 26384 5856
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 26608 4616 26660 4622
rect 26608 4558 26660 4564
rect 25872 4548 25924 4554
rect 25872 4490 25924 4496
rect 25780 3732 25832 3738
rect 25780 3674 25832 3680
rect 25884 3058 25912 4490
rect 26424 4480 26476 4486
rect 26424 4422 26476 4428
rect 26332 3936 26384 3942
rect 26332 3878 26384 3884
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 26344 3641 26372 3878
rect 26330 3632 26386 3641
rect 26330 3567 26386 3576
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 25872 3052 25924 3058
rect 25872 2994 25924 3000
rect 26160 2922 26188 3470
rect 26148 2916 26200 2922
rect 26148 2858 26200 2864
rect 26332 2848 26384 2854
rect 26332 2790 26384 2796
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 26344 2632 26372 2790
rect 25976 2604 26372 2632
rect 25976 1442 26004 2604
rect 26054 2544 26110 2553
rect 26330 2544 26386 2553
rect 26054 2479 26110 2488
rect 26148 2508 26200 2514
rect 26068 2446 26096 2479
rect 26330 2479 26386 2488
rect 26148 2450 26200 2456
rect 26056 2440 26108 2446
rect 26056 2382 26108 2388
rect 26056 2304 26108 2310
rect 26056 2246 26108 2252
rect 26068 1562 26096 2246
rect 26056 1556 26108 1562
rect 26056 1498 26108 1504
rect 25884 1414 26004 1442
rect 25688 468 25740 474
rect 25688 410 25740 416
rect 25884 56 25912 1414
rect 26160 56 26188 2450
rect 26240 2304 26292 2310
rect 26240 2246 26292 2252
rect 26252 1902 26280 2246
rect 26240 1896 26292 1902
rect 26240 1838 26292 1844
rect 26344 377 26372 2479
rect 26436 1426 26464 4422
rect 26514 3632 26570 3641
rect 26514 3567 26570 3576
rect 26528 3534 26556 3567
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 26516 2304 26568 2310
rect 26516 2246 26568 2252
rect 26424 1420 26476 1426
rect 26424 1362 26476 1368
rect 26528 1170 26556 2246
rect 26620 1873 26648 4558
rect 26792 4548 26844 4554
rect 26792 4490 26844 4496
rect 26700 2848 26752 2854
rect 26700 2790 26752 2796
rect 26606 1864 26662 1873
rect 26606 1799 26662 1808
rect 26436 1142 26556 1170
rect 26330 368 26386 377
rect 26330 303 26386 312
rect 26436 56 26464 1142
rect 26712 56 26740 2790
rect 26804 2689 26832 4490
rect 26790 2680 26846 2689
rect 26790 2615 26846 2624
rect 26896 2496 26924 6870
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 27356 2774 27384 7346
rect 27540 7206 27568 8978
rect 27712 7404 27764 7410
rect 27712 7346 27764 7352
rect 27528 7200 27580 7206
rect 27528 7142 27580 7148
rect 27724 6934 27752 7346
rect 27816 7206 27844 9046
rect 28080 8968 28132 8974
rect 28080 8910 28132 8916
rect 27988 7404 28040 7410
rect 27988 7346 28040 7352
rect 27804 7200 27856 7206
rect 27804 7142 27856 7148
rect 27712 6928 27764 6934
rect 27712 6870 27764 6876
rect 27436 5160 27488 5166
rect 27436 5102 27488 5108
rect 27620 5160 27672 5166
rect 27620 5102 27672 5108
rect 26804 2468 26924 2496
rect 27264 2746 27384 2774
rect 26804 1290 26832 2468
rect 27264 2394 27292 2746
rect 27448 2514 27476 5102
rect 27632 4826 27660 5102
rect 27620 4820 27672 4826
rect 27620 4762 27672 4768
rect 27896 3936 27948 3942
rect 27896 3878 27948 3884
rect 27908 3058 27936 3878
rect 28000 3097 28028 7346
rect 28092 7206 28120 8910
rect 28184 8634 28212 11194
rect 30116 8634 30144 11194
rect 30196 9240 30248 9246
rect 30196 9182 30248 9188
rect 28172 8628 28224 8634
rect 28172 8570 28224 8576
rect 30104 8628 30156 8634
rect 30104 8570 30156 8576
rect 30208 8498 30236 9182
rect 32048 8634 32076 11194
rect 33784 8832 33836 8838
rect 33784 8774 33836 8780
rect 33010 8732 33318 8741
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 33010 8667 33318 8676
rect 32036 8628 32088 8634
rect 32036 8570 32088 8576
rect 30196 8492 30248 8498
rect 30196 8434 30248 8440
rect 32588 8492 32640 8498
rect 32588 8434 32640 8440
rect 31024 8424 31076 8430
rect 31024 8366 31076 8372
rect 28356 7744 28408 7750
rect 28356 7686 28408 7692
rect 28264 7404 28316 7410
rect 28264 7346 28316 7352
rect 28080 7200 28132 7206
rect 28080 7142 28132 7148
rect 28080 5228 28132 5234
rect 28080 5170 28132 5176
rect 27986 3088 28042 3097
rect 27896 3052 27948 3058
rect 27986 3023 28042 3032
rect 27896 2994 27948 3000
rect 27712 2916 27764 2922
rect 27712 2858 27764 2864
rect 27620 2644 27672 2650
rect 27620 2586 27672 2592
rect 27436 2508 27488 2514
rect 27436 2450 27488 2456
rect 26884 2372 26936 2378
rect 27264 2366 27476 2394
rect 26884 2314 26936 2320
rect 26792 1284 26844 1290
rect 26792 1226 26844 1232
rect 26896 1170 26924 2314
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 27252 1896 27304 1902
rect 27252 1838 27304 1844
rect 26896 1142 27016 1170
rect 26988 56 27016 1142
rect 27264 56 27292 1838
rect 27448 1329 27476 2366
rect 27632 1902 27660 2586
rect 27620 1896 27672 1902
rect 27620 1838 27672 1844
rect 27528 1692 27580 1698
rect 27528 1634 27580 1640
rect 27434 1320 27490 1329
rect 27434 1255 27490 1264
rect 27540 56 27568 1634
rect 27724 406 27752 2858
rect 27804 2848 27856 2854
rect 27804 2790 27856 2796
rect 27712 400 27764 406
rect 27712 342 27764 348
rect 27816 56 27844 2790
rect 28092 2774 28120 5170
rect 28172 4140 28224 4146
rect 28172 4082 28224 4088
rect 28184 4049 28212 4082
rect 28170 4040 28226 4049
rect 28170 3975 28226 3984
rect 28276 3618 28304 7346
rect 28368 7206 28396 7686
rect 28448 7472 28500 7478
rect 28448 7414 28500 7420
rect 28460 7206 28488 7414
rect 28816 7404 28868 7410
rect 28816 7346 28868 7352
rect 28356 7200 28408 7206
rect 28356 7142 28408 7148
rect 28448 7200 28500 7206
rect 28448 7142 28500 7148
rect 28540 4480 28592 4486
rect 28540 4422 28592 4428
rect 28276 3590 28396 3618
rect 28368 3505 28396 3590
rect 28354 3496 28410 3505
rect 28354 3431 28410 3440
rect 28448 3120 28500 3126
rect 28448 3062 28500 3068
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 28000 2746 28120 2774
rect 27896 2440 27948 2446
rect 27896 2382 27948 2388
rect 27908 1698 27936 2382
rect 28000 1766 28028 2746
rect 28080 2576 28132 2582
rect 28080 2518 28132 2524
rect 27988 1760 28040 1766
rect 27988 1702 28040 1708
rect 27896 1692 27948 1698
rect 27896 1634 27948 1640
rect 28092 56 28120 2518
rect 28172 2440 28224 2446
rect 28172 2382 28224 2388
rect 28184 2106 28212 2382
rect 28172 2100 28224 2106
rect 28172 2042 28224 2048
rect 28368 56 28396 2790
rect 28460 2446 28488 3062
rect 28448 2440 28500 2446
rect 28448 2382 28500 2388
rect 28448 2032 28500 2038
rect 28448 1974 28500 1980
rect 28460 1834 28488 1974
rect 28552 1952 28580 4422
rect 28632 3936 28684 3942
rect 28632 3878 28684 3884
rect 28644 2446 28672 3878
rect 28632 2440 28684 2446
rect 28632 2382 28684 2388
rect 28724 2304 28776 2310
rect 28724 2246 28776 2252
rect 28632 1964 28684 1970
rect 28552 1924 28632 1952
rect 28632 1906 28684 1912
rect 28448 1828 28500 1834
rect 28448 1770 28500 1776
rect 28736 762 28764 2246
rect 28828 1358 28856 7346
rect 30840 4752 30892 4758
rect 30840 4694 30892 4700
rect 29552 4548 29604 4554
rect 29552 4490 29604 4496
rect 29000 4480 29052 4486
rect 29000 4422 29052 4428
rect 29012 4214 29040 4422
rect 29000 4208 29052 4214
rect 29000 4150 29052 4156
rect 29460 4140 29512 4146
rect 29460 4082 29512 4088
rect 29472 4026 29500 4082
rect 29288 4010 29500 4026
rect 29276 4004 29500 4010
rect 29328 3998 29500 4004
rect 29276 3946 29328 3952
rect 29000 3936 29052 3942
rect 29000 3878 29052 3884
rect 29184 3936 29236 3942
rect 29184 3878 29236 3884
rect 28908 2848 28960 2854
rect 28908 2790 28960 2796
rect 28816 1352 28868 1358
rect 28816 1294 28868 1300
rect 28644 734 28764 762
rect 28644 56 28672 734
rect 28920 56 28948 2790
rect 29012 2417 29040 3878
rect 29196 3058 29224 3878
rect 29184 3052 29236 3058
rect 29184 2994 29236 3000
rect 29184 2576 29236 2582
rect 29184 2518 29236 2524
rect 28998 2408 29054 2417
rect 28998 2343 29054 2352
rect 29196 56 29224 2518
rect 29460 2372 29512 2378
rect 29460 2314 29512 2320
rect 29472 56 29500 2314
rect 29564 241 29592 4490
rect 30380 4140 30432 4146
rect 30380 4082 30432 4088
rect 30104 4004 30156 4010
rect 30104 3946 30156 3952
rect 29828 3936 29880 3942
rect 29828 3878 29880 3884
rect 30012 3936 30064 3942
rect 30012 3878 30064 3884
rect 29736 2644 29788 2650
rect 29736 2586 29788 2592
rect 29550 232 29606 241
rect 29550 167 29606 176
rect 29748 56 29776 2586
rect 29840 270 29868 3878
rect 29920 3528 29972 3534
rect 29920 3470 29972 3476
rect 29932 338 29960 3470
rect 30024 2446 30052 3878
rect 30116 3058 30144 3946
rect 30196 3732 30248 3738
rect 30196 3674 30248 3680
rect 30104 3052 30156 3058
rect 30104 2994 30156 3000
rect 30104 2848 30156 2854
rect 30104 2790 30156 2796
rect 30012 2440 30064 2446
rect 30012 2382 30064 2388
rect 30116 1442 30144 2790
rect 30208 2446 30236 3674
rect 30288 2576 30340 2582
rect 30288 2518 30340 2524
rect 30196 2440 30248 2446
rect 30196 2382 30248 2388
rect 30024 1414 30144 1442
rect 29920 332 29972 338
rect 29920 274 29972 280
rect 29828 264 29880 270
rect 29828 206 29880 212
rect 30024 56 30052 1414
rect 30300 56 30328 2518
rect 30392 134 30420 4082
rect 30748 4004 30800 4010
rect 30748 3946 30800 3952
rect 30760 2774 30788 3946
rect 30852 3058 30880 4694
rect 31036 4486 31064 8366
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 32312 6860 32364 6866
rect 32312 6802 32364 6808
rect 31576 6724 31628 6730
rect 31576 6666 31628 6672
rect 31588 5778 31616 6666
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 31576 5772 31628 5778
rect 31576 5714 31628 5720
rect 31392 5228 31444 5234
rect 31392 5170 31444 5176
rect 31404 4826 31432 5170
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 31300 4820 31352 4826
rect 31300 4762 31352 4768
rect 31392 4820 31444 4826
rect 31392 4762 31444 4768
rect 30932 4480 30984 4486
rect 30932 4422 30984 4428
rect 31024 4480 31076 4486
rect 31024 4422 31076 4428
rect 30840 3052 30892 3058
rect 30840 2994 30892 3000
rect 30840 2848 30892 2854
rect 30840 2790 30892 2796
rect 30668 2746 30788 2774
rect 30668 2446 30696 2746
rect 30656 2440 30708 2446
rect 30656 2382 30708 2388
rect 30564 2304 30616 2310
rect 30564 2246 30616 2252
rect 30380 128 30432 134
rect 30380 70 30432 76
rect 30576 56 30604 2246
rect 30852 56 30880 2790
rect 30944 2774 30972 4422
rect 31024 3936 31076 3942
rect 31024 3878 31076 3884
rect 31116 3936 31168 3942
rect 31116 3878 31168 3884
rect 31036 3534 31064 3878
rect 31128 3738 31156 3878
rect 31116 3732 31168 3738
rect 31116 3674 31168 3680
rect 31024 3528 31076 3534
rect 31024 3470 31076 3476
rect 31312 3058 31340 4762
rect 31496 4690 31800 4706
rect 31496 4684 31812 4690
rect 31496 4678 31576 4684
rect 31300 3052 31352 3058
rect 31300 2994 31352 3000
rect 31208 2848 31260 2854
rect 31128 2796 31208 2802
rect 31128 2790 31260 2796
rect 31128 2774 31248 2790
rect 31496 2774 31524 4678
rect 31628 4678 31760 4684
rect 31576 4626 31628 4632
rect 31760 4626 31812 4632
rect 31852 4616 31904 4622
rect 31904 4564 31984 4570
rect 31852 4558 31984 4564
rect 31864 4542 31984 4558
rect 31760 4480 31812 4486
rect 31760 4422 31812 4428
rect 31852 4480 31904 4486
rect 31852 4422 31904 4428
rect 31576 4140 31628 4146
rect 31576 4082 31628 4088
rect 30944 2746 31064 2774
rect 31036 2650 31064 2746
rect 31024 2644 31076 2650
rect 31024 2586 31076 2592
rect 31128 56 31156 2774
rect 31312 2746 31524 2774
rect 31312 105 31340 2746
rect 31392 2644 31444 2650
rect 31392 2586 31444 2592
rect 31404 2446 31432 2586
rect 31484 2576 31536 2582
rect 31484 2518 31536 2524
rect 31392 2440 31444 2446
rect 31392 2382 31444 2388
rect 31496 1306 31524 2518
rect 31404 1278 31524 1306
rect 31298 96 31354 105
rect 22388 14 22508 42
rect 22558 0 22614 56
rect 22834 0 22890 56
rect 23110 0 23166 56
rect 23386 0 23442 56
rect 23662 0 23718 56
rect 23938 0 23994 56
rect 24214 0 24270 56
rect 24490 0 24546 56
rect 24766 0 24822 56
rect 25042 0 25098 56
rect 25318 0 25374 56
rect 25594 0 25650 56
rect 25870 0 25926 56
rect 26146 0 26202 56
rect 26422 0 26478 56
rect 26698 0 26754 56
rect 26974 0 27030 56
rect 27250 0 27306 56
rect 27526 0 27582 56
rect 27802 0 27858 56
rect 28078 0 28134 56
rect 28354 0 28410 56
rect 28630 0 28686 56
rect 28906 0 28962 56
rect 29182 0 29238 56
rect 29458 0 29514 56
rect 29734 0 29790 56
rect 30010 0 30066 56
rect 30286 0 30342 56
rect 30562 0 30618 56
rect 30838 0 30894 56
rect 31114 0 31170 56
rect 31404 56 31432 1278
rect 31588 202 31616 4082
rect 31772 2514 31800 4422
rect 31760 2508 31812 2514
rect 31760 2450 31812 2456
rect 31864 2378 31892 4422
rect 31956 4214 31984 4542
rect 31944 4208 31996 4214
rect 31944 4150 31996 4156
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 32324 2564 32352 6802
rect 32496 5160 32548 5166
rect 32496 5102 32548 5108
rect 32404 4480 32456 4486
rect 32404 4422 32456 4428
rect 32416 3126 32444 4422
rect 32404 3120 32456 3126
rect 32404 3062 32456 3068
rect 32232 2536 32352 2564
rect 32036 2508 32088 2514
rect 32036 2450 32088 2456
rect 31852 2372 31904 2378
rect 31852 2314 31904 2320
rect 31944 2372 31996 2378
rect 31944 2314 31996 2320
rect 31668 2304 31720 2310
rect 31668 2246 31720 2252
rect 31576 196 31628 202
rect 31576 138 31628 144
rect 31680 56 31708 2246
rect 31956 56 31984 2314
rect 32048 2038 32076 2450
rect 32128 2440 32180 2446
rect 32128 2382 32180 2388
rect 32036 2032 32088 2038
rect 32036 1974 32088 1980
rect 32140 1970 32168 2382
rect 32128 1964 32180 1970
rect 32128 1906 32180 1912
rect 32232 56 32260 2536
rect 32508 2446 32536 5102
rect 32600 3398 32628 8434
rect 33796 8362 33824 8774
rect 33980 8634 34008 11194
rect 35912 8634 35940 11194
rect 37738 9616 37794 9625
rect 37738 9551 37794 9560
rect 37004 8968 37056 8974
rect 37004 8910 37056 8916
rect 37016 8634 37044 8910
rect 37556 8900 37608 8906
rect 37556 8842 37608 8848
rect 33968 8628 34020 8634
rect 33968 8570 34020 8576
rect 35900 8628 35952 8634
rect 35900 8570 35952 8576
rect 37004 8628 37056 8634
rect 37004 8570 37056 8576
rect 37568 8498 37596 8842
rect 37752 8634 37780 9551
rect 37844 8634 37872 11194
rect 38382 9888 38438 9897
rect 38382 9823 38438 9832
rect 38290 9344 38346 9353
rect 38290 9279 38346 9288
rect 37740 8628 37792 8634
rect 37740 8570 37792 8576
rect 37832 8628 37884 8634
rect 37832 8570 37884 8576
rect 35992 8492 36044 8498
rect 35992 8434 36044 8440
rect 36820 8492 36872 8498
rect 36820 8434 36872 8440
rect 37556 8492 37608 8498
rect 37556 8434 37608 8440
rect 37648 8492 37700 8498
rect 37648 8434 37700 8440
rect 33784 8356 33836 8362
rect 33784 8298 33836 8304
rect 33010 7644 33318 7653
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 34704 7404 34756 7410
rect 34704 7346 34756 7352
rect 33876 6928 33928 6934
rect 33876 6870 33928 6876
rect 32772 6792 32824 6798
rect 32772 6734 32824 6740
rect 32680 4616 32732 4622
rect 32680 4558 32732 4564
rect 32588 3392 32640 3398
rect 32588 3334 32640 3340
rect 32496 2440 32548 2446
rect 32496 2382 32548 2388
rect 32496 1284 32548 1290
rect 32496 1226 32548 1232
rect 32508 56 32536 1226
rect 32692 66 32720 4558
rect 32784 1970 32812 6734
rect 33010 6556 33318 6565
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 33508 6180 33560 6186
rect 33508 6122 33560 6128
rect 33010 5468 33318 5477
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 33010 5403 33318 5412
rect 33010 4380 33318 4389
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 33010 3292 33318 3301
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 32772 1964 32824 1970
rect 32772 1906 32824 1912
rect 32770 1728 32826 1737
rect 32876 1698 32904 2382
rect 33010 2204 33318 2213
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 33428 2106 33456 2382
rect 33416 2100 33468 2106
rect 33416 2042 33468 2048
rect 33048 1964 33100 1970
rect 33048 1906 33100 1912
rect 32770 1663 32826 1672
rect 32864 1692 32916 1698
rect 32680 60 32732 66
rect 31298 31 31354 40
rect 31390 0 31446 56
rect 31666 0 31722 56
rect 31942 0 31998 56
rect 32218 0 32274 56
rect 32494 0 32550 56
rect 32784 56 32812 1663
rect 32864 1634 32916 1640
rect 33060 56 33088 1906
rect 33336 56 33456 82
rect 32680 2 32732 8
rect 32770 0 32826 56
rect 33046 0 33102 56
rect 33322 54 33456 56
rect 33322 0 33378 54
rect 33428 42 33456 54
rect 33520 42 33548 6122
rect 33784 5092 33836 5098
rect 33784 5034 33836 5040
rect 33796 4758 33824 5034
rect 33784 4752 33836 4758
rect 33784 4694 33836 4700
rect 33600 536 33652 542
rect 33600 478 33652 484
rect 33612 56 33640 478
rect 33888 56 33916 6870
rect 34426 3496 34482 3505
rect 34426 3431 34482 3440
rect 34150 3088 34206 3097
rect 34150 3023 34206 3032
rect 34164 56 34192 3023
rect 34440 56 34468 3431
rect 34716 56 34744 7346
rect 35532 6316 35584 6322
rect 35532 6258 35584 6264
rect 35256 1352 35308 1358
rect 34978 1320 35034 1329
rect 35256 1294 35308 1300
rect 34978 1255 35034 1264
rect 34992 56 35020 1255
rect 35268 56 35296 1294
rect 35544 56 35572 6258
rect 35808 5704 35860 5710
rect 35808 5646 35860 5652
rect 35820 56 35848 5646
rect 36004 4826 36032 8434
rect 36832 5370 36860 8434
rect 37660 8378 37688 8434
rect 37200 8350 37688 8378
rect 36820 5364 36872 5370
rect 36820 5306 36872 5312
rect 35992 4820 36044 4826
rect 35992 4762 36044 4768
rect 37096 4684 37148 4690
rect 37096 4626 37148 4632
rect 35900 4276 35952 4282
rect 35900 4218 35952 4224
rect 35912 4078 35940 4218
rect 36912 4208 36964 4214
rect 36912 4150 36964 4156
rect 35900 4072 35952 4078
rect 35900 4014 35952 4020
rect 36634 3632 36690 3641
rect 36634 3567 36690 3576
rect 36084 468 36136 474
rect 36084 410 36136 416
rect 36096 56 36124 410
rect 36360 400 36412 406
rect 36360 342 36412 348
rect 36372 56 36400 342
rect 36648 56 36676 3567
rect 36924 56 36952 4150
rect 37108 2394 37136 4626
rect 37200 4486 37228 8350
rect 37950 8188 38258 8197
rect 37950 8186 37956 8188
rect 38012 8186 38036 8188
rect 38092 8186 38116 8188
rect 38172 8186 38196 8188
rect 38252 8186 38258 8188
rect 38012 8134 38014 8186
rect 38194 8134 38196 8186
rect 37950 8132 37956 8134
rect 38012 8132 38036 8134
rect 38092 8132 38116 8134
rect 38172 8132 38196 8134
rect 38252 8132 38258 8134
rect 37950 8123 38258 8132
rect 38304 8090 38332 9279
rect 38292 8084 38344 8090
rect 38292 8026 38344 8032
rect 37740 7880 37792 7886
rect 37740 7822 37792 7828
rect 38108 7880 38160 7886
rect 38108 7822 38160 7828
rect 37752 7478 37780 7822
rect 37832 7812 37884 7818
rect 37832 7754 37884 7760
rect 38016 7812 38068 7818
rect 38016 7754 38068 7760
rect 37844 7478 37872 7754
rect 37740 7472 37792 7478
rect 37740 7414 37792 7420
rect 37832 7472 37884 7478
rect 37832 7414 37884 7420
rect 38028 7274 38056 7754
rect 38120 7342 38148 7822
rect 38396 7750 38424 9823
rect 39578 9072 39634 9081
rect 39578 9007 39634 9016
rect 39486 8800 39542 8809
rect 39010 8732 39318 8741
rect 39486 8735 39542 8744
rect 39010 8730 39016 8732
rect 39072 8730 39096 8732
rect 39152 8730 39176 8732
rect 39232 8730 39256 8732
rect 39312 8730 39318 8732
rect 39072 8678 39074 8730
rect 39254 8678 39256 8730
rect 39010 8676 39016 8678
rect 39072 8676 39096 8678
rect 39152 8676 39176 8678
rect 39232 8676 39256 8678
rect 39312 8676 39318 8678
rect 39010 8667 39318 8676
rect 38660 8628 38712 8634
rect 38660 8570 38712 8576
rect 38672 8537 38700 8570
rect 38658 8528 38714 8537
rect 38658 8463 38714 8472
rect 39028 8356 39080 8362
rect 39028 8298 39080 8304
rect 39396 8356 39448 8362
rect 39396 8298 39448 8304
rect 39040 8265 39068 8298
rect 39026 8256 39082 8265
rect 39026 8191 39082 8200
rect 39408 7993 39436 8298
rect 39500 8090 39528 8735
rect 39488 8084 39540 8090
rect 39488 8026 39540 8032
rect 39394 7984 39450 7993
rect 39394 7919 39450 7928
rect 38384 7744 38436 7750
rect 38384 7686 38436 7692
rect 38936 7744 38988 7750
rect 39396 7744 39448 7750
rect 38936 7686 38988 7692
rect 39394 7712 39396 7721
rect 39448 7712 39450 7721
rect 38948 7449 38976 7686
rect 39010 7644 39318 7653
rect 39394 7647 39450 7656
rect 39010 7642 39016 7644
rect 39072 7642 39096 7644
rect 39152 7642 39176 7644
rect 39232 7642 39256 7644
rect 39312 7642 39318 7644
rect 39072 7590 39074 7642
rect 39254 7590 39256 7642
rect 39010 7588 39016 7590
rect 39072 7588 39096 7590
rect 39152 7588 39176 7590
rect 39232 7588 39256 7590
rect 39312 7588 39318 7590
rect 39010 7579 39318 7588
rect 39592 7546 39620 9007
rect 39776 8974 39804 11194
rect 39764 8968 39816 8974
rect 39764 8910 39816 8916
rect 39580 7540 39632 7546
rect 39580 7482 39632 7488
rect 38934 7440 38990 7449
rect 38844 7404 38896 7410
rect 38934 7375 38990 7384
rect 38844 7346 38896 7352
rect 38108 7336 38160 7342
rect 38108 7278 38160 7284
rect 38016 7268 38068 7274
rect 38016 7210 38068 7216
rect 37950 7100 38258 7109
rect 37950 7098 37956 7100
rect 38012 7098 38036 7100
rect 38092 7098 38116 7100
rect 38172 7098 38196 7100
rect 38252 7098 38258 7100
rect 38012 7046 38014 7098
rect 38194 7046 38196 7098
rect 37950 7044 37956 7046
rect 38012 7044 38036 7046
rect 38092 7044 38116 7046
rect 38172 7044 38196 7046
rect 38252 7044 38258 7046
rect 37950 7035 38258 7044
rect 38856 7002 38884 7346
rect 39396 7200 39448 7206
rect 39394 7168 39396 7177
rect 39448 7168 39450 7177
rect 39394 7103 39450 7112
rect 38844 6996 38896 7002
rect 38844 6938 38896 6944
rect 39394 6896 39450 6905
rect 39394 6831 39450 6840
rect 39212 6792 39264 6798
rect 39210 6760 39212 6769
rect 39264 6760 39266 6769
rect 39210 6695 39266 6704
rect 39408 6662 39436 6831
rect 39948 6724 40000 6730
rect 39948 6666 40000 6672
rect 39396 6656 39448 6662
rect 39960 6633 39988 6666
rect 39396 6598 39448 6604
rect 39946 6624 40002 6633
rect 39010 6556 39318 6565
rect 39946 6559 40002 6568
rect 39010 6554 39016 6556
rect 39072 6554 39096 6556
rect 39152 6554 39176 6556
rect 39232 6554 39256 6556
rect 39312 6554 39318 6556
rect 39072 6502 39074 6554
rect 39254 6502 39256 6554
rect 39010 6500 39016 6502
rect 39072 6500 39096 6502
rect 39152 6500 39176 6502
rect 39232 6500 39256 6502
rect 39312 6500 39318 6502
rect 39010 6491 39318 6500
rect 39396 6452 39448 6458
rect 39396 6394 39448 6400
rect 39408 6361 39436 6394
rect 39394 6352 39450 6361
rect 38660 6316 38712 6322
rect 39394 6287 39450 6296
rect 38660 6258 38712 6264
rect 37950 6012 38258 6021
rect 37950 6010 37956 6012
rect 38012 6010 38036 6012
rect 38092 6010 38116 6012
rect 38172 6010 38196 6012
rect 38252 6010 38258 6012
rect 38012 5958 38014 6010
rect 38194 5958 38196 6010
rect 37950 5956 37956 5958
rect 38012 5956 38036 5958
rect 38092 5956 38116 5958
rect 38172 5956 38196 5958
rect 38252 5956 38258 5958
rect 37950 5947 38258 5956
rect 37740 5228 37792 5234
rect 37740 5170 37792 5176
rect 37464 4616 37516 4622
rect 37464 4558 37516 4564
rect 37188 4480 37240 4486
rect 37188 4422 37240 4428
rect 37108 2366 37228 2394
rect 37200 56 37228 2366
rect 37476 56 37504 4558
rect 37752 56 37780 5170
rect 38672 5030 38700 6258
rect 39028 6112 39080 6118
rect 39026 6080 39028 6089
rect 39080 6080 39082 6089
rect 39026 6015 39082 6024
rect 39396 5840 39448 5846
rect 39394 5808 39396 5817
rect 39448 5808 39450 5817
rect 39394 5743 39450 5752
rect 38844 5704 38896 5710
rect 38842 5672 38844 5681
rect 38896 5672 38898 5681
rect 38842 5607 38898 5616
rect 39948 5568 40000 5574
rect 39946 5536 39948 5545
rect 40000 5536 40002 5545
rect 39010 5468 39318 5477
rect 39946 5471 40002 5480
rect 39010 5466 39016 5468
rect 39072 5466 39096 5468
rect 39152 5466 39176 5468
rect 39232 5466 39256 5468
rect 39312 5466 39318 5468
rect 39072 5414 39074 5466
rect 39254 5414 39256 5466
rect 39010 5412 39016 5414
rect 39072 5412 39096 5414
rect 39152 5412 39176 5414
rect 39232 5412 39256 5414
rect 39312 5412 39318 5414
rect 39010 5403 39318 5412
rect 39396 5364 39448 5370
rect 39396 5306 39448 5312
rect 39408 5273 39436 5306
rect 39210 5264 39266 5273
rect 39210 5199 39212 5208
rect 39264 5199 39266 5208
rect 39394 5264 39450 5273
rect 39394 5199 39450 5208
rect 39212 5170 39264 5176
rect 38660 5024 38712 5030
rect 39028 5024 39080 5030
rect 38660 4966 38712 4972
rect 39026 4992 39028 5001
rect 39080 4992 39082 5001
rect 37950 4924 38258 4933
rect 39026 4927 39082 4936
rect 37950 4922 37956 4924
rect 38012 4922 38036 4924
rect 38092 4922 38116 4924
rect 38172 4922 38196 4924
rect 38252 4922 38258 4924
rect 38012 4870 38014 4922
rect 38194 4870 38196 4922
rect 37950 4868 37956 4870
rect 38012 4868 38036 4870
rect 38092 4868 38116 4870
rect 38172 4868 38196 4870
rect 38252 4868 38258 4870
rect 37950 4859 38258 4868
rect 39396 4752 39448 4758
rect 39394 4720 39396 4729
rect 39448 4720 39450 4729
rect 39394 4655 39450 4664
rect 39948 4480 40000 4486
rect 39946 4448 39948 4457
rect 40000 4448 40002 4457
rect 39010 4380 39318 4389
rect 39946 4383 40002 4392
rect 39010 4378 39016 4380
rect 39072 4378 39096 4380
rect 39152 4378 39176 4380
rect 39232 4378 39256 4380
rect 39312 4378 39318 4380
rect 39072 4326 39074 4378
rect 39254 4326 39256 4378
rect 39010 4324 39016 4326
rect 39072 4324 39096 4326
rect 39152 4324 39176 4326
rect 39232 4324 39256 4326
rect 39312 4324 39318 4326
rect 39010 4315 39318 4324
rect 39394 4176 39450 4185
rect 39394 4111 39450 4120
rect 39408 4010 39436 4111
rect 39212 4004 39264 4010
rect 39212 3946 39264 3952
rect 39396 4004 39448 4010
rect 39396 3946 39448 3952
rect 39028 3936 39080 3942
rect 39026 3904 39028 3913
rect 39080 3904 39082 3913
rect 37950 3836 38258 3845
rect 39026 3839 39082 3848
rect 37950 3834 37956 3836
rect 38012 3834 38036 3836
rect 38092 3834 38116 3836
rect 38172 3834 38196 3836
rect 38252 3834 38258 3836
rect 38012 3782 38014 3834
rect 38194 3782 38196 3834
rect 37950 3780 37956 3782
rect 38012 3780 38036 3782
rect 38092 3780 38116 3782
rect 38172 3780 38196 3782
rect 38252 3780 38258 3782
rect 37950 3771 38258 3780
rect 38844 3664 38896 3670
rect 38844 3606 38896 3612
rect 38856 3058 38884 3606
rect 39224 3534 39252 3946
rect 39396 3664 39448 3670
rect 39394 3632 39396 3641
rect 39448 3632 39450 3641
rect 39394 3567 39450 3576
rect 39212 3528 39264 3534
rect 39212 3470 39264 3476
rect 38936 3460 38988 3466
rect 38936 3402 38988 3408
rect 38948 3058 38976 3402
rect 39948 3392 40000 3398
rect 39946 3360 39948 3369
rect 40000 3360 40002 3369
rect 39010 3292 39318 3301
rect 39946 3295 40002 3304
rect 39010 3290 39016 3292
rect 39072 3290 39096 3292
rect 39152 3290 39176 3292
rect 39232 3290 39256 3292
rect 39312 3290 39318 3292
rect 39072 3238 39074 3290
rect 39254 3238 39256 3290
rect 39010 3236 39016 3238
rect 39072 3236 39096 3238
rect 39152 3236 39176 3238
rect 39232 3236 39256 3238
rect 39312 3236 39318 3238
rect 39010 3227 39318 3236
rect 39396 3188 39448 3194
rect 39396 3130 39448 3136
rect 39408 3097 39436 3130
rect 39394 3088 39450 3097
rect 38844 3052 38896 3058
rect 38844 2994 38896 3000
rect 38936 3052 38988 3058
rect 39394 3023 39450 3032
rect 38936 2994 38988 3000
rect 40408 2916 40460 2922
rect 40408 2858 40460 2864
rect 39028 2848 39080 2854
rect 39026 2816 39028 2825
rect 39080 2816 39082 2825
rect 37950 2748 38258 2757
rect 39026 2751 39082 2760
rect 37950 2746 37956 2748
rect 38012 2746 38036 2748
rect 38092 2746 38116 2748
rect 38172 2746 38196 2748
rect 38252 2746 38258 2748
rect 38012 2694 38014 2746
rect 38194 2694 38196 2746
rect 37950 2692 37956 2694
rect 38012 2692 38036 2694
rect 38092 2692 38116 2694
rect 38172 2692 38196 2694
rect 38252 2692 38258 2694
rect 37950 2683 38258 2692
rect 39396 2576 39448 2582
rect 39394 2544 39396 2553
rect 39448 2544 39450 2553
rect 39394 2479 39450 2488
rect 38476 2440 38528 2446
rect 38476 2382 38528 2388
rect 37924 2304 37976 2310
rect 37924 2246 37976 2252
rect 38292 2304 38344 2310
rect 38292 2246 38344 2252
rect 37936 2009 37964 2246
rect 37922 2000 37978 2009
rect 37922 1935 37978 1944
rect 38304 1737 38332 2246
rect 38488 2106 38516 2382
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 38936 2304 38988 2310
rect 40420 2281 40448 2858
rect 38936 2246 38988 2252
rect 40406 2272 40462 2281
rect 38476 2100 38528 2106
rect 38476 2042 38528 2048
rect 38290 1728 38346 1737
rect 38290 1663 38346 1672
rect 38672 1465 38700 2246
rect 38948 1970 38976 2246
rect 39010 2204 39318 2213
rect 40406 2207 40462 2216
rect 39010 2202 39016 2204
rect 39072 2202 39096 2204
rect 39152 2202 39176 2204
rect 39232 2202 39256 2204
rect 39312 2202 39318 2204
rect 39072 2150 39074 2202
rect 39254 2150 39256 2202
rect 39010 2148 39016 2150
rect 39072 2148 39096 2150
rect 39152 2148 39176 2150
rect 39232 2148 39256 2150
rect 39312 2148 39318 2150
rect 39010 2139 39318 2148
rect 38936 1964 38988 1970
rect 38936 1906 38988 1912
rect 38658 1456 38714 1465
rect 38658 1391 38714 1400
rect 33428 14 33548 42
rect 33598 0 33654 56
rect 33874 0 33930 56
rect 34150 0 34206 56
rect 34426 0 34482 56
rect 34702 0 34758 56
rect 34978 0 35034 56
rect 35254 0 35310 56
rect 35530 0 35586 56
rect 35806 0 35862 56
rect 36082 0 36138 56
rect 36358 0 36414 56
rect 36634 0 36690 56
rect 36910 0 36966 56
rect 37186 0 37242 56
rect 37462 0 37518 56
rect 37738 0 37794 56
<< via2 >>
rect 2778 8744 2834 8800
rect 1306 7384 1362 7440
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 14830 9560 14886 9616
rect 2778 8336 2834 8392
rect 1766 8200 1822 8256
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 1766 7792 1822 7848
rect 14922 9288 14978 9344
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 16486 8336 16542 8392
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 16394 7828 16396 7848
rect 16396 7828 16448 7848
rect 16448 7828 16450 7848
rect 16394 7792 16450 7828
rect 15106 7404 15162 7440
rect 15106 7384 15108 7404
rect 15108 7384 15160 7404
rect 15160 7384 15162 7404
rect 16486 7284 16488 7304
rect 16488 7284 16540 7304
rect 16540 7284 16542 7304
rect 16486 7248 16542 7284
rect 18694 9016 18750 9072
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 19062 7928 19118 7984
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 22558 9832 22614 9888
rect 22098 8472 22154 8528
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 570 5480 626 5536
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 2778 5072 2834 5128
rect 1766 4936 1822 4992
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 1766 4528 1822 4584
rect 2778 4392 2834 4448
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 5538 1400 5594 1456
rect 17498 6860 17554 6896
rect 17498 6840 17500 6860
rect 17500 6840 17552 6860
rect 17552 6840 17554 6860
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 9678 6432 9734 6488
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 8666 2488 8722 2544
rect 8758 1536 8814 1592
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 9862 2216 9918 2272
rect 9586 1672 9642 1728
rect 11058 6296 11114 6352
rect 11242 6296 11298 6352
rect 10966 5616 11022 5672
rect 17406 6704 17462 6760
rect 17866 6704 17922 6760
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 14830 6432 14886 6488
rect 11886 2352 11942 2408
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 13174 1808 13230 1864
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 14830 6024 14886 6080
rect 14554 5652 14556 5672
rect 14556 5652 14608 5672
rect 14608 5652 14610 5672
rect 14554 5616 14610 5652
rect 14370 2488 14426 2544
rect 13634 1672 13690 1728
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 15106 1944 15162 2000
rect 15290 1944 15346 2000
rect 17314 3304 17370 3360
rect 17038 3168 17094 3224
rect 16578 2352 16634 2408
rect 16762 2352 16818 2408
rect 15290 1672 15346 1728
rect 13726 312 13782 368
rect 14554 176 14610 232
rect 14830 40 14886 96
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 19338 6024 19394 6080
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 19614 5616 19670 5672
rect 19154 5208 19210 5264
rect 19338 5208 19394 5264
rect 18510 1536 18566 1592
rect 19798 5752 19854 5808
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 20626 3984 20682 4040
rect 20442 3848 20498 3904
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 20350 3712 20406 3768
rect 20350 3304 20406 3360
rect 20442 3168 20498 3224
rect 20626 2896 20682 2952
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 21546 4528 21602 4584
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 22098 2896 22154 2952
rect 22374 6160 22430 6216
rect 23570 6296 23626 6352
rect 23478 5072 23534 5128
rect 22834 4684 22890 4720
rect 22834 4664 22836 4684
rect 22836 4664 22888 4684
rect 22888 4664 22890 4684
rect 22466 2624 22522 2680
rect 22742 2624 22798 2680
rect 22742 1672 22798 1728
rect 24030 4120 24086 4176
rect 24214 3576 24270 3632
rect 24122 3032 24178 3088
rect 24398 3476 24400 3496
rect 24400 3476 24452 3496
rect 24452 3476 24454 3496
rect 24398 3440 24454 3476
rect 24950 2760 25006 2816
rect 24858 1944 24914 2000
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 26330 3576 26386 3632
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 26054 2488 26110 2544
rect 26330 2488 26386 2544
rect 26514 3576 26570 3632
rect 26606 1808 26662 1864
rect 26330 312 26386 368
rect 26790 2624 26846 2680
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 27986 3032 28042 3088
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 27434 1264 27490 1320
rect 28170 3984 28226 4040
rect 28354 3440 28410 3496
rect 28998 2352 29054 2408
rect 29550 176 29606 232
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 31298 40 31354 96
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 37738 9560 37794 9616
rect 38382 9832 38438 9888
rect 38290 9288 38346 9344
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 32770 1672 32826 1728
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
rect 34426 3440 34482 3496
rect 34150 3032 34206 3088
rect 34978 1264 35034 1320
rect 36634 3576 36690 3632
rect 37956 8186 38012 8188
rect 38036 8186 38092 8188
rect 38116 8186 38172 8188
rect 38196 8186 38252 8188
rect 37956 8134 38002 8186
rect 38002 8134 38012 8186
rect 38036 8134 38066 8186
rect 38066 8134 38078 8186
rect 38078 8134 38092 8186
rect 38116 8134 38130 8186
rect 38130 8134 38142 8186
rect 38142 8134 38172 8186
rect 38196 8134 38206 8186
rect 38206 8134 38252 8186
rect 37956 8132 38012 8134
rect 38036 8132 38092 8134
rect 38116 8132 38172 8134
rect 38196 8132 38252 8134
rect 39578 9016 39634 9072
rect 39486 8744 39542 8800
rect 39016 8730 39072 8732
rect 39096 8730 39152 8732
rect 39176 8730 39232 8732
rect 39256 8730 39312 8732
rect 39016 8678 39062 8730
rect 39062 8678 39072 8730
rect 39096 8678 39126 8730
rect 39126 8678 39138 8730
rect 39138 8678 39152 8730
rect 39176 8678 39190 8730
rect 39190 8678 39202 8730
rect 39202 8678 39232 8730
rect 39256 8678 39266 8730
rect 39266 8678 39312 8730
rect 39016 8676 39072 8678
rect 39096 8676 39152 8678
rect 39176 8676 39232 8678
rect 39256 8676 39312 8678
rect 38658 8472 38714 8528
rect 39026 8200 39082 8256
rect 39394 7928 39450 7984
rect 39394 7692 39396 7712
rect 39396 7692 39448 7712
rect 39448 7692 39450 7712
rect 39394 7656 39450 7692
rect 39016 7642 39072 7644
rect 39096 7642 39152 7644
rect 39176 7642 39232 7644
rect 39256 7642 39312 7644
rect 39016 7590 39062 7642
rect 39062 7590 39072 7642
rect 39096 7590 39126 7642
rect 39126 7590 39138 7642
rect 39138 7590 39152 7642
rect 39176 7590 39190 7642
rect 39190 7590 39202 7642
rect 39202 7590 39232 7642
rect 39256 7590 39266 7642
rect 39266 7590 39312 7642
rect 39016 7588 39072 7590
rect 39096 7588 39152 7590
rect 39176 7588 39232 7590
rect 39256 7588 39312 7590
rect 38934 7384 38990 7440
rect 37956 7098 38012 7100
rect 38036 7098 38092 7100
rect 38116 7098 38172 7100
rect 38196 7098 38252 7100
rect 37956 7046 38002 7098
rect 38002 7046 38012 7098
rect 38036 7046 38066 7098
rect 38066 7046 38078 7098
rect 38078 7046 38092 7098
rect 38116 7046 38130 7098
rect 38130 7046 38142 7098
rect 38142 7046 38172 7098
rect 38196 7046 38206 7098
rect 38206 7046 38252 7098
rect 37956 7044 38012 7046
rect 38036 7044 38092 7046
rect 38116 7044 38172 7046
rect 38196 7044 38252 7046
rect 39394 7148 39396 7168
rect 39396 7148 39448 7168
rect 39448 7148 39450 7168
rect 39394 7112 39450 7148
rect 39394 6840 39450 6896
rect 39210 6740 39212 6760
rect 39212 6740 39264 6760
rect 39264 6740 39266 6760
rect 39210 6704 39266 6740
rect 39946 6568 40002 6624
rect 39016 6554 39072 6556
rect 39096 6554 39152 6556
rect 39176 6554 39232 6556
rect 39256 6554 39312 6556
rect 39016 6502 39062 6554
rect 39062 6502 39072 6554
rect 39096 6502 39126 6554
rect 39126 6502 39138 6554
rect 39138 6502 39152 6554
rect 39176 6502 39190 6554
rect 39190 6502 39202 6554
rect 39202 6502 39232 6554
rect 39256 6502 39266 6554
rect 39266 6502 39312 6554
rect 39016 6500 39072 6502
rect 39096 6500 39152 6502
rect 39176 6500 39232 6502
rect 39256 6500 39312 6502
rect 39394 6296 39450 6352
rect 37956 6010 38012 6012
rect 38036 6010 38092 6012
rect 38116 6010 38172 6012
rect 38196 6010 38252 6012
rect 37956 5958 38002 6010
rect 38002 5958 38012 6010
rect 38036 5958 38066 6010
rect 38066 5958 38078 6010
rect 38078 5958 38092 6010
rect 38116 5958 38130 6010
rect 38130 5958 38142 6010
rect 38142 5958 38172 6010
rect 38196 5958 38206 6010
rect 38206 5958 38252 6010
rect 37956 5956 38012 5958
rect 38036 5956 38092 5958
rect 38116 5956 38172 5958
rect 38196 5956 38252 5958
rect 39026 6060 39028 6080
rect 39028 6060 39080 6080
rect 39080 6060 39082 6080
rect 39026 6024 39082 6060
rect 39394 5788 39396 5808
rect 39396 5788 39448 5808
rect 39448 5788 39450 5808
rect 39394 5752 39450 5788
rect 38842 5652 38844 5672
rect 38844 5652 38896 5672
rect 38896 5652 38898 5672
rect 38842 5616 38898 5652
rect 39946 5516 39948 5536
rect 39948 5516 40000 5536
rect 40000 5516 40002 5536
rect 39946 5480 40002 5516
rect 39016 5466 39072 5468
rect 39096 5466 39152 5468
rect 39176 5466 39232 5468
rect 39256 5466 39312 5468
rect 39016 5414 39062 5466
rect 39062 5414 39072 5466
rect 39096 5414 39126 5466
rect 39126 5414 39138 5466
rect 39138 5414 39152 5466
rect 39176 5414 39190 5466
rect 39190 5414 39202 5466
rect 39202 5414 39232 5466
rect 39256 5414 39266 5466
rect 39266 5414 39312 5466
rect 39016 5412 39072 5414
rect 39096 5412 39152 5414
rect 39176 5412 39232 5414
rect 39256 5412 39312 5414
rect 39210 5228 39266 5264
rect 39210 5208 39212 5228
rect 39212 5208 39264 5228
rect 39264 5208 39266 5228
rect 39394 5208 39450 5264
rect 39026 4972 39028 4992
rect 39028 4972 39080 4992
rect 39080 4972 39082 4992
rect 39026 4936 39082 4972
rect 37956 4922 38012 4924
rect 38036 4922 38092 4924
rect 38116 4922 38172 4924
rect 38196 4922 38252 4924
rect 37956 4870 38002 4922
rect 38002 4870 38012 4922
rect 38036 4870 38066 4922
rect 38066 4870 38078 4922
rect 38078 4870 38092 4922
rect 38116 4870 38130 4922
rect 38130 4870 38142 4922
rect 38142 4870 38172 4922
rect 38196 4870 38206 4922
rect 38206 4870 38252 4922
rect 37956 4868 38012 4870
rect 38036 4868 38092 4870
rect 38116 4868 38172 4870
rect 38196 4868 38252 4870
rect 39394 4700 39396 4720
rect 39396 4700 39448 4720
rect 39448 4700 39450 4720
rect 39394 4664 39450 4700
rect 39946 4428 39948 4448
rect 39948 4428 40000 4448
rect 40000 4428 40002 4448
rect 39946 4392 40002 4428
rect 39016 4378 39072 4380
rect 39096 4378 39152 4380
rect 39176 4378 39232 4380
rect 39256 4378 39312 4380
rect 39016 4326 39062 4378
rect 39062 4326 39072 4378
rect 39096 4326 39126 4378
rect 39126 4326 39138 4378
rect 39138 4326 39152 4378
rect 39176 4326 39190 4378
rect 39190 4326 39202 4378
rect 39202 4326 39232 4378
rect 39256 4326 39266 4378
rect 39266 4326 39312 4378
rect 39016 4324 39072 4326
rect 39096 4324 39152 4326
rect 39176 4324 39232 4326
rect 39256 4324 39312 4326
rect 39394 4120 39450 4176
rect 39026 3884 39028 3904
rect 39028 3884 39080 3904
rect 39080 3884 39082 3904
rect 39026 3848 39082 3884
rect 37956 3834 38012 3836
rect 38036 3834 38092 3836
rect 38116 3834 38172 3836
rect 38196 3834 38252 3836
rect 37956 3782 38002 3834
rect 38002 3782 38012 3834
rect 38036 3782 38066 3834
rect 38066 3782 38078 3834
rect 38078 3782 38092 3834
rect 38116 3782 38130 3834
rect 38130 3782 38142 3834
rect 38142 3782 38172 3834
rect 38196 3782 38206 3834
rect 38206 3782 38252 3834
rect 37956 3780 38012 3782
rect 38036 3780 38092 3782
rect 38116 3780 38172 3782
rect 38196 3780 38252 3782
rect 39394 3612 39396 3632
rect 39396 3612 39448 3632
rect 39448 3612 39450 3632
rect 39394 3576 39450 3612
rect 39946 3340 39948 3360
rect 39948 3340 40000 3360
rect 40000 3340 40002 3360
rect 39946 3304 40002 3340
rect 39016 3290 39072 3292
rect 39096 3290 39152 3292
rect 39176 3290 39232 3292
rect 39256 3290 39312 3292
rect 39016 3238 39062 3290
rect 39062 3238 39072 3290
rect 39096 3238 39126 3290
rect 39126 3238 39138 3290
rect 39138 3238 39152 3290
rect 39176 3238 39190 3290
rect 39190 3238 39202 3290
rect 39202 3238 39232 3290
rect 39256 3238 39266 3290
rect 39266 3238 39312 3290
rect 39016 3236 39072 3238
rect 39096 3236 39152 3238
rect 39176 3236 39232 3238
rect 39256 3236 39312 3238
rect 39394 3032 39450 3088
rect 39026 2796 39028 2816
rect 39028 2796 39080 2816
rect 39080 2796 39082 2816
rect 39026 2760 39082 2796
rect 37956 2746 38012 2748
rect 38036 2746 38092 2748
rect 38116 2746 38172 2748
rect 38196 2746 38252 2748
rect 37956 2694 38002 2746
rect 38002 2694 38012 2746
rect 38036 2694 38066 2746
rect 38066 2694 38078 2746
rect 38078 2694 38092 2746
rect 38116 2694 38130 2746
rect 38130 2694 38142 2746
rect 38142 2694 38172 2746
rect 38196 2694 38206 2746
rect 38206 2694 38252 2746
rect 37956 2692 38012 2694
rect 38036 2692 38092 2694
rect 38116 2692 38172 2694
rect 38196 2692 38252 2694
rect 39394 2524 39396 2544
rect 39396 2524 39448 2544
rect 39448 2524 39450 2544
rect 39394 2488 39450 2524
rect 37922 1944 37978 2000
rect 38290 1672 38346 1728
rect 40406 2216 40462 2272
rect 39016 2202 39072 2204
rect 39096 2202 39152 2204
rect 39176 2202 39232 2204
rect 39256 2202 39312 2204
rect 39016 2150 39062 2202
rect 39062 2150 39072 2202
rect 39096 2150 39126 2202
rect 39126 2150 39138 2202
rect 39138 2150 39152 2202
rect 39176 2150 39190 2202
rect 39190 2150 39202 2202
rect 39202 2150 39232 2202
rect 39256 2150 39266 2202
rect 39266 2150 39312 2202
rect 39016 2148 39072 2150
rect 39096 2148 39152 2150
rect 39176 2148 39232 2150
rect 39256 2148 39312 2150
rect 38658 1400 38714 1456
<< metal3 >>
rect 0 9890 120 9920
rect 22553 9890 22619 9893
rect 0 9888 22619 9890
rect 0 9832 22558 9888
rect 22614 9832 22619 9888
rect 0 9830 22619 9832
rect 0 9800 120 9830
rect 22553 9827 22619 9830
rect 38377 9890 38443 9893
rect 40880 9890 41000 9920
rect 38377 9888 41000 9890
rect 38377 9832 38382 9888
rect 38438 9832 41000 9888
rect 38377 9830 41000 9832
rect 38377 9827 38443 9830
rect 40880 9800 41000 9830
rect 0 9618 120 9648
rect 14825 9618 14891 9621
rect 0 9616 14891 9618
rect 0 9560 14830 9616
rect 14886 9560 14891 9616
rect 0 9558 14891 9560
rect 0 9528 120 9558
rect 14825 9555 14891 9558
rect 37733 9618 37799 9621
rect 40880 9618 41000 9648
rect 37733 9616 41000 9618
rect 37733 9560 37738 9616
rect 37794 9560 41000 9616
rect 37733 9558 41000 9560
rect 37733 9555 37799 9558
rect 40880 9528 41000 9558
rect 0 9346 120 9376
rect 14917 9346 14983 9349
rect 0 9344 14983 9346
rect 0 9288 14922 9344
rect 14978 9288 14983 9344
rect 0 9286 14983 9288
rect 0 9256 120 9286
rect 14917 9283 14983 9286
rect 38285 9346 38351 9349
rect 40880 9346 41000 9376
rect 38285 9344 41000 9346
rect 38285 9288 38290 9344
rect 38346 9288 41000 9344
rect 38285 9286 41000 9288
rect 38285 9283 38351 9286
rect 40880 9256 41000 9286
rect 0 9074 120 9104
rect 18689 9074 18755 9077
rect 0 9072 18755 9074
rect 0 9016 18694 9072
rect 18750 9016 18755 9072
rect 0 9014 18755 9016
rect 0 8984 120 9014
rect 18689 9011 18755 9014
rect 39573 9074 39639 9077
rect 40880 9074 41000 9104
rect 39573 9072 41000 9074
rect 39573 9016 39578 9072
rect 39634 9016 41000 9072
rect 39573 9014 41000 9016
rect 39573 9011 39639 9014
rect 40880 8984 41000 9014
rect 0 8802 120 8832
rect 2773 8802 2839 8805
rect 0 8800 2839 8802
rect 0 8744 2778 8800
rect 2834 8744 2839 8800
rect 0 8742 2839 8744
rect 0 8712 120 8742
rect 2773 8739 2839 8742
rect 39481 8802 39547 8805
rect 40880 8802 41000 8832
rect 39481 8800 41000 8802
rect 39481 8744 39486 8800
rect 39542 8744 41000 8800
rect 39481 8742 41000 8744
rect 39481 8739 39547 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 33006 8671 33322 8672
rect 39006 8736 39322 8737
rect 39006 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39322 8736
rect 40880 8712 41000 8742
rect 39006 8671 39322 8672
rect 0 8530 120 8560
rect 22093 8530 22159 8533
rect 0 8528 22159 8530
rect 0 8472 22098 8528
rect 22154 8472 22159 8528
rect 0 8470 22159 8472
rect 0 8440 120 8470
rect 22093 8467 22159 8470
rect 38653 8530 38719 8533
rect 40880 8530 41000 8560
rect 38653 8528 41000 8530
rect 38653 8472 38658 8528
rect 38714 8472 41000 8528
rect 38653 8470 41000 8472
rect 38653 8467 38719 8470
rect 40880 8440 41000 8470
rect 2773 8394 2839 8397
rect 16481 8394 16547 8397
rect 2773 8392 16547 8394
rect 2773 8336 2778 8392
rect 2834 8336 16486 8392
rect 16542 8336 16547 8392
rect 2773 8334 16547 8336
rect 2773 8331 2839 8334
rect 16481 8331 16547 8334
rect 0 8258 120 8288
rect 1761 8258 1827 8261
rect 0 8256 1827 8258
rect 0 8200 1766 8256
rect 1822 8200 1827 8256
rect 0 8198 1827 8200
rect 0 8168 120 8198
rect 1761 8195 1827 8198
rect 39021 8258 39087 8261
rect 40880 8258 41000 8288
rect 39021 8256 41000 8258
rect 39021 8200 39026 8256
rect 39082 8200 41000 8256
rect 39021 8198 41000 8200
rect 39021 8195 39087 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 37946 8192 38262 8193
rect 37946 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38262 8192
rect 40880 8168 41000 8198
rect 37946 8127 38262 8128
rect 0 7986 120 8016
rect 19057 7986 19123 7989
rect 0 7984 19123 7986
rect 0 7928 19062 7984
rect 19118 7928 19123 7984
rect 0 7926 19123 7928
rect 0 7896 120 7926
rect 19057 7923 19123 7926
rect 39389 7986 39455 7989
rect 40880 7986 41000 8016
rect 39389 7984 41000 7986
rect 39389 7928 39394 7984
rect 39450 7928 41000 7984
rect 39389 7926 41000 7928
rect 39389 7923 39455 7926
rect 40880 7896 41000 7926
rect 1761 7850 1827 7853
rect 16389 7850 16455 7853
rect 1761 7848 16455 7850
rect 1761 7792 1766 7848
rect 1822 7792 16394 7848
rect 16450 7792 16455 7848
rect 1761 7790 16455 7792
rect 1761 7787 1827 7790
rect 16389 7787 16455 7790
rect 0 7714 120 7744
rect 39389 7714 39455 7717
rect 40880 7714 41000 7744
rect 0 7654 2790 7714
rect 0 7624 120 7654
rect 0 7442 120 7472
rect 1301 7442 1367 7445
rect 0 7440 1367 7442
rect 0 7384 1306 7440
rect 1362 7384 1367 7440
rect 0 7382 1367 7384
rect 2730 7442 2790 7654
rect 39389 7712 41000 7714
rect 39389 7656 39394 7712
rect 39450 7656 41000 7712
rect 39389 7654 41000 7656
rect 39389 7651 39455 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 33006 7583 33322 7584
rect 39006 7648 39322 7649
rect 39006 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39322 7648
rect 40880 7624 41000 7654
rect 39006 7583 39322 7584
rect 15101 7442 15167 7445
rect 2730 7440 15167 7442
rect 2730 7384 15106 7440
rect 15162 7384 15167 7440
rect 2730 7382 15167 7384
rect 0 7352 120 7382
rect 1301 7379 1367 7382
rect 15101 7379 15167 7382
rect 38929 7442 38995 7445
rect 40880 7442 41000 7472
rect 38929 7440 41000 7442
rect 38929 7384 38934 7440
rect 38990 7384 41000 7440
rect 38929 7382 41000 7384
rect 38929 7379 38995 7382
rect 40880 7352 41000 7382
rect 16481 7306 16547 7309
rect 1718 7304 16547 7306
rect 1718 7248 16486 7304
rect 16542 7248 16547 7304
rect 1718 7246 16547 7248
rect 0 7170 120 7200
rect 1718 7170 1778 7246
rect 16481 7243 16547 7246
rect 0 7110 1778 7170
rect 39389 7170 39455 7173
rect 40880 7170 41000 7200
rect 39389 7168 41000 7170
rect 39389 7112 39394 7168
rect 39450 7112 41000 7168
rect 39389 7110 41000 7112
rect 0 7080 120 7110
rect 39389 7107 39455 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 37946 7104 38262 7105
rect 37946 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38262 7104
rect 40880 7080 41000 7110
rect 37946 7039 38262 7040
rect 0 6898 120 6928
rect 17493 6898 17559 6901
rect 0 6896 17559 6898
rect 0 6840 17498 6896
rect 17554 6840 17559 6896
rect 0 6838 17559 6840
rect 0 6808 120 6838
rect 17493 6835 17559 6838
rect 39389 6898 39455 6901
rect 40880 6898 41000 6928
rect 39389 6896 41000 6898
rect 39389 6840 39394 6896
rect 39450 6840 41000 6896
rect 39389 6838 41000 6840
rect 39389 6835 39455 6838
rect 40880 6808 41000 6838
rect 17401 6762 17467 6765
rect 2730 6760 17467 6762
rect 2730 6704 17406 6760
rect 17462 6704 17467 6760
rect 2730 6702 17467 6704
rect 0 6626 120 6656
rect 2730 6626 2790 6702
rect 17401 6699 17467 6702
rect 17861 6762 17927 6765
rect 39205 6762 39271 6765
rect 17861 6760 39271 6762
rect 17861 6704 17866 6760
rect 17922 6704 39210 6760
rect 39266 6704 39271 6760
rect 17861 6702 39271 6704
rect 17861 6699 17927 6702
rect 39205 6699 39271 6702
rect 0 6566 2790 6626
rect 39941 6626 40007 6629
rect 40880 6626 41000 6656
rect 39941 6624 41000 6626
rect 39941 6568 39946 6624
rect 40002 6568 41000 6624
rect 39941 6566 41000 6568
rect 0 6536 120 6566
rect 39941 6563 40007 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 33006 6495 33322 6496
rect 39006 6560 39322 6561
rect 39006 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39322 6560
rect 40880 6536 41000 6566
rect 39006 6495 39322 6496
rect 9673 6490 9739 6493
rect 14825 6490 14891 6493
rect 9673 6488 14891 6490
rect 9673 6432 9678 6488
rect 9734 6432 14830 6488
rect 14886 6432 14891 6488
rect 9673 6430 14891 6432
rect 9673 6427 9739 6430
rect 14825 6427 14891 6430
rect 0 6354 120 6384
rect 11053 6354 11119 6357
rect 0 6352 11119 6354
rect 0 6296 11058 6352
rect 11114 6296 11119 6352
rect 0 6294 11119 6296
rect 0 6264 120 6294
rect 11053 6291 11119 6294
rect 11237 6354 11303 6357
rect 23565 6354 23631 6357
rect 11237 6352 23631 6354
rect 11237 6296 11242 6352
rect 11298 6296 23570 6352
rect 23626 6296 23631 6352
rect 11237 6294 23631 6296
rect 11237 6291 11303 6294
rect 23565 6291 23631 6294
rect 39389 6354 39455 6357
rect 40880 6354 41000 6384
rect 39389 6352 41000 6354
rect 39389 6296 39394 6352
rect 39450 6296 41000 6352
rect 39389 6294 41000 6296
rect 39389 6291 39455 6294
rect 40880 6264 41000 6294
rect 22369 6218 22435 6221
rect 1718 6216 22435 6218
rect 1718 6160 22374 6216
rect 22430 6160 22435 6216
rect 1718 6158 22435 6160
rect 0 6082 120 6112
rect 1718 6082 1778 6158
rect 22369 6155 22435 6158
rect 0 6022 1778 6082
rect 14825 6082 14891 6085
rect 19333 6082 19399 6085
rect 14825 6080 19399 6082
rect 14825 6024 14830 6080
rect 14886 6024 19338 6080
rect 19394 6024 19399 6080
rect 14825 6022 19399 6024
rect 0 5992 120 6022
rect 14825 6019 14891 6022
rect 19333 6019 19399 6022
rect 39021 6082 39087 6085
rect 40880 6082 41000 6112
rect 39021 6080 41000 6082
rect 39021 6024 39026 6080
rect 39082 6024 41000 6080
rect 39021 6022 41000 6024
rect 39021 6019 39087 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 37946 6016 38262 6017
rect 37946 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38262 6016
rect 40880 5992 41000 6022
rect 37946 5951 38262 5952
rect 0 5810 120 5840
rect 19793 5810 19859 5813
rect 0 5808 19859 5810
rect 0 5752 19798 5808
rect 19854 5752 19859 5808
rect 0 5750 19859 5752
rect 0 5720 120 5750
rect 19793 5747 19859 5750
rect 39389 5810 39455 5813
rect 40880 5810 41000 5840
rect 39389 5808 41000 5810
rect 39389 5752 39394 5808
rect 39450 5752 41000 5808
rect 39389 5750 41000 5752
rect 39389 5747 39455 5750
rect 40880 5720 41000 5750
rect 10961 5674 11027 5677
rect 14549 5674 14615 5677
rect 10961 5672 14615 5674
rect 10961 5616 10966 5672
rect 11022 5616 14554 5672
rect 14610 5616 14615 5672
rect 10961 5614 14615 5616
rect 10961 5611 11027 5614
rect 14549 5611 14615 5614
rect 19609 5674 19675 5677
rect 38837 5674 38903 5677
rect 19609 5672 38903 5674
rect 19609 5616 19614 5672
rect 19670 5616 38842 5672
rect 38898 5616 38903 5672
rect 19609 5614 38903 5616
rect 19609 5611 19675 5614
rect 38837 5611 38903 5614
rect 0 5538 120 5568
rect 565 5538 631 5541
rect 0 5536 631 5538
rect 0 5480 570 5536
rect 626 5480 631 5536
rect 0 5478 631 5480
rect 0 5448 120 5478
rect 565 5475 631 5478
rect 39941 5538 40007 5541
rect 40880 5538 41000 5568
rect 39941 5536 41000 5538
rect 39941 5480 39946 5536
rect 40002 5480 41000 5536
rect 39941 5478 41000 5480
rect 39941 5475 40007 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 33006 5407 33322 5408
rect 39006 5472 39322 5473
rect 39006 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39322 5472
rect 40880 5448 41000 5478
rect 39006 5407 39322 5408
rect 0 5266 120 5296
rect 19149 5266 19215 5269
rect 0 5264 19215 5266
rect 0 5208 19154 5264
rect 19210 5208 19215 5264
rect 0 5206 19215 5208
rect 0 5176 120 5206
rect 19149 5203 19215 5206
rect 19333 5266 19399 5269
rect 39205 5266 39271 5269
rect 19333 5264 39271 5266
rect 19333 5208 19338 5264
rect 19394 5208 39210 5264
rect 39266 5208 39271 5264
rect 19333 5206 39271 5208
rect 19333 5203 19399 5206
rect 39205 5203 39271 5206
rect 39389 5266 39455 5269
rect 40880 5266 41000 5296
rect 39389 5264 41000 5266
rect 39389 5208 39394 5264
rect 39450 5208 41000 5264
rect 39389 5206 41000 5208
rect 39389 5203 39455 5206
rect 40880 5176 41000 5206
rect 2773 5130 2839 5133
rect 23473 5130 23539 5133
rect 2773 5128 23539 5130
rect 2773 5072 2778 5128
rect 2834 5072 23478 5128
rect 23534 5072 23539 5128
rect 2773 5070 23539 5072
rect 2773 5067 2839 5070
rect 23473 5067 23539 5070
rect 0 4994 120 5024
rect 1761 4994 1827 4997
rect 0 4992 1827 4994
rect 0 4936 1766 4992
rect 1822 4936 1827 4992
rect 0 4934 1827 4936
rect 0 4904 120 4934
rect 1761 4931 1827 4934
rect 39021 4994 39087 4997
rect 40880 4994 41000 5024
rect 39021 4992 41000 4994
rect 39021 4936 39026 4992
rect 39082 4936 41000 4992
rect 39021 4934 41000 4936
rect 39021 4931 39087 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 37946 4928 38262 4929
rect 37946 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38262 4928
rect 40880 4904 41000 4934
rect 37946 4863 38262 4864
rect 0 4722 120 4752
rect 22829 4722 22895 4725
rect 0 4720 22895 4722
rect 0 4664 22834 4720
rect 22890 4664 22895 4720
rect 0 4662 22895 4664
rect 0 4632 120 4662
rect 22829 4659 22895 4662
rect 39389 4722 39455 4725
rect 40880 4722 41000 4752
rect 39389 4720 41000 4722
rect 39389 4664 39394 4720
rect 39450 4664 41000 4720
rect 39389 4662 41000 4664
rect 39389 4659 39455 4662
rect 40880 4632 41000 4662
rect 1761 4586 1827 4589
rect 21541 4586 21607 4589
rect 1761 4584 21607 4586
rect 1761 4528 1766 4584
rect 1822 4528 21546 4584
rect 21602 4528 21607 4584
rect 1761 4526 21607 4528
rect 1761 4523 1827 4526
rect 21541 4523 21607 4526
rect 0 4450 120 4480
rect 2773 4450 2839 4453
rect 0 4448 2839 4450
rect 0 4392 2778 4448
rect 2834 4392 2839 4448
rect 0 4390 2839 4392
rect 0 4360 120 4390
rect 2773 4387 2839 4390
rect 39941 4450 40007 4453
rect 40880 4450 41000 4480
rect 39941 4448 41000 4450
rect 39941 4392 39946 4448
rect 40002 4392 41000 4448
rect 39941 4390 41000 4392
rect 39941 4387 40007 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 33006 4319 33322 4320
rect 39006 4384 39322 4385
rect 39006 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39322 4384
rect 40880 4360 41000 4390
rect 39006 4319 39322 4320
rect 0 4178 120 4208
rect 24025 4178 24091 4181
rect 0 4176 24091 4178
rect 0 4120 24030 4176
rect 24086 4120 24091 4176
rect 0 4118 24091 4120
rect 0 4088 120 4118
rect 24025 4115 24091 4118
rect 39389 4178 39455 4181
rect 40880 4178 41000 4208
rect 39389 4176 41000 4178
rect 39389 4120 39394 4176
rect 39450 4120 41000 4176
rect 39389 4118 41000 4120
rect 39389 4115 39455 4118
rect 40880 4088 41000 4118
rect 20621 4042 20687 4045
rect 28165 4042 28231 4045
rect 1718 4040 20687 4042
rect 1718 3984 20626 4040
rect 20682 3984 20687 4040
rect 1718 3982 20687 3984
rect 0 3906 120 3936
rect 1718 3906 1778 3982
rect 20621 3979 20687 3982
rect 22050 4040 28231 4042
rect 22050 3984 28170 4040
rect 28226 3984 28231 4040
rect 22050 3982 28231 3984
rect 0 3846 1778 3906
rect 20437 3906 20503 3909
rect 22050 3906 22110 3982
rect 28165 3979 28231 3982
rect 20437 3904 22110 3906
rect 20437 3848 20442 3904
rect 20498 3848 22110 3904
rect 20437 3846 22110 3848
rect 39021 3906 39087 3909
rect 40880 3906 41000 3936
rect 39021 3904 41000 3906
rect 39021 3848 39026 3904
rect 39082 3848 41000 3904
rect 39021 3846 41000 3848
rect 0 3816 120 3846
rect 20437 3843 20503 3846
rect 39021 3843 39087 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 37946 3840 38262 3841
rect 37946 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38262 3840
rect 40880 3816 41000 3846
rect 37946 3775 38262 3776
rect 20345 3770 20411 3773
rect 20345 3768 25882 3770
rect 20345 3712 20350 3768
rect 20406 3712 25882 3768
rect 20345 3710 25882 3712
rect 20345 3707 20411 3710
rect 0 3634 120 3664
rect 24209 3634 24275 3637
rect 0 3632 24275 3634
rect 0 3576 24214 3632
rect 24270 3576 24275 3632
rect 0 3574 24275 3576
rect 25822 3634 25882 3710
rect 26325 3634 26391 3637
rect 25822 3632 26391 3634
rect 25822 3576 26330 3632
rect 26386 3576 26391 3632
rect 25822 3574 26391 3576
rect 0 3544 120 3574
rect 24209 3571 24275 3574
rect 26325 3571 26391 3574
rect 26509 3634 26575 3637
rect 36629 3634 36695 3637
rect 26509 3632 36695 3634
rect 26509 3576 26514 3632
rect 26570 3576 36634 3632
rect 36690 3576 36695 3632
rect 26509 3574 36695 3576
rect 26509 3571 26575 3574
rect 36629 3571 36695 3574
rect 39389 3634 39455 3637
rect 40880 3634 41000 3664
rect 39389 3632 41000 3634
rect 39389 3576 39394 3632
rect 39450 3576 41000 3632
rect 39389 3574 41000 3576
rect 39389 3571 39455 3574
rect 40880 3544 41000 3574
rect 24393 3498 24459 3501
rect 2730 3496 24459 3498
rect 2730 3440 24398 3496
rect 24454 3440 24459 3496
rect 2730 3438 24459 3440
rect 0 3362 120 3392
rect 2730 3362 2790 3438
rect 24393 3435 24459 3438
rect 28349 3498 28415 3501
rect 34421 3498 34487 3501
rect 28349 3496 34487 3498
rect 28349 3440 28354 3496
rect 28410 3440 34426 3496
rect 34482 3440 34487 3496
rect 28349 3438 34487 3440
rect 28349 3435 28415 3438
rect 34421 3435 34487 3438
rect 0 3302 2790 3362
rect 17309 3362 17375 3365
rect 20345 3362 20411 3365
rect 17309 3360 20411 3362
rect 17309 3304 17314 3360
rect 17370 3304 20350 3360
rect 20406 3304 20411 3360
rect 17309 3302 20411 3304
rect 0 3272 120 3302
rect 17309 3299 17375 3302
rect 20345 3299 20411 3302
rect 39941 3362 40007 3365
rect 40880 3362 41000 3392
rect 39941 3360 41000 3362
rect 39941 3304 39946 3360
rect 40002 3304 41000 3360
rect 39941 3302 41000 3304
rect 39941 3299 40007 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 33006 3231 33322 3232
rect 39006 3296 39322 3297
rect 39006 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39322 3296
rect 40880 3272 41000 3302
rect 39006 3231 39322 3232
rect 17033 3226 17099 3229
rect 20437 3226 20503 3229
rect 17033 3224 20503 3226
rect 17033 3168 17038 3224
rect 17094 3168 20442 3224
rect 20498 3168 20503 3224
rect 17033 3166 20503 3168
rect 17033 3163 17099 3166
rect 20437 3163 20503 3166
rect 0 3090 120 3120
rect 24117 3090 24183 3093
rect 0 3088 24183 3090
rect 0 3032 24122 3088
rect 24178 3032 24183 3088
rect 0 3030 24183 3032
rect 0 3000 120 3030
rect 24117 3027 24183 3030
rect 27981 3090 28047 3093
rect 34145 3090 34211 3093
rect 27981 3088 34211 3090
rect 27981 3032 27986 3088
rect 28042 3032 34150 3088
rect 34206 3032 34211 3088
rect 27981 3030 34211 3032
rect 27981 3027 28047 3030
rect 34145 3027 34211 3030
rect 39389 3090 39455 3093
rect 40880 3090 41000 3120
rect 39389 3088 41000 3090
rect 39389 3032 39394 3088
rect 39450 3032 41000 3088
rect 39389 3030 41000 3032
rect 39389 3027 39455 3030
rect 40880 3000 41000 3030
rect 20621 2954 20687 2957
rect 22093 2954 22159 2957
rect 1718 2894 20546 2954
rect 0 2818 120 2848
rect 1718 2818 1778 2894
rect 0 2758 1778 2818
rect 20486 2818 20546 2894
rect 20621 2952 22159 2954
rect 20621 2896 20626 2952
rect 20682 2896 22098 2952
rect 22154 2896 22159 2952
rect 20621 2894 22159 2896
rect 20621 2891 20687 2894
rect 22093 2891 22159 2894
rect 24945 2818 25011 2821
rect 20486 2816 25011 2818
rect 20486 2760 24950 2816
rect 25006 2760 25011 2816
rect 20486 2758 25011 2760
rect 0 2728 120 2758
rect 24945 2755 25011 2758
rect 39021 2818 39087 2821
rect 40880 2818 41000 2848
rect 39021 2816 41000 2818
rect 39021 2760 39026 2816
rect 39082 2760 41000 2816
rect 39021 2758 41000 2760
rect 39021 2755 39087 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 37946 2752 38262 2753
rect 37946 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38262 2752
rect 40880 2728 41000 2758
rect 37946 2687 38262 2688
rect 22461 2682 22527 2685
rect 22737 2682 22803 2685
rect 26785 2682 26851 2685
rect 22461 2680 22803 2682
rect 22461 2624 22466 2680
rect 22522 2624 22742 2680
rect 22798 2624 22803 2680
rect 22461 2622 22803 2624
rect 22461 2619 22527 2622
rect 22737 2619 22803 2622
rect 26558 2680 26851 2682
rect 26558 2624 26790 2680
rect 26846 2624 26851 2680
rect 26558 2622 26851 2624
rect 0 2546 120 2576
rect 8661 2546 8727 2549
rect 0 2544 8727 2546
rect 0 2488 8666 2544
rect 8722 2488 8727 2544
rect 0 2486 8727 2488
rect 0 2456 120 2486
rect 8661 2483 8727 2486
rect 14365 2546 14431 2549
rect 26049 2546 26115 2549
rect 14365 2544 26115 2546
rect 14365 2488 14370 2544
rect 14426 2488 26054 2544
rect 26110 2488 26115 2544
rect 14365 2486 26115 2488
rect 14365 2483 14431 2486
rect 26049 2483 26115 2486
rect 26325 2546 26391 2549
rect 26558 2546 26618 2622
rect 26785 2619 26851 2622
rect 26325 2544 26618 2546
rect 26325 2488 26330 2544
rect 26386 2488 26618 2544
rect 26325 2486 26618 2488
rect 39389 2546 39455 2549
rect 40880 2546 41000 2576
rect 39389 2544 41000 2546
rect 39389 2488 39394 2544
rect 39450 2488 41000 2544
rect 39389 2486 41000 2488
rect 26325 2483 26391 2486
rect 39389 2483 39455 2486
rect 40880 2456 41000 2486
rect 11881 2410 11947 2413
rect 16573 2410 16639 2413
rect 2822 2408 11947 2410
rect 2822 2352 11886 2408
rect 11942 2352 11947 2408
rect 2822 2350 11947 2352
rect 0 2274 120 2304
rect 2822 2274 2882 2350
rect 11881 2347 11947 2350
rect 12022 2408 16639 2410
rect 12022 2352 16578 2408
rect 16634 2352 16639 2408
rect 12022 2350 16639 2352
rect 0 2214 2882 2274
rect 9857 2274 9923 2277
rect 12022 2274 12082 2350
rect 16573 2347 16639 2350
rect 16757 2410 16823 2413
rect 28993 2410 29059 2413
rect 16757 2408 29059 2410
rect 16757 2352 16762 2408
rect 16818 2352 28998 2408
rect 29054 2352 29059 2408
rect 16757 2350 29059 2352
rect 16757 2347 16823 2350
rect 28993 2347 29059 2350
rect 9857 2272 12082 2274
rect 9857 2216 9862 2272
rect 9918 2216 12082 2272
rect 9857 2214 12082 2216
rect 40401 2274 40467 2277
rect 40880 2274 41000 2304
rect 40401 2272 41000 2274
rect 40401 2216 40406 2272
rect 40462 2216 41000 2272
rect 40401 2214 41000 2216
rect 0 2184 120 2214
rect 9857 2211 9923 2214
rect 40401 2211 40467 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 33006 2143 33322 2144
rect 39006 2208 39322 2209
rect 39006 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39322 2208
rect 40880 2184 41000 2214
rect 39006 2143 39322 2144
rect 0 2002 120 2032
rect 15101 2002 15167 2005
rect 0 2000 15167 2002
rect 0 1944 15106 2000
rect 15162 1944 15167 2000
rect 0 1942 15167 1944
rect 0 1912 120 1942
rect 15101 1939 15167 1942
rect 15285 2002 15351 2005
rect 24853 2002 24919 2005
rect 15285 2000 24919 2002
rect 15285 1944 15290 2000
rect 15346 1944 24858 2000
rect 24914 1944 24919 2000
rect 15285 1942 24919 1944
rect 15285 1939 15351 1942
rect 24853 1939 24919 1942
rect 37917 2002 37983 2005
rect 40880 2002 41000 2032
rect 37917 2000 41000 2002
rect 37917 1944 37922 2000
rect 37978 1944 41000 2000
rect 37917 1942 41000 1944
rect 37917 1939 37983 1942
rect 40880 1912 41000 1942
rect 13169 1866 13235 1869
rect 26601 1866 26667 1869
rect 13169 1864 26667 1866
rect 13169 1808 13174 1864
rect 13230 1808 26606 1864
rect 26662 1808 26667 1864
rect 13169 1806 26667 1808
rect 13169 1803 13235 1806
rect 26601 1803 26667 1806
rect 0 1730 120 1760
rect 9581 1730 9647 1733
rect 0 1728 9647 1730
rect 0 1672 9586 1728
rect 9642 1672 9647 1728
rect 0 1670 9647 1672
rect 0 1640 120 1670
rect 9581 1667 9647 1670
rect 13629 1730 13695 1733
rect 15285 1730 15351 1733
rect 13629 1728 15351 1730
rect 13629 1672 13634 1728
rect 13690 1672 15290 1728
rect 15346 1672 15351 1728
rect 13629 1670 15351 1672
rect 13629 1667 13695 1670
rect 15285 1667 15351 1670
rect 22737 1730 22803 1733
rect 32765 1730 32831 1733
rect 22737 1728 32831 1730
rect 22737 1672 22742 1728
rect 22798 1672 32770 1728
rect 32826 1672 32831 1728
rect 22737 1670 32831 1672
rect 22737 1667 22803 1670
rect 32765 1667 32831 1670
rect 38285 1730 38351 1733
rect 40880 1730 41000 1760
rect 38285 1728 41000 1730
rect 38285 1672 38290 1728
rect 38346 1672 41000 1728
rect 38285 1670 41000 1672
rect 38285 1667 38351 1670
rect 40880 1640 41000 1670
rect 8753 1594 8819 1597
rect 18505 1594 18571 1597
rect 8753 1592 18571 1594
rect 8753 1536 8758 1592
rect 8814 1536 18510 1592
rect 18566 1536 18571 1592
rect 8753 1534 18571 1536
rect 8753 1531 8819 1534
rect 18505 1531 18571 1534
rect 0 1458 120 1488
rect 5533 1458 5599 1461
rect 0 1456 5599 1458
rect 0 1400 5538 1456
rect 5594 1400 5599 1456
rect 0 1398 5599 1400
rect 0 1368 120 1398
rect 5533 1395 5599 1398
rect 38653 1458 38719 1461
rect 40880 1458 41000 1488
rect 38653 1456 41000 1458
rect 38653 1400 38658 1456
rect 38714 1400 41000 1456
rect 38653 1398 41000 1400
rect 38653 1395 38719 1398
rect 40880 1368 41000 1398
rect 27429 1322 27495 1325
rect 34973 1322 35039 1325
rect 27429 1320 35039 1322
rect 27429 1264 27434 1320
rect 27490 1264 34978 1320
rect 35034 1264 35039 1320
rect 27429 1262 35039 1264
rect 27429 1259 27495 1262
rect 34973 1259 35039 1262
rect 13721 370 13787 373
rect 26325 370 26391 373
rect 13721 368 26391 370
rect 13721 312 13726 368
rect 13782 312 26330 368
rect 26386 312 26391 368
rect 13721 310 26391 312
rect 13721 307 13787 310
rect 26325 307 26391 310
rect 14549 234 14615 237
rect 29545 234 29611 237
rect 14549 232 29611 234
rect 14549 176 14554 232
rect 14610 176 29550 232
rect 29606 176 29611 232
rect 14549 174 29611 176
rect 14549 171 14615 174
rect 29545 171 29611 174
rect 14825 98 14891 101
rect 31293 98 31359 101
rect 14825 96 31359 98
rect 14825 40 14830 96
rect 14886 40 31298 96
rect 31354 40 31359 96
rect 14825 38 31359 40
rect 14825 35 14891 38
rect 31293 35 31359 38
<< via3 >>
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 39012 8732 39076 8736
rect 39012 8676 39016 8732
rect 39016 8676 39072 8732
rect 39072 8676 39076 8732
rect 39012 8672 39076 8676
rect 39092 8732 39156 8736
rect 39092 8676 39096 8732
rect 39096 8676 39152 8732
rect 39152 8676 39156 8732
rect 39092 8672 39156 8676
rect 39172 8732 39236 8736
rect 39172 8676 39176 8732
rect 39176 8676 39232 8732
rect 39232 8676 39236 8732
rect 39172 8672 39236 8676
rect 39252 8732 39316 8736
rect 39252 8676 39256 8732
rect 39256 8676 39312 8732
rect 39312 8676 39316 8732
rect 39252 8672 39316 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 37952 8188 38016 8192
rect 37952 8132 37956 8188
rect 37956 8132 38012 8188
rect 38012 8132 38016 8188
rect 37952 8128 38016 8132
rect 38032 8188 38096 8192
rect 38032 8132 38036 8188
rect 38036 8132 38092 8188
rect 38092 8132 38096 8188
rect 38032 8128 38096 8132
rect 38112 8188 38176 8192
rect 38112 8132 38116 8188
rect 38116 8132 38172 8188
rect 38172 8132 38176 8188
rect 38112 8128 38176 8132
rect 38192 8188 38256 8192
rect 38192 8132 38196 8188
rect 38196 8132 38252 8188
rect 38252 8132 38256 8188
rect 38192 8128 38256 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 39012 7644 39076 7648
rect 39012 7588 39016 7644
rect 39016 7588 39072 7644
rect 39072 7588 39076 7644
rect 39012 7584 39076 7588
rect 39092 7644 39156 7648
rect 39092 7588 39096 7644
rect 39096 7588 39152 7644
rect 39152 7588 39156 7644
rect 39092 7584 39156 7588
rect 39172 7644 39236 7648
rect 39172 7588 39176 7644
rect 39176 7588 39232 7644
rect 39232 7588 39236 7644
rect 39172 7584 39236 7588
rect 39252 7644 39316 7648
rect 39252 7588 39256 7644
rect 39256 7588 39312 7644
rect 39312 7588 39316 7644
rect 39252 7584 39316 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 37952 7100 38016 7104
rect 37952 7044 37956 7100
rect 37956 7044 38012 7100
rect 38012 7044 38016 7100
rect 37952 7040 38016 7044
rect 38032 7100 38096 7104
rect 38032 7044 38036 7100
rect 38036 7044 38092 7100
rect 38092 7044 38096 7100
rect 38032 7040 38096 7044
rect 38112 7100 38176 7104
rect 38112 7044 38116 7100
rect 38116 7044 38172 7100
rect 38172 7044 38176 7100
rect 38112 7040 38176 7044
rect 38192 7100 38256 7104
rect 38192 7044 38196 7100
rect 38196 7044 38252 7100
rect 38252 7044 38256 7100
rect 38192 7040 38256 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 39012 6556 39076 6560
rect 39012 6500 39016 6556
rect 39016 6500 39072 6556
rect 39072 6500 39076 6556
rect 39012 6496 39076 6500
rect 39092 6556 39156 6560
rect 39092 6500 39096 6556
rect 39096 6500 39152 6556
rect 39152 6500 39156 6556
rect 39092 6496 39156 6500
rect 39172 6556 39236 6560
rect 39172 6500 39176 6556
rect 39176 6500 39232 6556
rect 39232 6500 39236 6556
rect 39172 6496 39236 6500
rect 39252 6556 39316 6560
rect 39252 6500 39256 6556
rect 39256 6500 39312 6556
rect 39312 6500 39316 6556
rect 39252 6496 39316 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 37952 6012 38016 6016
rect 37952 5956 37956 6012
rect 37956 5956 38012 6012
rect 38012 5956 38016 6012
rect 37952 5952 38016 5956
rect 38032 6012 38096 6016
rect 38032 5956 38036 6012
rect 38036 5956 38092 6012
rect 38092 5956 38096 6012
rect 38032 5952 38096 5956
rect 38112 6012 38176 6016
rect 38112 5956 38116 6012
rect 38116 5956 38172 6012
rect 38172 5956 38176 6012
rect 38112 5952 38176 5956
rect 38192 6012 38256 6016
rect 38192 5956 38196 6012
rect 38196 5956 38252 6012
rect 38252 5956 38256 6012
rect 38192 5952 38256 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 39012 5468 39076 5472
rect 39012 5412 39016 5468
rect 39016 5412 39072 5468
rect 39072 5412 39076 5468
rect 39012 5408 39076 5412
rect 39092 5468 39156 5472
rect 39092 5412 39096 5468
rect 39096 5412 39152 5468
rect 39152 5412 39156 5468
rect 39092 5408 39156 5412
rect 39172 5468 39236 5472
rect 39172 5412 39176 5468
rect 39176 5412 39232 5468
rect 39232 5412 39236 5468
rect 39172 5408 39236 5412
rect 39252 5468 39316 5472
rect 39252 5412 39256 5468
rect 39256 5412 39312 5468
rect 39312 5412 39316 5468
rect 39252 5408 39316 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 37952 4924 38016 4928
rect 37952 4868 37956 4924
rect 37956 4868 38012 4924
rect 38012 4868 38016 4924
rect 37952 4864 38016 4868
rect 38032 4924 38096 4928
rect 38032 4868 38036 4924
rect 38036 4868 38092 4924
rect 38092 4868 38096 4924
rect 38032 4864 38096 4868
rect 38112 4924 38176 4928
rect 38112 4868 38116 4924
rect 38116 4868 38172 4924
rect 38172 4868 38176 4924
rect 38112 4864 38176 4868
rect 38192 4924 38256 4928
rect 38192 4868 38196 4924
rect 38196 4868 38252 4924
rect 38252 4868 38256 4924
rect 38192 4864 38256 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 39012 4380 39076 4384
rect 39012 4324 39016 4380
rect 39016 4324 39072 4380
rect 39072 4324 39076 4380
rect 39012 4320 39076 4324
rect 39092 4380 39156 4384
rect 39092 4324 39096 4380
rect 39096 4324 39152 4380
rect 39152 4324 39156 4380
rect 39092 4320 39156 4324
rect 39172 4380 39236 4384
rect 39172 4324 39176 4380
rect 39176 4324 39232 4380
rect 39232 4324 39236 4380
rect 39172 4320 39236 4324
rect 39252 4380 39316 4384
rect 39252 4324 39256 4380
rect 39256 4324 39312 4380
rect 39312 4324 39316 4380
rect 39252 4320 39316 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 37952 3836 38016 3840
rect 37952 3780 37956 3836
rect 37956 3780 38012 3836
rect 38012 3780 38016 3836
rect 37952 3776 38016 3780
rect 38032 3836 38096 3840
rect 38032 3780 38036 3836
rect 38036 3780 38092 3836
rect 38092 3780 38096 3836
rect 38032 3776 38096 3780
rect 38112 3836 38176 3840
rect 38112 3780 38116 3836
rect 38116 3780 38172 3836
rect 38172 3780 38176 3836
rect 38112 3776 38176 3780
rect 38192 3836 38256 3840
rect 38192 3780 38196 3836
rect 38196 3780 38252 3836
rect 38252 3780 38256 3836
rect 38192 3776 38256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 39012 3292 39076 3296
rect 39012 3236 39016 3292
rect 39016 3236 39072 3292
rect 39072 3236 39076 3292
rect 39012 3232 39076 3236
rect 39092 3292 39156 3296
rect 39092 3236 39096 3292
rect 39096 3236 39152 3292
rect 39152 3236 39156 3292
rect 39092 3232 39156 3236
rect 39172 3292 39236 3296
rect 39172 3236 39176 3292
rect 39176 3236 39232 3292
rect 39232 3236 39236 3292
rect 39172 3232 39236 3236
rect 39252 3292 39316 3296
rect 39252 3236 39256 3292
rect 39256 3236 39312 3292
rect 39312 3236 39316 3292
rect 39252 3232 39316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 37952 2748 38016 2752
rect 37952 2692 37956 2748
rect 37956 2692 38012 2748
rect 38012 2692 38016 2748
rect 37952 2688 38016 2692
rect 38032 2748 38096 2752
rect 38032 2692 38036 2748
rect 38036 2692 38092 2748
rect 38092 2692 38096 2748
rect 38032 2688 38096 2692
rect 38112 2748 38176 2752
rect 38112 2692 38116 2748
rect 38116 2692 38172 2748
rect 38172 2692 38176 2748
rect 38112 2688 38176 2692
rect 38192 2748 38256 2752
rect 38192 2692 38196 2748
rect 38196 2692 38252 2748
rect 38252 2692 38256 2748
rect 38192 2688 38256 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
rect 39012 2204 39076 2208
rect 39012 2148 39016 2204
rect 39016 2148 39072 2204
rect 39072 2148 39076 2204
rect 39012 2144 39076 2148
rect 39092 2204 39156 2208
rect 39092 2148 39096 2204
rect 39096 2148 39152 2204
rect 39152 2148 39156 2204
rect 39092 2144 39156 2148
rect 39172 2204 39236 2208
rect 39172 2148 39176 2204
rect 39176 2148 39232 2204
rect 39232 2148 39236 2204
rect 39172 2144 39236 2148
rect 39252 2204 39316 2208
rect 39252 2148 39256 2204
rect 39256 2148 39312 2204
rect 39312 2148 39316 2204
rect 39252 2144 39316 2148
<< metal4 >>
rect 1944 8192 2264 11250
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 8736 3324 11250
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11250
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 8736 9324 11250
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 8192 14264 11250
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13944 0 14264 2688
rect 15004 8736 15324 11250
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 8192 20264 11250
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19944 0 20264 2688
rect 21004 8736 21324 11250
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 21004 6560 21324 7584
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25944 8192 26264 11250
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25944 0 26264 2688
rect 27004 8736 27324 11250
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 31944 8192 32264 11250
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 0 32264 2688
rect 33004 8736 33324 11250
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
rect 37944 8192 38264 11250
rect 37944 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38264 8192
rect 37944 7104 38264 8128
rect 37944 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38264 7104
rect 37944 6016 38264 7040
rect 37944 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38264 6016
rect 37944 4928 38264 5952
rect 37944 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38264 4928
rect 37944 3840 38264 4864
rect 37944 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38264 3840
rect 37944 2752 38264 3776
rect 37944 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38264 2752
rect 37944 0 38264 2688
rect 39004 8736 39324 11250
rect 39004 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39324 8736
rect 39004 7648 39324 8672
rect 39004 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39324 7648
rect 39004 6560 39324 7584
rect 39004 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39324 6560
rect 39004 5472 39324 6496
rect 39004 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39324 5472
rect 39004 4384 39324 5408
rect 39004 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39324 4384
rect 39004 3296 39324 4320
rect 39004 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39324 3296
rect 39004 2208 39324 3232
rect 39004 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39324 2208
rect 39004 0 39324 2144
use sky130_fd_sc_hd__buf_1  _000_
timestamp -3599
transform 1 0 21712 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _001_
timestamp -3599
transform 1 0 22816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _002_
timestamp -3599
transform 1 0 23092 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _003_
timestamp -3599
transform 1 0 23368 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _004_
timestamp -3599
transform 1 0 22356 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _005_
timestamp -3599
transform 1 0 24932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _006_
timestamp -3599
transform 1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _007_
timestamp -3599
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _008_
timestamp -3599
transform 1 0 24380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _009_
timestamp -3599
transform 1 0 22172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _010_
timestamp -3599
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _011_
timestamp -3599
transform 1 0 23644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _012_
timestamp -3599
transform 1 0 23000 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _013_
timestamp -3599
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _014_
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _015_
timestamp -3599
transform 1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _016_
timestamp -3599
transform 1 0 20240 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _017_
timestamp -3599
transform 1 0 22356 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _018_
timestamp -3599
transform 1 0 17756 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _019_
timestamp -3599
transform 1 0 19688 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _020_
timestamp -3599
transform 1 0 17664 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _021_
timestamp -3599
transform 1 0 16928 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _022_
timestamp -3599
transform 1 0 23000 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _023_
timestamp -3599
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _024_
timestamp -3599
transform 1 0 20516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _025_
timestamp -3599
transform 1 0 19964 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _026_
timestamp -3599
transform 1 0 22172 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _027_
timestamp -3599
transform 1 0 19044 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _028_
timestamp -3599
transform 1 0 19596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _029_
timestamp -3599
transform -1 0 17480 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _030_
timestamp -3599
transform 1 0 17756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _031_
timestamp -3599
transform 1 0 22724 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _032_
timestamp -3599
transform -1 0 21068 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _033_
timestamp -3599
transform -1 0 18400 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _034_
timestamp -3599
transform -1 0 22448 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _035_
timestamp -3599
transform 1 0 19320 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _036_
timestamp -3599
transform -1 0 26220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _037_
timestamp -3599
transform -1 0 27784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _038_
timestamp -3599
transform -1 0 28060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _039_
timestamp -3599
transform -1 0 28336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp -3599
transform 1 0 28336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp -3599
transform 1 0 27140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp -3599
transform 1 0 28612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp -3599
transform 1 0 27416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp -3599
transform -1 0 26404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp -3599
transform -1 0 25668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp -3599
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp -3599
transform -1 0 26772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp -3599
transform -1 0 31096 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp -3599
transform -1 0 33396 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp -3599
transform -1 0 35972 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp -3599
transform 1 0 36892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _052_
timestamp -3599
transform 1 0 2944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _053_
timestamp -3599
transform 1 0 2668 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _054_
timestamp -3599
transform 1 0 3220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _055_
timestamp -3599
transform 1 0 2944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _056_
timestamp -3599
transform 1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _057_
timestamp -3599
transform 1 0 4232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _058_
timestamp -3599
transform 1 0 4692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _059_
timestamp -3599
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _060_
timestamp -3599
transform 1 0 7544 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _061_
timestamp -3599
transform 1 0 9016 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _062_
timestamp -3599
transform 1 0 10396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _063_
timestamp -3599
transform 1 0 11408 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _064_
timestamp -3599
transform 1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _065_
timestamp -3599
transform 1 0 9292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _066_
timestamp -3599
transform 1 0 9016 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _067_
timestamp -3599
transform 1 0 9568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _068_
timestamp -3599
transform 1 0 9936 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _069_
timestamp -3599
transform 1 0 10672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _070_
timestamp -3599
transform 1 0 11040 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _071_
timestamp -3599
transform 1 0 11684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp -3599
transform -1 0 15916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp -3599
transform -1 0 15180 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _074_
timestamp -3599
transform 1 0 14260 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _075_
timestamp -3599
transform 1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _076_
timestamp -3599
transform 1 0 13616 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _077_
timestamp -3599
transform 1 0 14168 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _078_
timestamp -3599
transform 1 0 13432 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _079_
timestamp -3599
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _080_
timestamp -3599
transform 1 0 14536 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _081_
timestamp -3599
transform 1 0 15364 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _082_
timestamp -3599
transform 1 0 15916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _083_
timestamp -3599
transform 1 0 16560 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp -3599
transform -1 0 17296 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp -3599
transform -1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp -3599
transform -1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp -3599
transform -1 0 18952 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp -3599
transform -1 0 27600 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp -3599
transform -1 0 28428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp -3599
transform 1 0 29164 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp -3599
transform 1 0 29992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp -3599
transform 1 0 30636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp -3599
transform 1 0 31096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp -3599
transform 1 0 31372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp -3599
transform 1 0 32016 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp -3599
transform 1 0 32292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp -3599
transform 1 0 31740 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp -3599
transform -1 0 30544 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp -3599
transform -1 0 29900 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp -3599
transform -1 0 29440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp -3599
transform -1 0 28980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp -3599
transform -1 0 27692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp -3599
transform -1 0 26772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp -3599
transform -1 0 22172 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform -1 0 24564 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform -1 0 23644 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform 1 0 22816 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform -1 0 21712 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform -1 0 19688 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform 1 0 20056 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 17756 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform 1 0 19504 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform -1 0 22816 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform 1 0 17480 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform -1 0 17664 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform -1 0 16560 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform -1 0 20516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform -1 0 21252 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform -1 0 22172 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform -1 0 19044 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp -3599
transform -1 0 18860 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp -3599
transform -1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp -3599
transform -1 0 23828 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp -3599
transform -1 0 18584 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp -3599
transform -1 0 22724 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp -3599
transform -1 0 24012 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp -3599
transform -1 0 22356 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp -3599
transform -1 0 25392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp -3599
transform -1 0 24288 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp -3599
transform -1 0 25576 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp -3599
transform 1 0 24196 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp -3599
transform -1 0 22632 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp -3599
transform 1 0 39008 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp -3599
transform 1 0 21252 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp -3599
transform -1 0 16192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp -3599
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp -3599
transform -1 0 18400 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp -3599
transform 1 0 30912 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp -3599
transform 1 0 29808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp -3599
transform 1 0 28980 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp -3599
transform 1 0 27140 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp -3599
transform -1 0 27416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp -3599
transform -1 0 29164 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp -3599
transform -1 0 30084 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp -3599
transform -1 0 30268 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp -3599
transform -1 0 31464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp -3599
transform -1 0 31740 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636964856
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636964856
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636964856
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636964856
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636964856
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636964856
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636964856
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636964856
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -3599
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636964856
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636964856
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -3599
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636964856
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636964856
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -3599
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp -3599
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_177
timestamp -3599
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp -3599
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp -3599
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -3599
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -3599
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -3599
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp -3599
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1636964856
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp -3599
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1636964856
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1636964856
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp -3599
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_393
timestamp -3599
transform 1 0 37260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_397
timestamp -3599
transform 1 0 37628 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_410
timestamp -3599
transform 1 0 38824 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636964856
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636964856
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636964856
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636964856
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp -3599
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -3599
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636964856
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636964856
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636964856
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636964856
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp -3599
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -3599
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636964856
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636964856
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636964856
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636964856
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp -3599
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -3599
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636964856
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp -3599
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_185
timestamp -3599
transform 1 0 18124 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_190
timestamp -3599
transform 1 0 18584 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_194
timestamp -3599
transform 1 0 18952 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_199
timestamp -3599
transform 1 0 19412 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636964856
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp -3599
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp -3599
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636964856
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_237
timestamp -3599
transform 1 0 22908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_248
timestamp -3599
transform 1 0 23920 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_254
timestamp -3599
transform 1 0 24472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_259
timestamp -3599
transform 1 0 24932 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_275
timestamp -3599
transform 1 0 26404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp -3599
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_285
timestamp -3599
transform 1 0 27324 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_295
timestamp -3599
transform 1 0 28244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_301
timestamp -3599
transform 1 0 28796 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_307
timestamp -3599
transform 1 0 29348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_319
timestamp -3599
transform 1 0 30452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_323
timestamp -3599
transform 1 0 30820 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp -3599
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636964856
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636964856
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636964856
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636964856
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp -3599
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp -3599
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636964856
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_405
timestamp -3599
transform 1 0 38364 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636964856
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636964856
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636964856
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636964856
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636964856
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636964856
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636964856
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636964856
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636964856
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636964856
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp -3599
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp -3599
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636964856
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636964856
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636964856
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_177
timestamp -3599
transform 1 0 17388 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_185
timestamp -3599
transform 1 0 18124 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp -3599
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_202
timestamp 1636964856
transform 1 0 19688 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_214
timestamp -3599
transform 1 0 20792 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_222
timestamp -3599
transform 1 0 21528 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_227
timestamp -3599
transform 1 0 21988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_249
timestamp -3599
transform 1 0 24012 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_269
timestamp -3599
transform 1 0 25852 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_275
timestamp -3599
transform 1 0 26404 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_279
timestamp 1636964856
transform 1 0 26772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_291
timestamp 1636964856
transform 1 0 27876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_303
timestamp -3599
transform 1 0 28980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp -3599
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636964856
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636964856
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636964856
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636964856
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp -3599
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp -3599
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636964856
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636964856
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636964856
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_401
timestamp -3599
transform 1 0 37996 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_409
timestamp -3599
transform 1 0 38732 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636964856
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636964856
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636964856
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_42
timestamp 1636964856
transform 1 0 4968 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp -3599
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636964856
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636964856
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636964856
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636964856
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp -3599
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -3599
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636964856
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636964856
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636964856
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636964856
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp -3599
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -3599
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp -3599
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_176
timestamp -3599
transform 1 0 17296 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636964856
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_193
timestamp -3599
transform 1 0 18860 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_202
timestamp 1636964856
transform 1 0 19688 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_214
timestamp -3599
transform 1 0 20792 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_228
timestamp -3599
transform 1 0 22080 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_234
timestamp 1636964856
transform 1 0 22632 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_246
timestamp -3599
transform 1 0 23736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_250
timestamp -3599
transform 1 0 24104 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_256
timestamp 1636964856
transform 1 0 24656 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_268
timestamp 1636964856
transform 1 0 25760 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp -3599
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_288
timestamp -3599
transform 1 0 27600 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_297
timestamp -3599
transform 1 0 28428 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_308
timestamp -3599
transform 1 0 29440 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_317
timestamp -3599
transform 1 0 30268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_332
timestamp -3599
transform 1 0 31648 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636964856
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636964856
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636964856
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636964856
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp -3599
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp -3599
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636964856
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_405
timestamp -3599
transform 1 0 38364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_409
timestamp -3599
transform 1 0 38732 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636964856
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp -3599
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_19
timestamp -3599
transform 1 0 2852 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp -3599
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp -3599
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_33
timestamp -3599
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_37
timestamp -3599
transform 1 0 4508 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_42
timestamp 1636964856
transform 1 0 4968 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_54
timestamp 1636964856
transform 1 0 6072 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_66
timestamp 1636964856
transform 1 0 7176 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_78
timestamp -3599
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636964856
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636964856
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636964856
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636964856
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp -3599
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp -3599
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636964856
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636964856
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_165
timestamp -3599
transform 1 0 16284 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_171
timestamp 1636964856
transform 1 0 16836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_183
timestamp 1636964856
transform 1 0 17940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp -3599
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_197
timestamp -3599
transform 1 0 19228 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_205
timestamp -3599
transform 1 0 19964 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_211
timestamp 1636964856
transform 1 0 20516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_223
timestamp 1636964856
transform 1 0 21620 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_235
timestamp -3599
transform 1 0 22724 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_241
timestamp -3599
transform 1 0 23276 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_248
timestamp -3599
transform 1 0 23920 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_255
timestamp -3599
transform 1 0 24564 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_263
timestamp -3599
transform 1 0 25300 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_267
timestamp -3599
transform 1 0 25668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_275
timestamp -3599
transform 1 0 26404 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_279
timestamp -3599
transform 1 0 26772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_283
timestamp -3599
transform 1 0 27140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_289
timestamp -3599
transform 1 0 27692 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_297
timestamp -3599
transform 1 0 28428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_309
timestamp -3599
transform 1 0 29532 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_320
timestamp -3599
transform 1 0 30544 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_326
timestamp -3599
transform 1 0 31096 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_330
timestamp -3599
transform 1 0 31464 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_342
timestamp -3599
transform 1 0 32568 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_351
timestamp 1636964856
transform 1 0 33396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp -3599
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_365
timestamp -3599
transform 1 0 34684 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_373
timestamp -3599
transform 1 0 35420 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_379
timestamp 1636964856
transform 1 0 35972 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_391
timestamp 1636964856
transform 1 0 37076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_403
timestamp -3599
transform 1 0 38180 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_409
timestamp -3599
transform 1 0 38732 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636964856
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_15
timestamp -3599
transform 1 0 2484 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_26
timestamp 1636964856
transform 1 0 3496 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_38
timestamp 1636964856
transform 1 0 4600 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_50
timestamp -3599
transform 1 0 5704 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636964856
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636964856
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636964856
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636964856
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp -3599
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp -3599
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636964856
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636964856
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636964856
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_149
timestamp -3599
transform 1 0 14812 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp -3599
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_177
timestamp -3599
transform 1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_184
timestamp 1636964856
transform 1 0 18032 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_196
timestamp 1636964856
transform 1 0 19136 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_208
timestamp 1636964856
transform 1 0 20240 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp -3599
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_225
timestamp -3599
transform 1 0 21804 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_234
timestamp 1636964856
transform 1 0 22632 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_246
timestamp 1636964856
transform 1 0 23736 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_258
timestamp 1636964856
transform 1 0 24840 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_270
timestamp -3599
transform 1 0 25944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp -3599
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636964856
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636964856
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636964856
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1636964856
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp -3599
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp -3599
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636964856
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636964856
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636964856
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636964856
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_385
timestamp -3599
transform 1 0 36524 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636964856
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_405
timestamp -3599
transform 1 0 38364 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_409
timestamp -3599
transform 1 0 38732 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636964856
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636964856
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636964856
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636964856
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636964856
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_65
timestamp -3599
transform 1 0 7084 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_69
timestamp -3599
transform 1 0 7452 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_73
timestamp -3599
transform 1 0 7820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp -3599
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp -3599
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_89
timestamp 1636964856
transform 1 0 9292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_101
timestamp 1636964856
transform 1 0 10396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_113
timestamp 1636964856
transform 1 0 11500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_125
timestamp -3599
transform 1 0 12604 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_133
timestamp -3599
transform 1 0 13340 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp -3599
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_149
timestamp -3599
transform 1 0 14812 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636964856
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636964856
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636964856
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp -3599
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp -3599
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_197
timestamp -3599
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_205
timestamp 1636964856
transform 1 0 19964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_217
timestamp 1636964856
transform 1 0 21068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_229
timestamp 1636964856
transform 1 0 22172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_241
timestamp -3599
transform 1 0 23276 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp -3599
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636964856
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_265
timestamp -3599
transform 1 0 25484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_271
timestamp -3599
transform 1 0 26036 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_275
timestamp 1636964856
transform 1 0 26404 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_287
timestamp 1636964856
transform 1 0 27508 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_299
timestamp -3599
transform 1 0 28612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp -3599
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636964856
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1636964856
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1636964856
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1636964856
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp -3599
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp -3599
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636964856
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1636964856
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1636964856
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_401
timestamp -3599
transform 1 0 37996 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_409
timestamp -3599
transform 1 0 38732 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636964856
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636964856
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636964856
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636964856
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp -3599
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -3599
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636964856
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636964856
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_81
timestamp -3599
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_87
timestamp 1636964856
transform 1 0 9108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_99
timestamp 1636964856
transform 1 0 10212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp -3599
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636964856
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_125
timestamp -3599
transform 1 0 12604 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_133
timestamp -3599
transform 1 0 13340 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_145
timestamp 1636964856
transform 1 0 14444 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_157
timestamp -3599
transform 1 0 15548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp -3599
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636964856
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636964856
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1636964856
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1636964856
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp -3599
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp -3599
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636964856
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636964856
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636964856
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1636964856
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp -3599
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp -3599
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_281
timestamp -3599
transform 1 0 26956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_285
timestamp -3599
transform 1 0 27324 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_289
timestamp 1636964856
transform 1 0 27692 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_301
timestamp 1636964856
transform 1 0 28796 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_313
timestamp 1636964856
transform 1 0 29900 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_325
timestamp -3599
transform 1 0 31004 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_333
timestamp -3599
transform 1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1636964856
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1636964856
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1636964856
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1636964856
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp -3599
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp -3599
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1636964856
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_405
timestamp -3599
transform 1 0 38364 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_409
timestamp -3599
transform 1 0 38732 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636964856
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636964856
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -3599
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636964856
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636964856
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636964856
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636964856
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp -3599
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp -3599
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_95
timestamp -3599
transform 1 0 9844 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_99
timestamp -3599
transform 1 0 10212 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_107
timestamp -3599
transform 1 0 10948 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_111
timestamp -3599
transform 1 0 11316 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_118
timestamp 1636964856
transform 1 0 11960 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_130
timestamp -3599
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp -3599
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636964856
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636964856
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636964856
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_177
timestamp -3599
transform 1 0 17388 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_183
timestamp 1636964856
transform 1 0 17940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp -3599
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636964856
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636964856
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_221
timestamp -3599
transform 1 0 21436 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_232
timestamp 1636964856
transform 1 0 22448 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_244
timestamp -3599
transform 1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636964856
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1636964856
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1636964856
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1636964856
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp -3599
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp -3599
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1636964856
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1636964856
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1636964856
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1636964856
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp -3599
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp -3599
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1636964856
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1636964856
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1636964856
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_401
timestamp -3599
transform 1 0 37996 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_409
timestamp -3599
transform 1 0 38732 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636964856
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636964856
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636964856
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1636964856
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp -3599
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -3599
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636964856
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636964856
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1636964856
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1636964856
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp -3599
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp -3599
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636964856
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1636964856
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1636964856
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1636964856
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_161
timestamp -3599
transform 1 0 15916 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_180
timestamp -3599
transform 1 0 17664 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_184
timestamp -3599
transform 1 0 18032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_190
timestamp -3599
transform 1 0 18584 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_204
timestamp -3599
transform 1 0 19872 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_208
timestamp -3599
transform 1 0 20240 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp -3599
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp -3599
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_232
timestamp -3599
transform 1 0 22448 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_241
timestamp 1636964856
transform 1 0 23276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_253
timestamp 1636964856
transform 1 0 24380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_265
timestamp -3599
transform 1 0 25484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_269
timestamp -3599
transform 1 0 25852 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp -3599
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp -3599
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp -3599
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_286
timestamp -3599
transform 1 0 27416 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_302
timestamp 1636964856
transform 1 0 28888 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_314
timestamp 1636964856
transform 1 0 29992 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_326
timestamp -3599
transform 1 0 31096 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp -3599
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1636964856
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1636964856
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1636964856
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1636964856
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp -3599
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp -3599
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1636964856
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_405
timestamp -3599
transform 1 0 38364 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_409
timestamp -3599
transform 1 0 38732 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636964856
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636964856
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -3599
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636964856
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636964856
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1636964856
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1636964856
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp -3599
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp -3599
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636964856
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1636964856
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1636964856
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1636964856
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp -3599
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp -3599
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1636964856
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1636964856
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1636964856
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1636964856
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp -3599
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp -3599
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1636964856
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1636964856
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1636964856
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1636964856
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp -3599
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp -3599
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1636964856
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1636964856
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1636964856
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1636964856
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp -3599
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp -3599
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1636964856
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1636964856
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1636964856
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1636964856
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp -3599
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp -3599
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1636964856
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1636964856
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_389
timestamp -3599
transform 1 0 36892 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_397
timestamp -3599
transform 1 0 37628 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_6
timestamp 1636964856
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_18
timestamp -3599
transform 1 0 2760 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_26
timestamp -3599
transform 1 0 3496 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_29
timestamp 1636964856
transform 1 0 3772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_41
timestamp -3599
transform 1 0 4876 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_47
timestamp -3599
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp -3599
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_63
timestamp -3599
transform 1 0 6900 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_68
timestamp 1636964856
transform 1 0 7360 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_80
timestamp -3599
transform 1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_89
timestamp 1636964856
transform 1 0 9292 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_101
timestamp -3599
transform 1 0 10396 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_105
timestamp -3599
transform 1 0 10764 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp -3599
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1636964856
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_125
timestamp -3599
transform 1 0 12604 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_131
timestamp -3599
transform 1 0 13156 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_139
timestamp -3599
transform 1 0 13892 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_141
timestamp -3599
transform 1 0 14076 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_147
timestamp -3599
transform 1 0 14628 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_152
timestamp 1636964856
transform 1 0 15088 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp -3599
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_173
timestamp 1636964856
transform 1 0 17020 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_185
timestamp -3599
transform 1 0 18124 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_189
timestamp -3599
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_194
timestamp -3599
transform 1 0 18952 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_197
timestamp 1636964856
transform 1 0 19228 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_209
timestamp -3599
transform 1 0 20332 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_215
timestamp -3599
transform 1 0 20884 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp -3599
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_225
timestamp -3599
transform 1 0 21804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_231
timestamp -3599
transform 1 0 22356 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_236
timestamp 1636964856
transform 1 0 22816 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_248
timestamp -3599
transform 1 0 23920 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_257
timestamp 1636964856
transform 1 0 24748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_269
timestamp -3599
transform 1 0 25852 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_273
timestamp -3599
transform 1 0 26220 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp -3599
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1636964856
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_293
timestamp -3599
transform 1 0 28060 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_299
timestamp -3599
transform 1 0 28612 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_307
timestamp -3599
transform 1 0 29348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_309
timestamp -3599
transform 1 0 29532 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_315
timestamp -3599
transform 1 0 30084 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_320
timestamp 1636964856
transform 1 0 30544 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_332
timestamp -3599
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_341
timestamp 1636964856
transform 1 0 32476 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_353
timestamp -3599
transform 1 0 33580 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_357
timestamp -3599
transform 1 0 33948 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_362
timestamp -3599
transform 1 0 34408 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_365
timestamp 1636964856
transform 1 0 34684 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_377
timestamp -3599
transform 1 0 35788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_383
timestamp -3599
transform 1 0 36340 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_387
timestamp -3599
transform 1 0 36708 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_393
timestamp -3599
transform 1 0 37260 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_404
timestamp -3599
transform 1 0 38272 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output1
timestamp -3599
transform 1 0 38456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform 1 0 39192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform 1 0 38824 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform 1 0 39192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform 1 0 38824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform 1 0 39192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 38824 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform 1 0 39192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 38824 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -3599
transform 1 0 39192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -3599
transform 1 0 38824 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -3599
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp -3599
transform 1 0 39192 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp -3599
transform 1 0 39192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp -3599
transform 1 0 38824 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp -3599
transform 1 0 39192 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp -3599
transform 1 0 39192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -3599
transform 1 0 38824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp -3599
transform 1 0 38456 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp -3599
transform 1 0 38456 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp -3599
transform 1 0 38824 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp -3599
transform 1 0 38088 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp -3599
transform 1 0 37720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp -3599
transform 1 0 37536 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp -3599
transform 1 0 37720 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp -3599
transform 1 0 38456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp -3599
transform 1 0 39192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp -3599
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp -3599
transform 1 0 39192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp -3599
transform 1 0 38824 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp -3599
transform 1 0 39192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp -3599
transform 1 0 38824 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp -3599
transform -1 0 3496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp -3599
transform -1 0 22816 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp -3599
transform -1 0 24748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp -3599
transform 1 0 26312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp -3599
transform 1 0 28244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp -3599
transform 1 0 30176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp -3599
transform 1 0 32108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp -3599
transform 1 0 34040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp -3599
transform 1 0 35972 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp -3599
transform 1 0 37904 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp -3599
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp -3599
transform -1 0 5428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp -3599
transform -1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp -3599
transform -1 0 9292 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp -3599
transform -1 0 11224 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp -3599
transform -1 0 13156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp -3599
transform -1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp -3599
transform -1 0 17020 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp -3599
transform -1 0 18952 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp -3599
transform -1 0 20884 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp -3599
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp -3599
transform 1 0 18216 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp -3599
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp -3599
transform 1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp -3599
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp -3599
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp -3599
transform 1 0 19596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp -3599
transform 1 0 19412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp -3599
transform 1 0 19780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp -3599
transform 1 0 20148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp -3599
transform 1 0 20516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp -3599
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp -3599
transform 1 0 21252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp -3599
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp -3599
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp -3599
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp -3599
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp -3599
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp -3599
transform 1 0 23644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp -3599
transform 1 0 23184 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp -3599
transform 1 0 23552 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp -3599
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp -3599
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp -3599
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform 1 0 27692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform 1 0 25116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform 1 0 24564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform 1 0 26220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform 1 0 25668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform 1 0 26036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform 1 0 27876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform 1 0 31372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform 1 0 30912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform 1 0 31280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform 1 0 32476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform 1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform 1 0 28796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform -1 0 28796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform -1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform -1 0 29348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform -1 0 30268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform -1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform -1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform -1 0 30452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform -1 0 31372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output105
timestamp -3599
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 39836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 39836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 39836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 39836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 39836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 39836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 39836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 39836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 39836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 39836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_38
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -3599
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_45
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_48
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_49
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_50
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -3599
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_52
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_53
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_54
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_55
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_56
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_57
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_58
timestamp -3599
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_59
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_60
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_61
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_62
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_63
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_65
timestamp -3599
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_66
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_67
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_68
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_69
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_70
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_71
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp -3599
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_73
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_74
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_75
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_76
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp -3599
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_83
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_84
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_85
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp -3599
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_87
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_88
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_92
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_93
timestamp -3599
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_95
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_96
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_97
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_98
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_99
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_100
timestamp -3599
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_101
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_102
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_103
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_104
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_105
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp -3599
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_108
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_109
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_110
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_111
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_112
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_113
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_114
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_115
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_116
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_117
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_118
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_119
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp -3599
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_121
timestamp -3599
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 17590 0 17646 56 0 FreeSans 224 0 0 0 Ci
port 0 nsew signal input
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[0]
port 1 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[10]
port 2 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[11]
port 3 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[12]
port 4 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[13]
port 5 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[14]
port 6 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[15]
port 7 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[16]
port 8 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[17]
port 9 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[18]
port 10 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[19]
port 11 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[1]
port 12 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[20]
port 13 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[21]
port 14 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[22]
port 15 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[23]
port 16 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[24]
port 17 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[25]
port 18 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[26]
port 19 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[27]
port 20 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[28]
port 21 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[29]
port 22 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[2]
port 23 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[30]
port 24 nsew signal input
flabel metal3 s 0 9800 120 9920 0 FreeSans 480 0 0 0 FrameData[31]
port 25 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[3]
port 26 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[4]
port 27 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[5]
port 28 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[6]
port 29 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[7]
port 30 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[8]
port 31 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[9]
port 32 nsew signal input
flabel metal3 s 40880 1368 41000 1488 0 FreeSans 480 0 0 0 FrameData_O[0]
port 33 nsew signal output
flabel metal3 s 40880 4088 41000 4208 0 FreeSans 480 0 0 0 FrameData_O[10]
port 34 nsew signal output
flabel metal3 s 40880 4360 41000 4480 0 FreeSans 480 0 0 0 FrameData_O[11]
port 35 nsew signal output
flabel metal3 s 40880 4632 41000 4752 0 FreeSans 480 0 0 0 FrameData_O[12]
port 36 nsew signal output
flabel metal3 s 40880 4904 41000 5024 0 FreeSans 480 0 0 0 FrameData_O[13]
port 37 nsew signal output
flabel metal3 s 40880 5176 41000 5296 0 FreeSans 480 0 0 0 FrameData_O[14]
port 38 nsew signal output
flabel metal3 s 40880 5448 41000 5568 0 FreeSans 480 0 0 0 FrameData_O[15]
port 39 nsew signal output
flabel metal3 s 40880 5720 41000 5840 0 FreeSans 480 0 0 0 FrameData_O[16]
port 40 nsew signal output
flabel metal3 s 40880 5992 41000 6112 0 FreeSans 480 0 0 0 FrameData_O[17]
port 41 nsew signal output
flabel metal3 s 40880 6264 41000 6384 0 FreeSans 480 0 0 0 FrameData_O[18]
port 42 nsew signal output
flabel metal3 s 40880 6536 41000 6656 0 FreeSans 480 0 0 0 FrameData_O[19]
port 43 nsew signal output
flabel metal3 s 40880 1640 41000 1760 0 FreeSans 480 0 0 0 FrameData_O[1]
port 44 nsew signal output
flabel metal3 s 40880 6808 41000 6928 0 FreeSans 480 0 0 0 FrameData_O[20]
port 45 nsew signal output
flabel metal3 s 40880 7080 41000 7200 0 FreeSans 480 0 0 0 FrameData_O[21]
port 46 nsew signal output
flabel metal3 s 40880 7352 41000 7472 0 FreeSans 480 0 0 0 FrameData_O[22]
port 47 nsew signal output
flabel metal3 s 40880 7624 41000 7744 0 FreeSans 480 0 0 0 FrameData_O[23]
port 48 nsew signal output
flabel metal3 s 40880 7896 41000 8016 0 FreeSans 480 0 0 0 FrameData_O[24]
port 49 nsew signal output
flabel metal3 s 40880 8168 41000 8288 0 FreeSans 480 0 0 0 FrameData_O[25]
port 50 nsew signal output
flabel metal3 s 40880 8440 41000 8560 0 FreeSans 480 0 0 0 FrameData_O[26]
port 51 nsew signal output
flabel metal3 s 40880 8712 41000 8832 0 FreeSans 480 0 0 0 FrameData_O[27]
port 52 nsew signal output
flabel metal3 s 40880 8984 41000 9104 0 FreeSans 480 0 0 0 FrameData_O[28]
port 53 nsew signal output
flabel metal3 s 40880 9256 41000 9376 0 FreeSans 480 0 0 0 FrameData_O[29]
port 54 nsew signal output
flabel metal3 s 40880 1912 41000 2032 0 FreeSans 480 0 0 0 FrameData_O[2]
port 55 nsew signal output
flabel metal3 s 40880 9528 41000 9648 0 FreeSans 480 0 0 0 FrameData_O[30]
port 56 nsew signal output
flabel metal3 s 40880 9800 41000 9920 0 FreeSans 480 0 0 0 FrameData_O[31]
port 57 nsew signal output
flabel metal3 s 40880 2184 41000 2304 0 FreeSans 480 0 0 0 FrameData_O[3]
port 58 nsew signal output
flabel metal3 s 40880 2456 41000 2576 0 FreeSans 480 0 0 0 FrameData_O[4]
port 59 nsew signal output
flabel metal3 s 40880 2728 41000 2848 0 FreeSans 480 0 0 0 FrameData_O[5]
port 60 nsew signal output
flabel metal3 s 40880 3000 41000 3120 0 FreeSans 480 0 0 0 FrameData_O[6]
port 61 nsew signal output
flabel metal3 s 40880 3272 41000 3392 0 FreeSans 480 0 0 0 FrameData_O[7]
port 62 nsew signal output
flabel metal3 s 40880 3544 41000 3664 0 FreeSans 480 0 0 0 FrameData_O[8]
port 63 nsew signal output
flabel metal3 s 40880 3816 41000 3936 0 FreeSans 480 0 0 0 FrameData_O[9]
port 64 nsew signal output
flabel metal2 s 32494 0 32550 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 65 nsew signal input
flabel metal2 s 35254 0 35310 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 66 nsew signal input
flabel metal2 s 35530 0 35586 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 67 nsew signal input
flabel metal2 s 35806 0 35862 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 68 nsew signal input
flabel metal2 s 36082 0 36138 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 69 nsew signal input
flabel metal2 s 36358 0 36414 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 70 nsew signal input
flabel metal2 s 36634 0 36690 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 71 nsew signal input
flabel metal2 s 36910 0 36966 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 72 nsew signal input
flabel metal2 s 37186 0 37242 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 73 nsew signal input
flabel metal2 s 37462 0 37518 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 74 nsew signal input
flabel metal2 s 37738 0 37794 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 75 nsew signal input
flabel metal2 s 32770 0 32826 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 76 nsew signal input
flabel metal2 s 33046 0 33102 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 77 nsew signal input
flabel metal2 s 33322 0 33378 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 78 nsew signal input
flabel metal2 s 33598 0 33654 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 79 nsew signal input
flabel metal2 s 33874 0 33930 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 80 nsew signal input
flabel metal2 s 34150 0 34206 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 81 nsew signal input
flabel metal2 s 34426 0 34482 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 82 nsew signal input
flabel metal2 s 34702 0 34758 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 83 nsew signal input
flabel metal2 s 34978 0 35034 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 84 nsew signal input
flabel metal2 s 3054 11194 3110 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 85 nsew signal output
flabel metal2 s 22374 11194 22430 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 86 nsew signal output
flabel metal2 s 24306 11194 24362 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 87 nsew signal output
flabel metal2 s 26238 11194 26294 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 88 nsew signal output
flabel metal2 s 28170 11194 28226 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 89 nsew signal output
flabel metal2 s 30102 11194 30158 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 90 nsew signal output
flabel metal2 s 32034 11194 32090 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 91 nsew signal output
flabel metal2 s 33966 11194 34022 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 92 nsew signal output
flabel metal2 s 35898 11194 35954 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 93 nsew signal output
flabel metal2 s 37830 11194 37886 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 94 nsew signal output
flabel metal2 s 39762 11194 39818 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 95 nsew signal output
flabel metal2 s 4986 11194 5042 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 96 nsew signal output
flabel metal2 s 6918 11194 6974 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 97 nsew signal output
flabel metal2 s 8850 11194 8906 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 98 nsew signal output
flabel metal2 s 10782 11194 10838 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 99 nsew signal output
flabel metal2 s 12714 11194 12770 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 100 nsew signal output
flabel metal2 s 14646 11194 14702 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 101 nsew signal output
flabel metal2 s 16578 11194 16634 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 102 nsew signal output
flabel metal2 s 18510 11194 18566 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 103 nsew signal output
flabel metal2 s 20442 11194 20498 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 104 nsew signal output
flabel metal2 s 3238 0 3294 56 0 FreeSans 224 0 0 0 N1END[0]
port 105 nsew signal input
flabel metal2 s 3514 0 3570 56 0 FreeSans 224 0 0 0 N1END[1]
port 106 nsew signal input
flabel metal2 s 3790 0 3846 56 0 FreeSans 224 0 0 0 N1END[2]
port 107 nsew signal input
flabel metal2 s 4066 0 4122 56 0 FreeSans 224 0 0 0 N1END[3]
port 108 nsew signal input
flabel metal2 s 6550 0 6606 56 0 FreeSans 224 0 0 0 N2END[0]
port 109 nsew signal input
flabel metal2 s 6826 0 6882 56 0 FreeSans 224 0 0 0 N2END[1]
port 110 nsew signal input
flabel metal2 s 7102 0 7158 56 0 FreeSans 224 0 0 0 N2END[2]
port 111 nsew signal input
flabel metal2 s 7378 0 7434 56 0 FreeSans 224 0 0 0 N2END[3]
port 112 nsew signal input
flabel metal2 s 7654 0 7710 56 0 FreeSans 224 0 0 0 N2END[4]
port 113 nsew signal input
flabel metal2 s 7930 0 7986 56 0 FreeSans 224 0 0 0 N2END[5]
port 114 nsew signal input
flabel metal2 s 8206 0 8262 56 0 FreeSans 224 0 0 0 N2END[6]
port 115 nsew signal input
flabel metal2 s 8482 0 8538 56 0 FreeSans 224 0 0 0 N2END[7]
port 116 nsew signal input
flabel metal2 s 4342 0 4398 56 0 FreeSans 224 0 0 0 N2MID[0]
port 117 nsew signal input
flabel metal2 s 4618 0 4674 56 0 FreeSans 224 0 0 0 N2MID[1]
port 118 nsew signal input
flabel metal2 s 4894 0 4950 56 0 FreeSans 224 0 0 0 N2MID[2]
port 119 nsew signal input
flabel metal2 s 5170 0 5226 56 0 FreeSans 224 0 0 0 N2MID[3]
port 120 nsew signal input
flabel metal2 s 5446 0 5502 56 0 FreeSans 224 0 0 0 N2MID[4]
port 121 nsew signal input
flabel metal2 s 5722 0 5778 56 0 FreeSans 224 0 0 0 N2MID[5]
port 122 nsew signal input
flabel metal2 s 5998 0 6054 56 0 FreeSans 224 0 0 0 N2MID[6]
port 123 nsew signal input
flabel metal2 s 6274 0 6330 56 0 FreeSans 224 0 0 0 N2MID[7]
port 124 nsew signal input
flabel metal2 s 8758 0 8814 56 0 FreeSans 224 0 0 0 N4END[0]
port 125 nsew signal input
flabel metal2 s 11518 0 11574 56 0 FreeSans 224 0 0 0 N4END[10]
port 126 nsew signal input
flabel metal2 s 11794 0 11850 56 0 FreeSans 224 0 0 0 N4END[11]
port 127 nsew signal input
flabel metal2 s 12070 0 12126 56 0 FreeSans 224 0 0 0 N4END[12]
port 128 nsew signal input
flabel metal2 s 12346 0 12402 56 0 FreeSans 224 0 0 0 N4END[13]
port 129 nsew signal input
flabel metal2 s 12622 0 12678 56 0 FreeSans 224 0 0 0 N4END[14]
port 130 nsew signal input
flabel metal2 s 12898 0 12954 56 0 FreeSans 224 0 0 0 N4END[15]
port 131 nsew signal input
flabel metal2 s 9034 0 9090 56 0 FreeSans 224 0 0 0 N4END[1]
port 132 nsew signal input
flabel metal2 s 9310 0 9366 56 0 FreeSans 224 0 0 0 N4END[2]
port 133 nsew signal input
flabel metal2 s 9586 0 9642 56 0 FreeSans 224 0 0 0 N4END[3]
port 134 nsew signal input
flabel metal2 s 9862 0 9918 56 0 FreeSans 224 0 0 0 N4END[4]
port 135 nsew signal input
flabel metal2 s 10138 0 10194 56 0 FreeSans 224 0 0 0 N4END[5]
port 136 nsew signal input
flabel metal2 s 10414 0 10470 56 0 FreeSans 224 0 0 0 N4END[6]
port 137 nsew signal input
flabel metal2 s 10690 0 10746 56 0 FreeSans 224 0 0 0 N4END[7]
port 138 nsew signal input
flabel metal2 s 10966 0 11022 56 0 FreeSans 224 0 0 0 N4END[8]
port 139 nsew signal input
flabel metal2 s 11242 0 11298 56 0 FreeSans 224 0 0 0 N4END[9]
port 140 nsew signal input
flabel metal2 s 13174 0 13230 56 0 FreeSans 224 0 0 0 NN4END[0]
port 141 nsew signal input
flabel metal2 s 15934 0 15990 56 0 FreeSans 224 0 0 0 NN4END[10]
port 142 nsew signal input
flabel metal2 s 16210 0 16266 56 0 FreeSans 224 0 0 0 NN4END[11]
port 143 nsew signal input
flabel metal2 s 16486 0 16542 56 0 FreeSans 224 0 0 0 NN4END[12]
port 144 nsew signal input
flabel metal2 s 16762 0 16818 56 0 FreeSans 224 0 0 0 NN4END[13]
port 145 nsew signal input
flabel metal2 s 17038 0 17094 56 0 FreeSans 224 0 0 0 NN4END[14]
port 146 nsew signal input
flabel metal2 s 17314 0 17370 56 0 FreeSans 224 0 0 0 NN4END[15]
port 147 nsew signal input
flabel metal2 s 13450 0 13506 56 0 FreeSans 224 0 0 0 NN4END[1]
port 148 nsew signal input
flabel metal2 s 13726 0 13782 56 0 FreeSans 224 0 0 0 NN4END[2]
port 149 nsew signal input
flabel metal2 s 14002 0 14058 56 0 FreeSans 224 0 0 0 NN4END[3]
port 150 nsew signal input
flabel metal2 s 14278 0 14334 56 0 FreeSans 224 0 0 0 NN4END[4]
port 151 nsew signal input
flabel metal2 s 14554 0 14610 56 0 FreeSans 224 0 0 0 NN4END[5]
port 152 nsew signal input
flabel metal2 s 14830 0 14886 56 0 FreeSans 224 0 0 0 NN4END[6]
port 153 nsew signal input
flabel metal2 s 15106 0 15162 56 0 FreeSans 224 0 0 0 NN4END[7]
port 154 nsew signal input
flabel metal2 s 15382 0 15438 56 0 FreeSans 224 0 0 0 NN4END[8]
port 155 nsew signal input
flabel metal2 s 15658 0 15714 56 0 FreeSans 224 0 0 0 NN4END[9]
port 156 nsew signal input
flabel metal2 s 17866 0 17922 56 0 FreeSans 224 0 0 0 S1BEG[0]
port 157 nsew signal output
flabel metal2 s 18142 0 18198 56 0 FreeSans 224 0 0 0 S1BEG[1]
port 158 nsew signal output
flabel metal2 s 18418 0 18474 56 0 FreeSans 224 0 0 0 S1BEG[2]
port 159 nsew signal output
flabel metal2 s 18694 0 18750 56 0 FreeSans 224 0 0 0 S1BEG[3]
port 160 nsew signal output
flabel metal2 s 18970 0 19026 56 0 FreeSans 224 0 0 0 S2BEG[0]
port 161 nsew signal output
flabel metal2 s 19246 0 19302 56 0 FreeSans 224 0 0 0 S2BEG[1]
port 162 nsew signal output
flabel metal2 s 19522 0 19578 56 0 FreeSans 224 0 0 0 S2BEG[2]
port 163 nsew signal output
flabel metal2 s 19798 0 19854 56 0 FreeSans 224 0 0 0 S2BEG[3]
port 164 nsew signal output
flabel metal2 s 20074 0 20130 56 0 FreeSans 224 0 0 0 S2BEG[4]
port 165 nsew signal output
flabel metal2 s 20350 0 20406 56 0 FreeSans 224 0 0 0 S2BEG[5]
port 166 nsew signal output
flabel metal2 s 20626 0 20682 56 0 FreeSans 224 0 0 0 S2BEG[6]
port 167 nsew signal output
flabel metal2 s 20902 0 20958 56 0 FreeSans 224 0 0 0 S2BEG[7]
port 168 nsew signal output
flabel metal2 s 21178 0 21234 56 0 FreeSans 224 0 0 0 S2BEGb[0]
port 169 nsew signal output
flabel metal2 s 21454 0 21510 56 0 FreeSans 224 0 0 0 S2BEGb[1]
port 170 nsew signal output
flabel metal2 s 21730 0 21786 56 0 FreeSans 224 0 0 0 S2BEGb[2]
port 171 nsew signal output
flabel metal2 s 22006 0 22062 56 0 FreeSans 224 0 0 0 S2BEGb[3]
port 172 nsew signal output
flabel metal2 s 22282 0 22338 56 0 FreeSans 224 0 0 0 S2BEGb[4]
port 173 nsew signal output
flabel metal2 s 22558 0 22614 56 0 FreeSans 224 0 0 0 S2BEGb[5]
port 174 nsew signal output
flabel metal2 s 22834 0 22890 56 0 FreeSans 224 0 0 0 S2BEGb[6]
port 175 nsew signal output
flabel metal2 s 23110 0 23166 56 0 FreeSans 224 0 0 0 S2BEGb[7]
port 176 nsew signal output
flabel metal2 s 23386 0 23442 56 0 FreeSans 224 0 0 0 S4BEG[0]
port 177 nsew signal output
flabel metal2 s 26146 0 26202 56 0 FreeSans 224 0 0 0 S4BEG[10]
port 178 nsew signal output
flabel metal2 s 26422 0 26478 56 0 FreeSans 224 0 0 0 S4BEG[11]
port 179 nsew signal output
flabel metal2 s 26698 0 26754 56 0 FreeSans 224 0 0 0 S4BEG[12]
port 180 nsew signal output
flabel metal2 s 26974 0 27030 56 0 FreeSans 224 0 0 0 S4BEG[13]
port 181 nsew signal output
flabel metal2 s 27250 0 27306 56 0 FreeSans 224 0 0 0 S4BEG[14]
port 182 nsew signal output
flabel metal2 s 27526 0 27582 56 0 FreeSans 224 0 0 0 S4BEG[15]
port 183 nsew signal output
flabel metal2 s 23662 0 23718 56 0 FreeSans 224 0 0 0 S4BEG[1]
port 184 nsew signal output
flabel metal2 s 23938 0 23994 56 0 FreeSans 224 0 0 0 S4BEG[2]
port 185 nsew signal output
flabel metal2 s 24214 0 24270 56 0 FreeSans 224 0 0 0 S4BEG[3]
port 186 nsew signal output
flabel metal2 s 24490 0 24546 56 0 FreeSans 224 0 0 0 S4BEG[4]
port 187 nsew signal output
flabel metal2 s 24766 0 24822 56 0 FreeSans 224 0 0 0 S4BEG[5]
port 188 nsew signal output
flabel metal2 s 25042 0 25098 56 0 FreeSans 224 0 0 0 S4BEG[6]
port 189 nsew signal output
flabel metal2 s 25318 0 25374 56 0 FreeSans 224 0 0 0 S4BEG[7]
port 190 nsew signal output
flabel metal2 s 25594 0 25650 56 0 FreeSans 224 0 0 0 S4BEG[8]
port 191 nsew signal output
flabel metal2 s 25870 0 25926 56 0 FreeSans 224 0 0 0 S4BEG[9]
port 192 nsew signal output
flabel metal2 s 27802 0 27858 56 0 FreeSans 224 0 0 0 SS4BEG[0]
port 193 nsew signal output
flabel metal2 s 30562 0 30618 56 0 FreeSans 224 0 0 0 SS4BEG[10]
port 194 nsew signal output
flabel metal2 s 30838 0 30894 56 0 FreeSans 224 0 0 0 SS4BEG[11]
port 195 nsew signal output
flabel metal2 s 31114 0 31170 56 0 FreeSans 224 0 0 0 SS4BEG[12]
port 196 nsew signal output
flabel metal2 s 31390 0 31446 56 0 FreeSans 224 0 0 0 SS4BEG[13]
port 197 nsew signal output
flabel metal2 s 31666 0 31722 56 0 FreeSans 224 0 0 0 SS4BEG[14]
port 198 nsew signal output
flabel metal2 s 31942 0 31998 56 0 FreeSans 224 0 0 0 SS4BEG[15]
port 199 nsew signal output
flabel metal2 s 28078 0 28134 56 0 FreeSans 224 0 0 0 SS4BEG[1]
port 200 nsew signal output
flabel metal2 s 28354 0 28410 56 0 FreeSans 224 0 0 0 SS4BEG[2]
port 201 nsew signal output
flabel metal2 s 28630 0 28686 56 0 FreeSans 224 0 0 0 SS4BEG[3]
port 202 nsew signal output
flabel metal2 s 28906 0 28962 56 0 FreeSans 224 0 0 0 SS4BEG[4]
port 203 nsew signal output
flabel metal2 s 29182 0 29238 56 0 FreeSans 224 0 0 0 SS4BEG[5]
port 204 nsew signal output
flabel metal2 s 29458 0 29514 56 0 FreeSans 224 0 0 0 SS4BEG[6]
port 205 nsew signal output
flabel metal2 s 29734 0 29790 56 0 FreeSans 224 0 0 0 SS4BEG[7]
port 206 nsew signal output
flabel metal2 s 30010 0 30066 56 0 FreeSans 224 0 0 0 SS4BEG[8]
port 207 nsew signal output
flabel metal2 s 30286 0 30342 56 0 FreeSans 224 0 0 0 SS4BEG[9]
port 208 nsew signal output
flabel metal2 s 32218 0 32274 56 0 FreeSans 224 0 0 0 UserCLK
port 209 nsew signal input
flabel metal2 s 1122 11194 1178 11250 0 FreeSans 224 0 0 0 UserCLKo
port 210 nsew signal output
flabel metal4 s 3004 0 3324 11250 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 3004 11190 3324 11250 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11250 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 9004 11190 9324 11250 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11250 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 15004 11190 15324 11250 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11250 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 21004 11190 21324 11250 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11250 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 27004 11190 27324 11250 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11250 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 33004 11190 33324 11250 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 39004 0 39324 11250 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 39004 0 39324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 39004 11190 39324 11250 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11250 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 1944 11190 2264 11250 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 7944 0 8264 11250 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 7944 11190 8264 11250 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 13944 0 14264 11250 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 13944 11190 14264 11250 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 19944 0 20264 11250 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 19944 11190 20264 11250 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 25944 0 26264 11250 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 25944 11190 26264 11250 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 31944 0 32264 11250 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 31944 11190 32264 11250 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 37944 0 38264 11250 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 37944 0 38264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 37944 11190 38264 11250 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
rlabel metal1 20470 8704 20470 8704 0 VGND
rlabel metal1 20470 8160 20470 8160 0 VPWR
rlabel metal3 2828 1428 2828 1428 0 FrameData[0]
rlabel metal2 24058 4369 24058 4369 0 FrameData[10]
rlabel metal2 2806 4760 2806 4760 0 FrameData[11]
rlabel via2 22862 4675 22862 4675 0 FrameData[12]
rlabel metal3 942 4964 942 4964 0 FrameData[13]
rlabel metal1 19228 3502 19228 3502 0 FrameData[14]
rlabel metal3 344 5508 344 5508 0 FrameData[15]
rlabel metal1 19964 4658 19964 4658 0 FrameData[16]
rlabel metal3 919 6052 919 6052 0 FrameData[17]
rlabel metal1 16836 5202 16836 5202 0 FrameData[18]
rlabel metal1 18492 5882 18492 5882 0 FrameData[19]
rlabel metal3 4852 1700 4852 1700 0 FrameData[1]
rlabel via2 17526 6851 17526 6851 0 FrameData[20]
rlabel metal3 919 7140 919 7140 0 FrameData[21]
rlabel metal3 712 7412 712 7412 0 FrameData[22]
rlabel metal1 15778 7378 15778 7378 0 FrameData[23]
rlabel metal2 20470 7616 20470 7616 0 FrameData[24]
rlabel metal3 942 8228 942 8228 0 FrameData[25]
rlabel metal2 22126 8007 22126 8007 0 FrameData[26]
rlabel metal2 18906 7786 18906 7786 0 FrameData[27]
rlabel metal2 18722 8279 18722 8279 0 FrameData[28]
rlabel metal1 15594 7514 15594 7514 0 FrameData[29]
rlabel metal2 15134 1649 15134 1649 0 FrameData[2]
rlabel metal2 17802 7548 17802 7548 0 FrameData[30]
rlabel metal2 22586 8687 22586 8687 0 FrameData[31]
rlabel metal3 1471 2244 1471 2244 0 FrameData[3]
rlabel metal3 4392 2516 4392 2516 0 FrameData[4]
rlabel metal3 919 2788 919 2788 0 FrameData[5]
rlabel metal2 24150 3213 24150 3213 0 FrameData[6]
rlabel metal3 1425 3332 1425 3332 0 FrameData[7]
rlabel metal2 24242 3757 24242 3757 0 FrameData[8]
rlabel metal3 919 3876 919 3876 0 FrameData[9]
rlabel metal3 39798 1428 39798 1428 0 FrameData_O[0]
rlabel metal3 40166 4148 40166 4148 0 FrameData_O[10]
rlabel metal3 40442 4420 40442 4420 0 FrameData_O[11]
rlabel metal3 40166 4692 40166 4692 0 FrameData_O[12]
rlabel metal3 39982 4964 39982 4964 0 FrameData_O[13]
rlabel metal3 40166 5236 40166 5236 0 FrameData_O[14]
rlabel metal3 40442 5508 40442 5508 0 FrameData_O[15]
rlabel metal3 40166 5780 40166 5780 0 FrameData_O[16]
rlabel metal3 39982 6052 39982 6052 0 FrameData_O[17]
rlabel metal3 40166 6324 40166 6324 0 FrameData_O[18]
rlabel metal3 40442 6596 40442 6596 0 FrameData_O[19]
rlabel metal3 39614 1700 39614 1700 0 FrameData_O[1]
rlabel metal3 40166 6868 40166 6868 0 FrameData_O[20]
rlabel metal3 40166 7140 40166 7140 0 FrameData_O[21]
rlabel metal3 39936 7412 39936 7412 0 FrameData_O[22]
rlabel metal3 40166 7684 40166 7684 0 FrameData_O[23]
rlabel metal3 40166 7956 40166 7956 0 FrameData_O[24]
rlabel metal3 39982 8228 39982 8228 0 FrameData_O[25]
rlabel metal3 39798 8500 39798 8500 0 FrameData_O[26]
rlabel metal1 39100 8058 39100 8058 0 FrameData_O[27]
rlabel metal1 39330 7514 39330 7514 0 FrameData_O[28]
rlabel metal2 38318 8687 38318 8687 0 FrameData_O[29]
rlabel metal3 39430 1972 39430 1972 0 FrameData_O[2]
rlabel metal2 37766 9095 37766 9095 0 FrameData_O[30]
rlabel metal1 38180 7718 38180 7718 0 FrameData_O[31]
rlabel metal3 40672 2244 40672 2244 0 FrameData_O[3]
rlabel metal3 40166 2516 40166 2516 0 FrameData_O[4]
rlabel metal3 39982 2788 39982 2788 0 FrameData_O[5]
rlabel metal3 40166 3060 40166 3060 0 FrameData_O[6]
rlabel metal3 40442 3332 40442 3332 0 FrameData_O[7]
rlabel metal3 40166 3604 40166 3604 0 FrameData_O[8]
rlabel metal3 39982 3876 39982 3876 0 FrameData_O[9]
rlabel metal2 32522 650 32522 650 0 FrameStrobe[0]
rlabel metal2 35282 684 35282 684 0 FrameStrobe[10]
rlabel metal2 35558 3166 35558 3166 0 FrameStrobe[11]
rlabel metal2 35834 2860 35834 2860 0 FrameStrobe[12]
rlabel metal2 36110 242 36110 242 0 FrameStrobe[13]
rlabel metal2 36386 208 36386 208 0 FrameStrobe[14]
rlabel metal2 36662 1823 36662 1823 0 FrameStrobe[15]
rlabel via1 31878 4573 31878 4573 0 FrameStrobe[16]
rlabel metal2 37214 1211 37214 1211 0 FrameStrobe[17]
rlabel metal1 36616 4590 36616 4590 0 FrameStrobe[18]
rlabel metal1 37444 5202 37444 5202 0 FrameStrobe[19]
rlabel metal2 32798 871 32798 871 0 FrameStrobe[1]
rlabel metal2 33074 990 33074 990 0 FrameStrobe[2]
rlabel metal2 33350 55 33350 55 0 FrameStrobe[3]
rlabel metal2 33626 276 33626 276 0 FrameStrobe[4]
rlabel metal2 33902 3472 33902 3472 0 FrameStrobe[5]
rlabel metal2 34178 1551 34178 1551 0 FrameStrobe[6]
rlabel metal2 34454 1755 34454 1755 0 FrameStrobe[7]
rlabel metal2 34730 3710 34730 3710 0 FrameStrobe[8]
rlabel metal2 35006 667 35006 667 0 FrameStrobe[9]
rlabel metal1 3082 8602 3082 8602 0 FrameStrobe_O[0]
rlabel metal1 22494 8602 22494 8602 0 FrameStrobe_O[10]
rlabel metal1 24426 8602 24426 8602 0 FrameStrobe_O[11]
rlabel metal1 26404 8602 26404 8602 0 FrameStrobe_O[12]
rlabel metal1 28336 8602 28336 8602 0 FrameStrobe_O[13]
rlabel metal1 30268 8602 30268 8602 0 FrameStrobe_O[14]
rlabel metal1 32200 8602 32200 8602 0 FrameStrobe_O[15]
rlabel metal1 34132 8602 34132 8602 0 FrameStrobe_O[16]
rlabel metal1 36064 8602 36064 8602 0 FrameStrobe_O[17]
rlabel metal1 37996 8602 37996 8602 0 FrameStrobe_O[18]
rlabel metal2 37030 8772 37030 8772 0 FrameStrobe_O[19]
rlabel metal1 5106 8602 5106 8602 0 FrameStrobe_O[1]
rlabel metal1 7038 8602 7038 8602 0 FrameStrobe_O[2]
rlabel metal1 8970 8602 8970 8602 0 FrameStrobe_O[3]
rlabel metal1 10902 8602 10902 8602 0 FrameStrobe_O[4]
rlabel metal1 12834 8602 12834 8602 0 FrameStrobe_O[5]
rlabel metal1 14766 8602 14766 8602 0 FrameStrobe_O[6]
rlabel metal1 16698 8602 16698 8602 0 FrameStrobe_O[7]
rlabel metal1 18630 8602 18630 8602 0 FrameStrobe_O[8]
rlabel metal1 20562 8602 20562 8602 0 FrameStrobe_O[9]
rlabel metal2 3266 55 3266 55 0 N1END[0]
rlabel metal1 3404 5202 3404 5202 0 N1END[1]
rlabel metal1 2714 5134 2714 5134 0 N1END[2]
rlabel metal1 3542 5134 3542 5134 0 N1END[3]
rlabel metal1 7774 6426 7774 6426 0 N2END[0]
rlabel metal1 8878 5542 8878 5542 0 N2END[1]
rlabel metal1 8832 5746 8832 5746 0 N2END[2]
rlabel metal1 8694 6222 8694 6222 0 N2END[3]
rlabel metal1 8418 6086 8418 6086 0 N2END[4]
rlabel metal2 7958 1279 7958 1279 0 N2END[5]
rlabel metal2 8234 1330 8234 1330 0 N2END[6]
rlabel metal1 8694 6290 8694 6290 0 N2END[7]
rlabel metal2 4370 55 4370 55 0 N2MID[0]
rlabel metal1 6900 6630 6900 6630 0 N2MID[1]
rlabel metal2 4922 1401 4922 1401 0 N2MID[2]
rlabel metal1 6394 5678 6394 5678 0 N2MID[3]
rlabel metal1 5750 5202 5750 5202 0 N2MID[4]
rlabel metal1 5244 4590 5244 4590 0 N2MID[5]
rlabel metal2 6026 650 6026 650 0 N2MID[6]
rlabel metal1 5520 4114 5520 4114 0 N2MID[7]
rlabel metal2 8786 803 8786 803 0 N4END[0]
rlabel metal1 14214 6324 14214 6324 0 N4END[10]
rlabel metal2 11822 3166 11822 3166 0 N4END[11]
rlabel metal1 13938 6256 13938 6256 0 N4END[12]
rlabel metal2 12558 4947 12558 4947 0 N4END[13]
rlabel metal1 13662 5610 13662 5610 0 N4END[14]
rlabel metal1 14306 5134 14306 5134 0 N4END[15]
rlabel metal2 9062 55 9062 55 0 N4END[1]
rlabel metal2 9338 1007 9338 1007 0 N4END[2]
rlabel metal2 9614 803 9614 803 0 N4END[3]
rlabel metal2 9890 1143 9890 1143 0 N4END[4]
rlabel metal1 15962 5236 15962 5236 0 N4END[5]
rlabel metal2 10442 2622 10442 2622 0 N4END[6]
rlabel via2 14582 5661 14582 5661 0 N4END[7]
rlabel metal2 10994 1330 10994 1330 0 N4END[8]
rlabel metal2 11270 2860 11270 2860 0 N4END[9]
rlabel metal2 13202 939 13202 939 0 NN4END[0]
rlabel metal2 15962 174 15962 174 0 NN4END[10]
rlabel metal2 16238 55 16238 55 0 NN4END[11]
rlabel metal2 16514 140 16514 140 0 NN4END[12]
rlabel metal2 16790 1211 16790 1211 0 NN4END[13]
rlabel metal3 18768 3196 18768 3196 0 NN4END[14]
rlabel metal3 18860 3332 18860 3332 0 NN4END[15]
rlabel metal2 13478 208 13478 208 0 NN4END[1]
rlabel metal2 13754 191 13754 191 0 NN4END[2]
rlabel metal2 14030 276 14030 276 0 NN4END[3]
rlabel metal2 14306 242 14306 242 0 NN4END[4]
rlabel metal2 14582 123 14582 123 0 NN4END[5]
rlabel via2 14858 55 14858 55 0 NN4END[6]
rlabel metal2 15134 106 15134 106 0 NN4END[7]
rlabel metal2 15410 854 15410 854 0 NN4END[8]
rlabel metal2 15686 106 15686 106 0 NN4END[9]
rlabel metal2 17894 1160 17894 1160 0 S1BEG[0]
rlabel metal1 18308 2822 18308 2822 0 S1BEG[1]
rlabel metal2 18446 1160 18446 1160 0 S1BEG[2]
rlabel metal2 18722 1160 18722 1160 0 S1BEG[3]
rlabel metal1 19136 2822 19136 2822 0 S2BEG[0]
rlabel metal2 19274 1160 19274 1160 0 S2BEG[1]
rlabel metal1 19688 2822 19688 2822 0 S2BEG[2]
rlabel metal2 19826 1160 19826 1160 0 S2BEG[3]
rlabel metal2 20102 1160 20102 1160 0 S2BEG[4]
rlabel metal2 20378 1160 20378 1160 0 S2BEG[5]
rlabel metal2 20654 1160 20654 1160 0 S2BEG[6]
rlabel metal2 20930 1160 20930 1160 0 S2BEG[7]
rlabel metal2 21206 55 21206 55 0 S2BEGb[0]
rlabel metal2 21482 1160 21482 1160 0 S2BEGb[1]
rlabel metal2 21758 1296 21758 1296 0 S2BEGb[2]
rlabel metal2 22034 1330 22034 1330 0 S2BEGb[3]
rlabel metal2 22310 55 22310 55 0 S2BEGb[4]
rlabel metal2 22586 1330 22586 1330 0 S2BEGb[5]
rlabel metal2 22862 1160 22862 1160 0 S2BEGb[6]
rlabel metal1 23276 2822 23276 2822 0 S2BEGb[7]
rlabel metal1 23598 3162 23598 3162 0 S4BEG[0]
rlabel metal2 26174 1262 26174 1262 0 S4BEG[10]
rlabel metal2 26450 599 26450 599 0 S4BEG[11]
rlabel metal1 26956 2822 26956 2822 0 S4BEG[12]
rlabel metal2 27002 599 27002 599 0 S4BEG[13]
rlabel metal2 27278 956 27278 956 0 S4BEG[14]
rlabel metal2 27554 854 27554 854 0 S4BEG[15]
rlabel metal2 23690 1296 23690 1296 0 S4BEG[1]
rlabel metal2 23966 1160 23966 1160 0 S4BEG[2]
rlabel metal2 24242 1330 24242 1330 0 S4BEG[3]
rlabel metal1 24656 2822 24656 2822 0 S4BEG[4]
rlabel metal2 24794 1296 24794 1296 0 S4BEG[5]
rlabel metal2 25070 786 25070 786 0 S4BEG[6]
rlabel metal2 25346 956 25346 956 0 S4BEG[7]
rlabel metal1 25760 2822 25760 2822 0 S4BEG[8]
rlabel metal2 25898 735 25898 735 0 S4BEG[9]
rlabel metal1 27968 2822 27968 2822 0 SS4BEG[0]
rlabel metal2 30590 1160 30590 1160 0 SS4BEG[10]
rlabel metal1 31004 2822 31004 2822 0 SS4BEG[11]
rlabel metal2 31188 2788 31188 2788 0 SS4BEG[12]
rlabel metal2 31418 667 31418 667 0 SS4BEG[13]
rlabel metal2 31694 1160 31694 1160 0 SS4BEG[14]
rlabel metal2 31970 1194 31970 1194 0 SS4BEG[15]
rlabel metal2 28106 1296 28106 1296 0 SS4BEG[1]
rlabel metal1 28474 2822 28474 2822 0 SS4BEG[2]
rlabel metal2 28658 395 28658 395 0 SS4BEG[3]
rlabel metal1 29026 2822 29026 2822 0 SS4BEG[4]
rlabel metal2 29210 1296 29210 1296 0 SS4BEG[5]
rlabel metal2 29486 1194 29486 1194 0 SS4BEG[6]
rlabel metal2 29762 1330 29762 1330 0 SS4BEG[7]
rlabel metal2 30038 735 30038 735 0 SS4BEG[8]
rlabel metal2 30314 1296 30314 1296 0 SS4BEG[9]
rlabel metal2 32246 1296 32246 1296 0 UserCLK
rlabel metal1 1288 8602 1288 8602 0 UserCLKo
rlabel metal2 38502 2244 38502 2244 0 net1
rlabel metal2 17986 5848 17986 5848 0 net10
rlabel metal1 30682 3706 30682 3706 0 net100
rlabel metal1 30636 2414 30636 2414 0 net101
rlabel metal1 31970 4454 31970 4454 0 net102
rlabel metal2 32430 3774 32430 3774 0 net103
rlabel metal2 31786 3468 31786 3468 0 net104
rlabel metal2 1610 7582 1610 7582 0 net105
rlabel metal1 20999 5814 20999 5814 0 net11
rlabel metal1 38134 2448 38134 2448 0 net12
rlabel metal2 17894 6817 17894 6817 0 net13
rlabel metal2 17158 7582 17158 7582 0 net14
rlabel metal1 38870 7922 38870 7922 0 net15
rlabel metal2 38042 7514 38042 7514 0 net16
rlabel metal2 20746 8398 20746 8398 0 net17
rlabel metal1 20286 7514 20286 7514 0 net18
rlabel metal1 23598 7174 23598 7174 0 net19
rlabel metal2 35926 4148 35926 4148 0 net2
rlabel metal2 19274 7786 19274 7786 0 net20
rlabel metal2 19826 7072 19826 7072 0 net21
rlabel metal2 38134 7582 38134 7582 0 net22
rlabel metal2 33442 2244 33442 2244 0 net23
rlabel metal2 17986 8194 17986 8194 0 net24
rlabel metal2 37766 7650 37766 7650 0 net25
rlabel metal1 38502 3094 38502 3094 0 net26
rlabel metal1 39008 2278 39008 2278 0 net27
rlabel metal2 38870 3332 38870 3332 0 net28
rlabel metal2 38962 3230 38962 3230 0 net29
rlabel metal1 38870 4556 38870 4556 0 net3
rlabel metal1 35305 3502 35305 3502 0 net30
rlabel metal2 39238 3740 39238 3740 0 net31
rlabel metal1 31694 4148 31694 4148 0 net32
rlabel metal2 20838 8364 20838 8364 0 net33
rlabel metal1 28566 7174 28566 7174 0 net34
rlabel metal1 26082 6426 26082 6426 0 net35
rlabel metal2 26358 7174 26358 7174 0 net36
rlabel metal2 25622 6426 25622 6426 0 net37
rlabel metal2 25806 6460 25806 6460 0 net38
rlabel metal2 32614 5916 32614 5916 0 net39
rlabel metal1 39238 4658 39238 4658 0 net4
rlabel metal1 34086 8432 34086 8432 0 net40
rlabel metal1 34684 4794 34684 4794 0 net41
rlabel metal1 36570 4454 36570 4454 0 net42
rlabel metal1 36892 5338 36892 5338 0 net43
rlabel metal2 5382 8636 5382 8636 0 net44
rlabel metal1 7314 8398 7314 8398 0 net45
rlabel metal2 19366 7650 19366 7650 0 net46
rlabel metal1 12420 8500 12420 8500 0 net47
rlabel metal2 13110 8738 13110 8738 0 net48
rlabel metal2 16882 8772 16882 8772 0 net49
rlabel metal1 38870 5236 38870 5236 0 net5
rlabel metal2 16974 8704 16974 8704 0 net50
rlabel metal2 18906 8806 18906 8806 0 net51
rlabel metal1 21459 8466 21459 8466 0 net52
rlabel metal1 17204 2414 17204 2414 0 net53
rlabel metal2 17986 3774 17986 3774 0 net54
rlabel metal1 17940 2414 17940 2414 0 net55
rlabel metal1 18446 2380 18446 2380 0 net56
rlabel metal1 19090 3060 19090 3060 0 net57
rlabel via1 18262 3485 18262 3485 0 net58
rlabel metal2 19642 3230 19642 3230 0 net59
rlabel metal2 19458 3417 19458 3417 0 net6
rlabel metal2 14858 6256 14858 6256 0 net60
rlabel metal1 19780 2414 19780 2414 0 net61
rlabel metal1 18722 2380 18722 2380 0 net62
rlabel metal1 19228 2550 19228 2550 0 net63
rlabel metal1 11937 1938 11937 1938 0 net64
rlabel metal1 21344 2414 21344 2414 0 net65
rlabel metal2 13662 5984 13662 5984 0 net66
rlabel metal1 22264 2414 22264 2414 0 net67
rlabel metal1 17250 1938 17250 1938 0 net68
rlabel metal1 10212 6630 10212 6630 0 net69
rlabel metal2 19642 4777 19642 4777 0 net7
rlabel metal1 17250 2584 17250 2584 0 net70
rlabel metal1 23644 2414 23644 2414 0 net71
rlabel metal2 12006 3485 12006 3485 0 net72
rlabel metal1 21666 5032 21666 5032 0 net73
rlabel metal1 16146 5304 16146 5304 0 net74
rlabel metal1 19274 4794 19274 4794 0 net75
rlabel metal1 19734 3468 19734 3468 0 net76
rlabel metal1 18515 3978 18515 3978 0 net77
rlabel metal2 18630 3264 18630 3264 0 net78
rlabel metal2 19366 3230 19366 3230 0 net79
rlabel metal2 20470 5032 20470 5032 0 net8
rlabel metal1 19090 5746 19090 5746 0 net80
rlabel metal1 15318 5814 15318 5814 0 net81
rlabel metal1 14214 6086 14214 6086 0 net82
rlabel metal2 20746 4896 20746 4896 0 net83
rlabel metal1 14674 6086 14674 6086 0 net84
rlabel metal3 14490 1700 14490 1700 0 net85
rlabel metal1 14168 5542 14168 5542 0 net86
rlabel metal1 20010 5576 20010 5576 0 net87
rlabel metal2 15594 4862 15594 4862 0 net88
rlabel metal2 27922 3468 27922 3468 0 net89
rlabel metal2 38686 5644 38686 5644 0 net9
rlabel metal1 31234 2618 31234 2618 0 net90
rlabel metal1 30912 3026 30912 3026 0 net91
rlabel metal2 31326 3910 31326 3910 0 net92
rlabel metal2 32154 2176 32154 2176 0 net93
rlabel metal2 32522 3774 32522 3774 0 net94
rlabel metal2 32890 2040 32890 2040 0 net95
rlabel metal1 28750 2414 28750 2414 0 net96
rlabel metal1 28980 3026 28980 3026 0 net97
rlabel metal1 29946 2414 29946 2414 0 net98
rlabel metal1 29716 3026 29716 3026 0 net99
<< properties >>
string FIXED_BBOX 0 0 41000 11250
<< end >>
