magic
tech ihp-sg13g2
magscale 1 2
timestamp 1743695212
<< metal1 >>
rect 1152 9848 38112 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 38112 9848
rect 1152 9784 38112 9808
rect 7323 9680 7365 9689
rect 7323 9640 7324 9680
rect 7364 9640 7365 9680
rect 7323 9631 7365 9640
rect 7707 9680 7749 9689
rect 7707 9640 7708 9680
rect 7748 9640 7749 9680
rect 7707 9631 7749 9640
rect 8091 9680 8133 9689
rect 8091 9640 8092 9680
rect 8132 9640 8133 9680
rect 8091 9631 8133 9640
rect 8475 9680 8517 9689
rect 8475 9640 8476 9680
rect 8516 9640 8517 9680
rect 8475 9631 8517 9640
rect 8859 9680 8901 9689
rect 8859 9640 8860 9680
rect 8900 9640 8901 9680
rect 8859 9631 8901 9640
rect 9243 9680 9285 9689
rect 9243 9640 9244 9680
rect 9284 9640 9285 9680
rect 9243 9631 9285 9640
rect 9627 9680 9669 9689
rect 9627 9640 9628 9680
rect 9668 9640 9669 9680
rect 9627 9631 9669 9640
rect 10011 9680 10053 9689
rect 10011 9640 10012 9680
rect 10052 9640 10053 9680
rect 10011 9631 10053 9640
rect 10395 9680 10437 9689
rect 10395 9640 10396 9680
rect 10436 9640 10437 9680
rect 10395 9631 10437 9640
rect 10779 9680 10821 9689
rect 10779 9640 10780 9680
rect 10820 9640 10821 9680
rect 10779 9631 10821 9640
rect 11163 9680 11205 9689
rect 11163 9640 11164 9680
rect 11204 9640 11205 9680
rect 11163 9631 11205 9640
rect 11547 9680 11589 9689
rect 11547 9640 11548 9680
rect 11588 9640 11589 9680
rect 11547 9631 11589 9640
rect 11931 9680 11973 9689
rect 11931 9640 11932 9680
rect 11972 9640 11973 9680
rect 11931 9631 11973 9640
rect 12315 9680 12357 9689
rect 12315 9640 12316 9680
rect 12356 9640 12357 9680
rect 12315 9631 12357 9640
rect 12699 9680 12741 9689
rect 12699 9640 12700 9680
rect 12740 9640 12741 9680
rect 12699 9631 12741 9640
rect 13083 9680 13125 9689
rect 13083 9640 13084 9680
rect 13124 9640 13125 9680
rect 13083 9631 13125 9640
rect 13467 9680 13509 9689
rect 13467 9640 13468 9680
rect 13508 9640 13509 9680
rect 13467 9631 13509 9640
rect 13851 9680 13893 9689
rect 13851 9640 13852 9680
rect 13892 9640 13893 9680
rect 13851 9631 13893 9640
rect 14235 9680 14277 9689
rect 14235 9640 14236 9680
rect 14276 9640 14277 9680
rect 14235 9631 14277 9640
rect 14619 9680 14661 9689
rect 14619 9640 14620 9680
rect 14660 9640 14661 9680
rect 14619 9631 14661 9640
rect 15003 9680 15045 9689
rect 15003 9640 15004 9680
rect 15044 9640 15045 9680
rect 15003 9631 15045 9640
rect 15387 9680 15429 9689
rect 15387 9640 15388 9680
rect 15428 9640 15429 9680
rect 15387 9631 15429 9640
rect 15771 9680 15813 9689
rect 15771 9640 15772 9680
rect 15812 9640 15813 9680
rect 15771 9631 15813 9640
rect 16539 9680 16581 9689
rect 16539 9640 16540 9680
rect 16580 9640 16581 9680
rect 16539 9631 16581 9640
rect 17019 9680 17061 9689
rect 17019 9640 17020 9680
rect 17060 9640 17061 9680
rect 17019 9631 17061 9640
rect 17403 9680 17445 9689
rect 17403 9640 17404 9680
rect 17444 9640 17445 9680
rect 17403 9631 17445 9640
rect 27579 9680 27621 9689
rect 27579 9640 27580 9680
rect 27620 9640 27621 9680
rect 27579 9631 27621 9640
rect 28347 9680 28389 9689
rect 28347 9640 28348 9680
rect 28388 9640 28389 9680
rect 28347 9631 28389 9640
rect 29115 9680 29157 9689
rect 29115 9640 29116 9680
rect 29156 9640 29157 9680
rect 29115 9631 29157 9640
rect 30651 9680 30693 9689
rect 30651 9640 30652 9680
rect 30692 9640 30693 9680
rect 30651 9631 30693 9640
rect 31035 9680 31077 9689
rect 31035 9640 31036 9680
rect 31076 9640 31077 9680
rect 31035 9631 31077 9640
rect 32187 9680 32229 9689
rect 32187 9640 32188 9680
rect 32228 9640 32229 9680
rect 32187 9631 32229 9640
rect 36123 9680 36165 9689
rect 36123 9640 36124 9680
rect 36164 9640 36165 9680
rect 36123 9631 36165 9640
rect 36507 9680 36549 9689
rect 36507 9640 36508 9680
rect 36548 9640 36549 9680
rect 36507 9631 36549 9640
rect 36891 9680 36933 9689
rect 36891 9640 36892 9680
rect 36932 9640 36933 9680
rect 36891 9631 36933 9640
rect 16635 9596 16677 9605
rect 16635 9556 16636 9596
rect 16676 9556 16677 9596
rect 16635 9547 16677 9556
rect 17787 9596 17829 9605
rect 17787 9556 17788 9596
rect 17828 9556 17829 9596
rect 17787 9547 17829 9556
rect 27963 9596 28005 9605
rect 27963 9556 27964 9596
rect 28004 9556 28005 9596
rect 27963 9547 28005 9556
rect 28731 9596 28773 9605
rect 28731 9556 28732 9596
rect 28772 9556 28773 9596
rect 28731 9547 28773 9556
rect 29883 9596 29925 9605
rect 29883 9556 29884 9596
rect 29924 9556 29925 9596
rect 29883 9547 29925 9556
rect 31803 9596 31845 9605
rect 31803 9556 31804 9596
rect 31844 9556 31845 9596
rect 31803 9547 31845 9556
rect 7083 9512 7125 9521
rect 7083 9472 7084 9512
rect 7124 9472 7125 9512
rect 7083 9463 7125 9472
rect 7467 9512 7509 9521
rect 7467 9472 7468 9512
rect 7508 9472 7509 9512
rect 7467 9463 7509 9472
rect 7851 9512 7893 9521
rect 7851 9472 7852 9512
rect 7892 9472 7893 9512
rect 7851 9463 7893 9472
rect 8235 9512 8277 9521
rect 8235 9472 8236 9512
rect 8276 9472 8277 9512
rect 8235 9463 8277 9472
rect 8619 9512 8661 9521
rect 8619 9472 8620 9512
rect 8660 9472 8661 9512
rect 8619 9463 8661 9472
rect 9003 9512 9045 9521
rect 9003 9472 9004 9512
rect 9044 9472 9045 9512
rect 9003 9463 9045 9472
rect 9387 9512 9429 9521
rect 9387 9472 9388 9512
rect 9428 9472 9429 9512
rect 9387 9463 9429 9472
rect 9771 9512 9813 9521
rect 9771 9472 9772 9512
rect 9812 9472 9813 9512
rect 9771 9463 9813 9472
rect 10155 9512 10197 9521
rect 10155 9472 10156 9512
rect 10196 9472 10197 9512
rect 10155 9463 10197 9472
rect 10539 9512 10581 9521
rect 10539 9472 10540 9512
rect 10580 9472 10581 9512
rect 10539 9463 10581 9472
rect 10923 9512 10965 9521
rect 10923 9472 10924 9512
rect 10964 9472 10965 9512
rect 10923 9463 10965 9472
rect 11307 9512 11349 9521
rect 11307 9472 11308 9512
rect 11348 9472 11349 9512
rect 11307 9463 11349 9472
rect 11691 9512 11733 9521
rect 11691 9472 11692 9512
rect 11732 9472 11733 9512
rect 11691 9463 11733 9472
rect 12075 9512 12117 9521
rect 12075 9472 12076 9512
rect 12116 9472 12117 9512
rect 12075 9463 12117 9472
rect 12459 9512 12501 9521
rect 12459 9472 12460 9512
rect 12500 9472 12501 9512
rect 12459 9463 12501 9472
rect 12843 9512 12885 9521
rect 12843 9472 12844 9512
rect 12884 9472 12885 9512
rect 12843 9463 12885 9472
rect 13227 9512 13269 9521
rect 13227 9472 13228 9512
rect 13268 9472 13269 9512
rect 13227 9463 13269 9472
rect 13611 9512 13653 9521
rect 13611 9472 13612 9512
rect 13652 9472 13653 9512
rect 13611 9463 13653 9472
rect 13995 9512 14037 9521
rect 13995 9472 13996 9512
rect 14036 9472 14037 9512
rect 13995 9463 14037 9472
rect 14379 9512 14421 9521
rect 14379 9472 14380 9512
rect 14420 9472 14421 9512
rect 14379 9463 14421 9472
rect 14763 9512 14805 9521
rect 14763 9472 14764 9512
rect 14804 9472 14805 9512
rect 14763 9463 14805 9472
rect 15147 9512 15189 9521
rect 15147 9472 15148 9512
rect 15188 9472 15189 9512
rect 15147 9463 15189 9472
rect 15531 9512 15573 9521
rect 15531 9472 15532 9512
rect 15572 9472 15573 9512
rect 15531 9463 15573 9472
rect 15915 9512 15957 9521
rect 15915 9472 15916 9512
rect 15956 9472 15957 9512
rect 15915 9463 15957 9472
rect 16155 9512 16197 9521
rect 16155 9472 16156 9512
rect 16196 9472 16197 9512
rect 16155 9463 16197 9472
rect 16299 9512 16341 9521
rect 16299 9472 16300 9512
rect 16340 9472 16341 9512
rect 16299 9463 16341 9472
rect 16875 9512 16917 9521
rect 16875 9472 16876 9512
rect 16916 9472 16917 9512
rect 16875 9463 16917 9472
rect 17259 9512 17301 9521
rect 17259 9472 17260 9512
rect 17300 9472 17301 9512
rect 17259 9463 17301 9472
rect 17643 9512 17685 9521
rect 17643 9472 17644 9512
rect 17684 9472 17685 9512
rect 17643 9463 17685 9472
rect 18027 9512 18069 9521
rect 18027 9472 18028 9512
rect 18068 9472 18069 9512
rect 18027 9463 18069 9472
rect 27819 9512 27861 9521
rect 27819 9472 27820 9512
rect 27860 9472 27861 9512
rect 27819 9463 27861 9472
rect 28203 9512 28245 9521
rect 28203 9472 28204 9512
rect 28244 9472 28245 9512
rect 28203 9463 28245 9472
rect 28587 9512 28629 9521
rect 28587 9472 28588 9512
rect 28628 9472 28629 9512
rect 28587 9463 28629 9472
rect 28971 9512 29013 9521
rect 28971 9472 28972 9512
rect 29012 9472 29013 9512
rect 28971 9463 29013 9472
rect 29355 9512 29397 9521
rect 29355 9472 29356 9512
rect 29396 9472 29397 9512
rect 29355 9463 29397 9472
rect 29739 9512 29781 9521
rect 29739 9472 29740 9512
rect 29780 9472 29781 9512
rect 29739 9463 29781 9472
rect 30123 9512 30165 9521
rect 30123 9472 30124 9512
rect 30164 9472 30165 9512
rect 30123 9463 30165 9472
rect 30507 9512 30549 9521
rect 30507 9472 30508 9512
rect 30548 9472 30549 9512
rect 30507 9463 30549 9472
rect 30891 9512 30933 9521
rect 30891 9472 30892 9512
rect 30932 9472 30933 9512
rect 30891 9463 30933 9472
rect 31275 9512 31317 9521
rect 31275 9472 31276 9512
rect 31316 9472 31317 9512
rect 31275 9463 31317 9472
rect 31659 9512 31701 9521
rect 31659 9472 31660 9512
rect 31700 9472 31701 9512
rect 31659 9463 31701 9472
rect 32043 9512 32085 9521
rect 32043 9472 32044 9512
rect 32084 9472 32085 9512
rect 32043 9463 32085 9472
rect 32427 9512 32469 9521
rect 32427 9472 32428 9512
rect 32468 9472 32469 9512
rect 32427 9463 32469 9472
rect 35883 9512 35925 9521
rect 35883 9472 35884 9512
rect 35924 9472 35925 9512
rect 35883 9463 35925 9472
rect 36267 9512 36309 9521
rect 36267 9472 36268 9512
rect 36308 9472 36309 9512
rect 36267 9463 36309 9472
rect 36651 9512 36693 9521
rect 36651 9472 36652 9512
rect 36692 9472 36693 9512
rect 36651 9463 36693 9472
rect 37035 9512 37077 9521
rect 37035 9472 37036 9512
rect 37076 9472 37077 9512
rect 37035 9463 37077 9472
rect 37419 9512 37461 9521
rect 37419 9472 37420 9512
rect 37460 9472 37461 9512
rect 37419 9463 37461 9472
rect 37803 9512 37845 9521
rect 37803 9472 37804 9512
rect 37844 9472 37845 9512
rect 37803 9463 37845 9472
rect 29499 9344 29541 9353
rect 29499 9304 29500 9344
rect 29540 9304 29541 9344
rect 29499 9295 29541 9304
rect 31419 9344 31461 9353
rect 31419 9304 31420 9344
rect 31460 9304 31461 9344
rect 31419 9295 31461 9304
rect 37275 9344 37317 9353
rect 37275 9304 37276 9344
rect 37316 9304 37317 9344
rect 37275 9295 37317 9304
rect 30267 9260 30309 9269
rect 30267 9220 30268 9260
rect 30308 9220 30309 9260
rect 30267 9211 30309 9220
rect 37659 9260 37701 9269
rect 37659 9220 37660 9260
rect 37700 9220 37701 9260
rect 37659 9211 37701 9220
rect 38043 9260 38085 9269
rect 38043 9220 38044 9260
rect 38084 9220 38085 9260
rect 38043 9211 38085 9220
rect 1152 9092 38112 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 38112 9092
rect 1152 9028 38112 9052
rect 7803 8924 7845 8933
rect 7803 8884 7804 8924
rect 7844 8884 7845 8924
rect 7803 8875 7845 8884
rect 8187 8924 8229 8933
rect 8187 8884 8188 8924
rect 8228 8884 8229 8924
rect 8187 8875 8229 8884
rect 8571 8924 8613 8933
rect 8571 8884 8572 8924
rect 8612 8884 8613 8924
rect 8571 8875 8613 8884
rect 8955 8924 8997 8933
rect 8955 8884 8956 8924
rect 8996 8884 8997 8924
rect 8955 8875 8997 8884
rect 9339 8924 9381 8933
rect 9339 8884 9340 8924
rect 9380 8884 9381 8924
rect 9339 8875 9381 8884
rect 9723 8924 9765 8933
rect 9723 8884 9724 8924
rect 9764 8884 9765 8924
rect 9723 8875 9765 8884
rect 10107 8924 10149 8933
rect 10107 8884 10108 8924
rect 10148 8884 10149 8924
rect 10107 8875 10149 8884
rect 10491 8924 10533 8933
rect 10491 8884 10492 8924
rect 10532 8884 10533 8924
rect 10491 8875 10533 8884
rect 10875 8924 10917 8933
rect 10875 8884 10876 8924
rect 10916 8884 10917 8924
rect 10875 8875 10917 8884
rect 11259 8924 11301 8933
rect 11259 8884 11260 8924
rect 11300 8884 11301 8924
rect 11259 8875 11301 8884
rect 11643 8924 11685 8933
rect 11643 8884 11644 8924
rect 11684 8884 11685 8924
rect 11643 8875 11685 8884
rect 12027 8924 12069 8933
rect 12027 8884 12028 8924
rect 12068 8884 12069 8924
rect 12027 8875 12069 8884
rect 12411 8924 12453 8933
rect 12411 8884 12412 8924
rect 12452 8884 12453 8924
rect 12411 8875 12453 8884
rect 12795 8924 12837 8933
rect 12795 8884 12796 8924
rect 12836 8884 12837 8924
rect 12795 8875 12837 8884
rect 13179 8924 13221 8933
rect 13179 8884 13180 8924
rect 13220 8884 13221 8924
rect 13179 8875 13221 8884
rect 13563 8924 13605 8933
rect 13563 8884 13564 8924
rect 13604 8884 13605 8924
rect 13563 8875 13605 8884
rect 13947 8924 13989 8933
rect 13947 8884 13948 8924
rect 13988 8884 13989 8924
rect 13947 8875 13989 8884
rect 14331 8924 14373 8933
rect 14331 8884 14332 8924
rect 14372 8884 14373 8924
rect 14331 8875 14373 8884
rect 14715 8924 14757 8933
rect 14715 8884 14716 8924
rect 14756 8884 14757 8924
rect 14715 8875 14757 8884
rect 15099 8924 15141 8933
rect 15099 8884 15100 8924
rect 15140 8884 15141 8924
rect 15099 8875 15141 8884
rect 15483 8924 15525 8933
rect 15483 8884 15484 8924
rect 15524 8884 15525 8924
rect 15483 8875 15525 8884
rect 15867 8924 15909 8933
rect 15867 8884 15868 8924
rect 15908 8884 15909 8924
rect 15867 8875 15909 8884
rect 16251 8924 16293 8933
rect 16251 8884 16252 8924
rect 16292 8884 16293 8924
rect 16251 8875 16293 8884
rect 28539 8924 28581 8933
rect 28539 8884 28540 8924
rect 28580 8884 28581 8924
rect 28539 8875 28581 8884
rect 28923 8924 28965 8933
rect 28923 8884 28924 8924
rect 28964 8884 28965 8924
rect 28923 8875 28965 8884
rect 29307 8924 29349 8933
rect 29307 8884 29308 8924
rect 29348 8884 29349 8924
rect 29307 8875 29349 8884
rect 29691 8924 29733 8933
rect 29691 8884 29692 8924
rect 29732 8884 29733 8924
rect 29691 8875 29733 8884
rect 30075 8924 30117 8933
rect 30075 8884 30076 8924
rect 30116 8884 30117 8924
rect 30075 8875 30117 8884
rect 30459 8924 30501 8933
rect 30459 8884 30460 8924
rect 30500 8884 30501 8924
rect 30459 8875 30501 8884
rect 30843 8924 30885 8933
rect 30843 8884 30844 8924
rect 30884 8884 30885 8924
rect 30843 8875 30885 8884
rect 31227 8924 31269 8933
rect 31227 8884 31228 8924
rect 31268 8884 31269 8924
rect 31227 8875 31269 8884
rect 36891 8924 36933 8933
rect 36891 8884 36892 8924
rect 36932 8884 36933 8924
rect 36891 8875 36933 8884
rect 37275 8924 37317 8933
rect 37275 8884 37276 8924
rect 37316 8884 37317 8924
rect 37275 8875 37317 8884
rect 8043 8672 8085 8681
rect 8043 8632 8044 8672
rect 8084 8632 8085 8672
rect 8043 8623 8085 8632
rect 8427 8672 8469 8681
rect 8427 8632 8428 8672
rect 8468 8632 8469 8672
rect 8427 8623 8469 8632
rect 8811 8672 8853 8681
rect 8811 8632 8812 8672
rect 8852 8632 8853 8672
rect 8811 8623 8853 8632
rect 9195 8672 9237 8681
rect 9195 8632 9196 8672
rect 9236 8632 9237 8672
rect 9195 8623 9237 8632
rect 9579 8672 9621 8681
rect 9579 8632 9580 8672
rect 9620 8632 9621 8672
rect 9579 8623 9621 8632
rect 9963 8672 10005 8681
rect 9963 8632 9964 8672
rect 10004 8632 10005 8672
rect 9963 8623 10005 8632
rect 10347 8672 10389 8681
rect 10347 8632 10348 8672
rect 10388 8632 10389 8672
rect 10347 8623 10389 8632
rect 10731 8672 10773 8681
rect 10731 8632 10732 8672
rect 10772 8632 10773 8672
rect 10731 8623 10773 8632
rect 11115 8672 11157 8681
rect 11115 8632 11116 8672
rect 11156 8632 11157 8672
rect 11115 8623 11157 8632
rect 11499 8672 11541 8681
rect 11499 8632 11500 8672
rect 11540 8632 11541 8672
rect 11499 8623 11541 8632
rect 11883 8672 11925 8681
rect 11883 8632 11884 8672
rect 11924 8632 11925 8672
rect 11883 8623 11925 8632
rect 12267 8672 12309 8681
rect 12267 8632 12268 8672
rect 12308 8632 12309 8672
rect 12267 8623 12309 8632
rect 12651 8672 12693 8681
rect 12651 8632 12652 8672
rect 12692 8632 12693 8672
rect 12651 8623 12693 8632
rect 13035 8672 13077 8681
rect 13035 8632 13036 8672
rect 13076 8632 13077 8672
rect 13035 8623 13077 8632
rect 13419 8672 13461 8681
rect 13419 8632 13420 8672
rect 13460 8632 13461 8672
rect 13419 8623 13461 8632
rect 13803 8672 13845 8681
rect 13803 8632 13804 8672
rect 13844 8632 13845 8672
rect 13803 8623 13845 8632
rect 14187 8672 14229 8681
rect 14187 8632 14188 8672
rect 14228 8632 14229 8672
rect 14187 8623 14229 8632
rect 14571 8672 14613 8681
rect 14571 8632 14572 8672
rect 14612 8632 14613 8672
rect 14571 8623 14613 8632
rect 14955 8672 14997 8681
rect 14955 8632 14956 8672
rect 14996 8632 14997 8672
rect 14955 8623 14997 8632
rect 15339 8672 15381 8681
rect 15339 8632 15340 8672
rect 15380 8632 15381 8672
rect 15339 8623 15381 8632
rect 15723 8672 15765 8681
rect 15723 8632 15724 8672
rect 15764 8632 15765 8672
rect 15723 8623 15765 8632
rect 16107 8672 16149 8681
rect 16107 8632 16108 8672
rect 16148 8632 16149 8672
rect 16107 8623 16149 8632
rect 16491 8672 16533 8681
rect 16491 8632 16492 8672
rect 16532 8632 16533 8672
rect 16491 8623 16533 8632
rect 28779 8672 28821 8681
rect 28779 8632 28780 8672
rect 28820 8632 28821 8672
rect 28779 8623 28821 8632
rect 29163 8672 29205 8681
rect 29163 8632 29164 8672
rect 29204 8632 29205 8672
rect 29163 8623 29205 8632
rect 29547 8672 29589 8681
rect 29547 8632 29548 8672
rect 29588 8632 29589 8672
rect 29547 8623 29589 8632
rect 29931 8672 29973 8681
rect 29931 8632 29932 8672
rect 29972 8632 29973 8672
rect 29931 8623 29973 8632
rect 30315 8672 30357 8681
rect 30315 8632 30316 8672
rect 30356 8632 30357 8672
rect 30315 8623 30357 8632
rect 30699 8672 30741 8681
rect 30699 8632 30700 8672
rect 30740 8632 30741 8672
rect 30699 8623 30741 8632
rect 31083 8672 31125 8681
rect 31083 8632 31084 8672
rect 31124 8632 31125 8672
rect 31083 8623 31125 8632
rect 31467 8672 31509 8681
rect 31467 8632 31468 8672
rect 31508 8632 31509 8672
rect 31467 8623 31509 8632
rect 32523 8672 32565 8681
rect 32523 8632 32524 8672
rect 32564 8632 32565 8672
rect 32523 8623 32565 8632
rect 32763 8672 32805 8681
rect 32763 8632 32764 8672
rect 32804 8632 32805 8672
rect 32763 8623 32805 8632
rect 36651 8672 36693 8681
rect 36651 8632 36652 8672
rect 36692 8632 36693 8672
rect 36651 8623 36693 8632
rect 37035 8672 37077 8681
rect 37035 8632 37036 8672
rect 37076 8632 37077 8672
rect 37035 8623 37077 8632
rect 37419 8672 37461 8681
rect 37419 8632 37420 8672
rect 37460 8632 37461 8672
rect 37419 8623 37461 8632
rect 37803 8672 37845 8681
rect 37803 8632 37804 8672
rect 37844 8632 37845 8672
rect 37803 8623 37845 8632
rect 37659 8504 37701 8513
rect 37659 8464 37660 8504
rect 37700 8464 37701 8504
rect 37659 8455 37701 8464
rect 38043 8504 38085 8513
rect 38043 8464 38044 8504
rect 38084 8464 38085 8504
rect 38043 8455 38085 8464
rect 1152 8336 38112 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 38112 8336
rect 1152 8272 38112 8296
rect 29883 8168 29925 8177
rect 29883 8128 29884 8168
rect 29924 8128 29925 8168
rect 29883 8119 29925 8128
rect 30651 8168 30693 8177
rect 30651 8128 30652 8168
rect 30692 8128 30693 8168
rect 30651 8119 30693 8128
rect 32379 8168 32421 8177
rect 32379 8128 32380 8168
rect 32420 8128 32421 8168
rect 32379 8119 32421 8128
rect 31419 8084 31461 8093
rect 31419 8044 31420 8084
rect 31460 8044 31461 8084
rect 31419 8035 31461 8044
rect 19611 8000 19653 8009
rect 19611 7960 19612 8000
rect 19652 7960 19653 8000
rect 19611 7951 19653 7960
rect 19851 8000 19893 8009
rect 19851 7960 19852 8000
rect 19892 7960 19893 8000
rect 19851 7951 19893 7960
rect 20235 8000 20277 8009
rect 20235 7960 20236 8000
rect 20276 7960 20277 8000
rect 20235 7951 20277 7960
rect 22155 8000 22197 8009
rect 22155 7960 22156 8000
rect 22196 7960 22197 8000
rect 22155 7951 22197 7960
rect 23019 8000 23061 8009
rect 23019 7960 23020 8000
rect 23060 7960 23061 8000
rect 23019 7951 23061 7960
rect 23931 8000 23973 8009
rect 23931 7960 23932 8000
rect 23972 7960 23973 8000
rect 23931 7951 23973 7960
rect 24171 8000 24213 8009
rect 24171 7960 24172 8000
rect 24212 7960 24213 8000
rect 24171 7951 24213 7960
rect 25515 8000 25557 8009
rect 25515 7960 25516 8000
rect 25556 7960 25557 8000
rect 25515 7951 25557 7960
rect 26187 8000 26229 8009
rect 26187 7960 26188 8000
rect 26228 7960 26229 8000
rect 26187 7951 26229 7960
rect 26763 8000 26805 8009
rect 26763 7960 26764 8000
rect 26804 7960 26805 8000
rect 26763 7951 26805 7960
rect 27579 8000 27621 8009
rect 27579 7960 27580 8000
rect 27620 7960 27621 8000
rect 27579 7951 27621 7960
rect 27819 8000 27861 8009
rect 27819 7960 27820 8000
rect 27860 7960 27861 8000
rect 27819 7951 27861 7960
rect 29643 8000 29685 8009
rect 29643 7960 29644 8000
rect 29684 7960 29685 8000
rect 29643 7951 29685 7960
rect 30027 8000 30069 8009
rect 30027 7960 30028 8000
rect 30068 7960 30069 8000
rect 30027 7951 30069 7960
rect 30411 8000 30453 8009
rect 30411 7960 30412 8000
rect 30452 7960 30453 8000
rect 30411 7951 30453 7960
rect 30795 8000 30837 8009
rect 30795 7960 30796 8000
rect 30836 7960 30837 8000
rect 30795 7951 30837 7960
rect 31179 8000 31221 8009
rect 31179 7960 31180 8000
rect 31220 7960 31221 8000
rect 31179 7951 31221 7960
rect 32139 8000 32181 8009
rect 32139 7960 32140 8000
rect 32180 7960 32181 8000
rect 32139 7951 32181 7960
rect 37419 8000 37461 8009
rect 37419 7960 37420 8000
rect 37460 7960 37461 8000
rect 37419 7951 37461 7960
rect 37803 8000 37845 8009
rect 37803 7960 37804 8000
rect 37844 7960 37845 8000
rect 37803 7951 37845 7960
rect 19995 7832 20037 7841
rect 19995 7792 19996 7832
rect 20036 7792 20037 7832
rect 19995 7783 20037 7792
rect 21915 7832 21957 7841
rect 21915 7792 21916 7832
rect 21956 7792 21957 7832
rect 21915 7783 21957 7792
rect 26427 7832 26469 7841
rect 26427 7792 26428 7832
rect 26468 7792 26469 7832
rect 26427 7783 26469 7792
rect 22779 7748 22821 7757
rect 22779 7708 22780 7748
rect 22820 7708 22821 7748
rect 22779 7699 22821 7708
rect 25275 7748 25317 7757
rect 25275 7708 25276 7748
rect 25316 7708 25317 7748
rect 25275 7699 25317 7708
rect 26523 7748 26565 7757
rect 26523 7708 26524 7748
rect 26564 7708 26565 7748
rect 26523 7699 26565 7708
rect 30267 7748 30309 7757
rect 30267 7708 30268 7748
rect 30308 7708 30309 7748
rect 30267 7699 30309 7708
rect 31035 7748 31077 7757
rect 31035 7708 31036 7748
rect 31076 7708 31077 7748
rect 31035 7699 31077 7708
rect 37659 7748 37701 7757
rect 37659 7708 37660 7748
rect 37700 7708 37701 7748
rect 37659 7699 37701 7708
rect 38043 7748 38085 7757
rect 38043 7708 38044 7748
rect 38084 7708 38085 7748
rect 38043 7699 38085 7708
rect 1152 7580 38112 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 38112 7580
rect 1152 7516 38112 7540
rect 19707 7412 19749 7421
rect 19707 7372 19708 7412
rect 19748 7372 19749 7412
rect 19707 7363 19749 7372
rect 30267 7412 30309 7421
rect 30267 7372 30268 7412
rect 30308 7372 30309 7412
rect 30267 7363 30309 7372
rect 18795 7160 18837 7169
rect 18795 7120 18796 7160
rect 18836 7120 18837 7160
rect 18795 7111 18837 7120
rect 19179 7160 19221 7169
rect 19179 7120 19180 7160
rect 19220 7120 19221 7160
rect 19179 7111 19221 7120
rect 19563 7160 19605 7169
rect 19563 7120 19564 7160
rect 19604 7120 19605 7160
rect 19563 7111 19605 7120
rect 19947 7160 19989 7169
rect 19947 7120 19948 7160
rect 19988 7120 19989 7160
rect 19947 7111 19989 7120
rect 20091 7160 20133 7169
rect 20091 7120 20092 7160
rect 20132 7120 20133 7160
rect 20091 7111 20133 7120
rect 20331 7160 20373 7169
rect 20331 7120 20332 7160
rect 20372 7120 20373 7160
rect 20331 7111 20373 7120
rect 20715 7160 20757 7169
rect 20715 7120 20716 7160
rect 20756 7120 20757 7160
rect 20715 7111 20757 7120
rect 21387 7160 21429 7169
rect 21387 7120 21388 7160
rect 21428 7120 21429 7160
rect 21387 7111 21429 7120
rect 25611 7160 25653 7169
rect 25611 7120 25612 7160
rect 25652 7120 25653 7160
rect 25611 7111 25653 7120
rect 29643 7160 29685 7169
rect 29643 7120 29644 7160
rect 29684 7120 29685 7160
rect 29643 7111 29685 7120
rect 30027 7160 30069 7169
rect 30027 7120 30028 7160
rect 30068 7120 30069 7160
rect 30027 7111 30069 7120
rect 31083 7160 31125 7169
rect 31083 7120 31084 7160
rect 31124 7120 31125 7160
rect 31083 7111 31125 7120
rect 31323 7160 31365 7169
rect 31323 7120 31324 7160
rect 31364 7120 31365 7160
rect 31323 7111 31365 7120
rect 37419 7160 37461 7169
rect 37419 7120 37420 7160
rect 37460 7120 37461 7160
rect 37419 7111 37461 7120
rect 37803 7160 37845 7169
rect 37803 7120 37804 7160
rect 37844 7120 37845 7160
rect 37803 7111 37845 7120
rect 18939 7076 18981 7085
rect 18939 7036 18940 7076
rect 18980 7036 18981 7076
rect 18939 7027 18981 7036
rect 29883 7076 29925 7085
rect 29883 7036 29884 7076
rect 29924 7036 29925 7076
rect 29883 7027 29925 7036
rect 18555 6992 18597 7001
rect 18555 6952 18556 6992
rect 18596 6952 18597 6992
rect 18555 6943 18597 6952
rect 19323 6992 19365 7001
rect 19323 6952 19324 6992
rect 19364 6952 19365 6992
rect 19323 6943 19365 6952
rect 20475 6992 20517 7001
rect 20475 6952 20476 6992
rect 20516 6952 20517 6992
rect 20475 6943 20517 6952
rect 21147 6992 21189 7001
rect 21147 6952 21148 6992
rect 21188 6952 21189 6992
rect 21147 6943 21189 6952
rect 25851 6992 25893 7001
rect 25851 6952 25852 6992
rect 25892 6952 25893 6992
rect 25851 6943 25893 6952
rect 37659 6992 37701 7001
rect 37659 6952 37660 6992
rect 37700 6952 37701 6992
rect 37659 6943 37701 6952
rect 38043 6992 38085 7001
rect 38043 6952 38044 6992
rect 38084 6952 38085 6992
rect 38043 6943 38085 6952
rect 1152 6824 38112 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 38112 6824
rect 1152 6760 38112 6784
rect 16731 6656 16773 6665
rect 16731 6616 16732 6656
rect 16772 6616 16773 6656
rect 16731 6607 16773 6616
rect 19803 6656 19845 6665
rect 19803 6616 19804 6656
rect 19844 6616 19845 6656
rect 19803 6607 19845 6616
rect 29691 6656 29733 6665
rect 29691 6616 29692 6656
rect 29732 6616 29733 6656
rect 29691 6607 29733 6616
rect 30075 6656 30117 6665
rect 30075 6616 30076 6656
rect 30116 6616 30117 6656
rect 30075 6607 30117 6616
rect 31899 6656 31941 6665
rect 31899 6616 31900 6656
rect 31940 6616 31941 6656
rect 31899 6607 31941 6616
rect 16971 6488 17013 6497
rect 16971 6448 16972 6488
rect 17012 6448 17013 6488
rect 16971 6439 17013 6448
rect 20043 6488 20085 6497
rect 20043 6448 20044 6488
rect 20084 6448 20085 6488
rect 20043 6439 20085 6448
rect 29451 6488 29493 6497
rect 29451 6448 29452 6488
rect 29492 6448 29493 6488
rect 29451 6439 29493 6448
rect 29835 6488 29877 6497
rect 29835 6448 29836 6488
rect 29876 6448 29877 6488
rect 29835 6439 29877 6448
rect 31659 6488 31701 6497
rect 31659 6448 31660 6488
rect 31700 6448 31701 6488
rect 31659 6439 31701 6448
rect 37419 6488 37461 6497
rect 37419 6448 37420 6488
rect 37460 6448 37461 6488
rect 37419 6439 37461 6448
rect 37803 6488 37845 6497
rect 37803 6448 37804 6488
rect 37844 6448 37845 6488
rect 37803 6439 37845 6448
rect 38043 6320 38085 6329
rect 38043 6280 38044 6320
rect 38084 6280 38085 6320
rect 38043 6271 38085 6280
rect 37659 6236 37701 6245
rect 37659 6196 37660 6236
rect 37700 6196 37701 6236
rect 37659 6187 37701 6196
rect 1152 6068 38112 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 38112 6068
rect 1152 6004 38112 6028
rect 6843 5900 6885 5909
rect 6843 5860 6844 5900
rect 6884 5860 6885 5900
rect 6843 5851 6885 5860
rect 15003 5900 15045 5909
rect 15003 5860 15004 5900
rect 15044 5860 15045 5900
rect 15003 5851 15045 5860
rect 16923 5816 16965 5825
rect 16923 5776 16924 5816
rect 16964 5776 16965 5816
rect 16923 5767 16965 5776
rect 5451 5648 5493 5657
rect 5451 5608 5452 5648
rect 5492 5608 5493 5648
rect 5451 5599 5493 5608
rect 5835 5648 5877 5657
rect 5835 5608 5836 5648
rect 5876 5608 5877 5648
rect 5835 5599 5877 5608
rect 6219 5648 6261 5657
rect 6219 5608 6220 5648
rect 6260 5608 6261 5648
rect 6219 5599 6261 5608
rect 6603 5648 6645 5657
rect 6603 5608 6604 5648
rect 6644 5608 6645 5648
rect 6603 5599 6645 5608
rect 6987 5648 7029 5657
rect 6987 5608 6988 5648
rect 7028 5608 7029 5648
rect 6987 5599 7029 5608
rect 7227 5648 7269 5657
rect 7227 5608 7228 5648
rect 7268 5608 7269 5648
rect 7227 5599 7269 5608
rect 15243 5648 15285 5657
rect 15243 5608 15244 5648
rect 15284 5608 15285 5648
rect 15243 5599 15285 5608
rect 15387 5648 15429 5657
rect 15387 5608 15388 5648
rect 15428 5608 15429 5648
rect 15387 5599 15429 5608
rect 15627 5648 15669 5657
rect 15627 5608 15628 5648
rect 15668 5608 15669 5648
rect 15627 5599 15669 5608
rect 16011 5648 16053 5657
rect 16011 5608 16012 5648
rect 16052 5608 16053 5648
rect 16011 5599 16053 5608
rect 16395 5648 16437 5657
rect 16395 5608 16396 5648
rect 16436 5608 16437 5648
rect 16395 5599 16437 5608
rect 16779 5648 16821 5657
rect 16779 5608 16780 5648
rect 16820 5608 16821 5648
rect 16779 5599 16821 5608
rect 17163 5648 17205 5657
rect 17163 5608 17164 5648
rect 17204 5608 17205 5648
rect 17163 5599 17205 5608
rect 17547 5648 17589 5657
rect 17547 5608 17548 5648
rect 17588 5608 17589 5648
rect 17547 5599 17589 5608
rect 17691 5648 17733 5657
rect 17691 5608 17692 5648
rect 17732 5608 17733 5648
rect 17691 5599 17733 5608
rect 17931 5648 17973 5657
rect 17931 5608 17932 5648
rect 17972 5608 17973 5648
rect 17931 5599 17973 5608
rect 29067 5648 29109 5657
rect 29067 5608 29068 5648
rect 29108 5608 29109 5648
rect 29067 5599 29109 5608
rect 29307 5648 29349 5657
rect 29307 5608 29308 5648
rect 29348 5608 29349 5648
rect 29307 5599 29349 5608
rect 37419 5648 37461 5657
rect 37419 5608 37420 5648
rect 37460 5608 37461 5648
rect 37419 5599 37461 5608
rect 37803 5648 37845 5657
rect 37803 5608 37804 5648
rect 37844 5608 37845 5648
rect 37803 5599 37845 5608
rect 38043 5648 38085 5657
rect 38043 5608 38044 5648
rect 38084 5608 38085 5648
rect 38043 5599 38085 5608
rect 5691 5564 5733 5573
rect 5691 5524 5692 5564
rect 5732 5524 5733 5564
rect 5691 5515 5733 5524
rect 6459 5564 6501 5573
rect 6459 5524 6460 5564
rect 6500 5524 6501 5564
rect 6459 5515 6501 5524
rect 15771 5564 15813 5573
rect 15771 5524 15772 5564
rect 15812 5524 15813 5564
rect 15771 5515 15813 5524
rect 17307 5564 17349 5573
rect 17307 5524 17308 5564
rect 17348 5524 17349 5564
rect 17307 5515 17349 5524
rect 6075 5480 6117 5489
rect 6075 5440 6076 5480
rect 6116 5440 6117 5480
rect 6075 5431 6117 5440
rect 16155 5480 16197 5489
rect 16155 5440 16156 5480
rect 16196 5440 16197 5480
rect 16155 5431 16197 5440
rect 16539 5480 16581 5489
rect 16539 5440 16540 5480
rect 16580 5440 16581 5480
rect 16539 5431 16581 5440
rect 37659 5480 37701 5489
rect 37659 5440 37660 5480
rect 37700 5440 37701 5480
rect 37659 5431 37701 5440
rect 1152 5312 38112 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 38112 5312
rect 1152 5248 38112 5272
rect 6075 5144 6117 5153
rect 6075 5104 6076 5144
rect 6116 5104 6117 5144
rect 6075 5095 6117 5104
rect 7131 5144 7173 5153
rect 7131 5104 7132 5144
rect 7172 5104 7173 5144
rect 7131 5095 7173 5104
rect 7515 5144 7557 5153
rect 7515 5104 7516 5144
rect 7556 5104 7557 5144
rect 7515 5095 7557 5104
rect 8283 5144 8325 5153
rect 8283 5104 8284 5144
rect 8324 5104 8325 5144
rect 8283 5095 8325 5104
rect 9051 5144 9093 5153
rect 9051 5104 9052 5144
rect 9092 5104 9093 5144
rect 9051 5095 9093 5104
rect 9435 5144 9477 5153
rect 9435 5104 9436 5144
rect 9476 5104 9477 5144
rect 9435 5095 9477 5104
rect 11739 5144 11781 5153
rect 11739 5104 11740 5144
rect 11780 5104 11781 5144
rect 11739 5095 11781 5104
rect 12507 5144 12549 5153
rect 12507 5104 12508 5144
rect 12548 5104 12549 5144
rect 12507 5095 12549 5104
rect 14523 5144 14565 5153
rect 14523 5104 14524 5144
rect 14564 5104 14565 5144
rect 14523 5095 14565 5104
rect 29211 5144 29253 5153
rect 29211 5104 29212 5144
rect 29252 5104 29253 5144
rect 29211 5095 29253 5104
rect 7899 5060 7941 5069
rect 7899 5020 7900 5060
rect 7940 5020 7941 5060
rect 7899 5011 7941 5020
rect 8667 5060 8709 5069
rect 8667 5020 8668 5060
rect 8708 5020 8709 5060
rect 8667 5011 8709 5020
rect 13659 5060 13701 5069
rect 13659 5020 13660 5060
rect 13700 5020 13701 5060
rect 13659 5011 13701 5020
rect 17115 5060 17157 5069
rect 17115 5020 17116 5060
rect 17156 5020 17157 5060
rect 17115 5011 17157 5020
rect 5835 4976 5877 4985
rect 5835 4936 5836 4976
rect 5876 4936 5877 4976
rect 5835 4927 5877 4936
rect 6891 4976 6933 4985
rect 6891 4936 6892 4976
rect 6932 4936 6933 4976
rect 6891 4927 6933 4936
rect 7275 4976 7317 4985
rect 7275 4936 7276 4976
rect 7316 4936 7317 4976
rect 7275 4927 7317 4936
rect 7659 4976 7701 4985
rect 7659 4936 7660 4976
rect 7700 4936 7701 4976
rect 7659 4927 7701 4936
rect 8043 4976 8085 4985
rect 8043 4936 8044 4976
rect 8084 4936 8085 4976
rect 8043 4927 8085 4936
rect 8427 4976 8469 4985
rect 8427 4936 8428 4976
rect 8468 4936 8469 4976
rect 8427 4927 8469 4936
rect 8811 4976 8853 4985
rect 8811 4936 8812 4976
rect 8852 4936 8853 4976
rect 8811 4927 8853 4936
rect 9195 4976 9237 4985
rect 9195 4936 9196 4976
rect 9236 4936 9237 4976
rect 9195 4927 9237 4936
rect 11979 4976 12021 4985
rect 11979 4936 11980 4976
rect 12020 4936 12021 4976
rect 11979 4927 12021 4936
rect 12123 4976 12165 4985
rect 12123 4936 12124 4976
rect 12164 4936 12165 4976
rect 12123 4927 12165 4936
rect 12363 4976 12405 4985
rect 12363 4936 12364 4976
rect 12404 4936 12405 4976
rect 12363 4927 12405 4936
rect 12747 4976 12789 4985
rect 12747 4936 12748 4976
rect 12788 4936 12789 4976
rect 12747 4927 12789 4936
rect 13131 4976 13173 4985
rect 13131 4936 13132 4976
rect 13172 4936 13173 4976
rect 13131 4927 13173 4936
rect 13515 4976 13557 4985
rect 13515 4936 13516 4976
rect 13556 4936 13557 4976
rect 13515 4927 13557 4936
rect 13899 4976 13941 4985
rect 13899 4936 13900 4976
rect 13940 4936 13941 4976
rect 13899 4927 13941 4936
rect 14763 4976 14805 4985
rect 14763 4936 14764 4976
rect 14804 4936 14805 4976
rect 14763 4927 14805 4936
rect 16971 4976 17013 4985
rect 16971 4936 16972 4976
rect 17012 4936 17013 4976
rect 16971 4927 17013 4936
rect 17355 4976 17397 4985
rect 17355 4936 17356 4976
rect 17396 4936 17397 4976
rect 17355 4927 17397 4936
rect 23979 4976 24021 4985
rect 23979 4936 23980 4976
rect 24020 4936 24021 4976
rect 23979 4927 24021 4936
rect 28971 4976 29013 4985
rect 28971 4936 28972 4976
rect 29012 4936 29013 4976
rect 28971 4927 29013 4936
rect 37419 4976 37461 4985
rect 37419 4936 37420 4976
rect 37460 4936 37461 4976
rect 37419 4927 37461 4936
rect 37803 4976 37845 4985
rect 37803 4936 37804 4976
rect 37844 4936 37845 4976
rect 37803 4927 37845 4936
rect 38043 4976 38085 4985
rect 38043 4936 38044 4976
rect 38084 4936 38085 4976
rect 38043 4927 38085 4936
rect 12891 4808 12933 4817
rect 12891 4768 12892 4808
rect 12932 4768 12933 4808
rect 12891 4759 12933 4768
rect 16731 4808 16773 4817
rect 16731 4768 16732 4808
rect 16772 4768 16773 4808
rect 16731 4759 16773 4768
rect 13275 4724 13317 4733
rect 13275 4684 13276 4724
rect 13316 4684 13317 4724
rect 13275 4675 13317 4684
rect 24219 4724 24261 4733
rect 24219 4684 24220 4724
rect 24260 4684 24261 4724
rect 24219 4675 24261 4684
rect 37659 4724 37701 4733
rect 37659 4684 37660 4724
rect 37700 4684 37701 4724
rect 37659 4675 37701 4684
rect 1152 4556 38112 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 38112 4556
rect 1152 4492 38112 4516
rect 3483 4304 3525 4313
rect 3483 4264 3484 4304
rect 3524 4264 3525 4304
rect 3483 4255 3525 4264
rect 8475 4304 8517 4313
rect 8475 4264 8476 4304
rect 8516 4264 8517 4304
rect 8475 4255 8517 4264
rect 9627 4304 9669 4313
rect 9627 4264 9628 4304
rect 9668 4264 9669 4304
rect 9627 4255 9669 4264
rect 11643 4304 11685 4313
rect 11643 4264 11644 4304
rect 11684 4264 11685 4304
rect 11643 4255 11685 4264
rect 24603 4304 24645 4313
rect 24603 4264 24604 4304
rect 24644 4264 24645 4304
rect 24603 4255 24645 4264
rect 29403 4304 29445 4313
rect 29403 4264 29404 4304
rect 29444 4264 29445 4304
rect 29403 4255 29445 4264
rect 38043 4304 38085 4313
rect 38043 4264 38044 4304
rect 38084 4264 38085 4304
rect 38043 4255 38085 4264
rect 3243 4136 3285 4145
rect 3243 4096 3244 4136
rect 3284 4096 3285 4136
rect 3243 4087 3285 4096
rect 3915 4136 3957 4145
rect 3915 4096 3916 4136
rect 3956 4096 3957 4136
rect 3915 4087 3957 4096
rect 8235 4136 8277 4145
rect 8235 4096 8236 4136
rect 8276 4096 8277 4136
rect 8235 4087 8277 4096
rect 9387 4136 9429 4145
rect 9387 4096 9388 4136
rect 9428 4096 9429 4136
rect 9387 4087 9429 4096
rect 10059 4136 10101 4145
rect 10059 4096 10060 4136
rect 10100 4096 10101 4136
rect 10059 4087 10101 4096
rect 10683 4136 10725 4145
rect 10683 4096 10684 4136
rect 10724 4096 10725 4136
rect 10683 4087 10725 4096
rect 10923 4136 10965 4145
rect 10923 4096 10924 4136
rect 10964 4096 10965 4136
rect 10923 4087 10965 4096
rect 11818 4136 11876 4137
rect 11818 4096 11827 4136
rect 11867 4096 11876 4136
rect 11818 4095 11876 4096
rect 24363 4136 24405 4145
rect 24363 4096 24364 4136
rect 24404 4096 24405 4136
rect 24363 4087 24405 4096
rect 29163 4136 29205 4145
rect 29163 4096 29164 4136
rect 29204 4096 29205 4136
rect 29163 4087 29205 4096
rect 37419 4136 37461 4145
rect 37419 4096 37420 4136
rect 37460 4096 37461 4136
rect 37419 4087 37461 4096
rect 37803 4136 37845 4145
rect 37803 4096 37804 4136
rect 37844 4096 37845 4136
rect 37803 4087 37845 4096
rect 4155 4052 4197 4061
rect 4155 4012 4156 4052
rect 4196 4012 4197 4052
rect 4155 4003 4197 4012
rect 37659 4052 37701 4061
rect 37659 4012 37660 4052
rect 37700 4012 37701 4052
rect 37659 4003 37701 4012
rect 10299 3968 10341 3977
rect 10299 3928 10300 3968
rect 10340 3928 10341 3968
rect 10299 3919 10341 3928
rect 1152 3800 38112 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 38112 3800
rect 1152 3736 38112 3760
rect 22587 3632 22629 3641
rect 22587 3592 22588 3632
rect 22628 3592 22629 3632
rect 22587 3583 22629 3592
rect 28827 3632 28869 3641
rect 28827 3592 28828 3632
rect 28868 3592 28869 3632
rect 28827 3583 28869 3592
rect 38043 3632 38085 3641
rect 38043 3592 38044 3632
rect 38084 3592 38085 3632
rect 38043 3583 38085 3592
rect 21819 3548 21861 3557
rect 21819 3508 21820 3548
rect 21860 3508 21861 3548
rect 21819 3499 21861 3508
rect 26523 3548 26565 3557
rect 26523 3508 26524 3548
rect 26564 3508 26565 3548
rect 26523 3499 26565 3508
rect 5355 3464 5397 3473
rect 5355 3424 5356 3464
rect 5396 3424 5397 3464
rect 5355 3415 5397 3424
rect 15627 3464 15669 3473
rect 15627 3424 15628 3464
rect 15668 3424 15669 3464
rect 15627 3415 15669 3424
rect 18507 3464 18549 3473
rect 18507 3424 18508 3464
rect 18548 3424 18549 3464
rect 18507 3415 18549 3424
rect 18891 3464 18933 3473
rect 18891 3424 18892 3464
rect 18932 3424 18933 3464
rect 18891 3415 18933 3424
rect 19563 3464 19605 3473
rect 19563 3424 19564 3464
rect 19604 3424 19605 3464
rect 19563 3415 19605 3424
rect 19947 3464 19989 3473
rect 19947 3424 19948 3464
rect 19988 3424 19989 3464
rect 19947 3415 19989 3424
rect 20331 3464 20373 3473
rect 20331 3424 20332 3464
rect 20372 3424 20373 3464
rect 20331 3415 20373 3424
rect 20715 3464 20757 3473
rect 20715 3424 20716 3464
rect 20756 3424 20757 3464
rect 20715 3415 20757 3424
rect 20955 3464 20997 3473
rect 20955 3424 20956 3464
rect 20996 3424 20997 3464
rect 20955 3415 20997 3424
rect 21195 3464 21237 3473
rect 21195 3424 21196 3464
rect 21236 3424 21237 3464
rect 21195 3415 21237 3424
rect 21435 3464 21477 3473
rect 21435 3424 21436 3464
rect 21476 3424 21477 3464
rect 21435 3415 21477 3424
rect 21579 3464 21621 3473
rect 21579 3424 21580 3464
rect 21620 3424 21621 3464
rect 21579 3415 21621 3424
rect 22347 3464 22389 3473
rect 22347 3424 22348 3464
rect 22388 3424 22389 3464
rect 22347 3415 22389 3424
rect 26283 3464 26325 3473
rect 26283 3424 26284 3464
rect 26324 3424 26325 3464
rect 26283 3415 26325 3424
rect 28587 3464 28629 3473
rect 28587 3424 28588 3464
rect 28628 3424 28629 3464
rect 28587 3415 28629 3424
rect 37419 3464 37461 3473
rect 37419 3424 37420 3464
rect 37460 3424 37461 3464
rect 37419 3415 37461 3424
rect 37803 3464 37845 3473
rect 37803 3424 37804 3464
rect 37844 3424 37845 3464
rect 37803 3415 37845 3424
rect 19131 3296 19173 3305
rect 19131 3256 19132 3296
rect 19172 3256 19173 3296
rect 19131 3247 19173 3256
rect 20187 3296 20229 3305
rect 20187 3256 20188 3296
rect 20228 3256 20229 3296
rect 20187 3247 20229 3256
rect 37659 3296 37701 3305
rect 37659 3256 37660 3296
rect 37700 3256 37701 3296
rect 37659 3247 37701 3256
rect 5595 3212 5637 3221
rect 5595 3172 5596 3212
rect 5636 3172 5637 3212
rect 5595 3163 5637 3172
rect 15867 3212 15909 3221
rect 15867 3172 15868 3212
rect 15908 3172 15909 3212
rect 15867 3163 15909 3172
rect 18747 3212 18789 3221
rect 18747 3172 18748 3212
rect 18788 3172 18789 3212
rect 18747 3163 18789 3172
rect 19803 3212 19845 3221
rect 19803 3172 19804 3212
rect 19844 3172 19845 3212
rect 19803 3163 19845 3172
rect 20571 3212 20613 3221
rect 20571 3172 20572 3212
rect 20612 3172 20613 3212
rect 20571 3163 20613 3172
rect 1152 3044 38112 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 38112 3044
rect 1152 2980 38112 3004
rect 8187 2876 8229 2885
rect 8187 2836 8188 2876
rect 8228 2836 8229 2876
rect 8187 2827 8229 2836
rect 8571 2876 8613 2885
rect 8571 2836 8572 2876
rect 8612 2836 8613 2876
rect 8571 2827 8613 2836
rect 14619 2876 14661 2885
rect 14619 2836 14620 2876
rect 14660 2836 14661 2876
rect 14619 2827 14661 2836
rect 15675 2876 15717 2885
rect 15675 2836 15676 2876
rect 15716 2836 15717 2876
rect 15675 2827 15717 2836
rect 17595 2876 17637 2885
rect 17595 2836 17596 2876
rect 17636 2836 17637 2876
rect 17595 2827 17637 2836
rect 21435 2876 21477 2885
rect 21435 2836 21436 2876
rect 21476 2836 21477 2876
rect 21435 2827 21477 2836
rect 27291 2876 27333 2885
rect 27291 2836 27292 2876
rect 27332 2836 27333 2876
rect 27291 2827 27333 2836
rect 29307 2876 29349 2885
rect 29307 2836 29308 2876
rect 29348 2836 29349 2876
rect 29307 2827 29349 2836
rect 30747 2876 30789 2885
rect 30747 2836 30748 2876
rect 30788 2836 30789 2876
rect 30747 2827 30789 2836
rect 38043 2876 38085 2885
rect 38043 2836 38044 2876
rect 38084 2836 38085 2876
rect 38043 2827 38085 2836
rect 25467 2792 25509 2801
rect 25467 2752 25468 2792
rect 25508 2752 25509 2792
rect 25467 2743 25509 2752
rect 25851 2792 25893 2801
rect 25851 2752 25852 2792
rect 25892 2752 25893 2792
rect 25851 2743 25893 2752
rect 28059 2792 28101 2801
rect 28059 2752 28060 2792
rect 28100 2752 28101 2792
rect 28059 2743 28101 2752
rect 7947 2624 7989 2633
rect 7947 2584 7948 2624
rect 7988 2584 7989 2624
rect 7947 2575 7989 2584
rect 8331 2624 8373 2633
rect 8331 2584 8332 2624
rect 8372 2584 8373 2624
rect 8331 2575 8373 2584
rect 11499 2624 11541 2633
rect 11499 2584 11500 2624
rect 11540 2584 11541 2624
rect 11499 2575 11541 2584
rect 13323 2624 13365 2633
rect 13323 2584 13324 2624
rect 13364 2584 13365 2624
rect 13323 2575 13365 2584
rect 14379 2624 14421 2633
rect 14379 2584 14380 2624
rect 14420 2584 14421 2624
rect 14379 2575 14421 2584
rect 14763 2624 14805 2633
rect 14763 2584 14764 2624
rect 14804 2584 14805 2624
rect 14763 2575 14805 2584
rect 15435 2624 15477 2633
rect 15435 2584 15436 2624
rect 15476 2584 15477 2624
rect 15435 2575 15477 2584
rect 15819 2624 15861 2633
rect 15819 2584 15820 2624
rect 15860 2584 15861 2624
rect 15819 2575 15861 2584
rect 17355 2624 17397 2633
rect 17355 2584 17356 2624
rect 17396 2584 17397 2624
rect 17355 2575 17397 2584
rect 21195 2624 21237 2633
rect 21195 2584 21196 2624
rect 21236 2584 21237 2624
rect 21195 2575 21237 2584
rect 21579 2624 21621 2633
rect 21579 2584 21580 2624
rect 21620 2584 21621 2624
rect 21579 2575 21621 2584
rect 25227 2624 25269 2633
rect 25227 2584 25228 2624
rect 25268 2584 25269 2624
rect 25227 2575 25269 2584
rect 25611 2624 25653 2633
rect 25611 2584 25612 2624
rect 25652 2584 25653 2624
rect 25611 2575 25653 2584
rect 27051 2624 27093 2633
rect 27051 2584 27052 2624
rect 27092 2584 27093 2624
rect 27051 2575 27093 2584
rect 27435 2624 27477 2633
rect 27435 2584 27436 2624
rect 27476 2584 27477 2624
rect 27435 2575 27477 2584
rect 27819 2624 27861 2633
rect 27819 2584 27820 2624
rect 27860 2584 27861 2624
rect 27819 2575 27861 2584
rect 29547 2624 29589 2633
rect 29547 2584 29548 2624
rect 29588 2584 29589 2624
rect 29547 2575 29589 2584
rect 30987 2624 31029 2633
rect 30987 2584 30988 2624
rect 31028 2584 31029 2624
rect 30987 2575 31029 2584
rect 37035 2624 37077 2633
rect 37035 2584 37036 2624
rect 37076 2584 37077 2624
rect 37035 2575 37077 2584
rect 37419 2624 37461 2633
rect 37419 2584 37420 2624
rect 37460 2584 37461 2624
rect 37419 2575 37461 2584
rect 37803 2624 37845 2633
rect 37803 2584 37804 2624
rect 37844 2584 37845 2624
rect 37803 2575 37845 2584
rect 15003 2540 15045 2549
rect 15003 2500 15004 2540
rect 15044 2500 15045 2540
rect 15003 2491 15045 2500
rect 37659 2540 37701 2549
rect 37659 2500 37660 2540
rect 37700 2500 37701 2540
rect 37659 2491 37701 2500
rect 11739 2456 11781 2465
rect 11739 2416 11740 2456
rect 11780 2416 11781 2456
rect 11739 2407 11781 2416
rect 13563 2456 13605 2465
rect 13563 2416 13564 2456
rect 13604 2416 13605 2456
rect 13563 2407 13605 2416
rect 16059 2456 16101 2465
rect 16059 2416 16060 2456
rect 16100 2416 16101 2456
rect 16059 2407 16101 2416
rect 21819 2456 21861 2465
rect 21819 2416 21820 2456
rect 21860 2416 21861 2456
rect 21819 2407 21861 2416
rect 27675 2456 27717 2465
rect 27675 2416 27676 2456
rect 27716 2416 27717 2456
rect 27675 2407 27717 2416
rect 37275 2456 37317 2465
rect 37275 2416 37276 2456
rect 37316 2416 37317 2456
rect 37275 2407 37317 2416
rect 1152 2288 38112 2312
rect 1152 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 38112 2288
rect 1152 2224 38112 2248
rect 38043 2120 38085 2129
rect 38043 2080 38044 2120
rect 38084 2080 38085 2120
rect 38043 2071 38085 2080
rect 36267 1952 36309 1961
rect 36267 1912 36268 1952
rect 36308 1912 36309 1952
rect 36267 1903 36309 1912
rect 36651 1952 36693 1961
rect 36651 1912 36652 1952
rect 36692 1912 36693 1952
rect 36651 1903 36693 1912
rect 37035 1952 37077 1961
rect 37035 1912 37036 1952
rect 37076 1912 37077 1952
rect 37035 1903 37077 1912
rect 37419 1952 37461 1961
rect 37419 1912 37420 1952
rect 37460 1912 37461 1952
rect 37419 1903 37461 1912
rect 37803 1952 37845 1961
rect 37803 1912 37804 1952
rect 37844 1912 37845 1952
rect 37803 1903 37845 1912
rect 36891 1784 36933 1793
rect 36891 1744 36892 1784
rect 36932 1744 36933 1784
rect 36891 1735 36933 1744
rect 36507 1700 36549 1709
rect 36507 1660 36508 1700
rect 36548 1660 36549 1700
rect 36507 1651 36549 1660
rect 37275 1700 37317 1709
rect 37275 1660 37276 1700
rect 37316 1660 37317 1700
rect 37275 1651 37317 1660
rect 37659 1700 37701 1709
rect 37659 1660 37660 1700
rect 37700 1660 37701 1700
rect 37659 1651 37701 1660
rect 1152 1532 38112 1556
rect 1152 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 38112 1532
rect 1152 1468 38112 1492
<< via1 >>
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 7324 9640 7364 9680
rect 7708 9640 7748 9680
rect 8092 9640 8132 9680
rect 8476 9640 8516 9680
rect 8860 9640 8900 9680
rect 9244 9640 9284 9680
rect 9628 9640 9668 9680
rect 10012 9640 10052 9680
rect 10396 9640 10436 9680
rect 10780 9640 10820 9680
rect 11164 9640 11204 9680
rect 11548 9640 11588 9680
rect 11932 9640 11972 9680
rect 12316 9640 12356 9680
rect 12700 9640 12740 9680
rect 13084 9640 13124 9680
rect 13468 9640 13508 9680
rect 13852 9640 13892 9680
rect 14236 9640 14276 9680
rect 14620 9640 14660 9680
rect 15004 9640 15044 9680
rect 15388 9640 15428 9680
rect 15772 9640 15812 9680
rect 16540 9640 16580 9680
rect 17020 9640 17060 9680
rect 17404 9640 17444 9680
rect 27580 9640 27620 9680
rect 28348 9640 28388 9680
rect 29116 9640 29156 9680
rect 30652 9640 30692 9680
rect 31036 9640 31076 9680
rect 32188 9640 32228 9680
rect 36124 9640 36164 9680
rect 36508 9640 36548 9680
rect 36892 9640 36932 9680
rect 16636 9556 16676 9596
rect 17788 9556 17828 9596
rect 27964 9556 28004 9596
rect 28732 9556 28772 9596
rect 29884 9556 29924 9596
rect 31804 9556 31844 9596
rect 7084 9472 7124 9512
rect 7468 9472 7508 9512
rect 7852 9472 7892 9512
rect 8236 9472 8276 9512
rect 8620 9472 8660 9512
rect 9004 9472 9044 9512
rect 9388 9472 9428 9512
rect 9772 9472 9812 9512
rect 10156 9472 10196 9512
rect 10540 9472 10580 9512
rect 10924 9472 10964 9512
rect 11308 9472 11348 9512
rect 11692 9472 11732 9512
rect 12076 9472 12116 9512
rect 12460 9472 12500 9512
rect 12844 9472 12884 9512
rect 13228 9472 13268 9512
rect 13612 9472 13652 9512
rect 13996 9472 14036 9512
rect 14380 9472 14420 9512
rect 14764 9472 14804 9512
rect 15148 9472 15188 9512
rect 15532 9472 15572 9512
rect 15916 9472 15956 9512
rect 16156 9472 16196 9512
rect 16300 9472 16340 9512
rect 16876 9472 16916 9512
rect 17260 9472 17300 9512
rect 17644 9472 17684 9512
rect 18028 9472 18068 9512
rect 27820 9472 27860 9512
rect 28204 9472 28244 9512
rect 28588 9472 28628 9512
rect 28972 9472 29012 9512
rect 29356 9472 29396 9512
rect 29740 9472 29780 9512
rect 30124 9472 30164 9512
rect 30508 9472 30548 9512
rect 30892 9472 30932 9512
rect 31276 9472 31316 9512
rect 31660 9472 31700 9512
rect 32044 9472 32084 9512
rect 32428 9472 32468 9512
rect 35884 9472 35924 9512
rect 36268 9472 36308 9512
rect 36652 9472 36692 9512
rect 37036 9472 37076 9512
rect 37420 9472 37460 9512
rect 37804 9472 37844 9512
rect 29500 9304 29540 9344
rect 31420 9304 31460 9344
rect 37276 9304 37316 9344
rect 30268 9220 30308 9260
rect 37660 9220 37700 9260
rect 38044 9220 38084 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 7804 8884 7844 8924
rect 8188 8884 8228 8924
rect 8572 8884 8612 8924
rect 8956 8884 8996 8924
rect 9340 8884 9380 8924
rect 9724 8884 9764 8924
rect 10108 8884 10148 8924
rect 10492 8884 10532 8924
rect 10876 8884 10916 8924
rect 11260 8884 11300 8924
rect 11644 8884 11684 8924
rect 12028 8884 12068 8924
rect 12412 8884 12452 8924
rect 12796 8884 12836 8924
rect 13180 8884 13220 8924
rect 13564 8884 13604 8924
rect 13948 8884 13988 8924
rect 14332 8884 14372 8924
rect 14716 8884 14756 8924
rect 15100 8884 15140 8924
rect 15484 8884 15524 8924
rect 15868 8884 15908 8924
rect 16252 8884 16292 8924
rect 28540 8884 28580 8924
rect 28924 8884 28964 8924
rect 29308 8884 29348 8924
rect 29692 8884 29732 8924
rect 30076 8884 30116 8924
rect 30460 8884 30500 8924
rect 30844 8884 30884 8924
rect 31228 8884 31268 8924
rect 36892 8884 36932 8924
rect 37276 8884 37316 8924
rect 8044 8632 8084 8672
rect 8428 8632 8468 8672
rect 8812 8632 8852 8672
rect 9196 8632 9236 8672
rect 9580 8632 9620 8672
rect 9964 8632 10004 8672
rect 10348 8632 10388 8672
rect 10732 8632 10772 8672
rect 11116 8632 11156 8672
rect 11500 8632 11540 8672
rect 11884 8632 11924 8672
rect 12268 8632 12308 8672
rect 12652 8632 12692 8672
rect 13036 8632 13076 8672
rect 13420 8632 13460 8672
rect 13804 8632 13844 8672
rect 14188 8632 14228 8672
rect 14572 8632 14612 8672
rect 14956 8632 14996 8672
rect 15340 8632 15380 8672
rect 15724 8632 15764 8672
rect 16108 8632 16148 8672
rect 16492 8632 16532 8672
rect 28780 8632 28820 8672
rect 29164 8632 29204 8672
rect 29548 8632 29588 8672
rect 29932 8632 29972 8672
rect 30316 8632 30356 8672
rect 30700 8632 30740 8672
rect 31084 8632 31124 8672
rect 31468 8632 31508 8672
rect 32524 8632 32564 8672
rect 32764 8632 32804 8672
rect 36652 8632 36692 8672
rect 37036 8632 37076 8672
rect 37420 8632 37460 8672
rect 37804 8632 37844 8672
rect 37660 8464 37700 8504
rect 38044 8464 38084 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 29884 8128 29924 8168
rect 30652 8128 30692 8168
rect 32380 8128 32420 8168
rect 31420 8044 31460 8084
rect 19612 7960 19652 8000
rect 19852 7960 19892 8000
rect 20236 7960 20276 8000
rect 22156 7960 22196 8000
rect 23020 7960 23060 8000
rect 23932 7960 23972 8000
rect 24172 7960 24212 8000
rect 25516 7960 25556 8000
rect 26188 7960 26228 8000
rect 26764 7960 26804 8000
rect 27580 7960 27620 8000
rect 27820 7960 27860 8000
rect 29644 7960 29684 8000
rect 30028 7960 30068 8000
rect 30412 7960 30452 8000
rect 30796 7960 30836 8000
rect 31180 7960 31220 8000
rect 32140 7960 32180 8000
rect 37420 7960 37460 8000
rect 37804 7960 37844 8000
rect 19996 7792 20036 7832
rect 21916 7792 21956 7832
rect 26428 7792 26468 7832
rect 22780 7708 22820 7748
rect 25276 7708 25316 7748
rect 26524 7708 26564 7748
rect 30268 7708 30308 7748
rect 31036 7708 31076 7748
rect 37660 7708 37700 7748
rect 38044 7708 38084 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 19708 7372 19748 7412
rect 30268 7372 30308 7412
rect 18796 7120 18836 7160
rect 19180 7120 19220 7160
rect 19564 7120 19604 7160
rect 19948 7120 19988 7160
rect 20092 7120 20132 7160
rect 20332 7120 20372 7160
rect 20716 7120 20756 7160
rect 21388 7120 21428 7160
rect 25612 7120 25652 7160
rect 29644 7120 29684 7160
rect 30028 7120 30068 7160
rect 31084 7120 31124 7160
rect 31324 7120 31364 7160
rect 37420 7120 37460 7160
rect 37804 7120 37844 7160
rect 18940 7036 18980 7076
rect 29884 7036 29924 7076
rect 18556 6952 18596 6992
rect 19324 6952 19364 6992
rect 20476 6952 20516 6992
rect 21148 6952 21188 6992
rect 25852 6952 25892 6992
rect 37660 6952 37700 6992
rect 38044 6952 38084 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 16732 6616 16772 6656
rect 19804 6616 19844 6656
rect 29692 6616 29732 6656
rect 30076 6616 30116 6656
rect 31900 6616 31940 6656
rect 16972 6448 17012 6488
rect 20044 6448 20084 6488
rect 29452 6448 29492 6488
rect 29836 6448 29876 6488
rect 31660 6448 31700 6488
rect 37420 6448 37460 6488
rect 37804 6448 37844 6488
rect 38044 6280 38084 6320
rect 37660 6196 37700 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 6844 5860 6884 5900
rect 15004 5860 15044 5900
rect 16924 5776 16964 5816
rect 5452 5608 5492 5648
rect 5836 5608 5876 5648
rect 6220 5608 6260 5648
rect 6604 5608 6644 5648
rect 6988 5608 7028 5648
rect 7228 5608 7268 5648
rect 15244 5608 15284 5648
rect 15388 5608 15428 5648
rect 15628 5608 15668 5648
rect 16012 5608 16052 5648
rect 16396 5608 16436 5648
rect 16780 5608 16820 5648
rect 17164 5608 17204 5648
rect 17548 5608 17588 5648
rect 17692 5608 17732 5648
rect 17932 5608 17972 5648
rect 29068 5608 29108 5648
rect 29308 5608 29348 5648
rect 37420 5608 37460 5648
rect 37804 5608 37844 5648
rect 38044 5608 38084 5648
rect 5692 5524 5732 5564
rect 6460 5524 6500 5564
rect 15772 5524 15812 5564
rect 17308 5524 17348 5564
rect 6076 5440 6116 5480
rect 16156 5440 16196 5480
rect 16540 5440 16580 5480
rect 37660 5440 37700 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 6076 5104 6116 5144
rect 7132 5104 7172 5144
rect 7516 5104 7556 5144
rect 8284 5104 8324 5144
rect 9052 5104 9092 5144
rect 9436 5104 9476 5144
rect 11740 5104 11780 5144
rect 12508 5104 12548 5144
rect 14524 5104 14564 5144
rect 29212 5104 29252 5144
rect 7900 5020 7940 5060
rect 8668 5020 8708 5060
rect 13660 5020 13700 5060
rect 17116 5020 17156 5060
rect 5836 4936 5876 4976
rect 6892 4936 6932 4976
rect 7276 4936 7316 4976
rect 7660 4936 7700 4976
rect 8044 4936 8084 4976
rect 8428 4936 8468 4976
rect 8812 4936 8852 4976
rect 9196 4936 9236 4976
rect 11980 4936 12020 4976
rect 12124 4936 12164 4976
rect 12364 4936 12404 4976
rect 12748 4936 12788 4976
rect 13132 4936 13172 4976
rect 13516 4936 13556 4976
rect 13900 4936 13940 4976
rect 14764 4936 14804 4976
rect 16972 4936 17012 4976
rect 17356 4936 17396 4976
rect 23980 4936 24020 4976
rect 28972 4936 29012 4976
rect 37420 4936 37460 4976
rect 37804 4936 37844 4976
rect 38044 4936 38084 4976
rect 12892 4768 12932 4808
rect 16732 4768 16772 4808
rect 13276 4684 13316 4724
rect 24220 4684 24260 4724
rect 37660 4684 37700 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 3484 4264 3524 4304
rect 8476 4264 8516 4304
rect 9628 4264 9668 4304
rect 11644 4264 11684 4304
rect 24604 4264 24644 4304
rect 29404 4264 29444 4304
rect 38044 4264 38084 4304
rect 3244 4096 3284 4136
rect 3916 4096 3956 4136
rect 8236 4096 8276 4136
rect 9388 4096 9428 4136
rect 10060 4096 10100 4136
rect 10684 4096 10724 4136
rect 10924 4096 10964 4136
rect 11827 4096 11867 4136
rect 24364 4096 24404 4136
rect 29164 4096 29204 4136
rect 37420 4096 37460 4136
rect 37804 4096 37844 4136
rect 4156 4012 4196 4052
rect 37660 4012 37700 4052
rect 10300 3928 10340 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 22588 3592 22628 3632
rect 28828 3592 28868 3632
rect 38044 3592 38084 3632
rect 21820 3508 21860 3548
rect 26524 3508 26564 3548
rect 5356 3424 5396 3464
rect 15628 3424 15668 3464
rect 18508 3424 18548 3464
rect 18892 3424 18932 3464
rect 19564 3424 19604 3464
rect 19948 3424 19988 3464
rect 20332 3424 20372 3464
rect 20716 3424 20756 3464
rect 20956 3424 20996 3464
rect 21196 3424 21236 3464
rect 21436 3424 21476 3464
rect 21580 3424 21620 3464
rect 22348 3424 22388 3464
rect 26284 3424 26324 3464
rect 28588 3424 28628 3464
rect 37420 3424 37460 3464
rect 37804 3424 37844 3464
rect 19132 3256 19172 3296
rect 20188 3256 20228 3296
rect 37660 3256 37700 3296
rect 5596 3172 5636 3212
rect 15868 3172 15908 3212
rect 18748 3172 18788 3212
rect 19804 3172 19844 3212
rect 20572 3172 20612 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 8188 2836 8228 2876
rect 8572 2836 8612 2876
rect 14620 2836 14660 2876
rect 15676 2836 15716 2876
rect 17596 2836 17636 2876
rect 21436 2836 21476 2876
rect 27292 2836 27332 2876
rect 29308 2836 29348 2876
rect 30748 2836 30788 2876
rect 38044 2836 38084 2876
rect 25468 2752 25508 2792
rect 25852 2752 25892 2792
rect 28060 2752 28100 2792
rect 7948 2584 7988 2624
rect 8332 2584 8372 2624
rect 11500 2584 11540 2624
rect 13324 2584 13364 2624
rect 14380 2584 14420 2624
rect 14764 2584 14804 2624
rect 15436 2584 15476 2624
rect 15820 2584 15860 2624
rect 17356 2584 17396 2624
rect 21196 2584 21236 2624
rect 21580 2584 21620 2624
rect 25228 2584 25268 2624
rect 25612 2584 25652 2624
rect 27052 2584 27092 2624
rect 27436 2584 27476 2624
rect 27820 2584 27860 2624
rect 29548 2584 29588 2624
rect 30988 2584 31028 2624
rect 37036 2584 37076 2624
rect 37420 2584 37460 2624
rect 37804 2584 37844 2624
rect 15004 2500 15044 2540
rect 37660 2500 37700 2540
rect 11740 2416 11780 2456
rect 13564 2416 13604 2456
rect 16060 2416 16100 2456
rect 21820 2416 21860 2456
rect 27676 2416 27716 2456
rect 37276 2416 37316 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 38044 2080 38084 2120
rect 36268 1912 36308 1952
rect 36652 1912 36692 1952
rect 37036 1912 37076 1952
rect 37420 1912 37460 1952
rect 37804 1912 37844 1952
rect 36892 1744 36932 1784
rect 36508 1660 36548 1700
rect 37276 1660 37316 1700
rect 37660 1660 37700 1700
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
<< metal2 >>
rect 7852 11740 24268 11780
rect 24308 11740 24317 11780
rect 7852 11696 7892 11740
rect 7843 11656 7852 11696
rect 7892 11656 7901 11696
rect 8803 11656 8812 11696
rect 8852 11656 17740 11696
rect 17780 11656 17789 11696
rect 9187 11572 9196 11612
rect 9236 11572 17932 11612
rect 17972 11572 17981 11612
rect 0 11024 90 11044
rect 39174 11024 39264 11044
rect 0 10984 460 11024
rect 500 10984 509 11024
rect 37027 10984 37036 11024
rect 37076 10984 39264 11024
rect 0 10964 90 10984
rect 39174 10964 39264 10984
rect 14179 10816 14188 10856
rect 14228 10816 21196 10856
rect 21236 10816 21245 10856
rect 0 10688 90 10708
rect 39174 10688 39264 10708
rect 0 10648 652 10688
rect 692 10648 701 10688
rect 36163 10648 36172 10688
rect 36212 10648 39264 10688
rect 0 10628 90 10648
rect 39174 10628 39264 10648
rect 10531 10564 10540 10604
rect 10580 10564 18700 10604
rect 18740 10564 18749 10604
rect 0 10352 90 10372
rect 39174 10352 39264 10372
rect 0 10312 1324 10352
rect 1364 10312 1373 10352
rect 36547 10312 36556 10352
rect 36596 10312 39264 10352
rect 0 10292 90 10312
rect 39174 10292 39264 10312
rect 19267 10144 19276 10184
rect 19316 10144 19325 10184
rect 19276 10100 19316 10144
rect 13411 10060 13420 10100
rect 13460 10060 19316 10100
rect 0 10016 90 10036
rect 39174 10016 39264 10036
rect 0 9976 1036 10016
rect 1076 9976 1085 10016
rect 11875 9976 11884 10016
rect 11924 9976 23884 10016
rect 23924 9976 23933 10016
rect 29827 9976 29836 10016
rect 29876 9976 30124 10016
rect 30164 9976 30173 10016
rect 37315 9976 37324 10016
rect 37364 9976 39264 10016
rect 0 9956 90 9976
rect 39174 9956 39264 9976
rect 13987 9892 13996 9932
rect 14036 9892 19564 9932
rect 19604 9892 19613 9932
rect 28771 9892 28780 9932
rect 28820 9892 31316 9932
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 13219 9808 13228 9848
rect 13268 9808 17740 9848
rect 17780 9808 17789 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 28003 9808 28012 9848
rect 28052 9808 30068 9848
rect 12940 9724 13036 9764
rect 13076 9724 13085 9764
rect 16108 9724 17452 9764
rect 17492 9724 17501 9764
rect 28291 9724 28300 9764
rect 28340 9724 28724 9764
rect 0 9680 90 9700
rect 12940 9680 12980 9724
rect 0 9640 940 9680
rect 980 9640 989 9680
rect 7315 9640 7324 9680
rect 7364 9640 7564 9680
rect 7604 9640 7613 9680
rect 7699 9640 7708 9680
rect 7748 9640 7948 9680
rect 7988 9640 7997 9680
rect 8083 9640 8092 9680
rect 8132 9640 8332 9680
rect 8372 9640 8381 9680
rect 8467 9640 8476 9680
rect 8516 9640 8716 9680
rect 8756 9640 8765 9680
rect 8851 9640 8860 9680
rect 8900 9640 9100 9680
rect 9140 9640 9149 9680
rect 9235 9640 9244 9680
rect 9284 9640 9484 9680
rect 9524 9640 9533 9680
rect 9619 9640 9628 9680
rect 9668 9640 9868 9680
rect 9908 9640 9917 9680
rect 10003 9640 10012 9680
rect 10052 9640 10252 9680
rect 10292 9640 10301 9680
rect 10387 9640 10396 9680
rect 10436 9640 10636 9680
rect 10676 9640 10685 9680
rect 10771 9640 10780 9680
rect 10820 9640 11020 9680
rect 11060 9640 11069 9680
rect 11155 9640 11164 9680
rect 11204 9640 11404 9680
rect 11444 9640 11453 9680
rect 11539 9640 11548 9680
rect 11588 9640 11788 9680
rect 11828 9640 11837 9680
rect 11923 9640 11932 9680
rect 11972 9640 12172 9680
rect 12212 9640 12221 9680
rect 12307 9640 12316 9680
rect 12356 9640 12556 9680
rect 12596 9640 12605 9680
rect 12691 9640 12700 9680
rect 12740 9640 12980 9680
rect 13075 9640 13084 9680
rect 13124 9640 13324 9680
rect 13364 9640 13373 9680
rect 13459 9640 13468 9680
rect 13508 9640 13708 9680
rect 13748 9640 13757 9680
rect 13843 9640 13852 9680
rect 13892 9640 14092 9680
rect 14132 9640 14141 9680
rect 14227 9640 14236 9680
rect 14276 9640 14476 9680
rect 14516 9640 14525 9680
rect 14611 9640 14620 9680
rect 14660 9640 14860 9680
rect 14900 9640 14909 9680
rect 14995 9640 15004 9680
rect 15044 9640 15244 9680
rect 15284 9640 15293 9680
rect 15379 9640 15388 9680
rect 15428 9640 15628 9680
rect 15668 9640 15677 9680
rect 15763 9640 15772 9680
rect 15812 9640 16012 9680
rect 16052 9640 16061 9680
rect 0 9620 90 9640
rect 16108 9596 16148 9724
rect 28684 9680 28724 9724
rect 16457 9640 16540 9680
rect 16580 9640 16588 9680
rect 16628 9640 16637 9680
rect 16963 9640 16972 9680
rect 17012 9640 17020 9680
rect 17060 9640 17143 9680
rect 17347 9640 17356 9680
rect 17396 9640 17404 9680
rect 17444 9640 17527 9680
rect 18883 9640 18892 9680
rect 18932 9640 19660 9680
rect 19700 9640 19709 9680
rect 27523 9640 27532 9680
rect 27572 9640 27580 9680
rect 27620 9640 27703 9680
rect 27907 9640 27916 9680
rect 27956 9640 28348 9680
rect 28388 9640 28397 9680
rect 28684 9640 29116 9680
rect 29156 9640 29165 9680
rect 30028 9596 30068 9808
rect 30211 9724 30220 9764
rect 30260 9724 30836 9764
rect 30796 9680 30836 9724
rect 30115 9640 30124 9680
rect 30164 9640 30652 9680
rect 30692 9640 30701 9680
rect 30796 9640 31036 9680
rect 31076 9640 31085 9680
rect 6115 9556 6124 9596
rect 6164 9556 7892 9596
rect 7852 9512 7892 9556
rect 10540 9556 11444 9596
rect 10540 9512 10580 9556
rect 5731 9472 5740 9512
rect 5780 9472 7084 9512
rect 7124 9472 7133 9512
rect 7337 9472 7468 9512
rect 7508 9472 7517 9512
rect 7843 9472 7852 9512
rect 7892 9472 7901 9512
rect 8227 9472 8236 9512
rect 8276 9472 8285 9512
rect 8489 9472 8620 9512
rect 8660 9472 8669 9512
rect 8873 9472 9004 9512
rect 9044 9472 9053 9512
rect 9379 9472 9388 9512
rect 9428 9472 9437 9512
rect 9763 9472 9772 9512
rect 9812 9472 9964 9512
rect 10004 9472 10013 9512
rect 10147 9472 10156 9512
rect 10196 9472 10327 9512
rect 10531 9472 10540 9512
rect 10580 9472 10589 9512
rect 10915 9472 10924 9512
rect 10964 9472 10973 9512
rect 11177 9472 11308 9512
rect 11348 9472 11357 9512
rect 8236 9428 8276 9472
rect 7171 9388 7180 9428
rect 7220 9388 8276 9428
rect 0 9344 90 9364
rect 9388 9344 9428 9472
rect 0 9304 1132 9344
rect 1172 9304 1181 9344
rect 7555 9304 7564 9344
rect 7604 9304 9428 9344
rect 0 9284 90 9304
rect 10924 9260 10964 9472
rect 11404 9428 11444 9556
rect 12940 9556 16148 9596
rect 16204 9556 16396 9596
rect 16436 9556 16445 9596
rect 16627 9556 16636 9596
rect 16676 9556 16780 9596
rect 16820 9556 16829 9596
rect 17155 9556 17164 9596
rect 17204 9556 17788 9596
rect 17828 9556 17837 9596
rect 27715 9556 27724 9596
rect 27764 9556 27964 9596
rect 28004 9556 28013 9596
rect 28099 9556 28108 9596
rect 28148 9556 28732 9596
rect 28772 9556 28781 9596
rect 29059 9556 29068 9596
rect 29108 9556 29884 9596
rect 29924 9556 29933 9596
rect 30028 9556 30548 9596
rect 12940 9512 12980 9556
rect 16204 9512 16244 9556
rect 30508 9512 30548 9556
rect 31276 9512 31316 9892
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 31459 9724 31468 9764
rect 31508 9724 32468 9764
rect 31363 9640 31372 9680
rect 31412 9640 32188 9680
rect 32228 9640 32237 9680
rect 31372 9556 31804 9596
rect 31844 9556 31853 9596
rect 11683 9472 11692 9512
rect 11732 9472 11741 9512
rect 11945 9472 12076 9512
rect 12116 9472 12125 9512
rect 12329 9472 12460 9512
rect 12500 9472 12509 9512
rect 12835 9472 12844 9512
rect 12884 9472 12980 9512
rect 13097 9472 13228 9512
rect 13268 9472 13277 9512
rect 13603 9472 13612 9512
rect 13652 9472 13708 9512
rect 13748 9472 13783 9512
rect 13987 9472 13996 9512
rect 14036 9472 14045 9512
rect 14371 9472 14380 9512
rect 14420 9472 14429 9512
rect 14755 9472 14764 9512
rect 14804 9472 14813 9512
rect 15017 9472 15148 9512
rect 15188 9472 15197 9512
rect 15401 9472 15532 9512
rect 15572 9472 15581 9512
rect 15785 9472 15916 9512
rect 15956 9472 15965 9512
rect 16147 9472 16156 9512
rect 16196 9472 16244 9512
rect 16291 9472 16300 9512
rect 16340 9472 16349 9512
rect 16867 9472 16876 9512
rect 16916 9472 16925 9512
rect 17129 9472 17260 9512
rect 17300 9472 17309 9512
rect 17513 9472 17644 9512
rect 17684 9472 17693 9512
rect 18019 9472 18028 9512
rect 18068 9472 18700 9512
rect 18740 9472 18749 9512
rect 27689 9472 27820 9512
rect 27860 9472 27869 9512
rect 28073 9472 28204 9512
rect 28244 9472 28253 9512
rect 28457 9472 28588 9512
rect 28628 9472 28637 9512
rect 28841 9472 28972 9512
rect 29012 9472 29021 9512
rect 29225 9472 29356 9512
rect 29396 9472 29405 9512
rect 29539 9472 29548 9512
rect 29588 9472 29740 9512
rect 29780 9472 29789 9512
rect 30115 9472 30124 9512
rect 30164 9472 30173 9512
rect 30499 9472 30508 9512
rect 30548 9472 30557 9512
rect 30883 9472 30892 9512
rect 30932 9472 30941 9512
rect 31267 9472 31276 9512
rect 31316 9472 31325 9512
rect 11692 9428 11732 9472
rect 11395 9388 11404 9428
rect 11444 9388 11453 9428
rect 11692 9388 12172 9428
rect 12212 9388 12221 9428
rect 8323 9220 8332 9260
rect 8372 9220 10964 9260
rect 13996 9092 14036 9472
rect 14380 9176 14420 9472
rect 14764 9260 14804 9472
rect 16300 9344 16340 9472
rect 16876 9428 16916 9472
rect 30124 9428 30164 9472
rect 30892 9428 30932 9472
rect 31372 9428 31412 9556
rect 32428 9512 32468 9724
rect 39174 9680 39264 9700
rect 36041 9640 36124 9680
rect 36164 9640 36172 9680
rect 36212 9640 36221 9680
rect 36425 9640 36508 9680
rect 36548 9640 36556 9680
rect 36596 9640 36605 9680
rect 36883 9640 36892 9680
rect 36932 9640 39264 9680
rect 39174 9620 39264 9640
rect 32611 9556 32620 9596
rect 32660 9556 37844 9596
rect 37804 9512 37844 9556
rect 31651 9472 31660 9512
rect 31700 9472 31709 9512
rect 32035 9472 32044 9512
rect 32084 9472 32093 9512
rect 32419 9472 32428 9512
rect 32468 9472 32477 9512
rect 35753 9472 35884 9512
rect 35924 9472 35933 9512
rect 36137 9472 36268 9512
rect 36308 9472 36317 9512
rect 36521 9472 36652 9512
rect 36692 9472 36701 9512
rect 37027 9472 37036 9512
rect 37076 9472 37085 9512
rect 37132 9472 37420 9512
rect 37460 9472 37469 9512
rect 37795 9472 37804 9512
rect 37844 9472 37853 9512
rect 16876 9388 19564 9428
rect 19604 9388 19613 9428
rect 29059 9388 29068 9428
rect 29108 9388 30164 9428
rect 30220 9388 30932 9428
rect 30979 9388 30988 9428
rect 31028 9388 31412 9428
rect 30220 9344 30260 9388
rect 16300 9304 19948 9344
rect 19988 9304 19997 9344
rect 28675 9304 28684 9344
rect 28724 9304 29500 9344
rect 29540 9304 29549 9344
rect 29731 9304 29740 9344
rect 29780 9304 30260 9344
rect 30595 9304 30604 9344
rect 30644 9304 31420 9344
rect 31460 9304 31469 9344
rect 14764 9220 19756 9260
rect 19796 9220 19805 9260
rect 29443 9220 29452 9260
rect 29492 9220 30268 9260
rect 30308 9220 30317 9260
rect 31660 9176 31700 9472
rect 14380 9136 24268 9176
rect 24308 9136 24317 9176
rect 30115 9136 30124 9176
rect 30164 9136 31700 9176
rect 32044 9092 32084 9472
rect 37036 9428 37076 9472
rect 33091 9388 33100 9428
rect 33140 9388 37076 9428
rect 37132 9344 37172 9472
rect 39174 9344 39264 9364
rect 32131 9304 32140 9344
rect 32180 9304 37172 9344
rect 37267 9304 37276 9344
rect 37316 9304 39264 9344
rect 39174 9284 39264 9304
rect 32227 9220 32236 9260
rect 32276 9220 36652 9260
rect 36692 9220 36701 9260
rect 37651 9220 37660 9260
rect 37700 9220 37709 9260
rect 38035 9220 38044 9260
rect 38084 9220 38668 9260
rect 38708 9220 38717 9260
rect 37660 9176 37700 9220
rect 37660 9136 39148 9176
rect 39188 9136 39197 9176
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 13996 9052 19124 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 29923 9052 29932 9092
rect 29972 9052 32084 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 0 9008 90 9028
rect 19084 9008 19124 9052
rect 39174 9008 39264 9028
rect 0 8968 1420 9008
rect 1460 8968 1469 9008
rect 14956 8968 19028 9008
rect 19084 8968 27244 9008
rect 27284 8968 27293 9008
rect 28963 8968 28972 9008
rect 29012 8968 29740 9008
rect 29780 8968 29789 9008
rect 30211 8968 30220 9008
rect 30260 8968 35884 9008
rect 35924 8968 35933 9008
rect 39139 8968 39148 9008
rect 39188 8968 39264 9008
rect 0 8948 90 8968
rect 7747 8884 7756 8924
rect 7796 8884 7804 8924
rect 7844 8884 7927 8924
rect 8131 8884 8140 8924
rect 8180 8884 8188 8924
rect 8228 8884 8311 8924
rect 8515 8884 8524 8924
rect 8564 8884 8572 8924
rect 8612 8884 8695 8924
rect 8899 8884 8908 8924
rect 8948 8884 8956 8924
rect 8996 8884 9079 8924
rect 9283 8884 9292 8924
rect 9332 8884 9340 8924
rect 9380 8884 9463 8924
rect 9667 8884 9676 8924
rect 9716 8884 9724 8924
rect 9764 8884 9847 8924
rect 10051 8884 10060 8924
rect 10100 8884 10108 8924
rect 10148 8884 10231 8924
rect 10435 8884 10444 8924
rect 10484 8884 10492 8924
rect 10532 8884 10615 8924
rect 10819 8884 10828 8924
rect 10868 8884 10876 8924
rect 10916 8884 10999 8924
rect 11203 8884 11212 8924
rect 11252 8884 11260 8924
rect 11300 8884 11383 8924
rect 11587 8884 11596 8924
rect 11636 8884 11644 8924
rect 11684 8884 11767 8924
rect 11971 8884 11980 8924
rect 12020 8884 12028 8924
rect 12068 8884 12151 8924
rect 12355 8884 12364 8924
rect 12404 8884 12412 8924
rect 12452 8884 12535 8924
rect 12739 8884 12748 8924
rect 12788 8884 12796 8924
rect 12836 8884 12919 8924
rect 13123 8884 13132 8924
rect 13172 8884 13180 8924
rect 13220 8884 13303 8924
rect 13507 8884 13516 8924
rect 13556 8884 13564 8924
rect 13604 8884 13687 8924
rect 13891 8884 13900 8924
rect 13940 8884 13948 8924
rect 13988 8884 14071 8924
rect 14275 8884 14284 8924
rect 14324 8884 14332 8924
rect 14372 8884 14455 8924
rect 14659 8884 14668 8924
rect 14708 8884 14716 8924
rect 14756 8884 14839 8924
rect 13027 8800 13036 8840
rect 13076 8800 14860 8840
rect 14900 8800 14909 8840
rect 6883 8716 6892 8756
rect 6932 8716 8468 8756
rect 8515 8716 8524 8756
rect 8564 8716 9236 8756
rect 9667 8716 9676 8756
rect 9716 8716 10388 8756
rect 10435 8716 10444 8756
rect 10484 8716 11924 8756
rect 0 8672 90 8692
rect 8428 8672 8468 8716
rect 9196 8672 9236 8716
rect 10348 8672 10388 8716
rect 11884 8672 11924 8716
rect 13036 8716 14380 8756
rect 14420 8716 14429 8756
rect 13036 8672 13076 8716
rect 14956 8672 14996 8968
rect 18988 8924 19028 8968
rect 39174 8948 39264 8968
rect 15043 8884 15052 8924
rect 15092 8884 15100 8924
rect 15140 8884 15223 8924
rect 15427 8884 15436 8924
rect 15476 8884 15484 8924
rect 15524 8884 15607 8924
rect 15811 8884 15820 8924
rect 15860 8884 15868 8924
rect 15908 8884 15991 8924
rect 16195 8884 16204 8924
rect 16244 8884 16252 8924
rect 16292 8884 16375 8924
rect 16483 8884 16492 8924
rect 16532 8884 18892 8924
rect 18932 8884 18941 8924
rect 18988 8884 24364 8924
rect 24404 8884 24413 8924
rect 28483 8884 28492 8924
rect 28532 8884 28540 8924
rect 28580 8884 28663 8924
rect 28867 8884 28876 8924
rect 28916 8884 28924 8924
rect 28964 8884 29047 8924
rect 29251 8884 29260 8924
rect 29300 8884 29308 8924
rect 29348 8884 29431 8924
rect 29635 8884 29644 8924
rect 29684 8884 29692 8924
rect 29732 8884 29815 8924
rect 30019 8884 30028 8924
rect 30068 8884 30076 8924
rect 30116 8884 30199 8924
rect 30403 8884 30412 8924
rect 30452 8884 30460 8924
rect 30500 8884 30583 8924
rect 30787 8884 30796 8924
rect 30836 8884 30844 8924
rect 30884 8884 30967 8924
rect 31171 8884 31180 8924
rect 31220 8884 31228 8924
rect 31268 8884 31351 8924
rect 36883 8884 36892 8924
rect 36932 8884 37036 8924
rect 37076 8884 37085 8924
rect 37193 8884 37276 8924
rect 37316 8884 37324 8924
rect 37364 8884 37373 8924
rect 15340 8800 23884 8840
rect 23924 8800 23933 8840
rect 29347 8800 29356 8840
rect 29396 8800 30740 8840
rect 31651 8800 31660 8840
rect 31700 8800 37076 8840
rect 15340 8672 15380 8800
rect 15724 8716 20140 8756
rect 20180 8716 20189 8756
rect 27427 8716 27436 8756
rect 27476 8716 29300 8756
rect 29443 8716 29452 8756
rect 29492 8716 30356 8756
rect 15724 8672 15764 8716
rect 29260 8672 29300 8716
rect 30316 8672 30356 8716
rect 30700 8672 30740 8800
rect 30787 8716 30796 8756
rect 30836 8716 31508 8756
rect 34531 8716 34540 8756
rect 34580 8716 36980 8756
rect 31468 8672 31508 8716
rect 0 8632 1228 8672
rect 1268 8632 1277 8672
rect 6499 8632 6508 8672
rect 6548 8632 8044 8672
rect 8084 8632 8093 8672
rect 8419 8632 8428 8672
rect 8468 8632 8477 8672
rect 8681 8632 8812 8672
rect 8852 8632 8861 8672
rect 9187 8632 9196 8672
rect 9236 8632 9245 8672
rect 9449 8632 9580 8672
rect 9620 8632 9629 8672
rect 9763 8632 9772 8672
rect 9812 8632 9964 8672
rect 10004 8632 10013 8672
rect 10339 8632 10348 8672
rect 10388 8632 10397 8672
rect 10601 8632 10732 8672
rect 10772 8632 10781 8672
rect 10985 8632 11116 8672
rect 11156 8632 11165 8672
rect 11369 8632 11500 8672
rect 11540 8632 11549 8672
rect 11875 8632 11884 8672
rect 11924 8632 11933 8672
rect 12259 8632 12268 8672
rect 12308 8632 12364 8672
rect 12404 8632 12439 8672
rect 12521 8632 12652 8672
rect 12692 8632 12701 8672
rect 13027 8632 13036 8672
rect 13076 8632 13085 8672
rect 13289 8632 13420 8672
rect 13460 8632 13469 8672
rect 13673 8632 13804 8672
rect 13844 8632 13853 8672
rect 14057 8632 14188 8672
rect 14228 8632 14237 8672
rect 14441 8632 14572 8672
rect 14612 8632 14621 8672
rect 14947 8632 14956 8672
rect 14996 8632 15005 8672
rect 15331 8632 15340 8672
rect 15380 8632 15389 8672
rect 15715 8632 15724 8672
rect 15764 8632 15773 8672
rect 15977 8632 16108 8672
rect 16148 8632 16157 8672
rect 16361 8632 16492 8672
rect 16532 8632 16541 8672
rect 25804 8632 26092 8672
rect 26132 8632 26141 8672
rect 27523 8632 27532 8672
rect 27572 8632 28780 8672
rect 28820 8632 28829 8672
rect 29033 8632 29164 8672
rect 29204 8632 29213 8672
rect 29260 8632 29548 8672
rect 29588 8632 29597 8672
rect 29644 8632 29932 8672
rect 29972 8632 29981 8672
rect 30307 8632 30316 8672
rect 30356 8632 30365 8672
rect 30691 8632 30700 8672
rect 30740 8632 30749 8672
rect 30796 8632 31084 8672
rect 31124 8632 31133 8672
rect 31459 8632 31468 8672
rect 31508 8632 31517 8672
rect 32393 8632 32524 8672
rect 32564 8632 32573 8672
rect 32755 8632 32764 8672
rect 32804 8632 36652 8672
rect 36692 8632 36701 8672
rect 0 8612 90 8632
rect 25804 8588 25844 8632
rect 29644 8588 29684 8632
rect 30796 8588 30836 8632
rect 1315 8548 1324 8588
rect 1364 8548 25844 8588
rect 25891 8548 25900 8588
rect 25940 8548 26956 8588
rect 26996 8548 27005 8588
rect 28867 8548 28876 8588
rect 28916 8548 29684 8588
rect 29731 8548 29740 8588
rect 29780 8548 30836 8588
rect 36940 8588 36980 8716
rect 37036 8672 37076 8800
rect 39174 8672 39264 8692
rect 37027 8632 37036 8672
rect 37076 8632 37085 8672
rect 37132 8632 37420 8672
rect 37460 8632 37469 8672
rect 37673 8632 37804 8672
rect 37844 8632 37853 8672
rect 38659 8632 38668 8672
rect 38708 8632 39264 8672
rect 37132 8588 37172 8632
rect 39174 8612 39264 8632
rect 36940 8548 37172 8588
rect 931 8464 940 8504
rect 980 8464 30028 8504
rect 30068 8464 30077 8504
rect 37651 8464 37660 8504
rect 37700 8464 37709 8504
rect 38035 8464 38044 8504
rect 38084 8464 38668 8504
rect 38708 8464 38717 8504
rect 643 8380 652 8420
rect 692 8380 29644 8420
rect 29684 8380 29693 8420
rect 0 8336 90 8356
rect 37660 8336 37700 8464
rect 39174 8336 39264 8356
rect 0 8296 1324 8336
rect 1364 8296 1373 8336
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 24163 8296 24172 8336
rect 24212 8296 26764 8336
rect 26804 8296 26813 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 37660 8296 39264 8336
rect 0 8276 90 8296
rect 39174 8276 39264 8296
rect 1027 8212 1036 8252
rect 1076 8212 25708 8252
rect 25748 8212 25757 8252
rect 1411 8128 1420 8168
rect 1460 8128 26380 8168
rect 26420 8128 26429 8168
rect 29875 8128 29884 8168
rect 29924 8128 30220 8168
rect 30260 8128 30269 8168
rect 30643 8128 30652 8168
rect 30692 8128 31660 8168
rect 31700 8128 31709 8168
rect 32371 8128 32380 8168
rect 32420 8128 33100 8168
rect 33140 8128 33149 8168
rect 1219 8044 1228 8084
rect 1268 8044 29300 8084
rect 31411 8044 31420 8084
rect 31460 8044 32620 8084
rect 32660 8044 32669 8084
rect 0 8000 90 8020
rect 0 7960 1420 8000
rect 1460 7960 1469 8000
rect 19555 7960 19564 8000
rect 19604 7960 19612 8000
rect 19652 7960 19735 8000
rect 19843 7960 19852 8000
rect 19892 7960 20023 8000
rect 20227 7960 20236 8000
rect 20276 7960 21676 8000
rect 21716 7960 21725 8000
rect 22147 7960 22156 8000
rect 22196 7960 22636 8000
rect 22676 7960 22685 8000
rect 22889 7960 22924 8000
rect 22964 7960 23020 8000
rect 23060 7960 23069 8000
rect 23801 7960 23884 8000
rect 23924 7960 23932 8000
rect 23972 7960 23981 8000
rect 24041 7960 24172 8000
rect 24212 7960 24221 8000
rect 25507 7960 25516 8000
rect 25556 7960 25900 8000
rect 25940 7960 25949 8000
rect 26057 7960 26092 8000
rect 26132 7960 26188 8000
rect 26228 7960 26237 8000
rect 26755 7960 26764 8000
rect 26804 7960 27148 8000
rect 27188 7960 27197 8000
rect 27331 7960 27340 8000
rect 27380 7960 27580 8000
rect 27620 7960 27629 8000
rect 27715 7960 27724 8000
rect 27764 7960 27820 8000
rect 27860 7960 27895 8000
rect 0 7940 90 7960
rect 29260 7916 29300 8044
rect 39174 8000 39264 8020
rect 29513 7960 29644 8000
rect 29684 7960 29693 8000
rect 29897 7960 30028 8000
rect 30068 7960 30077 8000
rect 30281 7960 30412 8000
rect 30452 7960 30461 8000
rect 30595 7960 30604 8000
rect 30644 7960 30796 8000
rect 30836 7960 30845 8000
rect 31171 7960 31180 8000
rect 31220 7960 31229 8000
rect 32131 7960 32140 8000
rect 32180 7960 32189 8000
rect 35971 7960 35980 8000
rect 36020 7960 37420 8000
rect 37460 7960 37469 8000
rect 37603 7960 37612 8000
rect 37652 7960 37804 8000
rect 37844 7960 37853 8000
rect 38659 7960 38668 8000
rect 38708 7960 39264 8000
rect 31180 7916 31220 7960
rect 1123 7876 1132 7916
rect 1172 7876 23060 7916
rect 19865 7792 19948 7832
rect 19988 7792 19996 7832
rect 20036 7792 20045 7832
rect 20131 7792 20140 7832
rect 20180 7792 21916 7832
rect 21956 7792 21965 7832
rect 23020 7748 23060 7876
rect 23884 7876 29204 7916
rect 29260 7876 31220 7916
rect 23884 7748 23924 7876
rect 29164 7832 29204 7876
rect 32140 7832 32180 7960
rect 39174 7940 39264 7960
rect 24355 7792 24364 7832
rect 24404 7792 25460 7832
rect 26419 7792 26428 7832
rect 26468 7792 27380 7832
rect 29164 7792 32180 7832
rect 25420 7748 25460 7792
rect 19747 7708 19756 7748
rect 19796 7708 22780 7748
rect 22820 7708 22829 7748
rect 23020 7708 23924 7748
rect 24259 7708 24268 7748
rect 24308 7708 25276 7748
rect 25316 7708 25325 7748
rect 25420 7708 26524 7748
rect 26564 7708 26573 7748
rect 0 7664 90 7684
rect 0 7624 1036 7664
rect 1076 7624 1085 7664
rect 0 7604 90 7624
rect 27340 7580 27380 7792
rect 30259 7708 30268 7748
rect 30308 7708 30932 7748
rect 31027 7708 31036 7748
rect 31076 7708 32140 7748
rect 32180 7708 32189 7748
rect 37651 7708 37660 7748
rect 37700 7708 37709 7748
rect 38035 7708 38044 7748
rect 38084 7708 38668 7748
rect 38708 7708 38717 7748
rect 30892 7664 30932 7708
rect 37660 7664 37700 7708
rect 39174 7664 39264 7684
rect 30892 7624 32236 7664
rect 32276 7624 32285 7664
rect 32332 7624 36268 7664
rect 36308 7624 36317 7664
rect 37660 7624 39264 7664
rect 32332 7580 32372 7624
rect 39174 7604 39264 7624
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 22627 7540 22636 7580
rect 22676 7540 26284 7580
rect 26324 7540 26333 7580
rect 27340 7540 32372 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 21667 7456 21676 7496
rect 21716 7456 25228 7496
rect 25268 7456 25277 7496
rect 18691 7372 18700 7412
rect 18740 7372 19708 7412
rect 19748 7372 19757 7412
rect 19843 7372 19852 7412
rect 19892 7372 25036 7412
rect 25076 7372 25085 7412
rect 30259 7372 30268 7412
rect 30308 7372 30796 7412
rect 30836 7372 30845 7412
rect 0 7328 90 7348
rect 39174 7328 39264 7348
rect 0 7288 844 7328
rect 884 7288 893 7328
rect 23011 7288 23020 7328
rect 23060 7288 26572 7328
rect 26612 7288 26621 7328
rect 38659 7288 38668 7328
rect 38708 7288 39264 7328
rect 0 7268 90 7288
rect 39174 7268 39264 7288
rect 18700 7204 20084 7244
rect 18700 7160 18740 7204
rect 20044 7160 20084 7204
rect 17635 7120 17644 7160
rect 17684 7120 18740 7160
rect 18787 7120 18796 7160
rect 18836 7120 18967 7160
rect 19171 7120 19180 7160
rect 19220 7120 19229 7160
rect 19555 7120 19564 7160
rect 19604 7120 19892 7160
rect 19939 7120 19948 7160
rect 19988 7120 19997 7160
rect 20044 7120 20092 7160
rect 20132 7120 20141 7160
rect 20323 7120 20332 7160
rect 20372 7120 20381 7160
rect 20707 7120 20716 7160
rect 20756 7120 21196 7160
rect 21236 7120 21245 7160
rect 21379 7120 21388 7160
rect 21428 7120 25556 7160
rect 25603 7120 25612 7160
rect 25652 7120 25783 7160
rect 29635 7120 29644 7160
rect 29684 7120 29693 7160
rect 30019 7120 30028 7160
rect 30068 7120 31028 7160
rect 31075 7120 31084 7160
rect 31124 7120 31255 7160
rect 31315 7120 31324 7160
rect 31364 7120 31372 7160
rect 31412 7120 31495 7160
rect 32707 7120 32716 7160
rect 32756 7120 37420 7160
rect 37460 7120 37469 7160
rect 37795 7120 37804 7160
rect 37844 7120 37853 7160
rect 19180 7076 19220 7120
rect 16483 7036 16492 7076
rect 16532 7036 18940 7076
rect 18980 7036 18989 7076
rect 19180 7036 19796 7076
rect 0 6992 90 7012
rect 0 6952 1132 6992
rect 1172 6952 1181 6992
rect 15907 6952 15916 6992
rect 15956 6952 18556 6992
rect 18596 6952 18605 6992
rect 18700 6952 19324 6992
rect 19364 6952 19373 6992
rect 0 6932 90 6952
rect 18700 6908 18740 6952
rect 15523 6868 15532 6908
rect 15572 6868 18740 6908
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 19756 6740 19796 7036
rect 19852 6824 19892 7120
rect 19948 6908 19988 7120
rect 20332 7076 20372 7120
rect 25516 7076 25556 7120
rect 20332 7036 24556 7076
rect 24596 7036 24605 7076
rect 25516 7036 26092 7076
rect 26132 7036 26141 7076
rect 20035 6952 20044 6992
rect 20084 6952 20476 6992
rect 20516 6952 20525 6992
rect 21017 6952 21100 6992
rect 21140 6952 21148 6992
rect 21188 6952 21197 6992
rect 21283 6952 21292 6992
rect 21332 6952 25748 6992
rect 25843 6952 25852 6992
rect 25892 6952 27380 6992
rect 25708 6908 25748 6952
rect 19948 6868 24652 6908
rect 24692 6868 24701 6908
rect 25708 6868 25996 6908
rect 26036 6868 26045 6908
rect 27340 6824 27380 6952
rect 29644 6908 29684 7120
rect 30988 7076 31028 7120
rect 37804 7076 37844 7120
rect 29801 7036 29884 7076
rect 29924 7036 29932 7076
rect 29972 7036 29981 7076
rect 30988 7036 34924 7076
rect 34964 7036 34973 7076
rect 36067 7036 36076 7076
rect 36116 7036 37844 7076
rect 39174 6992 39264 7012
rect 31075 6952 31084 6992
rect 31124 6952 36748 6992
rect 36788 6952 36797 6992
rect 37651 6952 37660 6992
rect 37700 6952 37940 6992
rect 38035 6952 38044 6992
rect 38084 6952 39264 6992
rect 29644 6868 33292 6908
rect 33332 6868 33341 6908
rect 33388 6868 34540 6908
rect 34580 6868 34589 6908
rect 33388 6824 33428 6868
rect 37900 6824 37940 6952
rect 39174 6932 39264 6952
rect 19852 6784 25708 6824
rect 25748 6784 25757 6824
rect 27340 6784 33428 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 37900 6784 39148 6824
rect 39188 6784 39197 6824
rect 19756 6700 23060 6740
rect 0 6656 90 6676
rect 23020 6656 23060 6700
rect 39174 6656 39264 6676
rect 0 6616 1228 6656
rect 1268 6616 1277 6656
rect 14563 6616 14572 6656
rect 14612 6616 16732 6656
rect 16772 6616 16781 6656
rect 17251 6616 17260 6656
rect 17300 6616 19804 6656
rect 19844 6616 19853 6656
rect 19948 6616 21388 6656
rect 21428 6616 21437 6656
rect 23020 6616 25516 6656
rect 25556 6616 25565 6656
rect 29609 6616 29692 6656
rect 29732 6616 29740 6656
rect 29780 6616 29789 6656
rect 30019 6616 30028 6656
rect 30068 6616 30076 6656
rect 30116 6616 30199 6656
rect 31891 6616 31900 6656
rect 31940 6616 37804 6656
rect 37844 6616 37853 6656
rect 39139 6616 39148 6656
rect 39188 6616 39264 6656
rect 0 6596 90 6616
rect 16099 6532 16108 6572
rect 16148 6532 19852 6572
rect 19892 6532 19901 6572
rect 19948 6488 19988 6616
rect 39174 6596 39264 6616
rect 20899 6532 20908 6572
rect 20948 6532 25420 6572
rect 25460 6532 25469 6572
rect 27340 6532 37460 6572
rect 16963 6448 16972 6488
rect 17012 6448 19988 6488
rect 20035 6448 20044 6488
rect 20084 6448 20215 6488
rect 21187 6448 21196 6488
rect 21236 6448 24844 6488
rect 24884 6448 24893 6488
rect 27340 6404 27380 6532
rect 37420 6488 37460 6532
rect 29443 6448 29452 6488
rect 29492 6448 29501 6488
rect 29705 6448 29836 6488
rect 29876 6448 29885 6488
rect 31651 6448 31660 6488
rect 31700 6448 31709 6488
rect 37411 6448 37420 6488
rect 37460 6448 37469 6488
rect 37795 6448 37804 6488
rect 37844 6448 37853 6488
rect 21475 6364 21484 6404
rect 21524 6364 27380 6404
rect 29452 6404 29492 6448
rect 29452 6364 31564 6404
rect 31604 6364 31613 6404
rect 0 6320 90 6340
rect 31660 6320 31700 6448
rect 37804 6404 37844 6448
rect 34531 6364 34540 6404
rect 34580 6364 37844 6404
rect 39174 6320 39264 6340
rect 0 6280 748 6320
rect 788 6280 797 6320
rect 1411 6280 1420 6320
rect 1460 6280 31700 6320
rect 38035 6280 38044 6320
rect 38084 6280 39264 6320
rect 0 6260 90 6280
rect 39174 6260 39264 6280
rect 15139 6196 15148 6236
rect 15188 6196 21100 6236
rect 21140 6196 21149 6236
rect 37651 6196 37660 6236
rect 37700 6196 38516 6236
rect 1315 6112 1324 6152
rect 1364 6112 25612 6152
rect 25652 6112 25661 6152
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 0 5984 90 6004
rect 38476 5984 38516 6196
rect 39174 5984 39264 6004
rect 0 5944 1420 5984
rect 1460 5944 1469 5984
rect 13507 5944 13516 5984
rect 13556 5944 23692 5984
rect 23732 5944 23741 5984
rect 38476 5944 39264 5984
rect 0 5924 90 5944
rect 39174 5924 39264 5944
rect 6761 5860 6844 5900
rect 6884 5860 6892 5900
rect 6932 5860 6941 5900
rect 13708 5860 15004 5900
rect 15044 5860 15053 5900
rect 6988 5776 8716 5816
rect 8756 5776 8765 5816
rect 12844 5776 13324 5816
rect 13364 5776 13373 5816
rect 2860 5692 6932 5732
rect 0 5648 90 5668
rect 2860 5648 2900 5692
rect 0 5608 2900 5648
rect 5443 5608 5452 5648
rect 5492 5608 5501 5648
rect 5827 5608 5836 5648
rect 5876 5608 5885 5648
rect 6211 5608 6220 5648
rect 6260 5608 6316 5648
rect 6356 5608 6391 5648
rect 6473 5608 6604 5648
rect 6644 5608 6653 5648
rect 0 5588 90 5608
rect 0 5312 90 5332
rect 5452 5312 5492 5608
rect 5609 5524 5692 5564
rect 5732 5524 5740 5564
rect 5780 5524 5789 5564
rect 5836 5396 5876 5608
rect 6892 5564 6932 5692
rect 6988 5648 7028 5776
rect 12844 5732 12884 5776
rect 7075 5692 7084 5732
rect 7124 5692 12884 5732
rect 12931 5692 12940 5732
rect 12980 5692 13612 5732
rect 13652 5692 13661 5732
rect 13708 5648 13748 5860
rect 14092 5776 16924 5816
rect 16964 5776 16973 5816
rect 14092 5732 14132 5776
rect 13795 5692 13804 5732
rect 13844 5692 14132 5732
rect 14284 5692 15428 5732
rect 6979 5608 6988 5648
rect 7028 5608 7037 5648
rect 7219 5608 7228 5648
rect 7268 5608 7468 5648
rect 7508 5608 7517 5648
rect 7564 5608 11788 5648
rect 11828 5608 11837 5648
rect 12067 5608 12076 5648
rect 12116 5608 12596 5648
rect 12643 5608 12652 5648
rect 12692 5608 13748 5648
rect 7564 5564 7604 5608
rect 12556 5564 12596 5608
rect 14284 5564 14324 5692
rect 15388 5648 15428 5692
rect 15628 5692 17356 5732
rect 17396 5692 17405 5732
rect 17548 5692 22348 5732
rect 22388 5692 22397 5732
rect 15628 5648 15668 5692
rect 17548 5648 17588 5692
rect 39174 5648 39264 5668
rect 15113 5608 15244 5648
rect 15284 5608 15293 5648
rect 15379 5608 15388 5648
rect 15428 5608 15437 5648
rect 15619 5608 15628 5648
rect 15668 5608 15677 5648
rect 15881 5608 16012 5648
rect 16052 5608 16061 5648
rect 16387 5608 16396 5648
rect 16436 5608 16445 5648
rect 16771 5608 16780 5648
rect 16820 5608 17108 5648
rect 17155 5608 17164 5648
rect 17204 5608 17213 5648
rect 17539 5608 17548 5648
rect 17588 5608 17597 5648
rect 17683 5608 17692 5648
rect 17732 5608 17740 5648
rect 17780 5608 17863 5648
rect 17923 5608 17932 5648
rect 17972 5608 21964 5648
rect 22004 5608 22013 5648
rect 28099 5608 28108 5648
rect 28148 5608 29068 5648
rect 29108 5608 29117 5648
rect 29251 5608 29260 5648
rect 29300 5608 29308 5648
rect 29348 5608 29431 5648
rect 37289 5608 37420 5648
rect 37460 5608 37469 5648
rect 37795 5608 37804 5648
rect 37844 5608 37853 5648
rect 38035 5608 38044 5648
rect 38084 5608 39264 5648
rect 16396 5564 16436 5608
rect 6377 5524 6460 5564
rect 6500 5524 6508 5564
rect 6548 5524 6557 5564
rect 6892 5524 7604 5564
rect 8419 5524 8428 5564
rect 8468 5524 12268 5564
rect 12308 5524 12317 5564
rect 12556 5524 14324 5564
rect 14380 5524 15772 5564
rect 15812 5524 15821 5564
rect 16396 5524 17012 5564
rect 14380 5480 14420 5524
rect 6067 5440 6076 5480
rect 6116 5440 8812 5480
rect 8852 5440 8861 5480
rect 12451 5440 12460 5480
rect 12500 5440 14420 5480
rect 15148 5440 16156 5480
rect 16196 5440 16205 5480
rect 16300 5440 16540 5480
rect 16580 5440 16589 5480
rect 15148 5396 15188 5440
rect 5836 5356 13996 5396
rect 14036 5356 14045 5396
rect 14179 5356 14188 5396
rect 14228 5356 15188 5396
rect 16300 5312 16340 5440
rect 0 5272 1652 5312
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 5452 5272 6988 5312
rect 7028 5272 7037 5312
rect 7276 5272 12940 5312
rect 12980 5272 12989 5312
rect 13411 5272 13420 5312
rect 13460 5272 16340 5312
rect 0 5252 90 5272
rect 1612 5228 1652 5272
rect 1612 5188 6836 5228
rect 5993 5104 6076 5144
rect 6116 5104 6124 5144
rect 6164 5104 6173 5144
rect 2860 5020 5972 5060
rect 0 4976 90 4996
rect 2860 4976 2900 5020
rect 0 4936 2900 4976
rect 5827 4936 5836 4976
rect 5876 4936 5885 4976
rect 0 4916 90 4936
rect 0 4640 90 4660
rect 0 4600 268 4640
rect 308 4600 317 4640
rect 0 4580 90 4600
rect 5836 4556 5876 4936
rect 5932 4640 5972 5020
rect 6796 4724 6836 5188
rect 7049 5104 7132 5144
rect 7172 5104 7180 5144
rect 7220 5104 7229 5144
rect 7276 4976 7316 5272
rect 16972 5228 17012 5524
rect 17068 5396 17108 5608
rect 17164 5480 17204 5608
rect 37804 5564 37844 5608
rect 39174 5588 39264 5608
rect 17299 5524 17308 5564
rect 17348 5524 17452 5564
rect 17492 5524 17501 5564
rect 17596 5524 22156 5564
rect 22196 5524 22205 5564
rect 37420 5524 37844 5564
rect 17596 5480 17636 5524
rect 17164 5440 17636 5480
rect 18691 5440 18700 5480
rect 18740 5440 19564 5480
rect 19604 5440 19613 5480
rect 17068 5356 22540 5396
rect 22580 5356 22589 5396
rect 17059 5272 17068 5312
rect 17108 5272 18700 5312
rect 18740 5272 18749 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 7660 5188 10676 5228
rect 11491 5188 11500 5228
rect 11540 5188 12020 5228
rect 12163 5188 12172 5228
rect 12212 5188 13748 5228
rect 16972 5188 21772 5228
rect 21812 5188 21821 5228
rect 7433 5104 7516 5144
rect 7556 5104 7564 5144
rect 7604 5104 7613 5144
rect 7660 4976 7700 5188
rect 8275 5104 8284 5144
rect 8324 5104 8620 5144
rect 8660 5104 8669 5144
rect 8995 5104 9004 5144
rect 9044 5104 9052 5144
rect 9092 5104 9175 5144
rect 9427 5104 9436 5144
rect 9476 5104 9580 5144
rect 9620 5104 9629 5144
rect 10636 5060 10676 5188
rect 11980 5144 12020 5188
rect 13708 5144 13748 5188
rect 10723 5104 10732 5144
rect 10772 5104 11740 5144
rect 11780 5104 11789 5144
rect 11980 5104 12508 5144
rect 12548 5104 12557 5144
rect 13708 5104 14524 5144
rect 14564 5104 14573 5144
rect 16003 5104 16012 5144
rect 16052 5104 22732 5144
rect 22772 5104 22781 5144
rect 28771 5104 28780 5144
rect 28820 5104 29212 5144
rect 29252 5104 29261 5144
rect 37420 5060 37460 5524
rect 37651 5440 37660 5480
rect 37700 5440 38516 5480
rect 38476 5312 38516 5440
rect 39174 5312 39264 5332
rect 38476 5272 39264 5312
rect 39174 5252 39264 5272
rect 7891 5020 7900 5060
rect 7940 5020 8524 5060
rect 8564 5020 8573 5060
rect 8659 5020 8668 5060
rect 8708 5020 9772 5060
rect 9812 5020 9821 5060
rect 10060 5020 10540 5060
rect 10580 5020 10589 5060
rect 10636 5020 11692 5060
rect 11732 5020 11741 5060
rect 11980 5020 12844 5060
rect 12884 5020 12893 5060
rect 12940 5020 13268 5060
rect 13603 5020 13612 5060
rect 13652 5020 13660 5060
rect 13700 5020 13783 5060
rect 14371 5020 14380 5060
rect 14420 5020 17116 5060
rect 17156 5020 17165 5060
rect 17260 5020 21580 5060
rect 21620 5020 21629 5060
rect 32332 5020 37460 5060
rect 10060 4976 10100 5020
rect 11980 4976 12020 5020
rect 12940 4976 12980 5020
rect 6883 4936 6892 4976
rect 6932 4936 7084 4976
rect 7124 4936 7133 4976
rect 7267 4936 7276 4976
rect 7316 4936 7325 4976
rect 7651 4936 7660 4976
rect 7700 4936 7709 4976
rect 8035 4936 8044 4976
rect 8084 4936 8093 4976
rect 8297 4936 8428 4976
rect 8468 4936 8477 4976
rect 8681 4936 8812 4976
rect 8852 4936 8861 4976
rect 9187 4936 9196 4976
rect 9236 4936 10100 4976
rect 10147 4936 10156 4976
rect 10196 4936 11732 4976
rect 11971 4936 11980 4976
rect 12020 4936 12029 4976
rect 12076 4936 12124 4976
rect 12164 4936 12173 4976
rect 12355 4936 12364 4976
rect 12404 4936 12556 4976
rect 12596 4936 12605 4976
rect 12739 4936 12748 4976
rect 12788 4936 12980 4976
rect 13123 4936 13132 4976
rect 13172 4936 13181 4976
rect 8044 4892 8084 4936
rect 11692 4892 11732 4936
rect 12076 4892 12116 4936
rect 8044 4852 11596 4892
rect 11636 4852 11645 4892
rect 11692 4852 12116 4892
rect 13132 4808 13172 4936
rect 13228 4892 13268 5020
rect 17260 4976 17300 5020
rect 13385 4936 13516 4976
rect 13556 4936 13565 4976
rect 13769 4936 13900 4976
rect 13940 4936 13949 4976
rect 14755 4936 14764 4976
rect 14804 4936 15052 4976
rect 15092 4936 15101 4976
rect 15148 4936 16780 4976
rect 16820 4936 16829 4976
rect 16963 4936 16972 4976
rect 17012 4936 17300 4976
rect 17347 4936 17356 4976
rect 17396 4936 22828 4976
rect 22868 4936 22877 4976
rect 23849 4936 23980 4976
rect 24020 4936 24029 4976
rect 26371 4936 26380 4976
rect 26420 4936 28972 4976
rect 29012 4936 29021 4976
rect 15148 4892 15188 4936
rect 13228 4852 15188 4892
rect 15235 4852 15244 4892
rect 15284 4852 23308 4892
rect 23348 4852 23357 4892
rect 32332 4808 32372 5020
rect 39174 4976 39264 4996
rect 34819 4936 34828 4976
rect 34868 4936 37420 4976
rect 37460 4936 37469 4976
rect 37795 4936 37804 4976
rect 37844 4936 37853 4976
rect 38035 4936 38044 4976
rect 38084 4936 39264 4976
rect 37804 4892 37844 4936
rect 39174 4916 39264 4936
rect 37507 4852 37516 4892
rect 37556 4852 37844 4892
rect 6979 4768 6988 4808
rect 7028 4768 10348 4808
rect 10388 4768 10397 4808
rect 11107 4768 11116 4808
rect 11156 4768 12892 4808
rect 12932 4768 12941 4808
rect 13132 4768 13652 4808
rect 13699 4768 13708 4808
rect 13748 4768 16732 4808
rect 16772 4768 16781 4808
rect 17635 4768 17644 4808
rect 17684 4768 32372 4808
rect 13612 4724 13652 4768
rect 6796 4684 12268 4724
rect 12308 4684 12317 4724
rect 12451 4684 12460 4724
rect 12500 4684 13276 4724
rect 13316 4684 13325 4724
rect 13603 4684 13612 4724
rect 13652 4684 13661 4724
rect 13891 4684 13900 4724
rect 13940 4684 19660 4724
rect 19700 4684 19709 4724
rect 19852 4684 20716 4724
rect 20756 4684 20765 4724
rect 24211 4684 24220 4724
rect 24260 4684 35884 4724
rect 35924 4684 35933 4724
rect 37651 4684 37660 4724
rect 37700 4684 38516 4724
rect 19852 4640 19892 4684
rect 38476 4640 38516 4684
rect 39174 4640 39264 4660
rect 5932 4600 12076 4640
rect 12116 4600 12125 4640
rect 12547 4600 12556 4640
rect 12596 4600 13516 4640
rect 13556 4600 13565 4640
rect 14947 4600 14956 4640
rect 14996 4600 18508 4640
rect 18548 4600 18557 4640
rect 18691 4600 18700 4640
rect 18740 4600 19892 4640
rect 19948 4600 20620 4640
rect 20660 4600 20669 4640
rect 38476 4600 39264 4640
rect 19948 4556 19988 4600
rect 39174 4580 39264 4600
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 5836 4516 12844 4556
rect 12884 4516 12893 4556
rect 12940 4516 17548 4556
rect 17588 4516 17597 4556
rect 17731 4516 17740 4556
rect 17780 4516 19988 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 12940 4472 12980 4516
rect 6595 4432 6604 4472
rect 6644 4432 12980 4472
rect 15043 4432 15052 4472
rect 15092 4432 23500 4472
rect 23540 4432 23549 4472
rect 8803 4348 8812 4388
rect 8852 4348 13556 4388
rect 13603 4348 13612 4388
rect 13652 4348 20524 4388
rect 20564 4348 20573 4388
rect 0 4304 90 4324
rect 13516 4304 13556 4348
rect 39174 4304 39264 4324
rect 0 4264 2900 4304
rect 3401 4264 3484 4304
rect 3524 4264 3532 4304
rect 3572 4264 3581 4304
rect 8323 4264 8332 4304
rect 8372 4264 8476 4304
rect 8516 4264 8525 4304
rect 9545 4264 9628 4304
rect 9668 4264 9676 4304
rect 9716 4264 9725 4304
rect 9772 4264 11020 4304
rect 11060 4264 11069 4304
rect 11299 4264 11308 4304
rect 11348 4264 11644 4304
rect 11684 4264 11693 4304
rect 11788 4264 12980 4304
rect 13516 4264 14956 4304
rect 14996 4264 15005 4304
rect 17836 4264 24076 4304
rect 24116 4264 24125 4304
rect 24595 4264 24604 4304
rect 24644 4264 29204 4304
rect 29321 4264 29404 4304
rect 29444 4264 29452 4304
rect 29492 4264 29501 4304
rect 38035 4264 38044 4304
rect 38084 4264 39264 4304
rect 0 4244 90 4264
rect 2860 4220 2900 4264
rect 9772 4220 9812 4264
rect 11788 4220 11828 4264
rect 12940 4220 12980 4264
rect 17836 4220 17876 4264
rect 29164 4220 29204 4264
rect 39174 4244 39264 4264
rect 2860 4180 9812 4220
rect 10060 4180 11828 4220
rect 11971 4180 11980 4220
rect 12020 4180 12116 4220
rect 12940 4180 13324 4220
rect 13364 4180 13373 4220
rect 13507 4180 13516 4220
rect 13556 4180 17876 4220
rect 17923 4180 17932 4220
rect 17972 4180 24404 4220
rect 24451 4180 24460 4220
rect 24500 4180 28780 4220
rect 28820 4180 28829 4220
rect 29164 4180 37612 4220
rect 37652 4180 37661 4220
rect 10060 4136 10100 4180
rect 12076 4136 12116 4180
rect 24364 4136 24404 4180
rect 3235 4096 3244 4136
rect 3284 4096 3340 4136
rect 3380 4096 3415 4136
rect 3907 4096 3916 4136
rect 3956 4096 3965 4136
rect 7843 4096 7852 4136
rect 7892 4096 8236 4136
rect 8276 4096 8285 4136
rect 9257 4096 9388 4136
rect 9428 4096 9437 4136
rect 10051 4096 10060 4136
rect 10100 4096 10109 4136
rect 10243 4096 10252 4136
rect 10292 4096 10684 4136
rect 10724 4096 10733 4136
rect 10793 4096 10924 4136
rect 10964 4096 10973 4136
rect 11683 4096 11692 4136
rect 11732 4096 11827 4136
rect 11867 4096 11876 4136
rect 12076 4096 21580 4136
rect 21620 4096 21629 4136
rect 24355 4096 24364 4136
rect 24404 4096 24413 4136
rect 24643 4096 24652 4136
rect 24692 4096 28244 4136
rect 29155 4096 29164 4136
rect 29204 4096 29213 4136
rect 37219 4096 37228 4136
rect 37268 4096 37420 4136
rect 37460 4096 37469 4136
rect 37516 4096 37804 4136
rect 37844 4096 37853 4136
rect 3916 4052 3956 4096
rect 28204 4052 28244 4096
rect 29164 4052 29204 4096
rect 2179 4012 2188 4052
rect 2228 4012 3956 4052
rect 4147 4012 4156 4052
rect 4196 4012 11060 4052
rect 12067 4012 12076 4052
rect 12116 4012 19948 4052
rect 19988 4012 19997 4052
rect 20419 4012 20428 4052
rect 20468 4012 21004 4052
rect 21044 4012 21053 4052
rect 24556 4012 27820 4052
rect 27860 4012 27869 4052
rect 28204 4012 29204 4052
rect 0 3968 90 3988
rect 11020 3968 11060 4012
rect 24556 3968 24596 4012
rect 0 3928 2900 3968
rect 10291 3928 10300 3968
rect 10340 3928 10444 3968
rect 10484 3928 10493 3968
rect 11020 3928 24596 3968
rect 24652 3928 27148 3968
rect 27188 3928 27197 3968
rect 27340 3928 36076 3968
rect 36116 3928 36125 3968
rect 0 3908 90 3928
rect 2860 3884 2900 3928
rect 2860 3844 21196 3884
rect 21236 3844 21245 3884
rect 21292 3844 24460 3884
rect 24500 3844 24509 3884
rect 21292 3800 21332 3844
rect 24652 3800 24692 3928
rect 27340 3884 27380 3928
rect 26755 3844 26764 3884
rect 26804 3844 27380 3884
rect 28771 3844 28780 3884
rect 28820 3844 37324 3884
rect 37364 3844 37373 3884
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 10915 3760 10924 3800
rect 10964 3760 18700 3800
rect 18740 3760 18749 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 19363 3760 19372 3800
rect 19412 3760 21332 3800
rect 21388 3760 22540 3800
rect 22580 3760 22589 3800
rect 22915 3760 22924 3800
rect 22964 3760 24692 3800
rect 27043 3760 27052 3800
rect 27092 3760 32716 3800
rect 32756 3760 32765 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 1219 3676 1228 3716
rect 1268 3676 2900 3716
rect 5443 3676 5452 3716
rect 5492 3676 20852 3716
rect 0 3632 90 3652
rect 2860 3632 2900 3676
rect 20812 3632 20852 3676
rect 21388 3632 21428 3760
rect 21667 3676 21676 3716
rect 21716 3676 28588 3716
rect 28628 3676 28637 3716
rect 28771 3676 28780 3716
rect 28820 3676 37420 3716
rect 37460 3676 37469 3716
rect 0 3592 76 3632
rect 116 3592 125 3632
rect 2860 3592 20756 3632
rect 20812 3592 21428 3632
rect 21484 3592 21716 3632
rect 22579 3592 22588 3632
rect 22628 3592 28724 3632
rect 28819 3592 28828 3632
rect 28868 3592 28972 3632
rect 29012 3592 29021 3632
rect 0 3572 90 3592
rect 259 3508 268 3548
rect 308 3508 20468 3548
rect 5347 3424 5356 3464
rect 5396 3424 5644 3464
rect 5684 3424 5693 3464
rect 5827 3424 5836 3464
rect 5876 3424 8660 3464
rect 12355 3424 12364 3464
rect 12404 3424 15628 3464
rect 15668 3424 15677 3464
rect 18377 3424 18508 3464
rect 18548 3424 18557 3464
rect 18761 3424 18892 3464
rect 18932 3424 18941 3464
rect 19267 3424 19276 3464
rect 19316 3424 19564 3464
rect 19604 3424 19613 3464
rect 19817 3424 19948 3464
rect 19988 3424 19997 3464
rect 20323 3424 20332 3464
rect 20372 3424 20381 3464
rect 8620 3380 8660 3424
rect 20332 3380 20372 3424
rect 8620 3340 20372 3380
rect 20428 3380 20468 3508
rect 20716 3464 20756 3592
rect 21484 3548 21524 3592
rect 20812 3508 21524 3548
rect 21571 3508 21580 3548
rect 21620 3508 21629 3548
rect 20707 3424 20716 3464
rect 20756 3424 20765 3464
rect 20812 3380 20852 3508
rect 21580 3464 21620 3508
rect 21676 3464 21716 3592
rect 21811 3508 21820 3548
rect 21860 3508 26420 3548
rect 26515 3508 26524 3548
rect 26564 3508 26764 3548
rect 26804 3508 26813 3548
rect 27052 3508 28588 3548
rect 28628 3508 28637 3548
rect 26380 3464 26420 3508
rect 27052 3464 27092 3508
rect 28684 3464 28724 3592
rect 37516 3548 37556 4096
rect 37651 4012 37660 4052
rect 37700 4012 38708 4052
rect 38668 3968 38708 4012
rect 39174 3968 39264 3988
rect 38668 3928 39264 3968
rect 39174 3908 39264 3928
rect 39174 3632 39264 3652
rect 38035 3592 38044 3632
rect 38084 3592 39264 3632
rect 39174 3572 39264 3592
rect 28771 3508 28780 3548
rect 28820 3508 37556 3548
rect 20947 3424 20956 3464
rect 20996 3424 21140 3464
rect 21187 3424 21196 3464
rect 21236 3424 21367 3464
rect 21427 3424 21436 3464
rect 21476 3424 21485 3464
rect 21533 3424 21580 3464
rect 21620 3424 21629 3464
rect 21676 3424 22348 3464
rect 22388 3424 22397 3464
rect 22531 3424 22540 3464
rect 22580 3424 26284 3464
rect 26324 3424 26333 3464
rect 26380 3424 27092 3464
rect 27139 3424 27148 3464
rect 27188 3424 28588 3464
rect 28628 3424 28637 3464
rect 28684 3424 34828 3464
rect 34868 3424 34877 3464
rect 35011 3424 35020 3464
rect 35060 3424 37420 3464
rect 37460 3424 37469 3464
rect 37795 3424 37804 3464
rect 37844 3424 37853 3464
rect 20428 3340 20852 3380
rect 0 3296 90 3316
rect 21100 3296 21140 3424
rect 21436 3380 21476 3424
rect 37804 3380 37844 3424
rect 21436 3340 22868 3380
rect 23011 3340 23020 3380
rect 23060 3340 37844 3380
rect 22828 3296 22868 3340
rect 39174 3296 39264 3316
rect 0 3256 5836 3296
rect 5876 3256 5885 3296
rect 14467 3256 14476 3296
rect 14516 3256 19028 3296
rect 19123 3256 19132 3296
rect 19172 3256 19372 3296
rect 19412 3256 19421 3296
rect 19660 3256 20084 3296
rect 20179 3256 20188 3296
rect 20228 3256 21004 3296
rect 21044 3256 21053 3296
rect 21100 3256 22004 3296
rect 22828 3256 37228 3296
rect 37268 3256 37277 3296
rect 37651 3256 37660 3296
rect 37700 3256 39264 3296
rect 0 3236 90 3256
rect 18988 3212 19028 3256
rect 19660 3212 19700 3256
rect 20044 3212 20084 3256
rect 21964 3212 22004 3256
rect 39174 3236 39264 3256
rect 1123 3172 1132 3212
rect 1172 3172 5452 3212
rect 5492 3172 5501 3212
rect 5587 3172 5596 3212
rect 5636 3172 5740 3212
rect 5780 3172 5789 3212
rect 8611 3172 8620 3212
rect 8660 3172 14284 3212
rect 14324 3172 14333 3212
rect 14380 3172 14660 3212
rect 15859 3172 15868 3212
rect 15908 3172 17740 3212
rect 17780 3172 17789 3212
rect 18739 3172 18748 3212
rect 18788 3172 18932 3212
rect 18988 3172 19700 3212
rect 19795 3172 19804 3212
rect 19844 3172 19948 3212
rect 19988 3172 19997 3212
rect 20044 3172 20428 3212
rect 20468 3172 20477 3212
rect 20563 3172 20572 3212
rect 20612 3172 21772 3212
rect 21812 3172 21821 3212
rect 21964 3172 27052 3212
rect 27092 3172 27101 3212
rect 37420 3172 37804 3212
rect 37844 3172 37853 3212
rect 14380 3128 14420 3172
rect 835 3088 844 3128
rect 884 3088 14420 3128
rect 14620 3128 14660 3172
rect 18892 3128 18932 3172
rect 37420 3128 37460 3172
rect 14620 3088 17932 3128
rect 17972 3088 17981 3128
rect 18892 3088 37460 3128
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 9379 3004 9388 3044
rect 9428 3004 14476 3044
rect 14516 3004 14525 3044
rect 14659 3004 14668 3044
rect 14708 3004 19852 3044
rect 19892 3004 19901 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 21763 3004 21772 3044
rect 21812 3004 35020 3044
rect 35060 3004 35069 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 0 2960 90 2980
rect 39174 2960 39264 2980
rect 0 2920 18508 2960
rect 18548 2920 18557 2960
rect 19939 2920 19948 2960
rect 19988 2920 37612 2960
rect 37652 2920 37661 2960
rect 38380 2920 39264 2960
rect 0 2900 90 2920
rect 38380 2876 38420 2920
rect 39174 2900 39264 2920
rect 1411 2836 1420 2876
rect 1460 2836 7220 2876
rect 8105 2836 8188 2876
rect 8228 2836 8236 2876
rect 8276 2836 8285 2876
rect 8419 2836 8428 2876
rect 8468 2836 8572 2876
rect 8612 2836 8621 2876
rect 14537 2836 14620 2876
rect 14660 2836 14668 2876
rect 14708 2836 14717 2876
rect 15593 2836 15676 2876
rect 15716 2836 15724 2876
rect 15764 2836 15773 2876
rect 17513 2836 17596 2876
rect 17636 2836 17644 2876
rect 17684 2836 17693 2876
rect 21353 2836 21436 2876
rect 21476 2836 21484 2876
rect 21524 2836 21533 2876
rect 23020 2836 25268 2876
rect 27283 2836 27292 2876
rect 27332 2836 28876 2876
rect 28916 2836 28925 2876
rect 29155 2836 29164 2876
rect 29204 2836 29308 2876
rect 29348 2836 29357 2876
rect 29539 2836 29548 2876
rect 29588 2836 30748 2876
rect 30788 2836 30797 2876
rect 38035 2836 38044 2876
rect 38084 2836 38420 2876
rect 7180 2792 7220 2836
rect 23020 2792 23060 2836
rect 7180 2752 11500 2792
rect 11540 2752 11549 2792
rect 13036 2752 18892 2792
rect 18932 2752 18941 2792
rect 19747 2752 19756 2792
rect 19796 2752 23060 2792
rect 13036 2708 13076 2752
rect 7948 2668 9100 2708
rect 9140 2668 9149 2708
rect 11404 2668 13076 2708
rect 15427 2668 15436 2708
rect 15476 2668 15523 2708
rect 0 2624 90 2644
rect 7948 2624 7988 2668
rect 0 2584 7220 2624
rect 7939 2584 7948 2624
rect 7988 2584 7997 2624
rect 8323 2584 8332 2624
rect 8372 2584 8381 2624
rect 0 2564 90 2584
rect 7180 2456 7220 2584
rect 8332 2540 8372 2584
rect 7363 2500 7372 2540
rect 7412 2500 8372 2540
rect 11404 2456 11444 2668
rect 15436 2624 15476 2668
rect 25228 2624 25268 2836
rect 25459 2752 25468 2792
rect 25508 2752 25748 2792
rect 25843 2752 25852 2792
rect 25892 2752 27436 2792
rect 27476 2752 27485 2792
rect 28051 2752 28060 2792
rect 28100 2752 29068 2792
rect 29108 2752 29117 2792
rect 25708 2708 25748 2752
rect 25708 2668 27628 2708
rect 27668 2668 27677 2708
rect 39174 2624 39264 2644
rect 11491 2584 11500 2624
rect 11540 2584 11671 2624
rect 13193 2584 13324 2624
rect 13364 2584 13373 2624
rect 14249 2584 14380 2624
rect 14420 2584 14429 2624
rect 14633 2584 14764 2624
rect 14804 2584 14813 2624
rect 15427 2584 15436 2624
rect 15476 2584 15485 2624
rect 15689 2584 15820 2624
rect 15860 2584 15869 2624
rect 17225 2584 17356 2624
rect 17396 2584 17405 2624
rect 17731 2584 17740 2624
rect 17780 2584 19660 2624
rect 19700 2584 19709 2624
rect 21065 2584 21196 2624
rect 21236 2584 21245 2624
rect 21449 2584 21580 2624
rect 21620 2584 21629 2624
rect 25219 2584 25228 2624
rect 25268 2584 25277 2624
rect 25481 2584 25612 2624
rect 25652 2584 25661 2624
rect 26921 2584 27052 2624
rect 27092 2584 27101 2624
rect 27427 2584 27436 2624
rect 27476 2584 27607 2624
rect 27811 2584 27820 2624
rect 27860 2584 27991 2624
rect 29417 2584 29548 2624
rect 29588 2584 29597 2624
rect 30857 2584 30988 2624
rect 31028 2584 31037 2624
rect 37027 2584 37036 2624
rect 37076 2584 37085 2624
rect 37356 2584 37420 2624
rect 37460 2584 37516 2624
rect 37556 2584 37591 2624
rect 37673 2584 37804 2624
rect 37844 2584 37853 2624
rect 38668 2584 39264 2624
rect 7180 2416 11444 2456
rect 11596 2500 13460 2540
rect 14995 2500 15004 2540
rect 15044 2500 36652 2540
rect 36692 2500 36701 2540
rect 11596 2372 11636 2500
rect 11731 2416 11740 2456
rect 11780 2416 13228 2456
rect 13268 2416 13277 2456
rect 3532 2332 11636 2372
rect 0 2288 90 2308
rect 3532 2288 3572 2332
rect 13420 2288 13460 2500
rect 13555 2416 13564 2456
rect 13604 2416 15956 2456
rect 16051 2416 16060 2456
rect 16100 2416 19508 2456
rect 21811 2416 21820 2456
rect 21860 2416 27532 2456
rect 27572 2416 27581 2456
rect 27667 2416 27676 2456
rect 27716 2416 34540 2456
rect 34580 2416 34589 2456
rect 15916 2372 15956 2416
rect 15916 2332 19316 2372
rect 19276 2288 19316 2332
rect 0 2248 3572 2288
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 13420 2248 17492 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 19276 2248 19372 2288
rect 19412 2248 19421 2288
rect 0 2228 90 2248
rect 17452 2204 17492 2248
rect 19468 2204 19508 2416
rect 37036 2372 37076 2584
rect 38668 2540 38708 2584
rect 39174 2564 39264 2584
rect 37651 2500 37660 2540
rect 37700 2500 38708 2540
rect 37267 2416 37276 2456
rect 37316 2416 37940 2456
rect 19555 2332 19564 2372
rect 19604 2332 37076 2372
rect 19651 2248 19660 2288
rect 19700 2248 25804 2288
rect 25844 2248 25853 2288
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 11779 2164 11788 2204
rect 11828 2164 17356 2204
rect 17396 2164 17405 2204
rect 17452 2164 19276 2204
rect 19316 2164 19325 2204
rect 19468 2164 36308 2204
rect 12547 2080 12556 2120
rect 12596 2080 30988 2120
rect 31028 2080 31037 2120
rect 14275 1996 14284 2036
rect 14324 1996 29548 2036
rect 29588 1996 29597 2036
rect 0 1952 90 1972
rect 36268 1952 36308 2164
rect 36364 1996 37460 2036
rect 0 1912 13324 1952
rect 13364 1912 13373 1952
rect 17731 1912 17740 1952
rect 17780 1912 25612 1952
rect 25652 1912 25661 1952
rect 25795 1912 25804 1952
rect 25844 1912 36212 1952
rect 36259 1912 36268 1952
rect 36308 1912 36317 1952
rect 0 1892 90 1912
rect 36172 1868 36212 1912
rect 36364 1868 36404 1996
rect 37420 1952 37460 1996
rect 37900 1952 37940 2416
rect 39174 2288 39264 2308
rect 38668 2248 39264 2288
rect 38668 2120 38708 2248
rect 39174 2228 39264 2248
rect 38035 2080 38044 2120
rect 38084 2080 38708 2120
rect 39174 1952 39264 1972
rect 36521 1912 36652 1952
rect 36692 1912 36701 1952
rect 36748 1912 37036 1952
rect 37076 1912 37085 1952
rect 37411 1912 37420 1952
rect 37460 1912 37469 1952
rect 37603 1912 37612 1952
rect 37652 1912 37804 1952
rect 37844 1912 37853 1952
rect 37900 1912 39264 1952
rect 16003 1828 16012 1868
rect 16052 1828 27820 1868
rect 27860 1828 27869 1868
rect 36172 1828 36404 1868
rect 36748 1784 36788 1912
rect 39174 1892 39264 1912
rect 10819 1744 10828 1784
rect 10868 1744 21580 1784
rect 21620 1744 21629 1784
rect 27340 1744 36788 1784
rect 36883 1744 36892 1784
rect 36932 1744 37804 1784
rect 37844 1744 37853 1784
rect 27340 1700 27380 1744
rect 13219 1660 13228 1700
rect 13268 1660 27380 1700
rect 36499 1660 36508 1700
rect 36548 1660 37172 1700
rect 37267 1660 37276 1700
rect 37316 1660 37516 1700
rect 37556 1660 37565 1700
rect 37651 1660 37660 1700
rect 37700 1660 37940 1700
rect 0 1616 90 1636
rect 0 1576 12364 1616
rect 12404 1576 12413 1616
rect 12940 1576 20564 1616
rect 21187 1576 21196 1616
rect 21236 1576 27052 1616
rect 27092 1576 27101 1616
rect 0 1556 90 1576
rect 12940 1532 12980 1576
rect 20524 1532 20564 1576
rect 37132 1532 37172 1660
rect 37900 1616 37940 1660
rect 39174 1616 39264 1636
rect 37900 1576 39264 1616
rect 39174 1556 39264 1576
rect 739 1492 748 1532
rect 788 1492 4820 1532
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 5356 1492 12980 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 20524 1492 27436 1532
rect 27476 1492 27485 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 37132 1492 37460 1532
rect 4780 1448 4820 1492
rect 5356 1448 5396 1492
rect 4780 1408 5396 1448
rect 0 1280 90 1300
rect 37420 1280 37460 1492
rect 39174 1280 39264 1300
rect 0 1240 15820 1280
rect 15860 1240 15869 1280
rect 37420 1240 39264 1280
rect 0 1220 90 1240
rect 39174 1220 39264 1240
rect 0 944 90 964
rect 39174 944 39264 964
rect 0 904 14764 944
rect 14804 904 14813 944
rect 37795 904 37804 944
rect 37844 904 39264 944
rect 0 884 90 904
rect 39174 884 39264 904
rect 0 608 90 628
rect 39174 608 39264 628
rect 0 568 11500 608
rect 11540 568 11549 608
rect 37507 568 37516 608
rect 37556 568 39264 608
rect 0 548 90 568
rect 39174 548 39264 568
<< via2 >>
rect 24268 11740 24308 11780
rect 7852 11656 7892 11696
rect 8812 11656 8852 11696
rect 17740 11656 17780 11696
rect 9196 11572 9236 11612
rect 17932 11572 17972 11612
rect 460 10984 500 11024
rect 37036 10984 37076 11024
rect 14188 10816 14228 10856
rect 21196 10816 21236 10856
rect 652 10648 692 10688
rect 36172 10648 36212 10688
rect 10540 10564 10580 10604
rect 18700 10564 18740 10604
rect 1324 10312 1364 10352
rect 36556 10312 36596 10352
rect 19276 10144 19316 10184
rect 13420 10060 13460 10100
rect 1036 9976 1076 10016
rect 11884 9976 11924 10016
rect 23884 9976 23924 10016
rect 29836 9976 29876 10016
rect 30124 9976 30164 10016
rect 37324 9976 37364 10016
rect 13996 9892 14036 9932
rect 19564 9892 19604 9932
rect 28780 9892 28820 9932
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 13228 9808 13268 9848
rect 17740 9808 17780 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 28012 9808 28052 9848
rect 13036 9724 13076 9764
rect 17452 9724 17492 9764
rect 28300 9724 28340 9764
rect 940 9640 980 9680
rect 7564 9640 7604 9680
rect 7948 9640 7988 9680
rect 8332 9640 8372 9680
rect 8716 9640 8756 9680
rect 9100 9640 9140 9680
rect 9484 9640 9524 9680
rect 9868 9640 9908 9680
rect 10252 9640 10292 9680
rect 10636 9640 10676 9680
rect 11020 9640 11060 9680
rect 11404 9640 11444 9680
rect 11788 9640 11828 9680
rect 12172 9640 12212 9680
rect 12556 9640 12596 9680
rect 13324 9640 13364 9680
rect 13708 9640 13748 9680
rect 14092 9640 14132 9680
rect 14476 9640 14516 9680
rect 14860 9640 14900 9680
rect 15244 9640 15284 9680
rect 15628 9640 15668 9680
rect 16012 9640 16052 9680
rect 16588 9640 16628 9680
rect 16972 9640 17012 9680
rect 17356 9640 17396 9680
rect 18892 9640 18932 9680
rect 19660 9640 19700 9680
rect 27532 9640 27572 9680
rect 27916 9640 27956 9680
rect 30220 9724 30260 9764
rect 30124 9640 30164 9680
rect 6124 9556 6164 9596
rect 5740 9472 5780 9512
rect 7468 9472 7508 9512
rect 8620 9472 8660 9512
rect 9004 9472 9044 9512
rect 9964 9472 10004 9512
rect 10156 9472 10196 9512
rect 11308 9472 11348 9512
rect 7180 9388 7220 9428
rect 1132 9304 1172 9344
rect 7564 9304 7604 9344
rect 16396 9556 16436 9596
rect 16780 9556 16820 9596
rect 17164 9556 17204 9596
rect 27724 9556 27764 9596
rect 28108 9556 28148 9596
rect 29068 9556 29108 9596
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 31468 9724 31508 9764
rect 31372 9640 31412 9680
rect 12076 9472 12116 9512
rect 12460 9472 12500 9512
rect 13228 9472 13268 9512
rect 13708 9472 13748 9512
rect 15148 9472 15188 9512
rect 15532 9472 15572 9512
rect 15916 9472 15956 9512
rect 17260 9472 17300 9512
rect 17644 9472 17684 9512
rect 18700 9472 18740 9512
rect 27820 9472 27860 9512
rect 28204 9472 28244 9512
rect 28588 9472 28628 9512
rect 28972 9472 29012 9512
rect 29356 9472 29396 9512
rect 29548 9472 29588 9512
rect 11404 9388 11444 9428
rect 12172 9388 12212 9428
rect 8332 9220 8372 9260
rect 36172 9640 36212 9680
rect 36556 9640 36596 9680
rect 32620 9556 32660 9596
rect 35884 9472 35924 9512
rect 36268 9472 36308 9512
rect 36652 9472 36692 9512
rect 19564 9388 19604 9428
rect 29068 9388 29108 9428
rect 30988 9388 31028 9428
rect 19948 9304 19988 9344
rect 28684 9304 28724 9344
rect 29740 9304 29780 9344
rect 30604 9304 30644 9344
rect 19756 9220 19796 9260
rect 29452 9220 29492 9260
rect 24268 9136 24308 9176
rect 30124 9136 30164 9176
rect 33100 9388 33140 9428
rect 32140 9304 32180 9344
rect 32236 9220 32276 9260
rect 36652 9220 36692 9260
rect 38668 9220 38708 9260
rect 39148 9136 39188 9176
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 29932 9052 29972 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 1420 8968 1460 9008
rect 27244 8968 27284 9008
rect 28972 8968 29012 9008
rect 29740 8968 29780 9008
rect 30220 8968 30260 9008
rect 35884 8968 35924 9008
rect 39148 8968 39188 9008
rect 7756 8884 7796 8924
rect 8140 8884 8180 8924
rect 8524 8884 8564 8924
rect 8908 8884 8948 8924
rect 9292 8884 9332 8924
rect 9676 8884 9716 8924
rect 10060 8884 10100 8924
rect 10444 8884 10484 8924
rect 10828 8884 10868 8924
rect 11212 8884 11252 8924
rect 11596 8884 11636 8924
rect 11980 8884 12020 8924
rect 12364 8884 12404 8924
rect 12748 8884 12788 8924
rect 13132 8884 13172 8924
rect 13516 8884 13556 8924
rect 13900 8884 13940 8924
rect 14284 8884 14324 8924
rect 14668 8884 14708 8924
rect 13036 8800 13076 8840
rect 14860 8800 14900 8840
rect 6892 8716 6932 8756
rect 8524 8716 8564 8756
rect 9676 8716 9716 8756
rect 10444 8716 10484 8756
rect 14380 8716 14420 8756
rect 15052 8884 15092 8924
rect 15436 8884 15476 8924
rect 15820 8884 15860 8924
rect 16204 8884 16244 8924
rect 16492 8884 16532 8924
rect 18892 8884 18932 8924
rect 24364 8884 24404 8924
rect 28492 8884 28532 8924
rect 28876 8884 28916 8924
rect 29260 8884 29300 8924
rect 29644 8884 29684 8924
rect 30028 8884 30068 8924
rect 30412 8884 30452 8924
rect 30796 8884 30836 8924
rect 31180 8884 31220 8924
rect 37036 8884 37076 8924
rect 37324 8884 37364 8924
rect 23884 8800 23924 8840
rect 29356 8800 29396 8840
rect 31660 8800 31700 8840
rect 20140 8716 20180 8756
rect 27436 8716 27476 8756
rect 29452 8716 29492 8756
rect 30796 8716 30836 8756
rect 34540 8716 34580 8756
rect 1228 8632 1268 8672
rect 6508 8632 6548 8672
rect 8812 8632 8852 8672
rect 9580 8632 9620 8672
rect 9772 8632 9812 8672
rect 10732 8632 10772 8672
rect 11116 8632 11156 8672
rect 11500 8632 11540 8672
rect 12364 8632 12404 8672
rect 12652 8632 12692 8672
rect 13420 8632 13460 8672
rect 13804 8632 13844 8672
rect 14188 8632 14228 8672
rect 14572 8632 14612 8672
rect 16108 8632 16148 8672
rect 16492 8632 16532 8672
rect 26092 8632 26132 8672
rect 27532 8632 27572 8672
rect 29164 8632 29204 8672
rect 32524 8632 32564 8672
rect 1324 8548 1364 8588
rect 25900 8548 25940 8588
rect 26956 8548 26996 8588
rect 28876 8548 28916 8588
rect 29740 8548 29780 8588
rect 37804 8632 37844 8672
rect 38668 8632 38708 8672
rect 940 8464 980 8504
rect 30028 8464 30068 8504
rect 38668 8464 38708 8504
rect 652 8380 692 8420
rect 29644 8380 29684 8420
rect 1324 8296 1364 8336
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 24172 8296 24212 8336
rect 26764 8296 26804 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 1036 8212 1076 8252
rect 25708 8212 25748 8252
rect 1420 8128 1460 8168
rect 26380 8128 26420 8168
rect 30220 8128 30260 8168
rect 31660 8128 31700 8168
rect 33100 8128 33140 8168
rect 1228 8044 1268 8084
rect 32620 8044 32660 8084
rect 1420 7960 1460 8000
rect 19564 7960 19604 8000
rect 19852 7960 19892 8000
rect 21676 7960 21716 8000
rect 22636 7960 22676 8000
rect 22924 7960 22964 8000
rect 23884 7960 23924 8000
rect 24172 7960 24212 8000
rect 25900 7960 25940 8000
rect 26092 7960 26132 8000
rect 27148 7960 27188 8000
rect 27340 7960 27380 8000
rect 27724 7960 27764 8000
rect 29644 7960 29684 8000
rect 30028 7960 30068 8000
rect 30412 7960 30452 8000
rect 30604 7960 30644 8000
rect 35980 7960 36020 8000
rect 37612 7960 37652 8000
rect 38668 7960 38708 8000
rect 1132 7876 1172 7916
rect 19948 7792 19988 7832
rect 20140 7792 20180 7832
rect 24364 7792 24404 7832
rect 19756 7708 19796 7748
rect 24268 7708 24308 7748
rect 1036 7624 1076 7664
rect 32140 7708 32180 7748
rect 38668 7708 38708 7748
rect 32236 7624 32276 7664
rect 36268 7624 36308 7664
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 22636 7540 22676 7580
rect 26284 7540 26324 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 21676 7456 21716 7496
rect 25228 7456 25268 7496
rect 18700 7372 18740 7412
rect 19852 7372 19892 7412
rect 25036 7372 25076 7412
rect 30796 7372 30836 7412
rect 844 7288 884 7328
rect 23020 7288 23060 7328
rect 26572 7288 26612 7328
rect 38668 7288 38708 7328
rect 17644 7120 17684 7160
rect 18796 7120 18836 7160
rect 21196 7120 21236 7160
rect 25612 7120 25652 7160
rect 31084 7120 31124 7160
rect 31372 7120 31412 7160
rect 32716 7120 32756 7160
rect 16492 7036 16532 7076
rect 1132 6952 1172 6992
rect 15916 6952 15956 6992
rect 15532 6868 15572 6908
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 24556 7036 24596 7076
rect 26092 7036 26132 7076
rect 20044 6952 20084 6992
rect 21100 6952 21140 6992
rect 21292 6952 21332 6992
rect 24652 6868 24692 6908
rect 25996 6868 26036 6908
rect 29932 7036 29972 7076
rect 34924 7036 34964 7076
rect 36076 7036 36116 7076
rect 31084 6952 31124 6992
rect 36748 6952 36788 6992
rect 33292 6868 33332 6908
rect 34540 6868 34580 6908
rect 25708 6784 25748 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 39148 6784 39188 6824
rect 1228 6616 1268 6656
rect 14572 6616 14612 6656
rect 17260 6616 17300 6656
rect 21388 6616 21428 6656
rect 25516 6616 25556 6656
rect 29740 6616 29780 6656
rect 30028 6616 30068 6656
rect 37804 6616 37844 6656
rect 39148 6616 39188 6656
rect 16108 6532 16148 6572
rect 19852 6532 19892 6572
rect 20908 6532 20948 6572
rect 25420 6532 25460 6572
rect 20044 6448 20084 6488
rect 21196 6448 21236 6488
rect 24844 6448 24884 6488
rect 29836 6448 29876 6488
rect 21484 6364 21524 6404
rect 31564 6364 31604 6404
rect 34540 6364 34580 6404
rect 748 6280 788 6320
rect 1420 6280 1460 6320
rect 15148 6196 15188 6236
rect 21100 6196 21140 6236
rect 1324 6112 1364 6152
rect 25612 6112 25652 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 1420 5944 1460 5984
rect 13516 5944 13556 5984
rect 23692 5944 23732 5984
rect 6892 5860 6932 5900
rect 8716 5776 8756 5816
rect 13324 5776 13364 5816
rect 6316 5608 6356 5648
rect 6604 5608 6644 5648
rect 5740 5524 5780 5564
rect 7084 5692 7124 5732
rect 12940 5692 12980 5732
rect 13612 5692 13652 5732
rect 13804 5692 13844 5732
rect 7468 5608 7508 5648
rect 11788 5608 11828 5648
rect 12076 5608 12116 5648
rect 12652 5608 12692 5648
rect 17356 5692 17396 5732
rect 22348 5692 22388 5732
rect 15244 5608 15284 5648
rect 16012 5608 16052 5648
rect 17740 5608 17780 5648
rect 21964 5608 22004 5648
rect 28108 5608 28148 5648
rect 29260 5608 29300 5648
rect 37420 5608 37460 5648
rect 6508 5524 6548 5564
rect 8428 5524 8468 5564
rect 12268 5524 12308 5564
rect 8812 5440 8852 5480
rect 12460 5440 12500 5480
rect 13996 5356 14036 5396
rect 14188 5356 14228 5396
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 6988 5272 7028 5312
rect 12940 5272 12980 5312
rect 13420 5272 13460 5312
rect 6124 5104 6164 5144
rect 268 4600 308 4640
rect 7180 5104 7220 5144
rect 17452 5524 17492 5564
rect 22156 5524 22196 5564
rect 18700 5440 18740 5480
rect 19564 5440 19604 5480
rect 22540 5356 22580 5396
rect 17068 5272 17108 5312
rect 18700 5272 18740 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 11500 5188 11540 5228
rect 12172 5188 12212 5228
rect 21772 5188 21812 5228
rect 7564 5104 7604 5144
rect 8620 5104 8660 5144
rect 9004 5104 9044 5144
rect 9580 5104 9620 5144
rect 10732 5104 10772 5144
rect 16012 5104 16052 5144
rect 22732 5104 22772 5144
rect 28780 5104 28820 5144
rect 8524 5020 8564 5060
rect 9772 5020 9812 5060
rect 10540 5020 10580 5060
rect 11692 5020 11732 5060
rect 12844 5020 12884 5060
rect 13612 5020 13652 5060
rect 14380 5020 14420 5060
rect 21580 5020 21620 5060
rect 7084 4936 7124 4976
rect 8428 4936 8468 4976
rect 8812 4936 8852 4976
rect 10156 4936 10196 4976
rect 12556 4936 12596 4976
rect 11596 4852 11636 4892
rect 13516 4936 13556 4976
rect 13900 4936 13940 4976
rect 15052 4936 15092 4976
rect 16780 4936 16820 4976
rect 22828 4936 22868 4976
rect 23980 4936 24020 4976
rect 26380 4936 26420 4976
rect 15244 4852 15284 4892
rect 23308 4852 23348 4892
rect 34828 4936 34868 4976
rect 37516 4852 37556 4892
rect 6988 4768 7028 4808
rect 10348 4768 10388 4808
rect 11116 4768 11156 4808
rect 13708 4768 13748 4808
rect 17644 4768 17684 4808
rect 12268 4684 12308 4724
rect 12460 4684 12500 4724
rect 13612 4684 13652 4724
rect 13900 4684 13940 4724
rect 19660 4684 19700 4724
rect 20716 4684 20756 4724
rect 35884 4684 35924 4724
rect 12076 4600 12116 4640
rect 12556 4600 12596 4640
rect 13516 4600 13556 4640
rect 14956 4600 14996 4640
rect 18508 4600 18548 4640
rect 18700 4600 18740 4640
rect 20620 4600 20660 4640
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 12844 4516 12884 4556
rect 17548 4516 17588 4556
rect 17740 4516 17780 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 6604 4432 6644 4472
rect 15052 4432 15092 4472
rect 23500 4432 23540 4472
rect 8812 4348 8852 4388
rect 13612 4348 13652 4388
rect 20524 4348 20564 4388
rect 3532 4264 3572 4304
rect 8332 4264 8372 4304
rect 9676 4264 9716 4304
rect 11020 4264 11060 4304
rect 11308 4264 11348 4304
rect 14956 4264 14996 4304
rect 24076 4264 24116 4304
rect 29452 4264 29492 4304
rect 11980 4180 12020 4220
rect 13324 4180 13364 4220
rect 13516 4180 13556 4220
rect 17932 4180 17972 4220
rect 24460 4180 24500 4220
rect 28780 4180 28820 4220
rect 37612 4180 37652 4220
rect 3340 4096 3380 4136
rect 7852 4096 7892 4136
rect 9388 4096 9428 4136
rect 10252 4096 10292 4136
rect 10924 4096 10964 4136
rect 11692 4096 11732 4136
rect 21580 4096 21620 4136
rect 24652 4096 24692 4136
rect 37228 4096 37268 4136
rect 2188 4012 2228 4052
rect 12076 4012 12116 4052
rect 19948 4012 19988 4052
rect 20428 4012 20468 4052
rect 21004 4012 21044 4052
rect 27820 4012 27860 4052
rect 10444 3928 10484 3968
rect 27148 3928 27188 3968
rect 36076 3928 36116 3968
rect 21196 3844 21236 3884
rect 24460 3844 24500 3884
rect 26764 3844 26804 3884
rect 28780 3844 28820 3884
rect 37324 3844 37364 3884
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 10924 3760 10964 3800
rect 18700 3760 18740 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 19372 3760 19412 3800
rect 22540 3760 22580 3800
rect 22924 3760 22964 3800
rect 27052 3760 27092 3800
rect 32716 3760 32756 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 1228 3676 1268 3716
rect 5452 3676 5492 3716
rect 21676 3676 21716 3716
rect 28588 3676 28628 3716
rect 28780 3676 28820 3716
rect 37420 3676 37460 3716
rect 76 3592 116 3632
rect 28972 3592 29012 3632
rect 268 3508 308 3548
rect 5644 3424 5684 3464
rect 5836 3424 5876 3464
rect 12364 3424 12404 3464
rect 18508 3424 18548 3464
rect 18892 3424 18932 3464
rect 19276 3424 19316 3464
rect 19948 3424 19988 3464
rect 21580 3508 21620 3548
rect 26764 3508 26804 3548
rect 28588 3508 28628 3548
rect 28780 3508 28820 3548
rect 21196 3424 21236 3464
rect 22540 3424 22580 3464
rect 27148 3424 27188 3464
rect 34828 3424 34868 3464
rect 35020 3424 35060 3464
rect 23020 3340 23060 3380
rect 5836 3256 5876 3296
rect 14476 3256 14516 3296
rect 19372 3256 19412 3296
rect 21004 3256 21044 3296
rect 37228 3256 37268 3296
rect 1132 3172 1172 3212
rect 5452 3172 5492 3212
rect 5740 3172 5780 3212
rect 8620 3172 8660 3212
rect 14284 3172 14324 3212
rect 17740 3172 17780 3212
rect 19948 3172 19988 3212
rect 20428 3172 20468 3212
rect 21772 3172 21812 3212
rect 27052 3172 27092 3212
rect 37804 3172 37844 3212
rect 844 3088 884 3128
rect 17932 3088 17972 3128
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 9388 3004 9428 3044
rect 14476 3004 14516 3044
rect 14668 3004 14708 3044
rect 19852 3004 19892 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 21772 3004 21812 3044
rect 35020 3004 35060 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 18508 2920 18548 2960
rect 19948 2920 19988 2960
rect 37612 2920 37652 2960
rect 1420 2836 1460 2876
rect 8236 2836 8276 2876
rect 8428 2836 8468 2876
rect 14668 2836 14708 2876
rect 15724 2836 15764 2876
rect 17644 2836 17684 2876
rect 21484 2836 21524 2876
rect 28876 2836 28916 2876
rect 29164 2836 29204 2876
rect 29548 2836 29588 2876
rect 11500 2752 11540 2792
rect 18892 2752 18932 2792
rect 19756 2752 19796 2792
rect 9100 2668 9140 2708
rect 15436 2668 15476 2708
rect 7372 2500 7412 2540
rect 27436 2752 27476 2792
rect 29068 2752 29108 2792
rect 27628 2668 27668 2708
rect 11500 2584 11540 2624
rect 13324 2584 13364 2624
rect 14380 2584 14420 2624
rect 14764 2584 14804 2624
rect 15820 2584 15860 2624
rect 17356 2584 17396 2624
rect 17740 2584 17780 2624
rect 19660 2584 19700 2624
rect 21196 2584 21236 2624
rect 21580 2584 21620 2624
rect 25612 2584 25652 2624
rect 27052 2584 27092 2624
rect 27436 2584 27476 2624
rect 27820 2584 27860 2624
rect 29548 2584 29588 2624
rect 30988 2584 31028 2624
rect 37516 2584 37556 2624
rect 37804 2584 37844 2624
rect 36652 2500 36692 2540
rect 13228 2416 13268 2456
rect 27532 2416 27572 2456
rect 34540 2416 34580 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 19372 2248 19412 2288
rect 19564 2332 19604 2372
rect 19660 2248 19700 2288
rect 25804 2248 25844 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 11788 2164 11828 2204
rect 17356 2164 17396 2204
rect 19276 2164 19316 2204
rect 12556 2080 12596 2120
rect 30988 2080 31028 2120
rect 14284 1996 14324 2036
rect 29548 1996 29588 2036
rect 13324 1912 13364 1952
rect 17740 1912 17780 1952
rect 25612 1912 25652 1952
rect 25804 1912 25844 1952
rect 36652 1912 36692 1952
rect 37612 1912 37652 1952
rect 16012 1828 16052 1868
rect 27820 1828 27860 1868
rect 10828 1744 10868 1784
rect 21580 1744 21620 1784
rect 37804 1744 37844 1784
rect 13228 1660 13268 1700
rect 37516 1660 37556 1700
rect 12364 1576 12404 1616
rect 21196 1576 21236 1616
rect 27052 1576 27092 1616
rect 748 1492 788 1532
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 27436 1492 27476 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 15820 1240 15860 1280
rect 14764 904 14804 944
rect 37804 904 37844 944
rect 11500 568 11540 608
rect 37516 568 37556 608
<< metal3 >>
rect 7544 11764 7624 11844
rect 7736 11764 7816 11844
rect 7928 11764 8008 11844
rect 8120 11764 8200 11844
rect 8312 11764 8392 11844
rect 8504 11764 8584 11844
rect 8696 11764 8776 11844
rect 8888 11764 8968 11844
rect 9080 11764 9160 11844
rect 9272 11764 9352 11844
rect 9464 11764 9544 11844
rect 9656 11764 9736 11844
rect 9848 11764 9928 11844
rect 10040 11764 10120 11844
rect 10232 11764 10312 11844
rect 10424 11764 10504 11844
rect 10616 11764 10696 11844
rect 10808 11764 10888 11844
rect 11000 11764 11080 11844
rect 11192 11764 11272 11844
rect 11384 11764 11464 11844
rect 11576 11764 11656 11844
rect 11768 11764 11848 11844
rect 11960 11764 12040 11844
rect 12152 11764 12232 11844
rect 12344 11764 12424 11844
rect 12536 11764 12616 11844
rect 12728 11764 12808 11844
rect 12920 11764 13000 11844
rect 13112 11764 13192 11844
rect 13304 11764 13384 11844
rect 13496 11764 13576 11844
rect 13688 11764 13768 11844
rect 13880 11764 13960 11844
rect 14072 11764 14152 11844
rect 14264 11764 14344 11844
rect 14456 11764 14536 11844
rect 14648 11764 14728 11844
rect 14840 11764 14920 11844
rect 15032 11764 15112 11844
rect 15224 11764 15304 11844
rect 15416 11764 15496 11844
rect 15608 11764 15688 11844
rect 15800 11764 15880 11844
rect 15992 11764 16072 11844
rect 16184 11764 16264 11844
rect 16376 11764 16456 11844
rect 16568 11764 16648 11844
rect 16760 11764 16840 11844
rect 16952 11764 17032 11844
rect 17144 11764 17224 11844
rect 17336 11764 17416 11844
rect 17528 11764 17608 11844
rect 17720 11764 17800 11844
rect 17912 11764 17992 11844
rect 18104 11764 18184 11844
rect 18296 11764 18376 11844
rect 18488 11764 18568 11844
rect 18680 11764 18760 11844
rect 18872 11764 18952 11844
rect 19064 11764 19144 11844
rect 19256 11764 19336 11844
rect 19448 11764 19528 11844
rect 19640 11764 19720 11844
rect 19832 11764 19912 11844
rect 20024 11764 20104 11844
rect 20216 11764 20296 11844
rect 20408 11764 20488 11844
rect 20600 11764 20680 11844
rect 20792 11764 20872 11844
rect 20984 11764 21064 11844
rect 21176 11764 21256 11844
rect 21368 11764 21448 11844
rect 21560 11764 21640 11844
rect 21752 11764 21832 11844
rect 21944 11764 22024 11844
rect 22136 11764 22216 11844
rect 22328 11764 22408 11844
rect 22520 11764 22600 11844
rect 22712 11764 22792 11844
rect 22904 11764 22984 11844
rect 23096 11764 23176 11844
rect 23288 11764 23368 11844
rect 23480 11764 23560 11844
rect 23672 11764 23752 11844
rect 23864 11764 23944 11844
rect 24056 11764 24136 11844
rect 24248 11780 24328 11844
rect 24248 11764 24268 11780
rect 460 11024 500 11033
rect 460 8672 500 10984
rect 460 8623 500 8632
rect 652 10688 692 10697
rect 652 8420 692 10648
rect 1324 10352 1364 10361
rect 1036 10016 1076 10025
rect 940 9680 980 9689
rect 940 8504 980 9640
rect 940 8455 980 8464
rect 652 8371 692 8380
rect 1036 8252 1076 9976
rect 1036 8203 1076 8212
rect 1132 9344 1172 9353
rect 1132 7916 1172 9304
rect 1228 8672 1268 8681
rect 1228 8084 1268 8632
rect 1324 8588 1364 10312
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 7564 9680 7604 11764
rect 7564 9631 7604 9640
rect 6124 9596 6164 9605
rect 3532 9512 3572 9521
rect 1324 8539 1364 8548
rect 1420 9008 1460 9017
rect 1228 8035 1268 8044
rect 1324 8336 1364 8345
rect 1132 7867 1172 7876
rect 1036 7664 1076 7673
rect 844 7328 884 7337
rect 748 6320 788 6329
rect 268 4640 308 4649
rect 76 3632 116 3641
rect 76 3212 116 3592
rect 268 3548 308 4600
rect 268 3499 308 3508
rect 76 3163 116 3172
rect 748 1532 788 6280
rect 844 3128 884 7288
rect 1036 4976 1076 7624
rect 1036 4927 1076 4936
rect 1132 6992 1172 7001
rect 1132 3212 1172 6952
rect 1228 6656 1268 6665
rect 1228 3716 1268 6616
rect 1324 6152 1364 8296
rect 1420 8168 1460 8968
rect 1420 8119 1460 8128
rect 1420 8000 1460 8009
rect 1420 6320 1460 7960
rect 1420 6271 1460 6280
rect 1324 6103 1364 6112
rect 1228 3667 1268 3676
rect 1420 5984 1460 5993
rect 1132 3163 1172 3172
rect 844 3079 884 3088
rect 1420 2876 1460 5944
rect 3532 4304 3572 9472
rect 5740 9512 5780 9521
rect 5644 9428 5684 9437
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 3532 4255 3572 4264
rect 3340 4136 3380 4145
rect 1420 2827 1460 2836
rect 2188 4052 2228 4061
rect 748 1483 788 1492
rect 2188 80 2228 4012
rect 2168 0 2248 80
rect 3340 60 3380 4096
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 5452 3716 5492 3725
rect 5452 3212 5492 3676
rect 5644 3632 5684 9388
rect 5740 5564 5780 9472
rect 5740 5515 5780 5524
rect 6124 5144 6164 9556
rect 7468 9512 7508 9521
rect 7180 9428 7220 9437
rect 6892 8756 6932 8765
rect 6508 8672 6548 8681
rect 6316 5648 6356 5657
rect 6316 5513 6356 5608
rect 6508 5564 6548 8632
rect 6892 5900 6932 8716
rect 6892 5851 6932 5860
rect 7084 5732 7124 5741
rect 6508 5515 6548 5524
rect 6604 5648 6644 5657
rect 6124 5095 6164 5104
rect 6604 4472 6644 5608
rect 6988 5312 7028 5321
rect 6988 4808 7028 5272
rect 7084 4976 7124 5692
rect 7180 5144 7220 9388
rect 7468 5648 7508 9472
rect 7468 5599 7508 5608
rect 7564 9344 7604 9353
rect 7180 5095 7220 5104
rect 7564 5144 7604 9304
rect 7756 8924 7796 11764
rect 7756 8875 7796 8884
rect 7852 11696 7892 11705
rect 7564 5095 7604 5104
rect 7084 4927 7124 4936
rect 6988 4759 7028 4768
rect 6604 4423 6644 4432
rect 7852 4136 7892 11656
rect 7948 9680 7988 11764
rect 7948 9631 7988 9640
rect 7852 4087 7892 4096
rect 8044 9260 8084 9269
rect 5644 3592 5780 3632
rect 5452 3163 5492 3172
rect 5644 3464 5684 3473
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 3688 2288 4056 2297
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 3688 2239 4056 2248
rect 4928 1532 5296 1541
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 4928 1483 5296 1492
rect 3724 148 3956 188
rect 3724 60 3764 148
rect 3916 80 3956 148
rect 5644 80 5684 3424
rect 5740 3212 5780 3592
rect 5836 3464 5876 3473
rect 5836 3296 5876 3424
rect 5836 3247 5876 3256
rect 5740 3163 5780 3172
rect 8044 2900 8084 9220
rect 8140 8924 8180 11764
rect 8332 9680 8372 11764
rect 8332 9631 8372 9640
rect 8140 8875 8180 8884
rect 8236 9344 8276 9353
rect 8236 4136 8276 9304
rect 8332 9260 8372 9269
rect 8332 4304 8372 9220
rect 8524 8924 8564 11764
rect 8716 9680 8756 11764
rect 8716 9631 8756 9640
rect 8812 11696 8852 11705
rect 8524 8875 8564 8884
rect 8620 9512 8660 9521
rect 8812 9512 8852 11656
rect 8524 8756 8564 8765
rect 8428 5564 8468 5573
rect 8428 4976 8468 5524
rect 8524 5060 8564 8716
rect 8620 5144 8660 9472
rect 8716 9472 8852 9512
rect 8716 5816 8756 9472
rect 8908 8924 8948 11764
rect 9100 9680 9140 11764
rect 9100 9631 9140 9640
rect 9196 11612 9236 11621
rect 8908 8875 8948 8884
rect 9004 9512 9044 9521
rect 8716 5767 8756 5776
rect 8812 8672 8852 8681
rect 8812 5480 8852 8632
rect 8812 5431 8852 5440
rect 8620 5095 8660 5104
rect 9004 5144 9044 9472
rect 9196 5648 9236 11572
rect 9292 8924 9332 11764
rect 9484 9680 9524 11764
rect 9484 9631 9524 9640
rect 9292 8875 9332 8884
rect 9676 8924 9716 11764
rect 9868 9680 9908 11764
rect 9868 9631 9908 9640
rect 9676 8875 9716 8884
rect 9964 9512 10004 9521
rect 9676 8756 9716 8765
rect 9196 5599 9236 5608
rect 9580 8672 9620 8681
rect 9004 5095 9044 5104
rect 9580 5144 9620 8632
rect 9580 5095 9620 5104
rect 8524 5011 8564 5020
rect 8428 4927 8468 4936
rect 8812 4976 8852 4985
rect 8812 4388 8852 4936
rect 8812 4339 8852 4348
rect 8332 4255 8372 4264
rect 9676 4304 9716 8716
rect 9772 8672 9812 8681
rect 9772 5060 9812 8632
rect 9772 5011 9812 5020
rect 9676 4255 9716 4264
rect 9388 4136 9428 4145
rect 8236 4096 8372 4136
rect 8044 2876 8276 2900
rect 8044 2860 8236 2876
rect 8332 2876 8372 4096
rect 9964 4136 10004 9472
rect 10060 8924 10100 11764
rect 10252 9680 10292 11764
rect 10252 9631 10292 9640
rect 10348 10688 10388 10697
rect 10060 8875 10100 8884
rect 10156 9512 10196 9521
rect 10156 4976 10196 9472
rect 10156 4927 10196 4936
rect 10348 4808 10388 10648
rect 10444 8924 10484 11764
rect 10444 8875 10484 8884
rect 10540 10604 10580 10613
rect 10348 4759 10388 4768
rect 10444 8756 10484 8765
rect 10252 4136 10292 4145
rect 9964 4096 10252 4136
rect 8620 3212 8660 3221
rect 8620 3077 8660 3172
rect 9388 3044 9428 4096
rect 10252 4087 10292 4096
rect 10444 3968 10484 8716
rect 10540 5060 10580 10564
rect 10636 9680 10676 11764
rect 10636 9631 10676 9640
rect 10828 8924 10868 11764
rect 11020 9680 11060 11764
rect 11020 9631 11060 9640
rect 10828 8875 10868 8884
rect 11212 8924 11252 11764
rect 11404 9680 11444 11764
rect 11404 9631 11444 9640
rect 11212 8875 11252 8884
rect 11308 9512 11348 9521
rect 10732 8672 10772 8681
rect 10732 5144 10772 8632
rect 10732 5095 10772 5104
rect 11116 8672 11156 8681
rect 10540 5011 10580 5020
rect 11116 4808 11156 8632
rect 11116 4759 11156 4768
rect 11020 4304 11060 4313
rect 11020 4169 11060 4264
rect 11308 4304 11348 9472
rect 11404 9428 11444 9437
rect 11404 5732 11444 9388
rect 11596 8924 11636 11764
rect 11788 9680 11828 11764
rect 11788 9631 11828 9640
rect 11884 10016 11924 10025
rect 11596 8875 11636 8884
rect 11404 5683 11444 5692
rect 11500 8672 11540 8681
rect 11500 5228 11540 8632
rect 11692 7160 11732 7169
rect 11500 5179 11540 5188
rect 11596 5816 11636 5825
rect 11596 4892 11636 5776
rect 11692 5060 11732 7120
rect 11692 5011 11732 5020
rect 11788 5648 11828 5657
rect 11596 4843 11636 4852
rect 11692 4892 11732 4901
rect 11308 4255 11348 4264
rect 10444 3919 10484 3928
rect 10924 4136 10964 4145
rect 10924 3800 10964 4096
rect 11692 4136 11732 4852
rect 11692 4087 11732 4096
rect 10924 3751 10964 3760
rect 9388 2995 9428 3004
rect 8428 2876 8468 2885
rect 8332 2836 8428 2876
rect 8236 2827 8276 2836
rect 8428 2827 8468 2836
rect 11500 2792 11540 2887
rect 11500 2743 11540 2752
rect 9100 2708 9140 2717
rect 7372 2540 7412 2549
rect 7372 80 7412 2500
rect 9100 80 9140 2668
rect 11500 2624 11540 2633
rect 10828 1784 10868 1793
rect 10828 80 10868 1744
rect 11500 608 11540 2584
rect 11788 2204 11828 5608
rect 11884 4892 11924 9976
rect 11980 8924 12020 11764
rect 12172 9680 12212 11764
rect 12172 9631 12212 9640
rect 11980 8875 12020 8884
rect 12076 9512 12116 9521
rect 12076 5648 12116 9472
rect 12076 5599 12116 5608
rect 12172 9428 12212 9437
rect 12172 5228 12212 9388
rect 12364 8924 12404 11764
rect 12556 9680 12596 11764
rect 12556 9631 12596 9640
rect 12364 8875 12404 8884
rect 12460 9512 12500 9521
rect 12364 8672 12404 8681
rect 12268 7664 12308 7673
rect 12268 5564 12308 7624
rect 12268 5515 12308 5524
rect 12172 5179 12212 5188
rect 11884 4843 11924 4852
rect 12268 4724 12308 4733
rect 12364 4724 12404 8632
rect 12460 5480 12500 9472
rect 12748 8924 12788 11764
rect 12940 11444 12980 11764
rect 12940 11404 13076 11444
rect 13036 9764 13076 11404
rect 13036 9715 13076 9724
rect 12748 8875 12788 8884
rect 13132 8924 13172 11764
rect 13228 9848 13268 9857
rect 13228 9512 13268 9808
rect 13324 9680 13364 11764
rect 13324 9631 13364 9640
rect 13420 10100 13460 10109
rect 13420 9512 13460 10060
rect 13228 9463 13268 9472
rect 13324 9472 13460 9512
rect 13132 8875 13172 8884
rect 13036 8840 13076 8849
rect 12652 8672 12692 8681
rect 12652 5648 12692 8632
rect 12652 5599 12692 5608
rect 12940 5732 12980 5741
rect 12940 5597 12980 5692
rect 12460 5431 12500 5440
rect 12940 5396 12980 5407
rect 12940 5312 12980 5356
rect 12940 5263 12980 5272
rect 12844 5060 12884 5069
rect 12556 4976 12596 4985
rect 12460 4724 12500 4733
rect 12364 4684 12460 4724
rect 12076 4640 12116 4649
rect 11980 4304 12020 4315
rect 11980 4220 12020 4264
rect 11980 4171 12020 4180
rect 12076 4052 12116 4600
rect 12076 4003 12116 4012
rect 12268 2708 12308 4684
rect 12460 4675 12500 4684
rect 12556 4640 12596 4936
rect 12844 4724 12884 5020
rect 12844 4675 12884 4684
rect 12556 4591 12596 4600
rect 12844 4556 12884 4565
rect 12844 4421 12884 4516
rect 13036 4556 13076 8800
rect 13324 5816 13364 9472
rect 13516 8924 13556 11764
rect 13708 9680 13748 11764
rect 13708 9631 13748 9640
rect 13516 8875 13556 8884
rect 13708 9512 13748 9521
rect 13324 5767 13364 5776
rect 13420 8672 13460 8681
rect 13420 5312 13460 8632
rect 13420 5263 13460 5272
rect 13516 5984 13556 5993
rect 13516 4976 13556 5944
rect 13612 5732 13652 5741
rect 13612 5060 13652 5692
rect 13612 5011 13652 5020
rect 13516 4927 13556 4936
rect 13708 4808 13748 9472
rect 13900 8924 13940 11764
rect 13900 8875 13940 8884
rect 13996 9932 14036 9941
rect 13804 8672 13844 8681
rect 13804 5732 13844 8632
rect 13804 5683 13844 5692
rect 13996 5396 14036 9892
rect 14092 9680 14132 11764
rect 14092 9631 14132 9640
rect 14188 10856 14228 10865
rect 14188 9512 14228 10816
rect 13996 5347 14036 5356
rect 14092 9472 14228 9512
rect 14092 5396 14132 9472
rect 14284 8924 14324 11764
rect 14476 9680 14516 11764
rect 14476 9631 14516 9640
rect 14284 8875 14324 8884
rect 14668 8924 14708 11764
rect 14860 9680 14900 11764
rect 14860 9631 14900 9640
rect 14668 8875 14708 8884
rect 15052 8924 15092 11764
rect 15244 9680 15284 11764
rect 15244 9631 15284 9640
rect 15052 8875 15092 8884
rect 15148 9512 15188 9521
rect 14860 8840 14900 8849
rect 14380 8756 14420 8765
rect 14092 5347 14132 5356
rect 14188 8672 14228 8681
rect 14188 5396 14228 8632
rect 14188 5347 14228 5356
rect 14380 5060 14420 8716
rect 14860 8705 14900 8800
rect 14572 8672 14612 8681
rect 14572 6656 14612 8632
rect 14572 6607 14612 6616
rect 15148 6236 15188 9472
rect 15436 8924 15476 11764
rect 15628 9680 15668 11764
rect 15628 9631 15668 9640
rect 15436 8875 15476 8884
rect 15532 9512 15572 9521
rect 15532 6908 15572 9472
rect 15820 8924 15860 11764
rect 16012 9680 16052 11764
rect 16012 9631 16052 9640
rect 15820 8875 15860 8884
rect 15916 9512 15956 9521
rect 15916 6992 15956 9472
rect 16204 8924 16244 11764
rect 16396 9596 16436 11764
rect 16588 9680 16628 11764
rect 16588 9631 16628 9640
rect 16396 9547 16436 9556
rect 16780 9596 16820 11764
rect 16972 9680 17012 11764
rect 16972 9631 17012 9640
rect 16780 9547 16820 9556
rect 17164 9596 17204 11764
rect 17356 9680 17396 11764
rect 17356 9631 17396 9640
rect 17452 9764 17492 9773
rect 17164 9547 17204 9556
rect 17260 9512 17300 9521
rect 16204 8875 16244 8884
rect 16492 8924 16532 8935
rect 16492 8840 16532 8884
rect 16492 8791 16532 8800
rect 15916 6943 15956 6952
rect 16108 8672 16148 8681
rect 15532 6859 15572 6868
rect 16108 6572 16148 8632
rect 16492 8672 16532 8681
rect 16492 7076 16532 8632
rect 16492 7027 16532 7036
rect 17260 6656 17300 9472
rect 17260 6607 17300 6616
rect 17356 8588 17396 8597
rect 16108 6523 16148 6532
rect 15148 6187 15188 6196
rect 17356 5732 17396 8548
rect 17356 5683 17396 5692
rect 14380 5011 14420 5020
rect 15244 5648 15284 5657
rect 13708 4759 13748 4768
rect 13900 4976 13940 4985
rect 13612 4724 13652 4733
rect 13036 4507 13076 4516
rect 13516 4640 13556 4649
rect 13516 4505 13556 4600
rect 13612 4388 13652 4684
rect 13900 4724 13940 4936
rect 13900 4675 13940 4684
rect 15052 4976 15092 4985
rect 13612 4339 13652 4348
rect 14956 4640 14996 4649
rect 14956 4304 14996 4600
rect 15052 4472 15092 4936
rect 15244 4892 15284 5608
rect 15244 4843 15284 4852
rect 15724 5648 15764 5657
rect 15052 4423 15092 4432
rect 14956 4255 14996 4264
rect 13324 4220 13364 4229
rect 13516 4220 13556 4229
rect 13364 4180 13516 4220
rect 13324 4171 13364 4180
rect 13516 4171 13556 4180
rect 12268 2659 12308 2668
rect 12364 3464 12404 3473
rect 11788 2155 11828 2164
rect 12364 1616 12404 3424
rect 14476 3296 14516 3305
rect 14284 3212 14324 3221
rect 14324 3172 14420 3212
rect 14284 3163 14324 3172
rect 13324 2624 13364 2633
rect 13228 2456 13268 2465
rect 12364 1567 12404 1576
rect 12556 2120 12596 2129
rect 11500 559 11540 568
rect 12556 80 12596 2080
rect 13228 1700 13268 2416
rect 13324 1952 13364 2584
rect 14380 2624 14420 3172
rect 14476 3044 14516 3256
rect 14476 2995 14516 3004
rect 14668 3044 14708 3053
rect 14668 2876 14708 3004
rect 14668 2827 14708 2836
rect 15724 2876 15764 5608
rect 16012 5648 16052 5657
rect 16012 5144 16052 5608
rect 17452 5564 17492 9724
rect 17452 5515 17492 5524
rect 16012 5095 16052 5104
rect 17068 5312 17108 5321
rect 16780 4976 16820 4985
rect 17068 4976 17108 5272
rect 16820 4936 17108 4976
rect 16780 4927 16820 4936
rect 17548 4556 17588 11764
rect 17740 11696 17780 11764
rect 17740 11647 17780 11656
rect 17932 11612 17972 11764
rect 17932 11563 17972 11572
rect 18124 10688 18164 11764
rect 18124 10639 18164 10648
rect 17740 9848 17780 9857
rect 17644 9512 17684 9521
rect 17644 7160 17684 9472
rect 17644 7111 17684 7120
rect 17740 5648 17780 9808
rect 18316 7664 18356 11764
rect 18316 7615 18356 7624
rect 17740 5599 17780 5608
rect 17548 4507 17588 4516
rect 17644 4808 17684 4817
rect 15724 2827 15764 2836
rect 17644 2876 17684 4768
rect 17740 4724 17780 4733
rect 17740 4556 17780 4684
rect 18508 4640 18548 11764
rect 18700 10604 18740 11764
rect 18700 10555 18740 10564
rect 18892 10016 18932 11764
rect 19084 10016 19124 11764
rect 19276 10184 19316 11764
rect 19468 10184 19508 11764
rect 19468 10144 19604 10184
rect 19276 10135 19316 10144
rect 19468 10016 19508 10025
rect 19084 9976 19412 10016
rect 18892 9967 18932 9976
rect 18808 9848 19176 9857
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 18808 9799 19176 9808
rect 18892 9680 18932 9689
rect 18700 9512 18740 9521
rect 18700 7412 18740 9472
rect 18892 8924 18932 9640
rect 18892 8875 18932 8884
rect 18808 8336 19176 8345
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 18808 8287 19176 8296
rect 18700 7363 18740 7372
rect 18796 7160 18836 7169
rect 18796 6992 18836 7120
rect 19372 7160 19412 9976
rect 19372 7111 19412 7120
rect 18796 6943 18836 6952
rect 18808 6824 19176 6833
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 18808 6775 19176 6784
rect 19468 5816 19508 9976
rect 19564 9932 19604 10144
rect 19564 9883 19604 9892
rect 19660 9680 19700 11764
rect 19660 9631 19700 9640
rect 19756 9596 19796 9605
rect 19756 9512 19796 9556
rect 19660 9472 19796 9512
rect 19564 9428 19604 9437
rect 19564 8000 19604 9388
rect 19564 7951 19604 7960
rect 19468 5767 19508 5776
rect 19564 7832 19604 7841
rect 18700 5480 18740 5489
rect 18700 5312 18740 5440
rect 19564 5480 19604 7792
rect 19564 5431 19604 5440
rect 18700 5263 18740 5272
rect 18808 5312 19176 5321
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 18808 5263 19176 5272
rect 19660 4724 19700 9472
rect 19756 9260 19796 9269
rect 19756 7748 19796 9220
rect 19852 8168 19892 11764
rect 20044 9596 20084 11764
rect 20044 9547 20084 9556
rect 19852 8119 19892 8128
rect 19948 9344 19988 9353
rect 19756 7699 19796 7708
rect 19852 8000 19892 8009
rect 19852 7412 19892 7960
rect 19948 7832 19988 9304
rect 20236 9260 20276 11764
rect 20428 9596 20468 11764
rect 20428 9547 20468 9556
rect 20236 9220 20564 9260
rect 20048 9092 20416 9101
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20048 9043 20416 9052
rect 19948 7783 19988 7792
rect 20140 8756 20180 8765
rect 20140 7832 20180 8716
rect 20140 7783 20180 7792
rect 20048 7580 20416 7589
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20048 7531 20416 7540
rect 19852 7363 19892 7372
rect 20044 6992 20084 7001
rect 19852 6952 20044 6992
rect 19852 6572 19892 6952
rect 20044 6943 20084 6952
rect 19852 6523 19892 6532
rect 20044 6488 20084 6497
rect 20044 6353 20084 6448
rect 20048 6068 20416 6077
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20048 6019 20416 6028
rect 19660 4675 19700 4684
rect 18508 4591 18548 4600
rect 18700 4640 18740 4649
rect 17740 4507 17780 4516
rect 18700 4505 18740 4600
rect 20048 4556 20416 4565
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20048 4507 20416 4516
rect 20524 4388 20564 9220
rect 20620 4640 20660 11764
rect 20716 9596 20756 9605
rect 20716 4724 20756 9556
rect 20716 4675 20756 4684
rect 20620 4591 20660 4600
rect 20524 4339 20564 4348
rect 17932 4220 17972 4229
rect 17644 2827 17684 2836
rect 17740 3212 17780 3221
rect 15436 2708 15476 2717
rect 14380 2575 14420 2584
rect 14764 2624 14804 2633
rect 13324 1903 13364 1912
rect 14284 2036 14324 2045
rect 13228 1651 13268 1660
rect 14284 80 14324 1996
rect 14764 944 14804 2584
rect 15436 2573 15476 2668
rect 15820 2624 15860 2633
rect 15820 1280 15860 2584
rect 17356 2624 17396 2633
rect 17356 2204 17396 2584
rect 17740 2624 17780 3172
rect 17932 3128 17972 4180
rect 19948 4052 19988 4061
rect 18700 3884 18740 3895
rect 18700 3800 18740 3844
rect 18700 3751 18740 3760
rect 18808 3800 19176 3809
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 18808 3751 19176 3760
rect 19372 3800 19412 3809
rect 17932 3079 17972 3088
rect 18508 3464 18548 3473
rect 18508 2960 18548 3424
rect 18508 2911 18548 2920
rect 18892 3464 18932 3473
rect 18892 2792 18932 3424
rect 18892 2743 18932 2752
rect 19276 3464 19316 3473
rect 17740 2575 17780 2584
rect 18808 2288 19176 2297
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 18808 2239 19176 2248
rect 17356 2155 17396 2164
rect 19276 2204 19316 3424
rect 19372 3296 19412 3760
rect 19948 3464 19988 4012
rect 19948 3415 19988 3424
rect 20428 4052 20468 4061
rect 19372 3247 19412 3256
rect 19852 3380 19892 3389
rect 19852 3044 19892 3340
rect 19852 2995 19892 3004
rect 19948 3212 19988 3221
rect 19948 2960 19988 3172
rect 20428 3212 20468 4012
rect 20812 3884 20852 11764
rect 20908 6992 20948 7001
rect 20908 6572 20948 6952
rect 20908 6523 20948 6532
rect 21004 4052 21044 11764
rect 21196 10856 21236 11764
rect 21196 10807 21236 10816
rect 21196 7160 21236 7169
rect 21100 6992 21140 7001
rect 21196 6992 21236 7120
rect 21292 6992 21332 7001
rect 21196 6952 21292 6992
rect 21100 6236 21140 6952
rect 21292 6943 21332 6952
rect 21388 6656 21428 11764
rect 21388 6607 21428 6616
rect 21196 6488 21236 6497
rect 21196 6353 21236 6448
rect 21484 6404 21524 6413
rect 21100 6187 21140 6196
rect 21004 4003 21044 4012
rect 20812 3835 20852 3844
rect 21196 3884 21236 3893
rect 21196 3464 21236 3844
rect 21196 3415 21236 3424
rect 20428 3163 20468 3172
rect 21004 3296 21044 3305
rect 21004 3161 21044 3256
rect 20048 3044 20416 3053
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20048 2995 20416 3004
rect 19948 2911 19988 2920
rect 21484 2876 21524 6364
rect 21580 5060 21620 11764
rect 21676 8000 21716 8009
rect 21676 7496 21716 7960
rect 21676 7447 21716 7456
rect 21772 5228 21812 11764
rect 21964 5648 22004 11764
rect 21964 5599 22004 5608
rect 22156 5564 22196 11764
rect 22348 5732 22388 11764
rect 22348 5683 22388 5692
rect 22156 5515 22196 5524
rect 22540 5396 22580 11764
rect 22636 8000 22676 8009
rect 22636 7580 22676 7960
rect 22636 7531 22676 7540
rect 22540 5347 22580 5356
rect 21772 5179 21812 5188
rect 22732 5144 22772 11764
rect 22924 9176 22964 11764
rect 22732 5095 22772 5104
rect 22828 9136 22964 9176
rect 21580 5011 21620 5020
rect 22828 4976 22868 9136
rect 23116 8588 23156 11764
rect 23116 8539 23156 8548
rect 22924 8000 22964 8009
rect 22924 7328 22964 7960
rect 23020 7328 23060 7337
rect 22924 7288 23020 7328
rect 23020 7279 23060 7288
rect 22828 4927 22868 4936
rect 23308 4892 23348 11764
rect 23308 4843 23348 4852
rect 23500 4472 23540 11764
rect 23692 5984 23732 11764
rect 23884 10016 23924 11764
rect 23884 9967 23924 9976
rect 23884 8840 23924 8849
rect 23884 8000 23924 8800
rect 23884 7951 23924 7960
rect 23692 5935 23732 5944
rect 23980 4976 24020 4985
rect 23980 4841 24020 4936
rect 23500 4423 23540 4432
rect 24076 4304 24116 11764
rect 24308 11764 24328 11780
rect 24440 11764 24520 11844
rect 24632 11764 24712 11844
rect 24824 11764 24904 11844
rect 25016 11764 25096 11844
rect 25208 11764 25288 11844
rect 25400 11764 25480 11844
rect 25592 11764 25672 11844
rect 25784 11764 25864 11844
rect 25976 11764 26056 11844
rect 26168 11764 26248 11844
rect 26360 11764 26440 11844
rect 26552 11764 26632 11844
rect 26744 11764 26824 11844
rect 26936 11764 27016 11844
rect 27128 11764 27208 11844
rect 27320 11764 27400 11844
rect 27512 11764 27592 11844
rect 27704 11764 27784 11844
rect 27896 11764 27976 11844
rect 28088 11764 28168 11844
rect 28280 11764 28360 11844
rect 28472 11764 28552 11844
rect 28664 11764 28744 11844
rect 28856 11764 28936 11844
rect 29048 11764 29128 11844
rect 29240 11764 29320 11844
rect 29432 11764 29512 11844
rect 29624 11764 29704 11844
rect 29816 11764 29896 11844
rect 30008 11764 30088 11844
rect 30200 11764 30280 11844
rect 30392 11764 30472 11844
rect 30584 11764 30664 11844
rect 30776 11764 30856 11844
rect 30968 11764 31048 11844
rect 31160 11764 31240 11844
rect 31352 11764 31432 11844
rect 24268 11731 24308 11740
rect 24268 9176 24308 9185
rect 24172 8336 24212 8345
rect 24172 8000 24212 8296
rect 24172 7951 24212 7960
rect 24268 7748 24308 9136
rect 24364 8924 24404 8933
rect 24364 7832 24404 8884
rect 24364 7783 24404 7792
rect 24268 7699 24308 7708
rect 24460 7220 24500 11764
rect 24460 7180 24596 7220
rect 24556 7076 24596 7180
rect 24556 7027 24596 7036
rect 24652 6908 24692 11764
rect 24652 6859 24692 6868
rect 24844 6488 24884 11764
rect 25036 7412 25076 11764
rect 25228 7496 25268 11764
rect 25228 7447 25268 7456
rect 25036 7363 25076 7372
rect 25420 6572 25460 11764
rect 25612 9512 25652 11764
rect 25516 9472 25652 9512
rect 25516 6656 25556 9472
rect 25708 8252 25748 8261
rect 25708 8117 25748 8212
rect 25804 7220 25844 11764
rect 25900 8588 25940 8597
rect 25900 8000 25940 8548
rect 25900 7951 25940 7960
rect 25708 7180 25844 7220
rect 25516 6607 25556 6616
rect 25612 7160 25652 7169
rect 25420 6523 25460 6532
rect 24844 6439 24884 6448
rect 25612 6152 25652 7120
rect 25708 6824 25748 7180
rect 25996 6908 26036 11764
rect 26092 8672 26132 8681
rect 26092 8000 26132 8632
rect 26092 7951 26132 7960
rect 26188 7220 26228 11764
rect 26380 9932 26420 11764
rect 26284 9892 26420 9932
rect 26284 7580 26324 9892
rect 26380 8168 26420 8177
rect 26380 8033 26420 8128
rect 26284 7531 26324 7540
rect 26572 7328 26612 11764
rect 26764 8336 26804 11764
rect 26956 8588 26996 11764
rect 26956 8539 26996 8548
rect 26764 8287 26804 8296
rect 27148 8000 27188 11764
rect 27340 11444 27380 11764
rect 27340 11404 27476 11444
rect 27436 9512 27476 11404
rect 27532 9680 27572 11764
rect 27532 9631 27572 9640
rect 27724 9596 27764 11764
rect 27916 9680 27956 11764
rect 27916 9631 27956 9640
rect 28012 9848 28052 9857
rect 27724 9547 27764 9556
rect 27820 9512 27860 9521
rect 27436 9472 27668 9512
rect 27244 9008 27284 9017
rect 27244 8000 27284 8968
rect 27436 8756 27476 8765
rect 27340 8000 27380 8009
rect 27244 7960 27340 8000
rect 27148 7951 27188 7960
rect 27340 7932 27380 7960
rect 26572 7279 26612 7288
rect 26092 7180 26228 7220
rect 26092 7076 26132 7180
rect 26092 7027 26132 7036
rect 25996 6859 26036 6868
rect 25708 6775 25748 6784
rect 25612 6103 25652 6112
rect 24076 4255 24116 4264
rect 26380 4976 26420 4985
rect 24460 4220 24500 4229
rect 21580 4136 21620 4145
rect 21580 3548 21620 4096
rect 24460 3884 24500 4180
rect 24460 3835 24500 3844
rect 24652 4136 24692 4145
rect 22540 3800 22580 3809
rect 21580 3499 21620 3508
rect 21676 3716 21716 3725
rect 21676 3296 21716 3676
rect 22540 3464 22580 3760
rect 22540 3415 22580 3424
rect 22924 3800 22964 3809
rect 21676 3247 21716 3256
rect 21772 3212 21812 3221
rect 21772 3044 21812 3172
rect 21772 2995 21812 3004
rect 21484 2827 21524 2836
rect 19756 2792 19796 2801
rect 19660 2624 19700 2633
rect 19564 2372 19604 2381
rect 19372 2332 19564 2372
rect 19372 2288 19412 2332
rect 19564 2323 19604 2332
rect 19372 2239 19412 2248
rect 19660 2288 19700 2584
rect 19660 2239 19700 2248
rect 19276 2155 19316 2164
rect 17740 1952 17780 1961
rect 15820 1231 15860 1240
rect 16012 1868 16052 1877
rect 14764 895 14804 904
rect 16012 80 16052 1828
rect 17740 80 17780 1912
rect 19756 188 19796 2752
rect 21196 2792 21236 2801
rect 21196 2624 21236 2752
rect 21196 2575 21236 2584
rect 21580 2624 21620 2633
rect 21580 1784 21620 2584
rect 21580 1735 21620 1744
rect 21196 1616 21236 1625
rect 20048 1532 20416 1541
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20048 1483 20416 1492
rect 19468 148 19796 188
rect 19468 80 19508 148
rect 21196 80 21236 1576
rect 22924 80 22964 3760
rect 23020 3380 23060 3389
rect 23020 3245 23060 3340
rect 24652 80 24692 4096
rect 25612 2624 25652 2633
rect 25612 1952 25652 2584
rect 25612 1903 25652 1912
rect 25804 2288 25844 2297
rect 25804 1952 25844 2248
rect 25804 1903 25844 1912
rect 26380 80 26420 4936
rect 27148 3968 27188 3977
rect 26764 3884 26804 3893
rect 26764 3548 26804 3844
rect 26764 3499 26804 3508
rect 27052 3800 27092 3809
rect 27052 3212 27092 3760
rect 27148 3464 27188 3928
rect 27148 3415 27188 3424
rect 27052 3163 27092 3172
rect 27436 2792 27476 8716
rect 27436 2743 27476 2752
rect 27532 8672 27572 8681
rect 27052 2624 27092 2633
rect 27052 1616 27092 2584
rect 27052 1567 27092 1576
rect 27436 2624 27476 2633
rect 27436 1532 27476 2584
rect 27532 2456 27572 8632
rect 27628 8000 27668 9472
rect 27724 8000 27764 8009
rect 27628 7960 27724 8000
rect 27724 7951 27764 7960
rect 27628 7832 27668 7841
rect 27628 2708 27668 7792
rect 27820 4052 27860 9472
rect 28012 7832 28052 9808
rect 28108 9596 28148 11764
rect 28300 9764 28340 11764
rect 28300 9715 28340 9724
rect 28108 9547 28148 9556
rect 28204 9512 28244 9521
rect 28204 9377 28244 9472
rect 28492 8924 28532 11764
rect 28588 9512 28628 9521
rect 28588 9428 28628 9472
rect 28588 9377 28628 9388
rect 28684 9344 28724 11764
rect 28684 9295 28724 9304
rect 28780 9932 28820 9941
rect 28492 8875 28532 8884
rect 28012 7783 28052 7792
rect 27820 4003 27860 4012
rect 28108 5648 28148 5657
rect 27628 2659 27668 2668
rect 27532 2407 27572 2416
rect 27820 2624 27860 2633
rect 27820 1868 27860 2584
rect 27820 1819 27860 1828
rect 27436 1483 27476 1492
rect 28108 80 28148 5608
rect 28780 5144 28820 9892
rect 28876 8924 28916 11764
rect 29068 9596 29108 11764
rect 29068 9547 29108 9556
rect 28972 9512 29012 9521
rect 28972 9344 29012 9472
rect 28972 9295 29012 9304
rect 29068 9428 29108 9437
rect 28876 8875 28916 8884
rect 28972 9008 29012 9017
rect 28780 5095 28820 5104
rect 28876 8588 28916 8597
rect 28780 4220 28820 4229
rect 28780 3884 28820 4180
rect 28780 3835 28820 3844
rect 28588 3716 28628 3725
rect 28780 3716 28820 3725
rect 28628 3676 28780 3716
rect 28588 3667 28628 3676
rect 28780 3667 28820 3676
rect 28588 3548 28628 3557
rect 28780 3548 28820 3557
rect 28628 3508 28780 3548
rect 28588 3499 28628 3508
rect 28780 3499 28820 3508
rect 28876 2876 28916 8548
rect 28972 3632 29012 8968
rect 28972 3583 29012 3592
rect 28876 2827 28916 2836
rect 29068 2792 29108 9388
rect 29260 8924 29300 11764
rect 29356 9512 29396 9521
rect 29356 9260 29396 9472
rect 29356 9211 29396 9220
rect 29452 9260 29492 11764
rect 29452 9211 29492 9220
rect 29548 9512 29588 9521
rect 29260 8875 29300 8884
rect 29356 8840 29396 8849
rect 29164 8672 29204 8681
rect 29164 2876 29204 8632
rect 29356 7220 29396 8800
rect 29260 7180 29396 7220
rect 29452 8756 29492 8765
rect 29260 5648 29300 7180
rect 29260 5599 29300 5608
rect 29452 4304 29492 8716
rect 29452 4255 29492 4264
rect 29164 2827 29204 2836
rect 29548 2876 29588 9472
rect 29644 8924 29684 11764
rect 29836 10016 29876 11764
rect 29836 9967 29876 9976
rect 29740 9344 29780 9353
rect 29740 9008 29780 9304
rect 29740 8959 29780 8968
rect 29932 9092 29972 9101
rect 29644 8875 29684 8884
rect 29740 8588 29780 8597
rect 29644 8420 29684 8429
rect 29644 8000 29684 8380
rect 29644 7951 29684 7960
rect 29740 6656 29780 8548
rect 29932 7076 29972 9052
rect 30028 8924 30068 11764
rect 30124 10016 30164 10025
rect 30124 9680 30164 9976
rect 30220 9764 30260 11764
rect 30220 9715 30260 9724
rect 30124 9631 30164 9640
rect 30028 8875 30068 8884
rect 30124 9176 30164 9185
rect 30028 8504 30068 8513
rect 30028 8000 30068 8464
rect 30028 7951 30068 7960
rect 30124 7220 30164 9136
rect 30220 9008 30260 9017
rect 30220 8168 30260 8968
rect 30412 8924 30452 11764
rect 30604 9344 30644 11764
rect 30604 9295 30644 9304
rect 30412 8875 30452 8884
rect 30796 8924 30836 11764
rect 30988 9428 31028 11764
rect 30988 9379 31028 9388
rect 30796 8875 30836 8884
rect 31180 8924 31220 11764
rect 31372 9680 31412 11764
rect 37036 11024 37076 11033
rect 36172 10688 36212 10697
rect 33928 9848 34296 9857
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 33928 9799 34296 9808
rect 31372 9631 31412 9640
rect 31468 9764 31508 9773
rect 31180 8875 31220 8884
rect 30796 8756 30836 8765
rect 30220 8119 30260 8128
rect 30412 8252 30452 8261
rect 30412 8000 30452 8212
rect 30412 7951 30452 7960
rect 30604 8168 30644 8177
rect 30604 8000 30644 8128
rect 30604 7951 30644 7960
rect 30796 7412 30836 8716
rect 30796 7363 30836 7372
rect 31468 7220 31508 9724
rect 36172 9680 36212 10648
rect 36172 9631 36212 9640
rect 36556 10352 36596 10361
rect 36556 9680 36596 10312
rect 36556 9631 36596 9640
rect 32620 9596 32660 9605
rect 32140 9344 32180 9353
rect 31660 8840 31700 8849
rect 31660 8168 31700 8800
rect 31660 8119 31700 8128
rect 32140 7748 32180 9304
rect 32140 7699 32180 7708
rect 32236 9260 32276 9269
rect 32236 7664 32276 9220
rect 32524 8672 32564 8681
rect 32524 8537 32564 8632
rect 32620 8084 32660 9556
rect 35884 9512 35924 9521
rect 33100 9428 33140 9437
rect 33100 8168 33140 9388
rect 35168 9092 35536 9101
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35168 9043 35536 9052
rect 35884 9008 35924 9472
rect 35884 8959 35924 8968
rect 36268 9512 36308 9521
rect 34540 8756 34580 8765
rect 33928 8336 34296 8345
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 33928 8287 34296 8296
rect 33100 8119 33140 8128
rect 32620 8035 32660 8044
rect 32236 7615 32276 7624
rect 29932 7027 29972 7036
rect 30028 7180 30164 7220
rect 31372 7180 31508 7220
rect 29740 6607 29780 6616
rect 30028 6656 30068 7180
rect 31084 7160 31124 7169
rect 31084 6992 31124 7120
rect 31372 7160 31412 7180
rect 31372 7111 31412 7120
rect 32716 7160 32756 7169
rect 31084 6943 31124 6952
rect 30028 6607 30068 6616
rect 29548 2827 29588 2836
rect 29836 6488 29876 6497
rect 29068 2743 29108 2752
rect 29548 2624 29588 2633
rect 29548 2036 29588 2584
rect 29548 1987 29588 1996
rect 29836 80 29876 6448
rect 31564 6404 31604 6413
rect 30988 2624 31028 2633
rect 30988 2120 31028 2584
rect 30988 2071 31028 2080
rect 31564 80 31604 6364
rect 32716 3800 32756 7120
rect 32716 3751 32756 3760
rect 33292 6908 33332 6917
rect 33292 80 33332 6868
rect 34540 6908 34580 8716
rect 35980 8000 36020 8009
rect 35168 7580 35536 7589
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35168 7531 35536 7540
rect 34540 6859 34580 6868
rect 34924 7076 34964 7085
rect 33928 6824 34296 6833
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 33928 6775 34296 6784
rect 34540 6404 34580 6413
rect 33928 5312 34296 5321
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 33928 5263 34296 5272
rect 33928 3800 34296 3809
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 33928 3751 34296 3760
rect 34540 2456 34580 6364
rect 34828 4976 34868 4985
rect 34828 3464 34868 4936
rect 34828 3415 34868 3424
rect 34924 2876 34964 7036
rect 35168 6068 35536 6077
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35168 6019 35536 6028
rect 35980 5144 36020 7960
rect 36268 7664 36308 9472
rect 36652 9512 36692 9521
rect 36652 9260 36692 9472
rect 36652 9211 36692 9220
rect 37036 8924 37076 10984
rect 37036 8875 37076 8884
rect 37324 10016 37364 10025
rect 37324 8924 37364 9976
rect 37324 8875 37364 8884
rect 38668 9260 38708 9269
rect 37804 8672 37844 8681
rect 36268 7615 36308 7624
rect 37612 8000 37652 8009
rect 35884 5104 36020 5144
rect 36076 7076 36116 7085
rect 35884 4724 35924 5104
rect 35884 4675 35924 4684
rect 35168 4556 35536 4565
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35168 4507 35536 4516
rect 36076 3968 36116 7036
rect 36076 3919 36116 3928
rect 36748 6992 36788 7001
rect 35020 3464 35060 3473
rect 35020 3044 35060 3424
rect 35020 2995 35060 3004
rect 35168 3044 35536 3053
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35168 2995 35536 3004
rect 34924 2836 35060 2876
rect 34540 2407 34580 2416
rect 33928 2288 34296 2297
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 33928 2239 34296 2248
rect 35020 80 35060 2836
rect 36652 2540 36692 2549
rect 36652 1952 36692 2500
rect 36652 1903 36692 1912
rect 35168 1532 35536 1541
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35168 1483 35536 1492
rect 36748 80 36788 6952
rect 37420 5648 37460 5657
rect 37420 5513 37460 5608
rect 37516 4892 37556 4901
rect 37228 4136 37268 4145
rect 37228 3296 37268 4096
rect 37324 3884 37364 3893
rect 37324 3548 37364 3844
rect 37420 3716 37460 3725
rect 37516 3716 37556 4852
rect 37612 4220 37652 7960
rect 37804 6656 37844 8632
rect 38668 8672 38708 9220
rect 39148 9176 39188 9185
rect 39148 9008 39188 9136
rect 39148 8959 39188 8968
rect 38668 8623 38708 8632
rect 38668 8504 38708 8513
rect 38668 8000 38708 8464
rect 38668 7951 38708 7960
rect 38668 7748 38708 7757
rect 38668 7328 38708 7708
rect 38668 7279 38708 7288
rect 37804 6607 37844 6616
rect 39148 6824 39188 6833
rect 39148 6656 39188 6784
rect 39148 6607 39188 6616
rect 37612 4171 37652 4180
rect 37460 3676 37556 3716
rect 37420 3648 37460 3676
rect 37324 3508 37556 3548
rect 37228 3247 37268 3256
rect 37516 2624 37556 3508
rect 37804 3212 37844 3221
rect 37516 2575 37556 2584
rect 37612 2960 37652 2969
rect 37612 1952 37652 2920
rect 37804 2624 37844 3172
rect 37804 2575 37844 2584
rect 37612 1903 37652 1912
rect 37804 1784 37844 1793
rect 37516 1700 37556 1709
rect 37516 608 37556 1660
rect 37804 944 37844 1744
rect 37804 895 37844 904
rect 37516 559 37556 568
rect 3340 20 3764 60
rect 3896 0 3976 80
rect 5624 0 5704 80
rect 7352 0 7432 80
rect 9080 0 9160 80
rect 10808 0 10888 80
rect 12536 0 12616 80
rect 14264 0 14344 80
rect 15992 0 16072 80
rect 17720 0 17800 80
rect 19448 0 19528 80
rect 21176 0 21256 80
rect 22904 0 22984 80
rect 24632 0 24712 80
rect 26360 0 26440 80
rect 28088 0 28168 80
rect 29816 0 29896 80
rect 31544 0 31624 80
rect 33272 0 33352 80
rect 35000 0 35080 80
rect 36728 0 36808 80
<< via3 >>
rect 460 8632 500 8672
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 3532 9472 3572 9512
rect 76 3172 116 3212
rect 1036 4936 1076 4976
rect 5644 9388 5684 9428
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 6316 5608 6356 5648
rect 8044 9220 8084 9260
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 8236 9304 8276 9344
rect 9196 5608 9236 5648
rect 10348 10648 10388 10688
rect 8620 3172 8660 3212
rect 11020 4264 11060 4304
rect 11404 5692 11444 5732
rect 11692 7120 11732 7160
rect 11596 5776 11636 5816
rect 11692 4852 11732 4892
rect 11500 2752 11540 2792
rect 12268 7624 12308 7664
rect 11884 4852 11924 4892
rect 12940 5692 12980 5732
rect 12940 5356 12980 5396
rect 11980 4264 12020 4304
rect 12844 4684 12884 4724
rect 12844 4516 12884 4556
rect 14860 8800 14900 8840
rect 14092 5356 14132 5396
rect 16492 8800 16532 8840
rect 17356 8548 17396 8588
rect 13036 4516 13076 4556
rect 13516 4600 13556 4640
rect 15724 5608 15764 5648
rect 12268 2668 12308 2708
rect 18124 10648 18164 10688
rect 18316 7624 18356 7664
rect 17740 4684 17780 4724
rect 18892 9976 18932 10016
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 19372 7120 19412 7160
rect 19468 9976 19508 10016
rect 18796 6952 18836 6992
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 19756 9556 19796 9596
rect 19468 5776 19508 5816
rect 19564 7792 19604 7832
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 20044 9556 20084 9596
rect 19852 8128 19892 8168
rect 20428 9556 20468 9596
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 20044 6448 20084 6488
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 18700 4600 18740 4640
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 20716 9556 20756 9596
rect 15436 2668 15476 2708
rect 18700 3844 18740 3884
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 19852 3340 19892 3380
rect 20908 6952 20948 6992
rect 21196 6448 21236 6488
rect 20812 3844 20852 3884
rect 21004 3256 21044 3296
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 23116 8548 23156 8588
rect 23980 4936 24020 4976
rect 25708 8212 25748 8252
rect 26380 8128 26420 8168
rect 21676 3256 21716 3296
rect 21196 2752 21236 2792
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 23020 3340 23060 3380
rect 27628 7792 27668 7832
rect 28204 9472 28244 9512
rect 28588 9388 28628 9428
rect 28012 7792 28052 7832
rect 28972 9304 29012 9344
rect 29356 9220 29396 9260
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 30412 8212 30452 8252
rect 30604 8128 30644 8168
rect 32524 8632 32564 8672
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 37420 5608 37460 5648
<< metal4 >>
rect 10339 10648 10348 10688
rect 10388 10648 18124 10688
rect 18164 10648 18173 10688
rect 18883 9976 18892 10016
rect 18932 9976 19468 10016
rect 19508 9976 19517 10016
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 19747 9556 19756 9596
rect 19796 9556 20044 9596
rect 20084 9556 20093 9596
rect 20419 9556 20428 9596
rect 20468 9556 20716 9596
rect 20756 9556 20765 9596
rect 3523 9472 3532 9512
rect 3572 9472 28204 9512
rect 28244 9472 28253 9512
rect 5635 9388 5644 9428
rect 5684 9388 28588 9428
rect 28628 9388 28637 9428
rect 8227 9304 8236 9344
rect 8276 9304 28972 9344
rect 29012 9304 29021 9344
rect 8035 9220 8044 9260
rect 8084 9220 29356 9260
rect 29396 9220 29405 9260
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 14851 8800 14860 8840
rect 14900 8800 16492 8840
rect 16532 8800 16541 8840
rect 451 8632 460 8672
rect 500 8632 32524 8672
rect 32564 8632 32573 8672
rect 17347 8548 17356 8588
rect 17396 8548 23116 8588
rect 23156 8548 23165 8588
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 25699 8212 25708 8252
rect 25748 8212 30412 8252
rect 30452 8212 30461 8252
rect 19564 8128 19852 8168
rect 19892 8128 19901 8168
rect 26371 8128 26380 8168
rect 26420 8128 30604 8168
rect 30644 8128 30653 8168
rect 19564 7832 19604 8128
rect 19555 7792 19564 7832
rect 19604 7792 19613 7832
rect 27619 7792 27628 7832
rect 27668 7792 28012 7832
rect 28052 7792 28061 7832
rect 12259 7624 12268 7664
rect 12308 7624 18316 7664
rect 18356 7624 18365 7664
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 11683 7120 11692 7160
rect 11732 7120 19372 7160
rect 19412 7120 19421 7160
rect 18787 6952 18796 6992
rect 18836 6952 20908 6992
rect 20948 6952 20957 6992
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 20035 6448 20044 6488
rect 20084 6448 21196 6488
rect 21236 6448 21245 6488
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 11587 5776 11596 5816
rect 11636 5776 19468 5816
rect 19508 5776 19517 5816
rect 11395 5692 11404 5732
rect 11444 5692 12940 5732
rect 12980 5692 12989 5732
rect 6307 5608 6316 5648
rect 6356 5608 9196 5648
rect 9236 5608 9245 5648
rect 15715 5608 15724 5648
rect 15764 5608 37420 5648
rect 37460 5608 37469 5648
rect 12931 5356 12940 5396
rect 12980 5356 14092 5396
rect 14132 5356 14141 5396
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 1027 4936 1036 4976
rect 1076 4936 23980 4976
rect 24020 4936 24029 4976
rect 11683 4852 11692 4892
rect 11732 4852 11884 4892
rect 11924 4852 11933 4892
rect 12835 4684 12844 4724
rect 12884 4684 17740 4724
rect 17780 4684 17789 4724
rect 13507 4600 13516 4640
rect 13556 4600 18700 4640
rect 18740 4600 18749 4640
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 12835 4516 12844 4556
rect 12884 4516 13036 4556
rect 13076 4516 13085 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 11011 4264 11020 4304
rect 11060 4264 11980 4304
rect 12020 4264 12029 4304
rect 18691 3844 18700 3884
rect 18740 3844 20812 3884
rect 20852 3844 20861 3884
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 19843 3340 19852 3380
rect 19892 3340 23020 3380
rect 23060 3340 23069 3380
rect 20995 3256 21004 3296
rect 21044 3256 21676 3296
rect 21716 3256 21725 3296
rect 67 3172 76 3212
rect 116 3172 8620 3212
rect 8660 3172 8669 3212
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 11491 2752 11500 2792
rect 11540 2752 21196 2792
rect 21236 2752 21245 2792
rect 12259 2668 12268 2708
rect 12308 2668 15436 2708
rect 15476 2668 15485 2708
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
<< via4 >>
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
<< metal5 >>
rect 3652 9848 4092 11844
rect 3652 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4092 9848
rect 3652 8336 4092 9808
rect 3652 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4092 8336
rect 3652 6824 4092 8296
rect 3652 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4092 6824
rect 3652 5312 4092 6784
rect 3652 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4092 5312
rect 3652 3800 4092 5272
rect 3652 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4092 3800
rect 3652 2288 4092 3760
rect 3652 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4092 2288
rect 3652 0 4092 2248
rect 4892 9092 5332 11844
rect 4892 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5332 9092
rect 4892 7580 5332 9052
rect 4892 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5332 7580
rect 4892 6068 5332 7540
rect 4892 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5332 6068
rect 4892 4556 5332 6028
rect 4892 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5332 4556
rect 4892 3044 5332 4516
rect 4892 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5332 3044
rect 4892 1532 5332 3004
rect 4892 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5332 1532
rect 4892 0 5332 1492
rect 18772 9848 19212 11844
rect 18772 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19212 9848
rect 18772 8336 19212 9808
rect 18772 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19212 8336
rect 18772 6824 19212 8296
rect 18772 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19212 6824
rect 18772 5312 19212 6784
rect 18772 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19212 5312
rect 18772 3800 19212 5272
rect 18772 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19212 3800
rect 18772 2288 19212 3760
rect 18772 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19212 2288
rect 18772 0 19212 2248
rect 20012 9092 20452 11844
rect 20012 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20452 9092
rect 20012 7580 20452 9052
rect 20012 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20452 7580
rect 20012 6068 20452 7540
rect 20012 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20452 6068
rect 20012 4556 20452 6028
rect 20012 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20452 4556
rect 20012 3044 20452 4516
rect 20012 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20452 3044
rect 20012 1532 20452 3004
rect 20012 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20452 1532
rect 20012 0 20452 1492
rect 33892 9848 34332 11844
rect 33892 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34332 9848
rect 33892 8336 34332 9808
rect 33892 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34332 8336
rect 33892 6824 34332 8296
rect 33892 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34332 6824
rect 33892 5312 34332 6784
rect 33892 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34332 5312
rect 33892 3800 34332 5272
rect 33892 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34332 3800
rect 33892 2288 34332 3760
rect 33892 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34332 2288
rect 33892 0 34332 2248
rect 35132 9092 35572 11844
rect 35132 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35572 9092
rect 35132 7580 35572 9052
rect 35132 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35572 7580
rect 35132 6068 35572 7540
rect 35132 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35572 6068
rect 35132 4556 35572 6028
rect 35132 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35572 4556
rect 35132 3044 35572 4516
rect 35132 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35572 3044
rect 35132 1532 35572 3004
rect 35132 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35572 1532
rect 35132 0 35572 1492
use sg13g2_buf_1  _000_
timestamp 1676381911
transform 1 0 11424 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _001_
timestamp 1676381911
transform 1 0 14688 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _002_
timestamp 1676381911
transform 1 0 15744 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _003_
timestamp 1676381911
transform 1 0 15552 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _004_
timestamp 1676381911
transform 1 0 13248 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _005_
timestamp 1676381911
transform 1 0 19488 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _006_
timestamp 1676381911
transform 1 0 18816 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _007_
timestamp 1676381911
transform 1 0 18432 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _008_
timestamp 1676381911
transform 1 0 20256 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _009_
timestamp 1676381911
transform 1 0 14304 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _010_
timestamp 1676381911
transform 1 0 21120 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _011_
timestamp 1676381911
transform 1 0 21504 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _012_
timestamp 1676381911
transform 1 0 22272 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _013_
timestamp 1676381911
transform 1 0 19872 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _014_
timestamp 1676381911
transform 1 0 15360 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _015_
timestamp 1676381911
transform 1 0 17280 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _016_
timestamp 1676381911
transform 1 0 21120 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _017_
timestamp 1676381911
transform 1 0 27360 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _018_
timestamp 1676381911
transform 1 0 20640 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _019_
timestamp 1676381911
transform 1 0 26208 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _020_
timestamp 1676381911
transform 1 0 24288 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _021_
timestamp 1676381911
transform 1 0 23904 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _022_
timestamp 1676381911
transform 1 0 31584 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _023_
timestamp 1676381911
transform 1 0 25536 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _024_
timestamp 1676381911
transform 1 0 31104 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _025_
timestamp 1676381911
transform 1 0 30720 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _026_
timestamp 1676381911
transform 1 0 32064 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _027_
timestamp 1676381911
transform 1 0 29952 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _028_
timestamp 1676381911
transform 1 0 30336 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _029_
timestamp 1676381911
transform 1 0 26112 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _030_
timestamp 1676381911
transform 1 0 29568 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _031_
timestamp 1676381911
transform 1 0 32448 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _032_
timestamp 1676381911
transform 1 0 3168 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _033_
timestamp 1676381911
transform 1 0 5280 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _034_
timestamp 1676381911
transform 1 0 8256 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _035_
timestamp 1676381911
transform 1 0 7872 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _036_
timestamp 1676381911
transform 1 0 21504 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _037_
timestamp 1676381911
transform -1 0 31104 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _038_
timestamp 1676381911
transform -1 0 29664 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _039_
timestamp 1676381911
transform 1 0 27744 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _040_
timestamp 1676381911
transform 1 0 25536 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _041_
timestamp 1676381911
transform 1 0 25152 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _042_
timestamp 1676381911
transform 1 0 26976 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _043_
timestamp 1676381911
transform 1 0 28512 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _044_
timestamp 1676381911
transform 1 0 29088 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _045_
timestamp 1676381911
transform 1 0 28896 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _046_
timestamp 1676381911
transform 1 0 28992 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _047_
timestamp 1676381911
transform 1 0 29760 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _048_
timestamp 1676381911
transform 1 0 29376 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _049_
timestamp 1676381911
transform 1 0 29568 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _050_
timestamp 1676381911
transform 1 0 29952 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _051_
timestamp 1676381911
transform 1 0 31008 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _052_
timestamp 1676381911
transform 1 0 5376 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _053_
timestamp 1676381911
transform 1 0 6144 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _054_
timestamp 1676381911
transform 1 0 6912 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _055_
timestamp 1676381911
transform 1 0 6528 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _056_
timestamp 1676381911
transform 1 0 5760 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _057_
timestamp 1676381911
transform 1 0 5760 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _058_
timestamp 1676381911
transform 1 0 6816 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _059_
timestamp 1676381911
transform 1 0 7584 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _060_
timestamp 1676381911
transform 1 0 7968 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _061_
timestamp 1676381911
transform 1 0 9120 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _062_
timestamp 1676381911
transform 1 0 8736 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _063_
timestamp 1676381911
transform 1 0 8352 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _064_
timestamp 1676381911
transform 1 0 7200 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _065_
timestamp 1676381911
transform 1 0 9312 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _066_
timestamp 1676381911
transform -1 0 11040 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _067_
timestamp 1676381911
transform -1 0 12096 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _068_
timestamp 1676381911
transform -1 0 12480 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _069_
timestamp 1676381911
transform -1 0 13248 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _070_
timestamp 1676381911
transform -1 0 14016 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _071_
timestamp 1676381911
transform -1 0 12864 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _072_
timestamp 1676381911
transform 1 0 8160 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _073_
timestamp 1676381911
transform 1 0 9984 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _074_
timestamp 1676381911
transform -1 0 12000 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _075_
timestamp 1676381911
transform -1 0 13632 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _076_
timestamp 1676381911
transform -1 0 14880 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _077_
timestamp 1676381911
transform -1 0 15360 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _078_
timestamp 1676381911
transform -1 0 15744 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _079_
timestamp 1676381911
transform -1 0 17472 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _080_
timestamp 1676381911
transform -1 0 16128 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _081_
timestamp 1676381911
transform -1 0 16896 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _082_
timestamp 1676381911
transform -1 0 17664 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _083_
timestamp 1676381911
transform -1 0 17280 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _084_
timestamp 1676381911
transform -1 0 18048 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _085_
timestamp 1676381911
transform -1 0 16512 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _086_
timestamp 1676381911
transform -1 0 17088 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _087_
timestamp 1676381911
transform -1 0 17088 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _088_
timestamp 1676381911
transform -1 0 27936 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _089_
timestamp 1676381911
transform -1 0 26880 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _090_
timestamp 1676381911
transform -1 0 25632 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _091_
timestamp 1676381911
transform -1 0 24288 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _092_
timestamp 1676381911
transform -1 0 23136 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _093_
timestamp 1676381911
transform -1 0 22272 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _094_
timestamp 1676381911
transform -1 0 21504 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _095_
timestamp 1676381911
transform -1 0 20832 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _096_
timestamp 1676381911
transform -1 0 19680 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _097_
timestamp 1676381911
transform -1 0 19296 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _098_
timestamp 1676381911
transform -1 0 18912 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _099_
timestamp 1676381911
transform -1 0 20352 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _100_
timestamp 1676381911
transform -1 0 19968 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _101_
timestamp 1676381911
transform -1 0 20160 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _102_
timestamp 1676381911
transform -1 0 20064 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _103_
timestamp 1676381911
transform -1 0 20448 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _104_
timestamp 1676381911
transform 1 0 3840 0 -1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 1152 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1824 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 2496 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 3168 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3840 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 4512 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 5184 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5856 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 6528 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 7200 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7872 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 8544 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 9216 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9888 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 10560 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 11232 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11904 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12576 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 13248 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13920 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14592 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 15264 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15936 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16608 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 17280 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 17952 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 18624 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 19296 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679581782
transform 1 0 19968 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679581782
transform 1 0 20640 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679581782
transform 1 0 21312 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679581782
transform 1 0 21984 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679581782
transform 1 0 22656 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679581782
transform 1 0 23328 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679581782
transform 1 0 24000 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679581782
transform 1 0 24672 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679581782
transform 1 0 25344 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1679581782
transform 1 0 26016 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1679581782
transform 1 0 26688 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1679581782
transform 1 0 27360 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1679581782
transform 1 0 28032 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1679581782
transform 1 0 28704 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1679581782
transform 1 0 29376 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1679581782
transform 1 0 30048 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1679581782
transform 1 0 30720 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_315
timestamp 1679581782
transform 1 0 31392 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_322
timestamp 1679581782
transform 1 0 32064 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_329
timestamp 1679581782
transform 1 0 32736 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_336
timestamp 1679581782
transform 1 0 33408 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_343
timestamp 1679581782
transform 1 0 34080 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_350
timestamp 1679581782
transform 1 0 34752 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_357
timestamp 1679581782
transform 1 0 35424 0 1 1512
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_364
timestamp 1677579658
transform 1 0 36096 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 1152 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1824 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 2496 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 3168 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3840 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 4512 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 5184 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5856 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 6528 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 7200 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_78
timestamp 1679581782
transform 1 0 8640 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_85
timestamp 1679581782
transform 1 0 9312 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_92
timestamp 1679581782
transform 1 0 9984 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_99
timestamp 1679581782
transform 1 0 10656 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_106
timestamp 1677579658
transform 1 0 11328 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_111
timestamp 1679581782
transform 1 0 11808 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_118
timestamp 1679581782
transform 1 0 12480 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_125
timestamp 1677579658
transform 1 0 13152 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_130
timestamp 1679581782
transform 1 0 13632 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_145
timestamp 1677580104
transform 1 0 15072 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_147
timestamp 1677579658
transform 1 0 15264 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_156
timestamp 1679581782
transform 1 0 16128 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_163
timestamp 1679577901
transform 1 0 16800 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_167
timestamp 1677579658
transform 1 0 17184 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_172
timestamp 1679581782
transform 1 0 17664 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_179
timestamp 1679581782
transform 1 0 18336 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_186
timestamp 1679581782
transform 1 0 19008 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_193
timestamp 1679581782
transform 1 0 19680 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_200
timestamp 1679581782
transform 1 0 20352 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_207
timestamp 1677579658
transform 1 0 21024 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_216
timestamp 1679581782
transform 1 0 21888 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_223
timestamp 1679581782
transform 1 0 22560 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_230
timestamp 1679581782
transform 1 0 23232 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_237
timestamp 1679581782
transform 1 0 23904 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_244
timestamp 1679577901
transform 1 0 24576 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_248
timestamp 1677580104
transform 1 0 24960 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_258
timestamp 1679581782
transform 1 0 25920 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_265
timestamp 1679577901
transform 1 0 26592 0 -1 3024
box -48 -56 432 834
use sg13g2_decap_8  FILLER_1_281
timestamp 1679581782
transform 1 0 28128 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_288
timestamp 1679577901
transform 1 0 28800 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_292
timestamp 1677579658
transform 1 0 29184 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_297
timestamp 1679581782
transform 1 0 29664 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_304
timestamp 1679577901
transform 1 0 30336 0 -1 3024
box -48 -56 432 834
use sg13g2_decap_8  FILLER_1_312
timestamp 1679581782
transform 1 0 31104 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_319
timestamp 1679581782
transform 1 0 31776 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_326
timestamp 1679581782
transform 1 0 32448 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_333
timestamp 1679581782
transform 1 0 33120 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_340
timestamp 1679581782
transform 1 0 33792 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_347
timestamp 1679581782
transform 1 0 34464 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_354
timestamp 1679581782
transform 1 0 35136 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_361
timestamp 1679581782
transform 1 0 35808 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_368
timestamp 1679577901
transform 1 0 36480 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_372
timestamp 1677579658
transform 1 0 36864 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679581782
transform 1 0 1152 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1679581782
transform 1 0 1824 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_14
timestamp 1679581782
transform 1 0 2496 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_21
timestamp 1679581782
transform 1 0 3168 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_28
timestamp 1679581782
transform 1 0 3840 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_35
timestamp 1679581782
transform 1 0 4512 0 1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_42
timestamp 1677579658
transform 1 0 5184 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_47
timestamp 1679581782
transform 1 0 5664 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_54
timestamp 1679581782
transform 1 0 6336 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_61
timestamp 1679581782
transform 1 0 7008 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_68
timestamp 1679581782
transform 1 0 7680 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_75
timestamp 1679581782
transform 1 0 8352 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_82
timestamp 1679581782
transform 1 0 9024 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_89
timestamp 1679581782
transform 1 0 9696 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_96
timestamp 1679581782
transform 1 0 10368 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_103
timestamp 1679581782
transform 1 0 11040 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_110
timestamp 1679581782
transform 1 0 11712 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_117
timestamp 1679581782
transform 1 0 12384 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_124
timestamp 1679581782
transform 1 0 13056 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_131
timestamp 1679581782
transform 1 0 13728 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_138
timestamp 1679581782
transform 1 0 14400 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_145
timestamp 1679577901
transform 1 0 15072 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_149
timestamp 1677579658
transform 1 0 15456 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_154
timestamp 1679581782
transform 1 0 15936 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_161
timestamp 1679581782
transform 1 0 16608 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_168
timestamp 1679581782
transform 1 0 17280 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_175
timestamp 1679577901
transform 1 0 17952 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_179
timestamp 1677579658
transform 1 0 18336 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_188
timestamp 1677580104
transform 1 0 19200 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_190
timestamp 1677579658
transform 1 0 19392 0 1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_207
timestamp 1677579658
transform 1 0 21024 0 1 3024
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_216
timestamp 1679577901
transform 1 0 21888 0 1 3024
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_224
timestamp 1679581782
transform 1 0 22656 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_231
timestamp 1679581782
transform 1 0 23328 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_238
timestamp 1679581782
transform 1 0 24000 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_245
timestamp 1679581782
transform 1 0 24672 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_252
timestamp 1679581782
transform 1 0 25344 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_259
timestamp 1677580104
transform 1 0 26016 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_265
timestamp 1679581782
transform 1 0 26592 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_272
timestamp 1679581782
transform 1 0 27264 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_279
timestamp 1679577901
transform 1 0 27936 0 1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_283
timestamp 1677580104
transform 1 0 28320 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_289
timestamp 1679581782
transform 1 0 28896 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_296
timestamp 1679581782
transform 1 0 29568 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_303
timestamp 1679581782
transform 1 0 30240 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_310
timestamp 1679581782
transform 1 0 30912 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_317
timestamp 1679581782
transform 1 0 31584 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_324
timestamp 1679581782
transform 1 0 32256 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_331
timestamp 1679581782
transform 1 0 32928 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_338
timestamp 1679581782
transform 1 0 33600 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_345
timestamp 1679581782
transform 1 0 34272 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_352
timestamp 1679581782
transform 1 0 34944 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_359
timestamp 1679581782
transform 1 0 35616 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_366
timestamp 1679581782
transform 1 0 36288 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_373
timestamp 1679577901
transform 1 0 36960 0 1 3024
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 1152 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_7
timestamp 1679581782
transform 1 0 1824 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1679581782
transform 1 0 2496 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_25
timestamp 1677580104
transform 1 0 3552 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_27
timestamp 1677579658
transform 1 0 3744 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_32
timestamp 1679581782
transform 1 0 4224 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_39
timestamp 1679581782
transform 1 0 4896 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_46
timestamp 1679581782
transform 1 0 5568 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_53
timestamp 1679581782
transform 1 0 6240 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_60
timestamp 1679581782
transform 1 0 6912 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_67
timestamp 1679577901
transform 1 0 7584 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_71
timestamp 1677580104
transform 1 0 7968 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_77
timestamp 1679581782
transform 1 0 8544 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_84
timestamp 1677579658
transform 1 0 9216 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_89
timestamp 1677580104
transform 1 0 9696 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_91
timestamp 1677579658
transform 1 0 9888 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_96
timestamp 1677580104
transform 1 0 10368 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_98
timestamp 1677579658
transform 1 0 10560 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_103
timestamp 1679577901
transform 1 0 11040 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_107
timestamp 1677580104
transform 1 0 11424 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_113
timestamp 1679581782
transform 1 0 12000 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_120
timestamp 1679581782
transform 1 0 12672 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_127
timestamp 1679581782
transform 1 0 13344 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_134
timestamp 1679581782
transform 1 0 14016 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_141
timestamp 1679581782
transform 1 0 14688 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_148
timestamp 1679581782
transform 1 0 15360 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_155
timestamp 1679581782
transform 1 0 16032 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_162
timestamp 1679581782
transform 1 0 16704 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_169
timestamp 1679581782
transform 1 0 17376 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_176
timestamp 1679581782
transform 1 0 18048 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_183
timestamp 1679581782
transform 1 0 18720 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_190
timestamp 1679581782
transform 1 0 19392 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_197
timestamp 1679581782
transform 1 0 20064 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_204
timestamp 1679581782
transform 1 0 20736 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_211
timestamp 1679581782
transform 1 0 21408 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_218
timestamp 1679581782
transform 1 0 22080 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_225
timestamp 1679581782
transform 1 0 22752 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_232
timestamp 1679581782
transform 1 0 23424 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_239
timestamp 1677580104
transform 1 0 24096 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_245
timestamp 1679581782
transform 1 0 24672 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_252
timestamp 1679581782
transform 1 0 25344 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_259
timestamp 1679581782
transform 1 0 26016 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_266
timestamp 1679581782
transform 1 0 26688 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_273
timestamp 1679581782
transform 1 0 27360 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_280
timestamp 1679581782
transform 1 0 28032 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_287
timestamp 1679577901
transform 1 0 28704 0 -1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_295
timestamp 1679581782
transform 1 0 29472 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_302
timestamp 1679581782
transform 1 0 30144 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_309
timestamp 1679581782
transform 1 0 30816 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_316
timestamp 1679581782
transform 1 0 31488 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_323
timestamp 1679581782
transform 1 0 32160 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_330
timestamp 1679581782
transform 1 0 32832 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_337
timestamp 1679581782
transform 1 0 33504 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_344
timestamp 1679581782
transform 1 0 34176 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_351
timestamp 1679581782
transform 1 0 34848 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_358
timestamp 1679581782
transform 1 0 35520 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_365
timestamp 1679581782
transform 1 0 36192 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_372
timestamp 1679577901
transform 1 0 36864 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_376
timestamp 1677579658
transform 1 0 37248 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679581782
transform 1 0 1152 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_7
timestamp 1679581782
transform 1 0 1824 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_14
timestamp 1679581782
transform 1 0 2496 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_21
timestamp 1679581782
transform 1 0 3168 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_28
timestamp 1679581782
transform 1 0 3840 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_35
timestamp 1679581782
transform 1 0 4512 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_42
timestamp 1679577901
transform 1 0 5184 0 1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_46
timestamp 1677580104
transform 1 0 5568 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_52
timestamp 1679581782
transform 1 0 6144 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_87
timestamp 1679581782
transform 1 0 9504 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_94
timestamp 1679581782
transform 1 0 10176 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_101
timestamp 1679581782
transform 1 0 10848 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_108
timestamp 1677580104
transform 1 0 11520 0 1 4536
box -48 -56 240 834
use sg13g2_decap_4  FILLER_4_134
timestamp 1679577901
transform 1 0 14016 0 1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_138
timestamp 1677579658
transform 1 0 14400 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_143
timestamp 1679581782
transform 1 0 14880 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_150
timestamp 1679581782
transform 1 0 15552 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_157
timestamp 1679577901
transform 1 0 16224 0 1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_161
timestamp 1677579658
transform 1 0 16608 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_170
timestamp 1679581782
transform 1 0 17472 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_177
timestamp 1679581782
transform 1 0 18144 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_184
timestamp 1679581782
transform 1 0 18816 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_191
timestamp 1679581782
transform 1 0 19488 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_198
timestamp 1679581782
transform 1 0 20160 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_205
timestamp 1679581782
transform 1 0 20832 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_212
timestamp 1679581782
transform 1 0 21504 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_219
timestamp 1679581782
transform 1 0 22176 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_226
timestamp 1679581782
transform 1 0 22848 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_233
timestamp 1679577901
transform 1 0 23520 0 1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_241
timestamp 1679581782
transform 1 0 24288 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_248
timestamp 1679581782
transform 1 0 24960 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_255
timestamp 1679581782
transform 1 0 25632 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_262
timestamp 1679581782
transform 1 0 26304 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_269
timestamp 1679581782
transform 1 0 26976 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_276
timestamp 1679581782
transform 1 0 27648 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_283
timestamp 1679577901
transform 1 0 28320 0 1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_287
timestamp 1677580104
transform 1 0 28704 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_293
timestamp 1679581782
transform 1 0 29280 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_300
timestamp 1679581782
transform 1 0 29952 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_307
timestamp 1679581782
transform 1 0 30624 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_314
timestamp 1679581782
transform 1 0 31296 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_321
timestamp 1679581782
transform 1 0 31968 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_328
timestamp 1679581782
transform 1 0 32640 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_335
timestamp 1679581782
transform 1 0 33312 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_342
timestamp 1679581782
transform 1 0 33984 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_349
timestamp 1679581782
transform 1 0 34656 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_356
timestamp 1679581782
transform 1 0 35328 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_363
timestamp 1679581782
transform 1 0 36000 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_370
timestamp 1679581782
transform 1 0 36672 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1679581782
transform 1 0 1152 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_7
timestamp 1679581782
transform 1 0 1824 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_14
timestamp 1679581782
transform 1 0 2496 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_21
timestamp 1679581782
transform 1 0 3168 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_28
timestamp 1679581782
transform 1 0 3840 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_35
timestamp 1679581782
transform 1 0 4512 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_42
timestamp 1677580104
transform 1 0 5184 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_64
timestamp 1679581782
transform 1 0 7296 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_71
timestamp 1679581782
transform 1 0 7968 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_78
timestamp 1679581782
transform 1 0 8640 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_85
timestamp 1679581782
transform 1 0 9312 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_92
timestamp 1679581782
transform 1 0 9984 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_99
timestamp 1679581782
transform 1 0 10656 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_106
timestamp 1679581782
transform 1 0 11328 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_113
timestamp 1679581782
transform 1 0 12000 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_120
timestamp 1679581782
transform 1 0 12672 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_127
timestamp 1679581782
transform 1 0 13344 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_134
timestamp 1679581782
transform 1 0 14016 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_141
timestamp 1677580104
transform 1 0 14688 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_143
timestamp 1677579658
transform 1 0 14880 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_176
timestamp 1679581782
transform 1 0 18048 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_183
timestamp 1679581782
transform 1 0 18720 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_190
timestamp 1679581782
transform 1 0 19392 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_197
timestamp 1679581782
transform 1 0 20064 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_204
timestamp 1679581782
transform 1 0 20736 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_211
timestamp 1679581782
transform 1 0 21408 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_218
timestamp 1679581782
transform 1 0 22080 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_225
timestamp 1679581782
transform 1 0 22752 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_232
timestamp 1679581782
transform 1 0 23424 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_239
timestamp 1679581782
transform 1 0 24096 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_246
timestamp 1679581782
transform 1 0 24768 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_253
timestamp 1679581782
transform 1 0 25440 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_260
timestamp 1679581782
transform 1 0 26112 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_267
timestamp 1679581782
transform 1 0 26784 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_274
timestamp 1679581782
transform 1 0 27456 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_281
timestamp 1679581782
transform 1 0 28128 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_288
timestamp 1677580104
transform 1 0 28800 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_294
timestamp 1679581782
transform 1 0 29376 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_301
timestamp 1679581782
transform 1 0 30048 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_308
timestamp 1679581782
transform 1 0 30720 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_315
timestamp 1679581782
transform 1 0 31392 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_322
timestamp 1679581782
transform 1 0 32064 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_329
timestamp 1679581782
transform 1 0 32736 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_336
timestamp 1679581782
transform 1 0 33408 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_343
timestamp 1679581782
transform 1 0 34080 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_350
timestamp 1679581782
transform 1 0 34752 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_357
timestamp 1679581782
transform 1 0 35424 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_364
timestamp 1679581782
transform 1 0 36096 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_371
timestamp 1679577901
transform 1 0 36768 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_375
timestamp 1677580104
transform 1 0 37152 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 1152 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1679581782
transform 1 0 1824 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_14
timestamp 1679581782
transform 1 0 2496 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_21
timestamp 1679581782
transform 1 0 3168 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_28
timestamp 1679581782
transform 1 0 3840 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_35
timestamp 1679581782
transform 1 0 4512 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_42
timestamp 1679581782
transform 1 0 5184 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_49
timestamp 1679581782
transform 1 0 5856 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_56
timestamp 1679581782
transform 1 0 6528 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_63
timestamp 1679581782
transform 1 0 7200 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_70
timestamp 1679581782
transform 1 0 7872 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_77
timestamp 1679581782
transform 1 0 8544 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_84
timestamp 1679581782
transform 1 0 9216 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_91
timestamp 1679581782
transform 1 0 9888 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_98
timestamp 1679581782
transform 1 0 10560 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_105
timestamp 1679581782
transform 1 0 11232 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_112
timestamp 1679581782
transform 1 0 11904 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_119
timestamp 1679581782
transform 1 0 12576 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_126
timestamp 1679581782
transform 1 0 13248 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_133
timestamp 1679581782
transform 1 0 13920 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_140
timestamp 1679581782
transform 1 0 14592 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_147
timestamp 1679581782
transform 1 0 15264 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_154
timestamp 1679581782
transform 1 0 15936 0 1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_161
timestamp 1677579658
transform 1 0 16608 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_166
timestamp 1679581782
transform 1 0 17088 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_173
timestamp 1679581782
transform 1 0 17760 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_180
timestamp 1679581782
transform 1 0 18432 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_187
timestamp 1679581782
transform 1 0 19104 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_198
timestamp 1679581782
transform 1 0 20160 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_205
timestamp 1679581782
transform 1 0 20832 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_212
timestamp 1679581782
transform 1 0 21504 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_219
timestamp 1679581782
transform 1 0 22176 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_226
timestamp 1679581782
transform 1 0 22848 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_233
timestamp 1679581782
transform 1 0 23520 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_240
timestamp 1679581782
transform 1 0 24192 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_247
timestamp 1679581782
transform 1 0 24864 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_254
timestamp 1679581782
transform 1 0 25536 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_261
timestamp 1679581782
transform 1 0 26208 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_268
timestamp 1679581782
transform 1 0 26880 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_275
timestamp 1679581782
transform 1 0 27552 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_282
timestamp 1679581782
transform 1 0 28224 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_289
timestamp 1679577901
transform 1 0 28896 0 1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_293
timestamp 1677579658
transform 1 0 29280 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_302
timestamp 1679581782
transform 1 0 30144 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_309
timestamp 1679581782
transform 1 0 30816 0 1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_316
timestamp 1677579658
transform 1 0 31488 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_321
timestamp 1679581782
transform 1 0 31968 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_328
timestamp 1679581782
transform 1 0 32640 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_335
timestamp 1679581782
transform 1 0 33312 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_342
timestamp 1679581782
transform 1 0 33984 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_349
timestamp 1679581782
transform 1 0 34656 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_356
timestamp 1679581782
transform 1 0 35328 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_363
timestamp 1679581782
transform 1 0 36000 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_370
timestamp 1679581782
transform 1 0 36672 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 1152 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1824 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 2496 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679581782
transform 1 0 3168 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679581782
transform 1 0 3840 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679581782
transform 1 0 4512 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679581782
transform 1 0 5184 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679581782
transform 1 0 5856 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_56
timestamp 1679581782
transform 1 0 6528 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_63
timestamp 1679581782
transform 1 0 7200 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_70
timestamp 1679581782
transform 1 0 7872 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_77
timestamp 1679581782
transform 1 0 8544 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_84
timestamp 1679581782
transform 1 0 9216 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_91
timestamp 1679581782
transform 1 0 9888 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_98
timestamp 1679581782
transform 1 0 10560 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_105
timestamp 1679581782
transform 1 0 11232 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_112
timestamp 1679581782
transform 1 0 11904 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_119
timestamp 1679581782
transform 1 0 12576 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_126
timestamp 1679581782
transform 1 0 13248 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_133
timestamp 1679581782
transform 1 0 13920 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_140
timestamp 1679581782
transform 1 0 14592 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_147
timestamp 1679581782
transform 1 0 15264 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_154
timestamp 1679581782
transform 1 0 15936 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_161
timestamp 1679581782
transform 1 0 16608 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_168
timestamp 1679581782
transform 1 0 17280 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_175
timestamp 1679577901
transform 1 0 17952 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_179
timestamp 1677580104
transform 1 0 18336 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_205
timestamp 1677580104
transform 1 0 20832 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_207
timestamp 1677579658
transform 1 0 21024 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_212
timestamp 1679581782
transform 1 0 21504 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_219
timestamp 1679581782
transform 1 0 22176 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_226
timestamp 1679581782
transform 1 0 22848 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_233
timestamp 1679581782
transform 1 0 23520 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_240
timestamp 1679581782
transform 1 0 24192 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_247
timestamp 1679581782
transform 1 0 24864 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_258
timestamp 1679581782
transform 1 0 25920 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_265
timestamp 1679581782
transform 1 0 26592 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_272
timestamp 1679581782
transform 1 0 27264 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_279
timestamp 1679581782
transform 1 0 27936 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_286
timestamp 1679581782
transform 1 0 28608 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_293
timestamp 1677580104
transform 1 0 29280 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_295
timestamp 1677579658
transform 1 0 29472 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_304
timestamp 1679581782
transform 1 0 30336 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_315
timestamp 1679581782
transform 1 0 31392 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_322
timestamp 1679581782
transform 1 0 32064 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_329
timestamp 1679581782
transform 1 0 32736 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_336
timestamp 1679581782
transform 1 0 33408 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_343
timestamp 1679581782
transform 1 0 34080 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_350
timestamp 1679581782
transform 1 0 34752 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_357
timestamp 1679581782
transform 1 0 35424 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_364
timestamp 1679581782
transform 1 0 36096 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_371
timestamp 1679577901
transform 1 0 36768 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_375
timestamp 1677580104
transform 1 0 37152 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1679581782
transform 1 0 1152 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_7
timestamp 1679581782
transform 1 0 1824 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_14
timestamp 1679581782
transform 1 0 2496 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_21
timestamp 1679581782
transform 1 0 3168 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_28
timestamp 1679581782
transform 1 0 3840 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_35
timestamp 1679581782
transform 1 0 4512 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_42
timestamp 1679581782
transform 1 0 5184 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_49
timestamp 1679581782
transform 1 0 5856 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_56
timestamp 1679581782
transform 1 0 6528 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_63
timestamp 1679581782
transform 1 0 7200 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_70
timestamp 1679581782
transform 1 0 7872 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_77
timestamp 1679581782
transform 1 0 8544 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_84
timestamp 1679581782
transform 1 0 9216 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_91
timestamp 1679581782
transform 1 0 9888 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_98
timestamp 1679581782
transform 1 0 10560 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_105
timestamp 1679581782
transform 1 0 11232 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_112
timestamp 1679581782
transform 1 0 11904 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_119
timestamp 1679581782
transform 1 0 12576 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_126
timestamp 1679581782
transform 1 0 13248 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_133
timestamp 1679581782
transform 1 0 13920 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_140
timestamp 1679581782
transform 1 0 14592 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_147
timestamp 1679581782
transform 1 0 15264 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_154
timestamp 1679581782
transform 1 0 15936 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_161
timestamp 1679581782
transform 1 0 16608 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_168
timestamp 1679581782
transform 1 0 17280 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_175
timestamp 1679581782
transform 1 0 17952 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_182
timestamp 1679581782
transform 1 0 18624 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_189
timestamp 1677580104
transform 1 0 19296 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_191
timestamp 1677579658
transform 1 0 19488 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_200
timestamp 1679581782
transform 1 0 20352 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_207
timestamp 1679581782
transform 1 0 21024 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_214
timestamp 1677580104
transform 1 0 21696 0 1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_220
timestamp 1679577901
transform 1 0 22272 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_224
timestamp 1677579658
transform 1 0 22656 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_229
timestamp 1679581782
transform 1 0 23136 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_236
timestamp 1677579658
transform 1 0 23808 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_241
timestamp 1679581782
transform 1 0 24288 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_248
timestamp 1677580104
transform 1 0 24960 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_250
timestamp 1677579658
transform 1 0 25152 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_255
timestamp 1679577901
transform 1 0 25632 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_259
timestamp 1677579658
transform 1 0 26016 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_268
timestamp 1679581782
transform 1 0 26880 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_279
timestamp 1679581782
transform 1 0 27936 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_286
timestamp 1679581782
transform 1 0 28608 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_293
timestamp 1677580104
transform 1 0 29280 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_295
timestamp 1677579658
transform 1 0 29472 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_316
timestamp 1679577901
transform 1 0 31488 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_320
timestamp 1677580104
transform 1 0 31872 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_326
timestamp 1679581782
transform 1 0 32448 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_333
timestamp 1679581782
transform 1 0 33120 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_340
timestamp 1679581782
transform 1 0 33792 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_347
timestamp 1679581782
transform 1 0 34464 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_354
timestamp 1679581782
transform 1 0 35136 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_361
timestamp 1679581782
transform 1 0 35808 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_368
timestamp 1679581782
transform 1 0 36480 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_375
timestamp 1677580104
transform 1 0 37152 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 1152 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_7
timestamp 1679581782
transform 1 0 1824 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_14
timestamp 1679581782
transform 1 0 2496 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_21
timestamp 1679581782
transform 1 0 3168 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_28
timestamp 1679581782
transform 1 0 3840 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_35
timestamp 1679581782
transform 1 0 4512 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_42
timestamp 1679581782
transform 1 0 5184 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_49
timestamp 1679581782
transform 1 0 5856 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_56
timestamp 1679581782
transform 1 0 6528 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_63
timestamp 1679577901
transform 1 0 7200 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_67
timestamp 1677580104
transform 1 0 7584 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_161
timestamp 1679581782
transform 1 0 16608 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_168
timestamp 1679581782
transform 1 0 17280 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_175
timestamp 1679581782
transform 1 0 17952 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_182
timestamp 1679581782
transform 1 0 18624 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_189
timestamp 1679581782
transform 1 0 19296 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_196
timestamp 1679581782
transform 1 0 19968 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_203
timestamp 1679581782
transform 1 0 20640 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_210
timestamp 1679581782
transform 1 0 21312 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_217
timestamp 1679581782
transform 1 0 21984 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_224
timestamp 1679581782
transform 1 0 22656 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_231
timestamp 1679581782
transform 1 0 23328 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_238
timestamp 1679581782
transform 1 0 24000 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_245
timestamp 1679581782
transform 1 0 24672 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_252
timestamp 1679581782
transform 1 0 25344 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_259
timestamp 1679581782
transform 1 0 26016 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_266
timestamp 1679581782
transform 1 0 26688 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_273
timestamp 1679581782
transform 1 0 27360 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_280
timestamp 1679577901
transform 1 0 28032 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_284
timestamp 1677579658
transform 1 0 28416 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_317
timestamp 1679581782
transform 1 0 31584 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_324
timestamp 1677580104
transform 1 0 32256 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_330
timestamp 1679581782
transform 1 0 32832 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_337
timestamp 1679581782
transform 1 0 33504 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_344
timestamp 1679581782
transform 1 0 34176 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_351
timestamp 1679581782
transform 1 0 34848 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_358
timestamp 1679581782
transform 1 0 35520 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_365
timestamp 1679577901
transform 1 0 36192 0 -1 9072
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_0
timestamp 1679581782
transform 1 0 1152 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_7
timestamp 1679581782
transform 1 0 1824 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_14
timestamp 1679581782
transform 1 0 2496 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_21
timestamp 1679581782
transform 1 0 3168 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_28
timestamp 1679581782
transform 1 0 3840 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_35
timestamp 1679581782
transform 1 0 4512 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_42
timestamp 1679581782
transform 1 0 5184 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_49
timestamp 1679581782
transform 1 0 5856 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_56
timestamp 1679577901
transform 1 0 6528 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_60
timestamp 1677579658
transform 1 0 6912 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_177
timestamp 1679581782
transform 1 0 18144 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_184
timestamp 1679581782
transform 1 0 18816 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_191
timestamp 1679581782
transform 1 0 19488 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_198
timestamp 1679581782
transform 1 0 20160 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_205
timestamp 1679581782
transform 1 0 20832 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_212
timestamp 1679581782
transform 1 0 21504 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_219
timestamp 1679581782
transform 1 0 22176 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_226
timestamp 1679581782
transform 1 0 22848 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_233
timestamp 1679581782
transform 1 0 23520 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_240
timestamp 1679581782
transform 1 0 24192 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_247
timestamp 1679581782
transform 1 0 24864 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_254
timestamp 1679581782
transform 1 0 25536 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_261
timestamp 1679581782
transform 1 0 26208 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_268
timestamp 1679581782
transform 1 0 26880 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_327
timestamp 1679581782
transform 1 0 32544 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_334
timestamp 1679581782
transform 1 0 33216 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_341
timestamp 1679581782
transform 1 0 33888 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_348
timestamp 1679581782
transform 1 0 34560 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_355
timestamp 1679577901
transform 1 0 35232 0 1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_359
timestamp 1677580104
transform 1 0 35616 0 1 9072
box -48 -56 240 834
use sg13g2_buf_1  output1
timestamp 1676381911
transform 1 0 36960 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output2
timestamp 1676381911
transform 1 0 37344 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output3
timestamp 1676381911
transform 1 0 37728 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output4
timestamp 1676381911
transform 1 0 37344 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output5
timestamp 1676381911
transform 1 0 37728 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output6
timestamp 1676381911
transform 1 0 37344 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676381911
transform 1 0 37728 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform 1 0 37344 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform 1 0 37728 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676381911
transform 1 0 37344 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676381911
transform 1 0 37728 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676381911
transform 1 0 36576 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676381911
transform 1 0 37728 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output14
timestamp 1676381911
transform 1 0 37344 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output15
timestamp 1676381911
transform 1 0 37728 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output16
timestamp 1676381911
transform 1 0 37344 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676381911
transform 1 0 37728 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676381911
transform 1 0 37344 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output19
timestamp 1676381911
transform 1 0 36960 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output20
timestamp 1676381911
transform 1 0 36576 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output21
timestamp 1676381911
transform 1 0 36960 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output22
timestamp 1676381911
transform 1 0 36192 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output23
timestamp 1676381911
transform 1 0 36192 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output24
timestamp 1676381911
transform 1 0 35808 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output25
timestamp 1676381911
transform 1 0 36576 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output26
timestamp 1676381911
transform 1 0 37344 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output27
timestamp 1676381911
transform 1 0 36960 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output28
timestamp 1676381911
transform 1 0 37728 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output29
timestamp 1676381911
transform 1 0 37344 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output30
timestamp 1676381911
transform 1 0 37728 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output31
timestamp 1676381911
transform 1 0 37344 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output32
timestamp 1676381911
transform 1 0 37728 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output33
timestamp 1676381911
transform -1 0 28320 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output34
timestamp 1676381911
transform -1 0 30048 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output35
timestamp 1676381911
transform -1 0 31008 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output36
timestamp 1676381911
transform -1 0 30432 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output37
timestamp 1676381911
transform -1 0 31392 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output38
timestamp 1676381911
transform -1 0 30816 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output39
timestamp 1676381911
transform -1 0 31776 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output40
timestamp 1676381911
transform -1 0 31200 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output41
timestamp 1676381911
transform -1 0 32160 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output42
timestamp 1676381911
transform -1 0 31584 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output43
timestamp 1676381911
transform -1 0 32544 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output44
timestamp 1676381911
transform -1 0 28704 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output45
timestamp 1676381911
transform -1 0 29088 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output46
timestamp 1676381911
transform -1 0 29472 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output47
timestamp 1676381911
transform -1 0 28896 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output48
timestamp 1676381911
transform -1 0 29856 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output49
timestamp 1676381911
transform -1 0 29280 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output50
timestamp 1676381911
transform -1 0 30240 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output51
timestamp 1676381911
transform -1 0 29664 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output52
timestamp 1676381911
transform -1 0 30624 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output53
timestamp 1676381911
transform 1 0 7008 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output54
timestamp 1676381911
transform -1 0 8160 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output55
timestamp 1676381911
transform 1 0 7392 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output56
timestamp 1676381911
transform -1 0 8544 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output57
timestamp 1676381911
transform 1 0 7776 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output58
timestamp 1676381911
transform -1 0 8928 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output59
timestamp 1676381911
transform 1 0 8160 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output60
timestamp 1676381911
transform -1 0 9312 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output61
timestamp 1676381911
transform 1 0 8544 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output62
timestamp 1676381911
transform -1 0 9696 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output63
timestamp 1676381911
transform 1 0 8928 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output64
timestamp 1676381911
transform -1 0 10080 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output65
timestamp 1676381911
transform 1 0 9312 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output66
timestamp 1676381911
transform -1 0 10464 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output67
timestamp 1676381911
transform 1 0 9696 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output68
timestamp 1676381911
transform -1 0 10848 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output69
timestamp 1676381911
transform 1 0 10080 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output70
timestamp 1676381911
transform -1 0 11232 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output71
timestamp 1676381911
transform 1 0 10464 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output72
timestamp 1676381911
transform -1 0 11616 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output73
timestamp 1676381911
transform 1 0 10848 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output74
timestamp 1676381911
transform 1 0 12768 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output75
timestamp 1676381911
transform -1 0 13920 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output76
timestamp 1676381911
transform 1 0 13152 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output77
timestamp 1676381911
transform -1 0 14304 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output78
timestamp 1676381911
transform 1 0 13536 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output79
timestamp 1676381911
transform -1 0 14688 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output80
timestamp 1676381911
transform -1 0 12000 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output81
timestamp 1676381911
transform 1 0 11232 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output82
timestamp 1676381911
transform -1 0 12384 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output83
timestamp 1676381911
transform 1 0 11616 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output84
timestamp 1676381911
transform -1 0 12768 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output85
timestamp 1676381911
transform 1 0 12000 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output86
timestamp 1676381911
transform -1 0 13152 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output87
timestamp 1676381911
transform 1 0 12384 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output88
timestamp 1676381911
transform -1 0 13536 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output89
timestamp 1676381911
transform 1 0 13920 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output90
timestamp 1676381911
transform 1 0 15840 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output91
timestamp 1676381911
transform 1 0 16224 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output92
timestamp 1676381911
transform -1 0 16992 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output93
timestamp 1676381911
transform -1 0 17376 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output94
timestamp 1676381911
transform -1 0 18144 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output95
timestamp 1676381911
transform -1 0 17760 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output96
timestamp 1676381911
transform -1 0 15072 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output97
timestamp 1676381911
transform 1 0 14304 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output98
timestamp 1676381911
transform -1 0 15456 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output99
timestamp 1676381911
transform 1 0 14688 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output100
timestamp 1676381911
transform -1 0 15840 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output101
timestamp 1676381911
transform 1 0 15072 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output102
timestamp 1676381911
transform -1 0 16224 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output103
timestamp 1676381911
transform 1 0 15456 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output104
timestamp 1676381911
transform -1 0 16608 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output105
timestamp 1676381911
transform -1 0 27936 0 1 9072
box -48 -56 432 834
<< labels >>
flabel metal2 s 0 548 90 628 0 FreeSans 320 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal2 s 0 3908 90 3988 0 FreeSans 320 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal2 s 0 4244 90 4324 0 FreeSans 320 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal2 s 0 4580 90 4660 0 FreeSans 320 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal2 s 0 4916 90 4996 0 FreeSans 320 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal2 s 0 5252 90 5332 0 FreeSans 320 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal2 s 0 5588 90 5668 0 FreeSans 320 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal2 s 0 5924 90 6004 0 FreeSans 320 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal2 s 0 6260 90 6340 0 FreeSans 320 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal2 s 0 6596 90 6676 0 FreeSans 320 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal2 s 0 6932 90 7012 0 FreeSans 320 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal2 s 0 884 90 964 0 FreeSans 320 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal2 s 0 7268 90 7348 0 FreeSans 320 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal2 s 0 7604 90 7684 0 FreeSans 320 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal2 s 0 7940 90 8020 0 FreeSans 320 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal2 s 0 8276 90 8356 0 FreeSans 320 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal2 s 0 8612 90 8692 0 FreeSans 320 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal2 s 0 8948 90 9028 0 FreeSans 320 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal2 s 0 9284 90 9364 0 FreeSans 320 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal2 s 0 9620 90 9700 0 FreeSans 320 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal2 s 0 9956 90 10036 0 FreeSans 320 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal2 s 0 10292 90 10372 0 FreeSans 320 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal2 s 0 1220 90 1300 0 FreeSans 320 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal2 s 0 10628 90 10708 0 FreeSans 320 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal2 s 0 10964 90 11044 0 FreeSans 320 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal2 s 0 1556 90 1636 0 FreeSans 320 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal2 s 0 1892 90 1972 0 FreeSans 320 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal2 s 0 2228 90 2308 0 FreeSans 320 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal2 s 0 2564 90 2644 0 FreeSans 320 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal2 s 0 2900 90 2980 0 FreeSans 320 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal2 s 0 3236 90 3316 0 FreeSans 320 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal2 s 0 3572 90 3652 0 FreeSans 320 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal2 s 39174 548 39264 628 0 FreeSans 320 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal2 s 39174 3908 39264 3988 0 FreeSans 320 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal2 s 39174 4244 39264 4324 0 FreeSans 320 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal2 s 39174 4580 39264 4660 0 FreeSans 320 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal2 s 39174 4916 39264 4996 0 FreeSans 320 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal2 s 39174 5252 39264 5332 0 FreeSans 320 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal2 s 39174 5588 39264 5668 0 FreeSans 320 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal2 s 39174 5924 39264 6004 0 FreeSans 320 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal2 s 39174 6260 39264 6340 0 FreeSans 320 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal2 s 39174 6596 39264 6676 0 FreeSans 320 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal2 s 39174 6932 39264 7012 0 FreeSans 320 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal2 s 39174 884 39264 964 0 FreeSans 320 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal2 s 39174 7268 39264 7348 0 FreeSans 320 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal2 s 39174 7604 39264 7684 0 FreeSans 320 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal2 s 39174 7940 39264 8020 0 FreeSans 320 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal2 s 39174 8276 39264 8356 0 FreeSans 320 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal2 s 39174 8612 39264 8692 0 FreeSans 320 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal2 s 39174 8948 39264 9028 0 FreeSans 320 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal2 s 39174 9284 39264 9364 0 FreeSans 320 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal2 s 39174 9620 39264 9700 0 FreeSans 320 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal2 s 39174 9956 39264 10036 0 FreeSans 320 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal2 s 39174 10292 39264 10372 0 FreeSans 320 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal2 s 39174 1220 39264 1300 0 FreeSans 320 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal2 s 39174 10628 39264 10708 0 FreeSans 320 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal2 s 39174 10964 39264 11044 0 FreeSans 320 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal2 s 39174 1556 39264 1636 0 FreeSans 320 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal2 s 39174 1892 39264 1972 0 FreeSans 320 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal2 s 39174 2228 39264 2308 0 FreeSans 320 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal2 s 39174 2564 39264 2644 0 FreeSans 320 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal2 s 39174 2900 39264 2980 0 FreeSans 320 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal2 s 39174 3236 39264 3316 0 FreeSans 320 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal2 s 39174 3572 39264 3652 0 FreeSans 320 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal3 s 3896 0 3976 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal3 s 21176 0 21256 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal3 s 22904 0 22984 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal3 s 24632 0 24712 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal3 s 26360 0 26440 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal3 s 28088 0 28168 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal3 s 29816 0 29896 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal3 s 31544 0 31624 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal3 s 33272 0 33352 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal3 s 35000 0 35080 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal3 s 36728 0 36808 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal3 s 5624 0 5704 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal3 s 7352 0 7432 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal3 s 9080 0 9160 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal3 s 10808 0 10888 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal3 s 12536 0 12616 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal3 s 14264 0 14344 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal3 s 15992 0 16072 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal3 s 17720 0 17800 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal3 s 19448 0 19528 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal3 s 27704 11764 27784 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal3 s 29624 11764 29704 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal3 s 29816 11764 29896 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal3 s 30008 11764 30088 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal3 s 30200 11764 30280 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal3 s 30392 11764 30472 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal3 s 30584 11764 30664 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal3 s 30776 11764 30856 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal3 s 30968 11764 31048 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal3 s 31160 11764 31240 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal3 s 31352 11764 31432 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal3 s 27896 11764 27976 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal3 s 28088 11764 28168 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal3 s 28280 11764 28360 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal3 s 28472 11764 28552 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal3 s 28664 11764 28744 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal3 s 28856 11764 28936 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal3 s 29048 11764 29128 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal3 s 29240 11764 29320 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal3 s 29432 11764 29512 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal3 s 7544 11764 7624 11844 0 FreeSans 320 0 0 0 N1BEG[0]
port 104 nsew signal output
flabel metal3 s 7736 11764 7816 11844 0 FreeSans 320 0 0 0 N1BEG[1]
port 105 nsew signal output
flabel metal3 s 7928 11764 8008 11844 0 FreeSans 320 0 0 0 N1BEG[2]
port 106 nsew signal output
flabel metal3 s 8120 11764 8200 11844 0 FreeSans 320 0 0 0 N1BEG[3]
port 107 nsew signal output
flabel metal3 s 8312 11764 8392 11844 0 FreeSans 320 0 0 0 N2BEG[0]
port 108 nsew signal output
flabel metal3 s 8504 11764 8584 11844 0 FreeSans 320 0 0 0 N2BEG[1]
port 109 nsew signal output
flabel metal3 s 8696 11764 8776 11844 0 FreeSans 320 0 0 0 N2BEG[2]
port 110 nsew signal output
flabel metal3 s 8888 11764 8968 11844 0 FreeSans 320 0 0 0 N2BEG[3]
port 111 nsew signal output
flabel metal3 s 9080 11764 9160 11844 0 FreeSans 320 0 0 0 N2BEG[4]
port 112 nsew signal output
flabel metal3 s 9272 11764 9352 11844 0 FreeSans 320 0 0 0 N2BEG[5]
port 113 nsew signal output
flabel metal3 s 9464 11764 9544 11844 0 FreeSans 320 0 0 0 N2BEG[6]
port 114 nsew signal output
flabel metal3 s 9656 11764 9736 11844 0 FreeSans 320 0 0 0 N2BEG[7]
port 115 nsew signal output
flabel metal3 s 9848 11764 9928 11844 0 FreeSans 320 0 0 0 N2BEGb[0]
port 116 nsew signal output
flabel metal3 s 10040 11764 10120 11844 0 FreeSans 320 0 0 0 N2BEGb[1]
port 117 nsew signal output
flabel metal3 s 10232 11764 10312 11844 0 FreeSans 320 0 0 0 N2BEGb[2]
port 118 nsew signal output
flabel metal3 s 10424 11764 10504 11844 0 FreeSans 320 0 0 0 N2BEGb[3]
port 119 nsew signal output
flabel metal3 s 10616 11764 10696 11844 0 FreeSans 320 0 0 0 N2BEGb[4]
port 120 nsew signal output
flabel metal3 s 10808 11764 10888 11844 0 FreeSans 320 0 0 0 N2BEGb[5]
port 121 nsew signal output
flabel metal3 s 11000 11764 11080 11844 0 FreeSans 320 0 0 0 N2BEGb[6]
port 122 nsew signal output
flabel metal3 s 11192 11764 11272 11844 0 FreeSans 320 0 0 0 N2BEGb[7]
port 123 nsew signal output
flabel metal3 s 11384 11764 11464 11844 0 FreeSans 320 0 0 0 N4BEG[0]
port 124 nsew signal output
flabel metal3 s 13304 11764 13384 11844 0 FreeSans 320 0 0 0 N4BEG[10]
port 125 nsew signal output
flabel metal3 s 13496 11764 13576 11844 0 FreeSans 320 0 0 0 N4BEG[11]
port 126 nsew signal output
flabel metal3 s 13688 11764 13768 11844 0 FreeSans 320 0 0 0 N4BEG[12]
port 127 nsew signal output
flabel metal3 s 13880 11764 13960 11844 0 FreeSans 320 0 0 0 N4BEG[13]
port 128 nsew signal output
flabel metal3 s 14072 11764 14152 11844 0 FreeSans 320 0 0 0 N4BEG[14]
port 129 nsew signal output
flabel metal3 s 14264 11764 14344 11844 0 FreeSans 320 0 0 0 N4BEG[15]
port 130 nsew signal output
flabel metal3 s 11576 11764 11656 11844 0 FreeSans 320 0 0 0 N4BEG[1]
port 131 nsew signal output
flabel metal3 s 11768 11764 11848 11844 0 FreeSans 320 0 0 0 N4BEG[2]
port 132 nsew signal output
flabel metal3 s 11960 11764 12040 11844 0 FreeSans 320 0 0 0 N4BEG[3]
port 133 nsew signal output
flabel metal3 s 12152 11764 12232 11844 0 FreeSans 320 0 0 0 N4BEG[4]
port 134 nsew signal output
flabel metal3 s 12344 11764 12424 11844 0 FreeSans 320 0 0 0 N4BEG[5]
port 135 nsew signal output
flabel metal3 s 12536 11764 12616 11844 0 FreeSans 320 0 0 0 N4BEG[6]
port 136 nsew signal output
flabel metal3 s 12728 11764 12808 11844 0 FreeSans 320 0 0 0 N4BEG[7]
port 137 nsew signal output
flabel metal3 s 12920 11764 13000 11844 0 FreeSans 320 0 0 0 N4BEG[8]
port 138 nsew signal output
flabel metal3 s 13112 11764 13192 11844 0 FreeSans 320 0 0 0 N4BEG[9]
port 139 nsew signal output
flabel metal3 s 14456 11764 14536 11844 0 FreeSans 320 0 0 0 NN4BEG[0]
port 140 nsew signal output
flabel metal3 s 16376 11764 16456 11844 0 FreeSans 320 0 0 0 NN4BEG[10]
port 141 nsew signal output
flabel metal3 s 16568 11764 16648 11844 0 FreeSans 320 0 0 0 NN4BEG[11]
port 142 nsew signal output
flabel metal3 s 16760 11764 16840 11844 0 FreeSans 320 0 0 0 NN4BEG[12]
port 143 nsew signal output
flabel metal3 s 16952 11764 17032 11844 0 FreeSans 320 0 0 0 NN4BEG[13]
port 144 nsew signal output
flabel metal3 s 17144 11764 17224 11844 0 FreeSans 320 0 0 0 NN4BEG[14]
port 145 nsew signal output
flabel metal3 s 17336 11764 17416 11844 0 FreeSans 320 0 0 0 NN4BEG[15]
port 146 nsew signal output
flabel metal3 s 14648 11764 14728 11844 0 FreeSans 320 0 0 0 NN4BEG[1]
port 147 nsew signal output
flabel metal3 s 14840 11764 14920 11844 0 FreeSans 320 0 0 0 NN4BEG[2]
port 148 nsew signal output
flabel metal3 s 15032 11764 15112 11844 0 FreeSans 320 0 0 0 NN4BEG[3]
port 149 nsew signal output
flabel metal3 s 15224 11764 15304 11844 0 FreeSans 320 0 0 0 NN4BEG[4]
port 150 nsew signal output
flabel metal3 s 15416 11764 15496 11844 0 FreeSans 320 0 0 0 NN4BEG[5]
port 151 nsew signal output
flabel metal3 s 15608 11764 15688 11844 0 FreeSans 320 0 0 0 NN4BEG[6]
port 152 nsew signal output
flabel metal3 s 15800 11764 15880 11844 0 FreeSans 320 0 0 0 NN4BEG[7]
port 153 nsew signal output
flabel metal3 s 15992 11764 16072 11844 0 FreeSans 320 0 0 0 NN4BEG[8]
port 154 nsew signal output
flabel metal3 s 16184 11764 16264 11844 0 FreeSans 320 0 0 0 NN4BEG[9]
port 155 nsew signal output
flabel metal3 s 17528 11764 17608 11844 0 FreeSans 320 0 0 0 S1END[0]
port 156 nsew signal input
flabel metal3 s 17720 11764 17800 11844 0 FreeSans 320 0 0 0 S1END[1]
port 157 nsew signal input
flabel metal3 s 17912 11764 17992 11844 0 FreeSans 320 0 0 0 S1END[2]
port 158 nsew signal input
flabel metal3 s 18104 11764 18184 11844 0 FreeSans 320 0 0 0 S1END[3]
port 159 nsew signal input
flabel metal3 s 19832 11764 19912 11844 0 FreeSans 320 0 0 0 S2END[0]
port 160 nsew signal input
flabel metal3 s 20024 11764 20104 11844 0 FreeSans 320 0 0 0 S2END[1]
port 161 nsew signal input
flabel metal3 s 20216 11764 20296 11844 0 FreeSans 320 0 0 0 S2END[2]
port 162 nsew signal input
flabel metal3 s 20408 11764 20488 11844 0 FreeSans 320 0 0 0 S2END[3]
port 163 nsew signal input
flabel metal3 s 20600 11764 20680 11844 0 FreeSans 320 0 0 0 S2END[4]
port 164 nsew signal input
flabel metal3 s 20792 11764 20872 11844 0 FreeSans 320 0 0 0 S2END[5]
port 165 nsew signal input
flabel metal3 s 20984 11764 21064 11844 0 FreeSans 320 0 0 0 S2END[6]
port 166 nsew signal input
flabel metal3 s 21176 11764 21256 11844 0 FreeSans 320 0 0 0 S2END[7]
port 167 nsew signal input
flabel metal3 s 18296 11764 18376 11844 0 FreeSans 320 0 0 0 S2MID[0]
port 168 nsew signal input
flabel metal3 s 18488 11764 18568 11844 0 FreeSans 320 0 0 0 S2MID[1]
port 169 nsew signal input
flabel metal3 s 18680 11764 18760 11844 0 FreeSans 320 0 0 0 S2MID[2]
port 170 nsew signal input
flabel metal3 s 18872 11764 18952 11844 0 FreeSans 320 0 0 0 S2MID[3]
port 171 nsew signal input
flabel metal3 s 19064 11764 19144 11844 0 FreeSans 320 0 0 0 S2MID[4]
port 172 nsew signal input
flabel metal3 s 19256 11764 19336 11844 0 FreeSans 320 0 0 0 S2MID[5]
port 173 nsew signal input
flabel metal3 s 19448 11764 19528 11844 0 FreeSans 320 0 0 0 S2MID[6]
port 174 nsew signal input
flabel metal3 s 19640 11764 19720 11844 0 FreeSans 320 0 0 0 S2MID[7]
port 175 nsew signal input
flabel metal3 s 21368 11764 21448 11844 0 FreeSans 320 0 0 0 S4END[0]
port 176 nsew signal input
flabel metal3 s 23288 11764 23368 11844 0 FreeSans 320 0 0 0 S4END[10]
port 177 nsew signal input
flabel metal3 s 23480 11764 23560 11844 0 FreeSans 320 0 0 0 S4END[11]
port 178 nsew signal input
flabel metal3 s 23672 11764 23752 11844 0 FreeSans 320 0 0 0 S4END[12]
port 179 nsew signal input
flabel metal3 s 23864 11764 23944 11844 0 FreeSans 320 0 0 0 S4END[13]
port 180 nsew signal input
flabel metal3 s 24056 11764 24136 11844 0 FreeSans 320 0 0 0 S4END[14]
port 181 nsew signal input
flabel metal3 s 24248 11764 24328 11844 0 FreeSans 320 0 0 0 S4END[15]
port 182 nsew signal input
flabel metal3 s 21560 11764 21640 11844 0 FreeSans 320 0 0 0 S4END[1]
port 183 nsew signal input
flabel metal3 s 21752 11764 21832 11844 0 FreeSans 320 0 0 0 S4END[2]
port 184 nsew signal input
flabel metal3 s 21944 11764 22024 11844 0 FreeSans 320 0 0 0 S4END[3]
port 185 nsew signal input
flabel metal3 s 22136 11764 22216 11844 0 FreeSans 320 0 0 0 S4END[4]
port 186 nsew signal input
flabel metal3 s 22328 11764 22408 11844 0 FreeSans 320 0 0 0 S4END[5]
port 187 nsew signal input
flabel metal3 s 22520 11764 22600 11844 0 FreeSans 320 0 0 0 S4END[6]
port 188 nsew signal input
flabel metal3 s 22712 11764 22792 11844 0 FreeSans 320 0 0 0 S4END[7]
port 189 nsew signal input
flabel metal3 s 22904 11764 22984 11844 0 FreeSans 320 0 0 0 S4END[8]
port 190 nsew signal input
flabel metal3 s 23096 11764 23176 11844 0 FreeSans 320 0 0 0 S4END[9]
port 191 nsew signal input
flabel metal3 s 24440 11764 24520 11844 0 FreeSans 320 0 0 0 SS4END[0]
port 192 nsew signal input
flabel metal3 s 26360 11764 26440 11844 0 FreeSans 320 0 0 0 SS4END[10]
port 193 nsew signal input
flabel metal3 s 26552 11764 26632 11844 0 FreeSans 320 0 0 0 SS4END[11]
port 194 nsew signal input
flabel metal3 s 26744 11764 26824 11844 0 FreeSans 320 0 0 0 SS4END[12]
port 195 nsew signal input
flabel metal3 s 26936 11764 27016 11844 0 FreeSans 320 0 0 0 SS4END[13]
port 196 nsew signal input
flabel metal3 s 27128 11764 27208 11844 0 FreeSans 320 0 0 0 SS4END[14]
port 197 nsew signal input
flabel metal3 s 27320 11764 27400 11844 0 FreeSans 320 0 0 0 SS4END[15]
port 198 nsew signal input
flabel metal3 s 24632 11764 24712 11844 0 FreeSans 320 0 0 0 SS4END[1]
port 199 nsew signal input
flabel metal3 s 24824 11764 24904 11844 0 FreeSans 320 0 0 0 SS4END[2]
port 200 nsew signal input
flabel metal3 s 25016 11764 25096 11844 0 FreeSans 320 0 0 0 SS4END[3]
port 201 nsew signal input
flabel metal3 s 25208 11764 25288 11844 0 FreeSans 320 0 0 0 SS4END[4]
port 202 nsew signal input
flabel metal3 s 25400 11764 25480 11844 0 FreeSans 320 0 0 0 SS4END[5]
port 203 nsew signal input
flabel metal3 s 25592 11764 25672 11844 0 FreeSans 320 0 0 0 SS4END[6]
port 204 nsew signal input
flabel metal3 s 25784 11764 25864 11844 0 FreeSans 320 0 0 0 SS4END[7]
port 205 nsew signal input
flabel metal3 s 25976 11764 26056 11844 0 FreeSans 320 0 0 0 SS4END[8]
port 206 nsew signal input
flabel metal3 s 26168 11764 26248 11844 0 FreeSans 320 0 0 0 SS4END[9]
port 207 nsew signal input
flabel metal3 s 2168 0 2248 80 0 FreeSans 320 0 0 0 UserCLK
port 208 nsew signal input
flabel metal3 s 27512 11764 27592 11844 0 FreeSans 320 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal5 s 4892 0 5332 11844 0 FreeSans 2560 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 4892 0 5332 40 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 4892 11804 5332 11844 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 20012 0 20452 11844 0 FreeSans 2560 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 20012 0 20452 40 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 20012 11804 20452 11844 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 35132 0 35572 11844 0 FreeSans 2560 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 35132 0 35572 40 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 35132 11804 35572 11844 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 3652 0 4092 11844 0 FreeSans 2560 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 3652 0 4092 40 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 3652 11804 4092 11844 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 18772 0 19212 11844 0 FreeSans 2560 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 18772 0 19212 40 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 18772 11804 19212 11844 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 33892 0 34332 11844 0 FreeSans 2560 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 33892 0 34332 40 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 33892 11804 34332 11844 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
rlabel metal1 19632 9072 19632 9072 0 VGND
rlabel metal1 19632 9828 19632 9828 0 VPWR
rlabel metal3 11520 1596 11520 1596 0 FrameData[0]
rlabel metal3 21216 3654 21216 3654 0 FrameData[10]
rlabel metal3 21600 3822 21600 3822 0 FrameData[11]
rlabel metal2 176 4620 176 4620 0 FrameData[12]
rlabel metal3 19968 3738 19968 3738 0 FrameData[13]
rlabel metal2 848 5292 848 5292 0 FrameData[14]
rlabel metal3 17376 2394 17376 2394 0 FrameData[15]
rlabel metal2 752 5964 752 5964 0 FrameData[16]
rlabel metal2 416 6300 416 6300 0 FrameData[17]
rlabel metal2 656 6636 656 6636 0 FrameData[18]
rlabel metal2 608 6972 608 6972 0 FrameData[19]
rlabel metal3 14784 1764 14784 1764 0 FrameData[1]
rlabel metal2 24384 4158 24384 4158 0 FrameData[20]
rlabel metal2 560 7644 560 7644 0 FrameData[21]
rlabel metal2 752 7980 752 7980 0 FrameData[22]
rlabel metal3 25632 6636 25632 6636 0 FrameData[23]
rlabel metal2 656 8652 656 8652 0 FrameData[24]
rlabel metal2 752 8988 752 8988 0 FrameData[25]
rlabel metal2 608 9324 608 9324 0 FrameData[26]
rlabel metal2 512 9660 512 9660 0 FrameData[27]
rlabel metal2 560 9996 560 9996 0 FrameData[28]
rlabel metal2 704 10332 704 10332 0 FrameData[29]
rlabel metal3 15840 1932 15840 1932 0 FrameData[2]
rlabel metal2 368 10668 368 10668 0 FrameData[30]
rlabel metal2 272 11004 272 11004 0 FrameData[31]
rlabel metal2 6224 1596 6224 1596 0 FrameData[3]
rlabel metal3 13344 2268 13344 2268 0 FrameData[4]
rlabel metal2 1808 2268 1808 2268 0 FrameData[5]
rlabel metal2 3632 2604 3632 2604 0 FrameData[6]
rlabel metal3 18528 3192 18528 3192 0 FrameData[7]
rlabel metal2 20352 3402 20352 3402 0 FrameData[8]
rlabel metal3 14352 3192 14352 3192 0 FrameData[9]
rlabel metal3 37536 1134 37536 1134 0 FrameData_O[0]
rlabel metal2 38943 3948 38943 3948 0 FrameData_O[10]
rlabel metal2 38631 4284 38631 4284 0 FrameData_O[11]
rlabel metal2 38847 4620 38847 4620 0 FrameData_O[12]
rlabel metal2 38631 4956 38631 4956 0 FrameData_O[13]
rlabel metal2 38847 5292 38847 5292 0 FrameData_O[14]
rlabel metal2 38631 5628 38631 5628 0 FrameData_O[15]
rlabel metal2 38847 5964 38847 5964 0 FrameData_O[16]
rlabel metal2 38631 6300 38631 6300 0 FrameData_O[17]
rlabel via2 39183 6636 39183 6636 0 FrameData_O[18]
rlabel metal2 38631 6972 38631 6972 0 FrameData_O[19]
rlabel metal3 37824 1344 37824 1344 0 FrameData_O[1]
rlabel metal2 38943 7308 38943 7308 0 FrameData_O[20]
rlabel metal2 38439 7644 38439 7644 0 FrameData_O[21]
rlabel metal2 38943 7980 38943 7980 0 FrameData_O[22]
rlabel metal2 38439 8316 38439 8316 0 FrameData_O[23]
rlabel metal2 38943 8652 38943 8652 0 FrameData_O[24]
rlabel via2 39183 8988 39183 8988 0 FrameData_O[25]
rlabel metal2 38247 9324 38247 9324 0 FrameData_O[26]
rlabel metal2 38055 9660 38055 9660 0 FrameData_O[27]
rlabel metal2 37320 8904 37320 8904 0 FrameData_O[28]
rlabel metal2 36552 9660 36552 9660 0 FrameData_O[29]
rlabel metal2 38319 1260 38319 1260 0 FrameData_O[2]
rlabel metal2 36168 9660 36168 9660 0 FrameData_O[30]
rlabel metal2 36984 8904 36984 8904 0 FrameData_O[31]
rlabel metal2 38559 1596 38559 1596 0 FrameData_O[3]
rlabel metal2 37920 2184 37920 2184 0 FrameData_O[4]
rlabel metal2 38376 2100 38376 2100 0 FrameData_O[5]
rlabel metal2 38943 2604 38943 2604 0 FrameData_O[6]
rlabel metal2 38232 2856 38232 2856 0 FrameData_O[7]
rlabel metal2 38439 3276 38439 3276 0 FrameData_O[8]
rlabel metal2 38631 3612 38631 3612 0 FrameData_O[9]
rlabel metal3 3936 114 3936 114 0 FrameStrobe[0]
rlabel metal3 27072 2100 27072 2100 0 FrameStrobe[10]
rlabel metal2 24672 3864 24672 3864 0 FrameStrobe[11]
rlabel metal3 24672 2088 24672 2088 0 FrameStrobe[12]
rlabel metal3 26400 2508 26400 2508 0 FrameStrobe[13]
rlabel metal3 28128 2844 28128 2844 0 FrameStrobe[14]
rlabel metal3 29856 3264 29856 3264 0 FrameStrobe[15]
rlabel metal3 31584 3222 31584 3222 0 FrameStrobe[16]
rlabel metal3 33312 3474 33312 3474 0 FrameStrobe[17]
rlabel metal3 35040 1458 35040 1458 0 FrameStrobe[18]
rlabel metal3 36768 3516 36768 3516 0 FrameStrobe[19]
rlabel metal2 5520 3444 5520 3444 0 FrameStrobe[1]
rlabel metal3 7392 1290 7392 1290 0 FrameStrobe[2]
rlabel metal3 9120 1374 9120 1374 0 FrameStrobe[3]
rlabel metal3 10848 912 10848 912 0 FrameStrobe[4]
rlabel metal3 12576 1080 12576 1080 0 FrameStrobe[5]
rlabel metal3 29568 2310 29568 2310 0 FrameStrobe[6]
rlabel metal3 27840 2226 27840 2226 0 FrameStrobe[7]
rlabel metal3 25632 2268 25632 2268 0 FrameStrobe[8]
rlabel metal2 25248 2730 25248 2730 0 FrameStrobe[9]
rlabel metal2 27864 9576 27864 9576 0 FrameStrobe_O[0]
rlabel metal2 29688 8904 29688 8904 0 FrameStrobe_O[10]
rlabel metal2 30408 9660 30408 9660 0 FrameStrobe_O[11]
rlabel metal2 30072 8904 30072 8904 0 FrameStrobe_O[12]
rlabel metal2 30936 9660 30936 9660 0 FrameStrobe_O[13]
rlabel metal2 30456 8904 30456 8904 0 FrameStrobe_O[14]
rlabel metal2 31032 9324 31032 9324 0 FrameStrobe_O[15]
rlabel metal2 30840 8904 30840 8904 0 FrameStrobe_O[16]
rlabel metal2 31608 9576 31608 9576 0 FrameStrobe_O[17]
rlabel metal2 31224 8904 31224 8904 0 FrameStrobe_O[18]
rlabel metal2 31800 9660 31800 9660 0 FrameStrobe_O[19]
rlabel metal2 28152 9660 28152 9660 0 FrameStrobe_O[1]
rlabel metal2 28440 9576 28440 9576 0 FrameStrobe_O[2]
rlabel metal2 28920 9660 28920 9660 0 FrameStrobe_O[3]
rlabel metal2 28536 8904 28536 8904 0 FrameStrobe_O[4]
rlabel metal2 29112 9324 29112 9324 0 FrameStrobe_O[5]
rlabel metal2 28920 8904 28920 8904 0 FrameStrobe_O[6]
rlabel metal2 29496 9576 29496 9576 0 FrameStrobe_O[7]
rlabel metal2 29304 8904 29304 8904 0 FrameStrobe_O[8]
rlabel metal2 29880 9240 29880 9240 0 FrameStrobe_O[9]
rlabel metal2 7464 9660 7464 9660 0 N1BEG[0]
rlabel metal2 7800 8904 7800 8904 0 N1BEG[1]
rlabel metal2 7848 9660 7848 9660 0 N1BEG[2]
rlabel metal2 8184 8904 8184 8904 0 N1BEG[3]
rlabel metal2 8232 9660 8232 9660 0 N2BEG[0]
rlabel metal2 8568 8904 8568 8904 0 N2BEG[1]
rlabel metal2 8616 9660 8616 9660 0 N2BEG[2]
rlabel metal2 8952 8904 8952 8904 0 N2BEG[3]
rlabel metal2 9000 9660 9000 9660 0 N2BEG[4]
rlabel metal2 9336 8904 9336 8904 0 N2BEG[5]
rlabel metal2 9384 9660 9384 9660 0 N2BEG[6]
rlabel metal2 9720 8904 9720 8904 0 N2BEG[7]
rlabel metal2 9768 9660 9768 9660 0 N2BEGb[0]
rlabel metal2 10104 8904 10104 8904 0 N2BEGb[1]
rlabel metal2 10152 9660 10152 9660 0 N2BEGb[2]
rlabel metal2 10488 8904 10488 8904 0 N2BEGb[3]
rlabel metal2 10536 9660 10536 9660 0 N2BEGb[4]
rlabel metal2 10872 8904 10872 8904 0 N2BEGb[5]
rlabel metal2 10920 9660 10920 9660 0 N2BEGb[6]
rlabel metal2 11256 8904 11256 8904 0 N2BEGb[7]
rlabel metal2 11304 9660 11304 9660 0 N4BEG[0]
rlabel metal2 13224 9660 13224 9660 0 N4BEG[10]
rlabel metal2 13560 8904 13560 8904 0 N4BEG[11]
rlabel metal2 13608 9660 13608 9660 0 N4BEG[12]
rlabel metal2 13944 8904 13944 8904 0 N4BEG[13]
rlabel metal2 13992 9660 13992 9660 0 N4BEG[14]
rlabel metal2 14328 8904 14328 8904 0 N4BEG[15]
rlabel metal2 11640 8904 11640 8904 0 N4BEG[1]
rlabel metal2 11688 9660 11688 9660 0 N4BEG[2]
rlabel metal2 12024 8904 12024 8904 0 N4BEG[3]
rlabel metal2 12072 9660 12072 9660 0 N4BEG[4]
rlabel metal2 12408 8904 12408 8904 0 N4BEG[5]
rlabel metal2 12456 9660 12456 9660 0 N4BEG[6]
rlabel metal2 12792 8904 12792 8904 0 N4BEG[7]
rlabel metal3 13056 10584 13056 10584 0 N4BEG[8]
rlabel metal2 13176 8904 13176 8904 0 N4BEG[9]
rlabel metal2 14376 9660 14376 9660 0 NN4BEG[0]
rlabel metal2 16200 9492 16200 9492 0 NN4BEG[10]
rlabel metal2 16584 9660 16584 9660 0 NN4BEG[11]
rlabel metal2 16728 9576 16728 9576 0 NN4BEG[12]
rlabel metal2 17016 9660 17016 9660 0 NN4BEG[13]
rlabel metal2 17496 9576 17496 9576 0 NN4BEG[14]
rlabel metal2 17400 9660 17400 9660 0 NN4BEG[15]
rlabel metal2 14712 8904 14712 8904 0 NN4BEG[1]
rlabel metal2 14760 9660 14760 9660 0 NN4BEG[2]
rlabel metal2 15096 8904 15096 8904 0 NN4BEG[3]
rlabel metal2 15144 9660 15144 9660 0 NN4BEG[4]
rlabel metal2 15480 8904 15480 8904 0 NN4BEG[5]
rlabel metal2 15528 9660 15528 9660 0 NN4BEG[6]
rlabel metal2 15864 8904 15864 8904 0 NN4BEG[7]
rlabel metal2 15912 9660 15912 9660 0 NN4BEG[8]
rlabel metal2 16248 8904 16248 8904 0 NN4BEG[9]
rlabel metal3 17568 8160 17568 8160 0 S1END[0]
rlabel metal3 17760 11730 17760 11730 0 S1END[1]
rlabel metal3 17952 11688 17952 11688 0 S1END[2]
rlabel metal3 18144 11226 18144 11226 0 S1END[3]
rlabel metal3 19872 9966 19872 9966 0 S2END[0]
rlabel metal3 20064 10680 20064 10680 0 S2END[1]
rlabel metal3 20256 10512 20256 10512 0 S2END[2]
rlabel metal3 20448 10680 20448 10680 0 S2END[3]
rlabel metal3 20640 8202 20640 8202 0 S2END[4]
rlabel metal3 20832 7824 20832 7824 0 S2END[5]
rlabel metal3 21024 7908 21024 7908 0 S2END[6]
rlabel metal3 21216 11310 21216 11310 0 S2END[7]
rlabel metal3 18336 9714 18336 9714 0 S2MID[0]
rlabel metal3 18528 8202 18528 8202 0 S2MID[1]
rlabel metal3 18720 11184 18720 11184 0 S2MID[2]
rlabel metal3 18912 10890 18912 10890 0 S2MID[3]
rlabel metal3 19104 10890 19104 10890 0 S2MID[4]
rlabel metal3 19296 10974 19296 10974 0 S2MID[5]
rlabel metal3 19488 10974 19488 10974 0 S2MID[6]
rlabel metal3 19680 10722 19680 10722 0 S2MID[7]
rlabel metal3 21408 9210 21408 9210 0 S4END[0]
rlabel metal3 23328 8328 23328 8328 0 S4END[10]
rlabel metal3 23520 8118 23520 8118 0 S4END[11]
rlabel metal3 23712 8874 23712 8874 0 S4END[12]
rlabel metal3 23904 10890 23904 10890 0 S4END[13]
rlabel metal3 24096 8034 24096 8034 0 S4END[14]
rlabel via2 24288 11772 24288 11772 0 S4END[15]
rlabel metal3 21600 8412 21600 8412 0 S4END[1]
rlabel metal3 21792 8496 21792 8496 0 S4END[2]
rlabel metal3 21984 8706 21984 8706 0 S4END[3]
rlabel metal3 22176 8664 22176 8664 0 S4END[4]
rlabel metal3 22368 8748 22368 8748 0 S4END[5]
rlabel metal3 22560 8580 22560 8580 0 S4END[6]
rlabel metal3 22752 8454 22752 8454 0 S4END[7]
rlabel metal3 22944 10470 22944 10470 0 S4END[8]
rlabel metal3 23136 10176 23136 10176 0 S4END[9]
rlabel metal3 24576 7128 24576 7128 0 SS4END[0]
rlabel metal3 26400 10848 26400 10848 0 SS4END[10]
rlabel metal3 26592 9546 26592 9546 0 SS4END[11]
rlabel metal3 26784 10050 26784 10050 0 SS4END[12]
rlabel metal3 26976 10176 26976 10176 0 SS4END[13]
rlabel metal3 27168 9882 27168 9882 0 SS4END[14]
rlabel metal3 27360 11604 27360 11604 0 SS4END[15]
rlabel metal3 24672 9336 24672 9336 0 SS4END[1]
rlabel metal3 24864 9126 24864 9126 0 SS4END[2]
rlabel metal3 25056 9588 25056 9588 0 SS4END[3]
rlabel metal3 25248 9630 25248 9630 0 SS4END[4]
rlabel metal3 25440 9168 25440 9168 0 SS4END[5]
rlabel metal3 25632 10638 25632 10638 0 SS4END[6]
rlabel metal3 25728 7002 25728 7002 0 SS4END[7]
rlabel metal2 25872 6888 25872 6888 0 SS4END[8]
rlabel metal2 25824 7056 25824 7056 0 SS4END[9]
rlabel metal3 2208 2046 2208 2046 0 UserCLK
rlabel metal2 27576 9660 27576 9660 0 UserCLKo
rlabel metal2 27360 1722 27360 1722 0 net1
rlabel metal3 27072 3486 27072 3486 0 net10
rlabel metal2 21048 7812 21048 7812 0 net100
rlabel metal2 21144 6972 21144 6972 0 net101
rlabel metal2 20280 6972 20280 6972 0 net102
rlabel metal2 19032 6972 19032 6972 0 net103
rlabel metal2 17736 7056 17736 7056 0 net104
rlabel metal2 24576 3990 24576 3990 0 net105
rlabel metal2 26664 3528 26664 3528 0 net11
rlabel metal3 36672 2226 36672 2226 0 net12
rlabel metal2 37728 7980 37728 7980 0 net13
rlabel metal3 35904 4914 35904 4914 0 net14
rlabel metal3 37824 7644 37824 7644 0 net15
rlabel metal2 26616 6972 26616 6972 0 net16
rlabel metal2 37824 9534 37824 9534 0 net17
rlabel metal2 31608 7728 31608 7728 0 net18
rlabel metal2 32760 8148 32760 8148 0 net19
rlabel metal2 37344 4116 37344 4116 0 net2
rlabel metal2 30600 7728 30600 7728 0 net20
rlabel metal2 31176 8148 31176 8148 0 net21
rlabel metal2 26904 7812 26904 7812 0 net22
rlabel metal2 36288 2058 36288 2058 0 net23
rlabel metal2 30072 8148 30072 8148 0 net24
rlabel metal2 34728 8652 34728 8652 0 net25
rlabel metal3 25824 2100 25824 2100 0 net26
rlabel metal2 37056 2478 37056 2478 0 net27
rlabel metal3 37632 2436 37632 2436 0 net28
rlabel metal3 24480 4032 24480 4032 0 net29
rlabel metal2 27072 3486 27072 3486 0 net3
rlabel metal3 37824 2898 37824 2898 0 net30
rlabel metal2 36240 3444 36240 3444 0 net31
rlabel metal2 37824 3402 37824 3402 0 net32
rlabel metal2 3528 4284 3528 4284 0 net33
rlabel metal2 28104 2856 28104 2856 0 net34
rlabel metal2 28920 3612 28920 3612 0 net35
rlabel metal2 29448 4284 29448 4284 0 net36
rlabel metal2 29016 5124 29016 5124 0 net37
rlabel metal2 29304 5628 29304 5628 0 net38
rlabel metal2 30072 6636 30072 6636 0 net39
rlabel metal2 36144 4956 36144 4956 0 net4
rlabel metal2 29736 6636 29736 6636 0 net40
rlabel metal2 29928 7056 29928 7056 0 net41
rlabel metal2 30552 7392 30552 7392 0 net42
rlabel metal2 31368 7140 31368 7140 0 net43
rlabel metal3 28608 9450 28608 9450 0 net44
rlabel metal2 8520 2856 8520 2856 0 net45
rlabel metal2 8232 2856 8232 2856 0 net46
rlabel metal2 28176 8652 28176 8652 0 net47
rlabel metal2 30168 2856 30168 2856 0 net48
rlabel metal2 29256 2856 29256 2856 0 net49
rlabel metal3 37536 4284 37536 4284 0 net5
rlabel metal2 28584 2772 28584 2772 0 net50
rlabel metal2 26664 2772 26664 2772 0 net51
rlabel metal2 25728 2730 25728 2730 0 net52
rlabel metal2 5736 5544 5736 5544 0 net53
rlabel metal2 6504 5544 6504 5544 0 net54
rlabel metal2 7368 5628 7368 5628 0 net55
rlabel metal2 6888 5880 6888 5880 0 net56
rlabel metal2 6120 5124 6120 5124 0 net57
rlabel metal2 7464 5460 7464 5460 0 net58
rlabel metal2 7176 5124 7176 5124 0 net59
rlabel metal2 15720 2856 15720 2856 0 net6
rlabel metal2 8232 5040 8232 5040 0 net60
rlabel metal2 8472 5124 8472 5124 0 net61
rlabel metal2 9528 5124 9528 5124 0 net62
rlabel metal2 9048 5124 9048 5124 0 net63
rlabel metal2 9240 5040 9240 5040 0 net64
rlabel metal2 7560 5124 7560 5124 0 net65
rlabel metal2 9672 4284 9672 4284 0 net66
rlabel metal2 10488 4116 10488 4116 0 net67
rlabel metal2 11256 5124 11256 5124 0 net68
rlabel metal2 12120 4956 12120 4956 0 net69
rlabel metal2 37824 5586 37824 5586 0 net7
rlabel metal2 12024 4788 12024 4788 0 net70
rlabel metal2 13656 5040 13656 5040 0 net71
rlabel metal2 12264 5124 12264 5124 0 net72
rlabel metal2 8424 4284 8424 4284 0 net73
rlabel metal2 17400 5544 17400 5544 0 net74
rlabel metal2 15528 5796 15528 5796 0 net75
rlabel metal2 17736 5628 17736 5628 0 net76
rlabel metal2 15672 5460 15672 5460 0 net77
rlabel metal2 15240 4788 15240 4788 0 net78
rlabel metal2 15672 6636 15672 6636 0 net79
rlabel metal2 37440 6510 37440 6510 0 net8
rlabel metal2 10392 3948 10392 3948 0 net80
rlabel metal2 11496 4284 11496 4284 0 net81
rlabel metal3 12432 4704 12432 4704 0 net82
rlabel metal2 14136 5124 14136 5124 0 net83
rlabel metal2 13728 5754 13728 5754 0 net84
rlabel metal2 14304 5628 14304 5628 0 net85
rlabel metal2 15768 5040 15768 5040 0 net86
rlabel metal2 14400 5502 14400 5502 0 net87
rlabel metal2 16440 5460 16440 5460 0 net88
rlabel metal3 27264 8484 27264 8484 0 net89
rlabel metal2 37824 6426 37824 6426 0 net9
rlabel metal2 17256 6972 17256 6972 0 net90
rlabel metal2 19992 7812 19992 7812 0 net91
rlabel metal2 19608 7980 19608 7980 0 net92
rlabel metal2 18552 6636 18552 6636 0 net93
rlabel metal2 19224 7392 19224 7392 0 net94
rlabel metal2 20088 7140 20088 7140 0 net95
rlabel metal2 25992 7728 25992 7728 0 net96
rlabel metal2 24792 7728 24792 7728 0 net97
rlabel metal2 23928 7980 23928 7980 0 net98
rlabel metal2 21288 7728 21288 7728 0 net99
<< properties >>
string FIXED_BBOX 0 0 39264 11844
<< end >>
