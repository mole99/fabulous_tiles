* NGSPICE file created from DSP.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlhq_1 abstract view
.subckt sg13g2_dlhq_1 D GATE Q VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd1_1 abstract view
.subckt sg13g2_dlygate4sd1_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_dfrbp_1 abstract view
.subckt sg13g2_dfrbp_1 CLK RESET_B D Q_N Q VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_16 abstract view
.subckt sg13g2_buf_16 X A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VSS VDD B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_mux2_2 abstract view
.subckt sg13g2_mux2_2 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_inv_16 abstract view
.subckt sg13g2_inv_16 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

.subckt DSP Tile_X0Y0_E1BEG[0] Tile_X0Y0_E1BEG[1] Tile_X0Y0_E1BEG[2] Tile_X0Y0_E1BEG[3]
+ Tile_X0Y0_E1END[0] Tile_X0Y0_E1END[1] Tile_X0Y0_E1END[2] Tile_X0Y0_E1END[3] Tile_X0Y0_E2BEG[0]
+ Tile_X0Y0_E2BEG[1] Tile_X0Y0_E2BEG[2] Tile_X0Y0_E2BEG[3] Tile_X0Y0_E2BEG[4] Tile_X0Y0_E2BEG[5]
+ Tile_X0Y0_E2BEG[6] Tile_X0Y0_E2BEG[7] Tile_X0Y0_E2BEGb[0] Tile_X0Y0_E2BEGb[1] Tile_X0Y0_E2BEGb[2]
+ Tile_X0Y0_E2BEGb[3] Tile_X0Y0_E2BEGb[4] Tile_X0Y0_E2BEGb[5] Tile_X0Y0_E2BEGb[6]
+ Tile_X0Y0_E2BEGb[7] Tile_X0Y0_E2END[0] Tile_X0Y0_E2END[1] Tile_X0Y0_E2END[2] Tile_X0Y0_E2END[3]
+ Tile_X0Y0_E2END[4] Tile_X0Y0_E2END[5] Tile_X0Y0_E2END[6] Tile_X0Y0_E2END[7] Tile_X0Y0_E2MID[0]
+ Tile_X0Y0_E2MID[1] Tile_X0Y0_E2MID[2] Tile_X0Y0_E2MID[3] Tile_X0Y0_E2MID[4] Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_E2MID[6] Tile_X0Y0_E2MID[7] Tile_X0Y0_E6BEG[0] Tile_X0Y0_E6BEG[10] Tile_X0Y0_E6BEG[11]
+ Tile_X0Y0_E6BEG[1] Tile_X0Y0_E6BEG[2] Tile_X0Y0_E6BEG[3] Tile_X0Y0_E6BEG[4] Tile_X0Y0_E6BEG[5]
+ Tile_X0Y0_E6BEG[6] Tile_X0Y0_E6BEG[7] Tile_X0Y0_E6BEG[8] Tile_X0Y0_E6BEG[9] Tile_X0Y0_E6END[0]
+ Tile_X0Y0_E6END[10] Tile_X0Y0_E6END[11] Tile_X0Y0_E6END[1] Tile_X0Y0_E6END[2] Tile_X0Y0_E6END[3]
+ Tile_X0Y0_E6END[4] Tile_X0Y0_E6END[5] Tile_X0Y0_E6END[6] Tile_X0Y0_E6END[7] Tile_X0Y0_E6END[8]
+ Tile_X0Y0_E6END[9] Tile_X0Y0_EE4BEG[0] Tile_X0Y0_EE4BEG[10] Tile_X0Y0_EE4BEG[11]
+ Tile_X0Y0_EE4BEG[12] Tile_X0Y0_EE4BEG[13] Tile_X0Y0_EE4BEG[14] Tile_X0Y0_EE4BEG[15]
+ Tile_X0Y0_EE4BEG[1] Tile_X0Y0_EE4BEG[2] Tile_X0Y0_EE4BEG[3] Tile_X0Y0_EE4BEG[4]
+ Tile_X0Y0_EE4BEG[5] Tile_X0Y0_EE4BEG[6] Tile_X0Y0_EE4BEG[7] Tile_X0Y0_EE4BEG[8]
+ Tile_X0Y0_EE4BEG[9] Tile_X0Y0_EE4END[0] Tile_X0Y0_EE4END[10] Tile_X0Y0_EE4END[11]
+ Tile_X0Y0_EE4END[12] Tile_X0Y0_EE4END[13] Tile_X0Y0_EE4END[14] Tile_X0Y0_EE4END[15]
+ Tile_X0Y0_EE4END[1] Tile_X0Y0_EE4END[2] Tile_X0Y0_EE4END[3] Tile_X0Y0_EE4END[4]
+ Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[6] Tile_X0Y0_EE4END[7] Tile_X0Y0_EE4END[8]
+ Tile_X0Y0_EE4END[9] Tile_X0Y0_FrameData[0] Tile_X0Y0_FrameData[10] Tile_X0Y0_FrameData[11]
+ Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData[13] Tile_X0Y0_FrameData[14] Tile_X0Y0_FrameData[15]
+ Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData[17] Tile_X0Y0_FrameData[18] Tile_X0Y0_FrameData[19]
+ Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData[20] Tile_X0Y0_FrameData[21] Tile_X0Y0_FrameData[22]
+ Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData[24] Tile_X0Y0_FrameData[25] Tile_X0Y0_FrameData[26]
+ Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData[28] Tile_X0Y0_FrameData[29] Tile_X0Y0_FrameData[2]
+ Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData[31] Tile_X0Y0_FrameData[3] Tile_X0Y0_FrameData[4]
+ Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData[6] Tile_X0Y0_FrameData[7] Tile_X0Y0_FrameData[8]
+ Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[0] Tile_X0Y0_FrameData_O[10] Tile_X0Y0_FrameData_O[11]
+ Tile_X0Y0_FrameData_O[12] Tile_X0Y0_FrameData_O[13] Tile_X0Y0_FrameData_O[14] Tile_X0Y0_FrameData_O[15]
+ Tile_X0Y0_FrameData_O[16] Tile_X0Y0_FrameData_O[17] Tile_X0Y0_FrameData_O[18] Tile_X0Y0_FrameData_O[19]
+ Tile_X0Y0_FrameData_O[1] Tile_X0Y0_FrameData_O[20] Tile_X0Y0_FrameData_O[21] Tile_X0Y0_FrameData_O[22]
+ Tile_X0Y0_FrameData_O[23] Tile_X0Y0_FrameData_O[24] Tile_X0Y0_FrameData_O[25] Tile_X0Y0_FrameData_O[26]
+ Tile_X0Y0_FrameData_O[27] Tile_X0Y0_FrameData_O[28] Tile_X0Y0_FrameData_O[29] Tile_X0Y0_FrameData_O[2]
+ Tile_X0Y0_FrameData_O[30] Tile_X0Y0_FrameData_O[31] Tile_X0Y0_FrameData_O[3] Tile_X0Y0_FrameData_O[4]
+ Tile_X0Y0_FrameData_O[5] Tile_X0Y0_FrameData_O[6] Tile_X0Y0_FrameData_O[7] Tile_X0Y0_FrameData_O[8]
+ Tile_X0Y0_FrameData_O[9] Tile_X0Y0_FrameStrobe_O[0] Tile_X0Y0_FrameStrobe_O[10]
+ Tile_X0Y0_FrameStrobe_O[11] Tile_X0Y0_FrameStrobe_O[12] Tile_X0Y0_FrameStrobe_O[13]
+ Tile_X0Y0_FrameStrobe_O[14] Tile_X0Y0_FrameStrobe_O[15] Tile_X0Y0_FrameStrobe_O[16]
+ Tile_X0Y0_FrameStrobe_O[17] Tile_X0Y0_FrameStrobe_O[18] Tile_X0Y0_FrameStrobe_O[19]
+ Tile_X0Y0_FrameStrobe_O[1] Tile_X0Y0_FrameStrobe_O[2] Tile_X0Y0_FrameStrobe_O[3]
+ Tile_X0Y0_FrameStrobe_O[4] Tile_X0Y0_FrameStrobe_O[5] Tile_X0Y0_FrameStrobe_O[6]
+ Tile_X0Y0_FrameStrobe_O[7] Tile_X0Y0_FrameStrobe_O[8] Tile_X0Y0_FrameStrobe_O[9]
+ Tile_X0Y0_N1BEG[0] Tile_X0Y0_N1BEG[1] Tile_X0Y0_N1BEG[2] Tile_X0Y0_N1BEG[3] Tile_X0Y0_N2BEG[0]
+ Tile_X0Y0_N2BEG[1] Tile_X0Y0_N2BEG[2] Tile_X0Y0_N2BEG[3] Tile_X0Y0_N2BEG[4] Tile_X0Y0_N2BEG[5]
+ Tile_X0Y0_N2BEG[6] Tile_X0Y0_N2BEG[7] Tile_X0Y0_N2BEGb[0] Tile_X0Y0_N2BEGb[1] Tile_X0Y0_N2BEGb[2]
+ Tile_X0Y0_N2BEGb[3] Tile_X0Y0_N2BEGb[4] Tile_X0Y0_N2BEGb[5] Tile_X0Y0_N2BEGb[6]
+ Tile_X0Y0_N2BEGb[7] Tile_X0Y0_N4BEG[0] Tile_X0Y0_N4BEG[10] Tile_X0Y0_N4BEG[11] Tile_X0Y0_N4BEG[12]
+ Tile_X0Y0_N4BEG[13] Tile_X0Y0_N4BEG[14] Tile_X0Y0_N4BEG[15] Tile_X0Y0_N4BEG[1] Tile_X0Y0_N4BEG[2]
+ Tile_X0Y0_N4BEG[3] Tile_X0Y0_N4BEG[4] Tile_X0Y0_N4BEG[5] Tile_X0Y0_N4BEG[6] Tile_X0Y0_N4BEG[7]
+ Tile_X0Y0_N4BEG[8] Tile_X0Y0_N4BEG[9] Tile_X0Y0_NN4BEG[0] Tile_X0Y0_NN4BEG[10] Tile_X0Y0_NN4BEG[11]
+ Tile_X0Y0_NN4BEG[12] Tile_X0Y0_NN4BEG[13] Tile_X0Y0_NN4BEG[14] Tile_X0Y0_NN4BEG[15]
+ Tile_X0Y0_NN4BEG[1] Tile_X0Y0_NN4BEG[2] Tile_X0Y0_NN4BEG[3] Tile_X0Y0_NN4BEG[4]
+ Tile_X0Y0_NN4BEG[5] Tile_X0Y0_NN4BEG[6] Tile_X0Y0_NN4BEG[7] Tile_X0Y0_NN4BEG[8]
+ Tile_X0Y0_NN4BEG[9] Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[1] Tile_X0Y0_S1END[2] Tile_X0Y0_S1END[3]
+ Tile_X0Y0_S2END[0] Tile_X0Y0_S2END[1] Tile_X0Y0_S2END[2] Tile_X0Y0_S2END[3] Tile_X0Y0_S2END[4]
+ Tile_X0Y0_S2END[5] Tile_X0Y0_S2END[6] Tile_X0Y0_S2END[7] Tile_X0Y0_S2MID[0] Tile_X0Y0_S2MID[1]
+ Tile_X0Y0_S2MID[2] Tile_X0Y0_S2MID[3] Tile_X0Y0_S2MID[4] Tile_X0Y0_S2MID[5] Tile_X0Y0_S2MID[6]
+ Tile_X0Y0_S2MID[7] Tile_X0Y0_S4END[0] Tile_X0Y0_S4END[10] Tile_X0Y0_S4END[11] Tile_X0Y0_S4END[12]
+ Tile_X0Y0_S4END[13] Tile_X0Y0_S4END[14] Tile_X0Y0_S4END[15] Tile_X0Y0_S4END[1] Tile_X0Y0_S4END[2]
+ Tile_X0Y0_S4END[3] Tile_X0Y0_S4END[4] Tile_X0Y0_S4END[5] Tile_X0Y0_S4END[6] Tile_X0Y0_S4END[7]
+ Tile_X0Y0_S4END[8] Tile_X0Y0_S4END[9] Tile_X0Y0_SS4END[0] Tile_X0Y0_SS4END[10] Tile_X0Y0_SS4END[11]
+ Tile_X0Y0_SS4END[12] Tile_X0Y0_SS4END[13] Tile_X0Y0_SS4END[14] Tile_X0Y0_SS4END[15]
+ Tile_X0Y0_SS4END[1] Tile_X0Y0_SS4END[2] Tile_X0Y0_SS4END[3] Tile_X0Y0_SS4END[4]
+ Tile_X0Y0_SS4END[5] Tile_X0Y0_SS4END[6] Tile_X0Y0_SS4END[7] Tile_X0Y0_SS4END[8]
+ Tile_X0Y0_SS4END[9] Tile_X0Y0_UserCLKo Tile_X0Y0_W1BEG[0] Tile_X0Y0_W1BEG[1] Tile_X0Y0_W1BEG[2]
+ Tile_X0Y0_W1BEG[3] Tile_X0Y0_W1END[0] Tile_X0Y0_W1END[1] Tile_X0Y0_W1END[2] Tile_X0Y0_W1END[3]
+ Tile_X0Y0_W2BEG[0] Tile_X0Y0_W2BEG[1] Tile_X0Y0_W2BEG[2] Tile_X0Y0_W2BEG[3] Tile_X0Y0_W2BEG[4]
+ Tile_X0Y0_W2BEG[5] Tile_X0Y0_W2BEG[6] Tile_X0Y0_W2BEG[7] Tile_X0Y0_W2BEGb[0] Tile_X0Y0_W2BEGb[1]
+ Tile_X0Y0_W2BEGb[2] Tile_X0Y0_W2BEGb[3] Tile_X0Y0_W2BEGb[4] Tile_X0Y0_W2BEGb[5]
+ Tile_X0Y0_W2BEGb[6] Tile_X0Y0_W2BEGb[7] Tile_X0Y0_W2END[0] Tile_X0Y0_W2END[1] Tile_X0Y0_W2END[2]
+ Tile_X0Y0_W2END[3] Tile_X0Y0_W2END[4] Tile_X0Y0_W2END[5] Tile_X0Y0_W2END[6] Tile_X0Y0_W2END[7]
+ Tile_X0Y0_W2MID[0] Tile_X0Y0_W2MID[1] Tile_X0Y0_W2MID[2] Tile_X0Y0_W2MID[3] Tile_X0Y0_W2MID[4]
+ Tile_X0Y0_W2MID[5] Tile_X0Y0_W2MID[6] Tile_X0Y0_W2MID[7] Tile_X0Y0_W6BEG[0] Tile_X0Y0_W6BEG[10]
+ Tile_X0Y0_W6BEG[11] Tile_X0Y0_W6BEG[1] Tile_X0Y0_W6BEG[2] Tile_X0Y0_W6BEG[3] Tile_X0Y0_W6BEG[4]
+ Tile_X0Y0_W6BEG[5] Tile_X0Y0_W6BEG[6] Tile_X0Y0_W6BEG[7] Tile_X0Y0_W6BEG[8] Tile_X0Y0_W6BEG[9]
+ Tile_X0Y0_W6END[0] Tile_X0Y0_W6END[10] Tile_X0Y0_W6END[11] Tile_X0Y0_W6END[1] Tile_X0Y0_W6END[2]
+ Tile_X0Y0_W6END[3] Tile_X0Y0_W6END[4] Tile_X0Y0_W6END[5] Tile_X0Y0_W6END[6] Tile_X0Y0_W6END[7]
+ Tile_X0Y0_W6END[8] Tile_X0Y0_W6END[9] Tile_X0Y0_WW4BEG[0] Tile_X0Y0_WW4BEG[10] Tile_X0Y0_WW4BEG[11]
+ Tile_X0Y0_WW4BEG[12] Tile_X0Y0_WW4BEG[13] Tile_X0Y0_WW4BEG[14] Tile_X0Y0_WW4BEG[15]
+ Tile_X0Y0_WW4BEG[1] Tile_X0Y0_WW4BEG[2] Tile_X0Y0_WW4BEG[3] Tile_X0Y0_WW4BEG[4]
+ Tile_X0Y0_WW4BEG[5] Tile_X0Y0_WW4BEG[6] Tile_X0Y0_WW4BEG[7] Tile_X0Y0_WW4BEG[8]
+ Tile_X0Y0_WW4BEG[9] Tile_X0Y0_WW4END[0] Tile_X0Y0_WW4END[10] Tile_X0Y0_WW4END[11]
+ Tile_X0Y0_WW4END[12] Tile_X0Y0_WW4END[13] Tile_X0Y0_WW4END[14] Tile_X0Y0_WW4END[15]
+ Tile_X0Y0_WW4END[1] Tile_X0Y0_WW4END[2] Tile_X0Y0_WW4END[3] Tile_X0Y0_WW4END[4]
+ Tile_X0Y0_WW4END[5] Tile_X0Y0_WW4END[6] Tile_X0Y0_WW4END[7] Tile_X0Y0_WW4END[8]
+ Tile_X0Y0_WW4END[9] Tile_X0Y1_E1BEG[0] Tile_X0Y1_E1BEG[1] Tile_X0Y1_E1BEG[2] Tile_X0Y1_E1BEG[3]
+ Tile_X0Y1_E1END[0] Tile_X0Y1_E1END[1] Tile_X0Y1_E1END[2] Tile_X0Y1_E1END[3] Tile_X0Y1_E2BEG[0]
+ Tile_X0Y1_E2BEG[1] Tile_X0Y1_E2BEG[2] Tile_X0Y1_E2BEG[3] Tile_X0Y1_E2BEG[4] Tile_X0Y1_E2BEG[5]
+ Tile_X0Y1_E2BEG[6] Tile_X0Y1_E2BEG[7] Tile_X0Y1_E2BEGb[0] Tile_X0Y1_E2BEGb[1] Tile_X0Y1_E2BEGb[2]
+ Tile_X0Y1_E2BEGb[3] Tile_X0Y1_E2BEGb[4] Tile_X0Y1_E2BEGb[5] Tile_X0Y1_E2BEGb[6]
+ Tile_X0Y1_E2BEGb[7] Tile_X0Y1_E2END[0] Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2] Tile_X0Y1_E2END[3]
+ Tile_X0Y1_E2END[4] Tile_X0Y1_E2END[5] Tile_X0Y1_E2END[6] Tile_X0Y1_E2END[7] Tile_X0Y1_E2MID[0]
+ Tile_X0Y1_E2MID[1] Tile_X0Y1_E2MID[2] Tile_X0Y1_E2MID[3] Tile_X0Y1_E2MID[4] Tile_X0Y1_E2MID[5]
+ Tile_X0Y1_E2MID[6] Tile_X0Y1_E2MID[7] Tile_X0Y1_E6BEG[0] Tile_X0Y1_E6BEG[10] Tile_X0Y1_E6BEG[11]
+ Tile_X0Y1_E6BEG[1] Tile_X0Y1_E6BEG[2] Tile_X0Y1_E6BEG[3] Tile_X0Y1_E6BEG[4] Tile_X0Y1_E6BEG[5]
+ Tile_X0Y1_E6BEG[6] Tile_X0Y1_E6BEG[7] Tile_X0Y1_E6BEG[8] Tile_X0Y1_E6BEG[9] Tile_X0Y1_E6END[0]
+ Tile_X0Y1_E6END[10] Tile_X0Y1_E6END[11] Tile_X0Y1_E6END[1] Tile_X0Y1_E6END[2] Tile_X0Y1_E6END[3]
+ Tile_X0Y1_E6END[4] Tile_X0Y1_E6END[5] Tile_X0Y1_E6END[6] Tile_X0Y1_E6END[7] Tile_X0Y1_E6END[8]
+ Tile_X0Y1_E6END[9] Tile_X0Y1_EE4BEG[0] Tile_X0Y1_EE4BEG[10] Tile_X0Y1_EE4BEG[11]
+ Tile_X0Y1_EE4BEG[12] Tile_X0Y1_EE4BEG[13] Tile_X0Y1_EE4BEG[14] Tile_X0Y1_EE4BEG[15]
+ Tile_X0Y1_EE4BEG[1] Tile_X0Y1_EE4BEG[2] Tile_X0Y1_EE4BEG[3] Tile_X0Y1_EE4BEG[4]
+ Tile_X0Y1_EE4BEG[5] Tile_X0Y1_EE4BEG[6] Tile_X0Y1_EE4BEG[7] Tile_X0Y1_EE4BEG[8]
+ Tile_X0Y1_EE4BEG[9] Tile_X0Y1_EE4END[0] Tile_X0Y1_EE4END[10] Tile_X0Y1_EE4END[11]
+ Tile_X0Y1_EE4END[12] Tile_X0Y1_EE4END[13] Tile_X0Y1_EE4END[14] Tile_X0Y1_EE4END[15]
+ Tile_X0Y1_EE4END[1] Tile_X0Y1_EE4END[2] Tile_X0Y1_EE4END[3] Tile_X0Y1_EE4END[4]
+ Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[6] Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[8]
+ Tile_X0Y1_EE4END[9] Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData[11]
+ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData[15]
+ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData[19]
+ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData[22]
+ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData[26]
+ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData[2]
+ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData[4]
+ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData[8]
+ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[0] Tile_X0Y1_FrameData_O[10] Tile_X0Y1_FrameData_O[11]
+ Tile_X0Y1_FrameData_O[12] Tile_X0Y1_FrameData_O[13] Tile_X0Y1_FrameData_O[14] Tile_X0Y1_FrameData_O[15]
+ Tile_X0Y1_FrameData_O[16] Tile_X0Y1_FrameData_O[17] Tile_X0Y1_FrameData_O[18] Tile_X0Y1_FrameData_O[19]
+ Tile_X0Y1_FrameData_O[1] Tile_X0Y1_FrameData_O[20] Tile_X0Y1_FrameData_O[21] Tile_X0Y1_FrameData_O[22]
+ Tile_X0Y1_FrameData_O[23] Tile_X0Y1_FrameData_O[24] Tile_X0Y1_FrameData_O[25] Tile_X0Y1_FrameData_O[26]
+ Tile_X0Y1_FrameData_O[27] Tile_X0Y1_FrameData_O[28] Tile_X0Y1_FrameData_O[29] Tile_X0Y1_FrameData_O[2]
+ Tile_X0Y1_FrameData_O[30] Tile_X0Y1_FrameData_O[31] Tile_X0Y1_FrameData_O[3] Tile_X0Y1_FrameData_O[4]
+ Tile_X0Y1_FrameData_O[5] Tile_X0Y1_FrameData_O[6] Tile_X0Y1_FrameData_O[7] Tile_X0Y1_FrameData_O[8]
+ Tile_X0Y1_FrameData_O[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_FrameStrobe[11]
+ Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_FrameStrobe[13] Tile_X0Y1_FrameStrobe[14] Tile_X0Y1_FrameStrobe[15]
+ Tile_X0Y1_FrameStrobe[16] Tile_X0Y1_FrameStrobe[17] Tile_X0Y1_FrameStrobe[18] Tile_X0Y1_FrameStrobe[19]
+ Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_FrameStrobe[4]
+ Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_FrameStrobe[8]
+ Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_N1END[0] Tile_X0Y1_N1END[1] Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[0] Tile_X0Y1_N2END[1] Tile_X0Y1_N2END[2] Tile_X0Y1_N2END[3]
+ Tile_X0Y1_N2END[4] Tile_X0Y1_N2END[5] Tile_X0Y1_N2END[6] Tile_X0Y1_N2END[7] Tile_X0Y1_N2MID[0]
+ Tile_X0Y1_N2MID[1] Tile_X0Y1_N2MID[2] Tile_X0Y1_N2MID[3] Tile_X0Y1_N2MID[4] Tile_X0Y1_N2MID[5]
+ Tile_X0Y1_N2MID[6] Tile_X0Y1_N2MID[7] Tile_X0Y1_N4END[0] Tile_X0Y1_N4END[10] Tile_X0Y1_N4END[11]
+ Tile_X0Y1_N4END[12] Tile_X0Y1_N4END[13] Tile_X0Y1_N4END[14] Tile_X0Y1_N4END[15]
+ Tile_X0Y1_N4END[1] Tile_X0Y1_N4END[2] Tile_X0Y1_N4END[3] Tile_X0Y1_N4END[4] Tile_X0Y1_N4END[5]
+ Tile_X0Y1_N4END[6] Tile_X0Y1_N4END[7] Tile_X0Y1_N4END[8] Tile_X0Y1_N4END[9] Tile_X0Y1_NN4END[0]
+ Tile_X0Y1_NN4END[10] Tile_X0Y1_NN4END[11] Tile_X0Y1_NN4END[12] Tile_X0Y1_NN4END[13]
+ Tile_X0Y1_NN4END[14] Tile_X0Y1_NN4END[15] Tile_X0Y1_NN4END[1] Tile_X0Y1_NN4END[2]
+ Tile_X0Y1_NN4END[3] Tile_X0Y1_NN4END[4] Tile_X0Y1_NN4END[5] Tile_X0Y1_NN4END[6]
+ Tile_X0Y1_NN4END[7] Tile_X0Y1_NN4END[8] Tile_X0Y1_NN4END[9] Tile_X0Y1_S1BEG[0] Tile_X0Y1_S1BEG[1]
+ Tile_X0Y1_S1BEG[2] Tile_X0Y1_S1BEG[3] Tile_X0Y1_S2BEG[0] Tile_X0Y1_S2BEG[1] Tile_X0Y1_S2BEG[2]
+ Tile_X0Y1_S2BEG[3] Tile_X0Y1_S2BEG[4] Tile_X0Y1_S2BEG[5] Tile_X0Y1_S2BEG[6] Tile_X0Y1_S2BEG[7]
+ Tile_X0Y1_S2BEGb[0] Tile_X0Y1_S2BEGb[1] Tile_X0Y1_S2BEGb[2] Tile_X0Y1_S2BEGb[3]
+ Tile_X0Y1_S2BEGb[4] Tile_X0Y1_S2BEGb[5] Tile_X0Y1_S2BEGb[6] Tile_X0Y1_S2BEGb[7]
+ Tile_X0Y1_S4BEG[0] Tile_X0Y1_S4BEG[10] Tile_X0Y1_S4BEG[11] Tile_X0Y1_S4BEG[12] Tile_X0Y1_S4BEG[13]
+ Tile_X0Y1_S4BEG[14] Tile_X0Y1_S4BEG[15] Tile_X0Y1_S4BEG[1] Tile_X0Y1_S4BEG[2] Tile_X0Y1_S4BEG[3]
+ Tile_X0Y1_S4BEG[4] Tile_X0Y1_S4BEG[5] Tile_X0Y1_S4BEG[6] Tile_X0Y1_S4BEG[7] Tile_X0Y1_S4BEG[8]
+ Tile_X0Y1_S4BEG[9] Tile_X0Y1_SS4BEG[0] Tile_X0Y1_SS4BEG[10] Tile_X0Y1_SS4BEG[11]
+ Tile_X0Y1_SS4BEG[12] Tile_X0Y1_SS4BEG[13] Tile_X0Y1_SS4BEG[14] Tile_X0Y1_SS4BEG[15]
+ Tile_X0Y1_SS4BEG[1] Tile_X0Y1_SS4BEG[2] Tile_X0Y1_SS4BEG[3] Tile_X0Y1_SS4BEG[4]
+ Tile_X0Y1_SS4BEG[5] Tile_X0Y1_SS4BEG[6] Tile_X0Y1_SS4BEG[7] Tile_X0Y1_SS4BEG[8]
+ Tile_X0Y1_SS4BEG[9] Tile_X0Y1_UserCLK Tile_X0Y1_W1BEG[0] Tile_X0Y1_W1BEG[1] Tile_X0Y1_W1BEG[2]
+ Tile_X0Y1_W1BEG[3] Tile_X0Y1_W1END[0] Tile_X0Y1_W1END[1] Tile_X0Y1_W1END[2] Tile_X0Y1_W1END[3]
+ Tile_X0Y1_W2BEG[0] Tile_X0Y1_W2BEG[1] Tile_X0Y1_W2BEG[2] Tile_X0Y1_W2BEG[3] Tile_X0Y1_W2BEG[4]
+ Tile_X0Y1_W2BEG[5] Tile_X0Y1_W2BEG[6] Tile_X0Y1_W2BEG[7] Tile_X0Y1_W2BEGb[0] Tile_X0Y1_W2BEGb[1]
+ Tile_X0Y1_W2BEGb[2] Tile_X0Y1_W2BEGb[3] Tile_X0Y1_W2BEGb[4] Tile_X0Y1_W2BEGb[5]
+ Tile_X0Y1_W2BEGb[6] Tile_X0Y1_W2BEGb[7] Tile_X0Y1_W2END[0] Tile_X0Y1_W2END[1] Tile_X0Y1_W2END[2]
+ Tile_X0Y1_W2END[3] Tile_X0Y1_W2END[4] Tile_X0Y1_W2END[5] Tile_X0Y1_W2END[6] Tile_X0Y1_W2END[7]
+ Tile_X0Y1_W2MID[0] Tile_X0Y1_W2MID[1] Tile_X0Y1_W2MID[2] Tile_X0Y1_W2MID[3] Tile_X0Y1_W2MID[4]
+ Tile_X0Y1_W2MID[5] Tile_X0Y1_W2MID[6] Tile_X0Y1_W2MID[7] Tile_X0Y1_W6BEG[0] Tile_X0Y1_W6BEG[10]
+ Tile_X0Y1_W6BEG[11] Tile_X0Y1_W6BEG[1] Tile_X0Y1_W6BEG[2] Tile_X0Y1_W6BEG[3] Tile_X0Y1_W6BEG[4]
+ Tile_X0Y1_W6BEG[5] Tile_X0Y1_W6BEG[6] Tile_X0Y1_W6BEG[7] Tile_X0Y1_W6BEG[8] Tile_X0Y1_W6BEG[9]
+ Tile_X0Y1_W6END[0] Tile_X0Y1_W6END[10] Tile_X0Y1_W6END[11] Tile_X0Y1_W6END[1] Tile_X0Y1_W6END[2]
+ Tile_X0Y1_W6END[3] Tile_X0Y1_W6END[4] Tile_X0Y1_W6END[5] Tile_X0Y1_W6END[6] Tile_X0Y1_W6END[7]
+ Tile_X0Y1_W6END[8] Tile_X0Y1_W6END[9] Tile_X0Y1_WW4BEG[0] Tile_X0Y1_WW4BEG[10] Tile_X0Y1_WW4BEG[11]
+ Tile_X0Y1_WW4BEG[12] Tile_X0Y1_WW4BEG[13] Tile_X0Y1_WW4BEG[14] Tile_X0Y1_WW4BEG[15]
+ Tile_X0Y1_WW4BEG[1] Tile_X0Y1_WW4BEG[2] Tile_X0Y1_WW4BEG[3] Tile_X0Y1_WW4BEG[4]
+ Tile_X0Y1_WW4BEG[5] Tile_X0Y1_WW4BEG[6] Tile_X0Y1_WW4BEG[7] Tile_X0Y1_WW4BEG[8]
+ Tile_X0Y1_WW4BEG[9] Tile_X0Y1_WW4END[0] Tile_X0Y1_WW4END[10] Tile_X0Y1_WW4END[11]
+ Tile_X0Y1_WW4END[12] Tile_X0Y1_WW4END[13] Tile_X0Y1_WW4END[14] Tile_X0Y1_WW4END[15]
+ Tile_X0Y1_WW4END[1] Tile_X0Y1_WW4END[2] Tile_X0Y1_WW4END[3] Tile_X0Y1_WW4END[4]
+ Tile_X0Y1_WW4END[5] Tile_X0Y1_WW4END[6] Tile_X0Y1_WW4END[7] Tile_X0Y1_WW4END[8]
+ Tile_X0Y1_WW4END[9] VGND VPWR
X_3155_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q VPWR _1211_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q _1210_ sg13g2_o21ai_1
X_3086_ _1144_ VPWR _1145_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q
+ _1143_ sg13g2_o21ai_1
X_3988_ net1701 net681 net1709 net1 net4 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q
+ _1993_ VPWR VGND sg13g2_mux4_1
X_5727_ net1859 net1739 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_2939_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6
+ net79 net44 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q
+ _1004_ VPWR VGND sg13g2_mux4_1
X_5658_ net1910 net1758 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_117_11 VPWR VGND sg13g2_fill_1
X_4609_ VPWR _0166_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q
+ VGND sg13g2_inv_1
X_5589_ net1901 net1782 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
Xfanout1807 net1808 net1807 VPWR VGND sg13g2_buf_1
Xfanout1829 net1830 net1829 VPWR VGND sg13g2_buf_1
Xfanout1818 net1819 net1818 VPWR VGND sg13g2_buf_1
Xrebuffer7 net634 net616 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_76_350 VPWR VGND sg13g2_fill_2
XFILLER_36_214 VPWR VGND sg13g2_fill_2
XFILLER_36_236 VPWR VGND sg13g2_fill_1
X_4960_ _0502_ VPWR _0503_ VGND net1695 net32 sg13g2_o21ai_1
X_4891_ _0436_ VPWR _0437_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 sg13g2_o21ai_1
X_3911_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q _1921_ _1922_
+ net1576 _1923_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X
+ VPWR VGND sg13g2_mux4_1
X_3842_ _1173_ net697 _1869_ VPWR VGND sg13g2_nor2_2
X_3773_ net1643 _1801_ _1802_ VPWR VGND sg13g2_nor2_2
X_5512_ net1871 net1811 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_2724_ VGND VPWR net1924 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q
+ _0802_ _0801_ sg13g2_a21oi_1
XFILLER_66_0 VPWR VGND sg13g2_fill_2
Xoutput401 net401 Tile_X0Y1_E6BEG[5] VPWR VGND sg13g2_buf_1
X_2655_ _0735_ VPWR _0736_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ net1531 sg13g2_o21ai_1
X_5443_ Tile_X0Y1_UserCLK net575 _0057_ _5443_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[19\]
+ VPWR VGND sg13g2_dfrbp_1
Xoutput412 net412 Tile_X0Y1_EE4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput434 net434 Tile_X0Y1_FrameData_O[20] VPWR VGND sg13g2_buf_1
Xoutput423 net423 Tile_X0Y1_FrameData_O[10] VPWR VGND sg13g2_buf_1
X_5374_ net1961 net1828 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_2586_ _0670_ VPWR _0671_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q
+ _0667_ sg13g2_o21ai_1
X_4325_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q net1711 net89
+ net149 net1544 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q _2259_
+ VPWR VGND sg13g2_mux4_1
Xoutput456 net456 Tile_X0Y1_S1BEG[2] VPWR VGND sg13g2_buf_1
Xoutput467 net467 Tile_X0Y1_S2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput478 net478 Tile_X0Y1_S4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput445 net445 Tile_X0Y1_FrameData_O[30] VPWR VGND sg13g2_buf_1
XFILLER_113_252 VPWR VGND sg13g2_fill_2
Xoutput489 net489 Tile_X0Y1_S4BEG[9] VPWR VGND sg13g2_buf_1
X_4256_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q net1589 net1523
+ net1519 net1541 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q _2215_
+ VPWR VGND sg13g2_mux4_1
XFILLER_47_18 VPWR VGND sg13g2_fill_1
X_3207_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q net1712 net120
+ net1927 net96 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q _1262_
+ VPWR VGND sg13g2_mux4_1
X_4187_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q net3 net1600
+ net1932 net1613 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q _2155_
+ VPWR VGND sg13g2_mux4_1
X_3138_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q _1194_
+ _1195_ _0120_ sg13g2_a21oi_1
XFILLER_27_225 VPWR VGND sg13g2_decap_4
XFILLER_27_203 VPWR VGND sg13g2_decap_4
XFILLER_67_383 VPWR VGND sg13g2_fill_2
X_3069_ _0127_ VPWR _1129_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q
+ _1128_ sg13g2_o21ai_1
XFILLER_63_28 VPWR VGND sg13g2_decap_8
XFILLER_50_250 VPWR VGND sg13g2_fill_2
XFILLER_50_283 VPWR VGND sg13g2_fill_1
XFILLER_10_169 VPWR VGND sg13g2_fill_1
Xfanout1615 net1615 net1616 VPWR VGND sg13g2_buf_16
Xfanout1648 net1651 net1648 VPWR VGND sg13g2_buf_1
Xfanout1637 net1639 net1637 VPWR VGND sg13g2_buf_1
Xfanout1626 net1627 net1626 VPWR VGND sg13g2_buf_1
XFILLER_104_285 VPWR VGND sg13g2_fill_1
Xfanout1659 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q net1659 VPWR
+ VGND sg13g2_buf_1
X_5090_ net1970 net1799 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_4110_ VGND VPWR net5 net1672 _2099_ _2098_ sg13g2_a21oi_1
X_4041_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q _2044_
+ _2045_ _0157_ sg13g2_a21oi_1
XFILLER_68_158 VPWR VGND sg13g2_fill_2
X_5992_ Tile_X0Y0_EE4END[12] net219 VPWR VGND sg13g2_buf_1
X_4943_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q _0484_
+ _0486_ _0485_ sg13g2_a21oi_1
X_4874_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q _0420_
+ _0421_ _0078_ sg13g2_a21oi_1
X_3825_ VGND VPWR net37 net1678 _1854_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q
+ sg13g2_a21oi_1
X_3756_ _1427_ VPWR _1786_ VGND _1214_ net1548 sg13g2_o21ai_1
XFILLER_118_344 VPWR VGND sg13g2_fill_2
X_2707_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q net1528 net1542
+ net1549 net1556 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q _0786_
+ VPWR VGND sg13g2_mux4_1
X_5426_ Tile_X0Y1_UserCLK net572 _0040_ _0020_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[2\]
+ VPWR VGND sg13g2_dfrbp_1
X_3687_ VGND VPWR net125 _0153_ _1722_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q
+ sg13g2_a21oi_1
Xoutput231 net231 Tile_X0Y0_FrameData_O[19] VPWR VGND sg13g2_buf_1
Xoutput253 net253 Tile_X0Y0_FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
Xoutput242 net242 Tile_X0Y0_FrameData_O[29] VPWR VGND sg13g2_buf_1
X_2638_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q _0719_ _0717_
+ _0713_ _0715_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q _0720_
+ VPWR VGND sg13g2_mux4_1
Xoutput220 net220 Tile_X0Y0_EE4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput264 net264 Tile_X0Y0_FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
Xoutput275 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 Tile_X0Y0_N1BEG[2]
+ VPWR VGND sg13g2_buf_1
Xoutput286 net286 Tile_X0Y0_N2BEGb[1] VPWR VGND sg13g2_buf_1
X_5357_ net1994 net1839 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_2569_ net1682 net137 _0655_ VPWR VGND sg13g2_nor2b_1
Xoutput297 net297 Tile_X0Y0_N4BEG[13] VPWR VGND sg13g2_buf_1
X_4308_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q net1564 net693
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 _0308_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 VPWR VGND sg13g2_mux4_1
XFILLER_59_136 VPWR VGND sg13g2_decap_8
X_5288_ net1984 net1729 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_99_294 VPWR VGND sg13g2_fill_1
XFILLER_101_266 VPWR VGND sg13g2_decap_4
X_4239_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q _2199_
+ _2200_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q sg13g2_a21oi_1
XFILLER_114_67 VPWR VGND sg13g2_fill_1
XFILLER_74_106 VPWR VGND sg13g2_fill_2
X_5456__588 VPWR VGND net588 sg13g2_tiehi
XFILLER_30_209 VPWR VGND sg13g2_decap_4
XFILLER_99_46 VPWR VGND sg13g2_fill_1
XFILLER_99_68 VPWR VGND sg13g2_fill_1
XFILLER_46_331 VPWR VGND sg13g2_fill_1
XFILLER_58_191 VPWR VGND sg13g2_fill_1
XFILLER_61_312 VPWR VGND sg13g2_fill_2
XFILLER_9_44 VPWR VGND sg13g2_fill_2
X_4590_ VPWR _0147_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q VGND
+ sg13g2_inv_1
X_3610_ VGND VPWR _1648_ _1649_ _1647_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q
+ sg13g2_a21oi_2
X_3541_ _1586_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q net1619
+ VPWR VGND sg13g2_nand2b_1
X_6260_ Tile_X0Y0_S4END[15] net487 VPWR VGND sg13g2_buf_1
X_3472_ VGND VPWR _0086_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q
+ _1521_ _1520_ sg13g2_a21oi_1
X_6191_ Tile_X0Y1_EE4END[10] net418 VPWR VGND sg13g2_buf_1
X_5211_ net1953 net1756 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_5142_ net1949 net1789 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_29_0 VPWR VGND sg13g2_fill_2
X_5073_ net1939 net1810 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_5479__555 VPWR VGND net555 sg13g2_tiehi
X_4024_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5
+ _2028_ VPWR VGND sg13g2_nor2b_1
Xfanout1990 Tile_X0Y0_FrameData[14] net1990 VPWR VGND sg13g2_buf_1
X_5975_ Tile_X0Y0_E6END[5] net198 VPWR VGND sg13g2_buf_1
X_4926_ _0469_ VPWR _0470_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q
+ net1577 sg13g2_o21ai_1
X_4857_ _0405_ net1685 net34 VPWR VGND sg13g2_nand2_1
X_3808_ _1836_ VPWR _1837_ VGND net49 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q
+ sg13g2_o21ai_1
XFILLER_118_141 VPWR VGND sg13g2_fill_2
X_4788_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q VPWR _0339_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q _0337_ sg13g2_o21ai_1
XFILLER_109_23 VPWR VGND sg13g2_fill_2
X_3739_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q net141 net52
+ net93 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q
+ _1770_ VPWR VGND sg13g2_mux4_1
XFILLER_109_67 VPWR VGND sg13g2_fill_2
X_5409_ net1968 net1817 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_70_175 VPWR VGND sg13g2_decap_8
XFILLER_70_197 VPWR VGND sg13g2_decap_8
XFILLER_46_194 VPWR VGND sg13g2_decap_4
XFILLER_34_345 VPWR VGND sg13g2_fill_1
X_5760_ net1861 net1726 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_2972_ VGND VPWR _1035_ _1032_ _1034_ sg13g2_or2_1
X_5691_ net1913 net1747 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_4711_ _0263_ VPWR _0264_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q
+ _0261_ sg13g2_o21ai_1
X_4642_ VGND VPWR net1657 net1569 _0199_ _0198_ sg13g2_a21oi_1
X_4573_ VPWR _0130_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q VGND
+ sg13g2_inv_1
X_6312_ Tile_X0Y1_W6END[9] net535 VPWR VGND sg13g2_buf_1
X_3524_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q VPWR _1570_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q net1571 sg13g2_o21ai_1
X_6243_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 net464 VPWR VGND sg13g2_buf_2
X_3455_ _1504_ _1502_ _1503_ _0002_ net1650 VPWR VGND sg13g2_a22oi_1
XFILLER_115_188 VPWR VGND sg13g2_fill_1
X_6174_ Tile_X0Y1_E6END[3] net397 VPWR VGND sg13g2_buf_1
X_3386_ _1431_ _1426_ _1438_ VPWR VGND sg13g2_xor2_1
X_5125_ net1975 net1785 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_29_117 VPWR VGND sg13g2_decap_4
X_5056_ net1965 net1809 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_4007_ _0230_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q _2012_
+ VPWR VGND sg13g2_nor2_2
XFILLER_71_17 VPWR VGND sg13g2_fill_1
XFILLER_71_28 VPWR VGND sg13g2_fill_2
X_5958_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 net179 VPWR VGND sg13g2_buf_1
X_4909_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q _0112_
+ _0454_ _0451_ _0455_ _0452_ sg13g2_a221oi_1
XFILLER_40_359 VPWR VGND sg13g2_fill_2
XFILLER_71_39 VPWR VGND sg13g2_fill_1
X_5889_ net1862 net1813 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_75_234 VPWR VGND sg13g2_fill_2
XFILLER_102_383 VPWR VGND sg13g2_fill_2
X_5471__603 VPWR VGND net603 sg13g2_tiehi
XFILLER_43_164 VPWR VGND sg13g2_decap_8
XFILLER_61_61 VPWR VGND sg13g2_fill_1
XFILLER_6_45 VPWR VGND sg13g2_fill_1
XFILLER_112_136 VPWR VGND sg13g2_decap_4
X_3240_ VGND VPWR _1241_ _1293_ _1292_ _1290_ sg13g2_a21oi_2
X_3171_ net1628 _0702_ _1224_ _1226_ VPWR VGND sg13g2_a21o_1
XFILLER_19_183 VPWR VGND sg13g2_fill_1
XFILLER_19_161 VPWR VGND sg13g2_fill_2
Xrebuffer28 net636 net637 VPWR VGND sg13g2_buf_2
Xrebuffer39 net648 net1607 VPWR VGND sg13g2_buf_16
XFILLER_34_142 VPWR VGND sg13g2_fill_2
X_5812_ net1898 net1836 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_5743_ net1886 net1726 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_2955_ _1016_ _1018_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q
+ _1019_ VPWR VGND sg13g2_nand3_1
X_2886_ _0955_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q _0953_
+ VPWR VGND sg13g2_nand2b_1
X_5674_ net1876 net1747 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
Xrebuffer129 net739 net738 VPWR VGND sg13g2_buf_2
Xrebuffer107 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 net716 VPWR VGND
+ sg13g2_buf_2
Xrebuffer118 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 net727 VPWR VGND
+ sg13g2_dlygate4sd1_1
X_4625_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q net1591 net1587
+ net1522 net1539 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q _0182_
+ VPWR VGND sg13g2_mux4_1
X_4556_ VPWR _0113_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q VGND
+ sg13g2_inv_1
X_3507_ VGND VPWR net1705 net1670 _1554_ _1553_ sg13g2_a21oi_1
X_4487_ net1512 _1890_ _0044_ VPWR VGND sg13g2_nor2_1
X_3438_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q VPWR _1489_ VGND
+ _1485_ _1487_ sg13g2_o21ai_1
X_6226_ net1885 net439 VPWR VGND sg13g2_buf_1
X_6157_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 net378 VPWR VGND sg13g2_buf_1
X_3369_ _1421_ _1419_ _1420_ VPWR VGND sg13g2_xnor2_1
X_5108_ net1945 net1796 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_6088_ Tile_X0Y1_NN4END[8] net309 VPWR VGND sg13g2_buf_1
XFILLER_72_237 VPWR VGND sg13g2_fill_2
X_5039_ net1997 net1852 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_122_67 VPWR VGND sg13g2_fill_2
XFILLER_25_131 VPWR VGND sg13g2_fill_1
XFILLER_13_315 VPWR VGND sg13g2_fill_1
XFILLER_31_20 VPWR VGND sg13g2_fill_1
XFILLER_31_31 VPWR VGND sg13g2_fill_2
Xinput120 Tile_X0Y1_N2END[5] net120 VPWR VGND sg13g2_buf_1
Xinput131 Tile_X0Y1_N4END[0] net131 VPWR VGND sg13g2_buf_1
Xinput153 Tile_X0Y1_W2END[2] net153 VPWR VGND sg13g2_buf_1
Xinput142 Tile_X0Y1_NN4END[3] net142 VPWR VGND sg13g2_buf_1
Xinput164 Tile_X0Y1_W2MID[5] net164 VPWR VGND sg13g2_buf_1
XFILLER_63_259 VPWR VGND sg13g2_fill_1
XFILLER_72_82 VPWR VGND sg13g2_fill_2
X_2740_ VGND VPWR _0074_ net1697 _0817_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q
+ sg13g2_a21oi_1
X_2671_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 _0749_ _0751_ _0747_
+ _0745_ VPWR VGND sg13g2_a22oi_1
X_4410_ _2332_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q _1780_
+ VPWR VGND sg13g2_nand2_1
X_5390_ net1996 net1827 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_4341_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q _2272_ _2273_
+ VPWR VGND sg13g2_nor2_1
X_4272_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q net117 net1921
+ net132 net1556 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A
+ VPWR VGND sg13g2_mux4_1
X_6011_ net1996 net223 VPWR VGND sg13g2_buf_1
X_3223_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q net126 net102
+ net639 net162 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q _1277_
+ VPWR VGND sg13g2_mux4_1
XFILLER_100_106 VPWR VGND sg13g2_fill_2
XFILLER_11_0 VPWR VGND sg13g2_fill_2
X_3154_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q net121 net97 net61
+ net157 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q _1210_ VPWR VGND
+ sg13g2_mux4_1
X_3085_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q _1142_ _1144_
+ VPWR VGND sg13g2_nor2_1
X_3987_ _1991_ VPWR _1992_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q
+ _0594_ sg13g2_o21ai_1
X_2938_ _0995_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 VGND _1003_
+ _1001_ sg13g2_o21ai_1
X_5726_ net1857 net1739 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_5657_ net1908 net1760 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_2869_ net1686 net1593 net1588 net1524 net1519 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q
+ _0939_ VPWR VGND sg13g2_mux4_1
X_5588_ net1898 net1784 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_4608_ VPWR _0165_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q VGND
+ sg13g2_inv_1
XFILLER_116_283 VPWR VGND sg13g2_fill_1
X_4539_ VPWR _0096_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q VGND
+ sg13g2_inv_1
X_6209_ net1858 net452 VPWR VGND sg13g2_buf_1
Xfanout1819 net1820 net1819 VPWR VGND sg13g2_buf_1
Xfanout1808 net1811 net1808 VPWR VGND sg13g2_buf_1
XFILLER_85_384 VPWR VGND sg13g2_fill_1
XFILLER_26_97 VPWR VGND sg13g2_fill_1
XFILLER_42_41 VPWR VGND sg13g2_fill_2
Xrebuffer8 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 net617 VPWR VGND sg13g2_buf_2
XFILLER_68_318 VPWR VGND sg13g2_fill_2
XFILLER_67_60 VPWR VGND sg13g2_fill_1
XFILLER_95_148 VPWR VGND sg13g2_decap_4
X_4890_ VGND VPWR _0080_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q
+ _0436_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q sg13g2_a21oi_1
X_3910_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q net137 net56
+ net67 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q
+ _1923_ VPWR VGND sg13g2_mux4_1
X_3841_ _1868_ _1463_ _1176_ VPWR VGND sg13g2_nand2b_1
X_3772_ VPWR Tile_X0Y1_DSP_bot.C0 net704 VGND sg13g2_inv_1
X_2723_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q net131 _0801_
+ VPWR VGND sg13g2_nor2b_1
X_5511_ net1919 net1845 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput402 net402 Tile_X0Y1_E6BEG[6] VPWR VGND sg13g2_buf_1
X_2654_ _0735_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q _0180_
+ VPWR VGND sg13g2_nand2_1
X_5442_ Tile_X0Y1_UserCLK net556 _0056_ _0036_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[18\]
+ VPWR VGND sg13g2_dfrbp_1
X_2585_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q _0669_
+ _0670_ _0089_ sg13g2_a21oi_1
Xoutput413 net413 Tile_X0Y1_EE4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput424 net424 Tile_X0Y1_FrameData_O[11] VPWR VGND sg13g2_buf_1
Xoutput435 net435 Tile_X0Y1_FrameData_O[21] VPWR VGND sg13g2_buf_1
X_5373_ net1960 net1830 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_4324_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q net1529 _0596_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 _0566_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 VPWR VGND sg13g2_mux4_1
Xoutput468 net468 Tile_X0Y1_S2BEGb[2] VPWR VGND sg13g2_buf_1
Xoutput457 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 Tile_X0Y1_S1BEG[3]
+ VPWR VGND sg13g2_buf_1
Xoutput446 net446 Tile_X0Y1_FrameData_O[31] VPWR VGND sg13g2_buf_1
Xoutput479 net479 Tile_X0Y1_S4BEG[14] VPWR VGND sg13g2_buf_1
X_4255_ _2213_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q _2214_
+ VPWR VGND sg13g2_nor2b_1
X_3206_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q net645 _0724_
+ _0099_ _0105_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q _1261_
+ VPWR VGND sg13g2_mux4_1
XFILLER_67_351 VPWR VGND sg13g2_fill_2
X_4186_ _2150_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 VGND _2152_
+ _2154_ sg13g2_o21ai_1
X_3137_ _1193_ VPWR _1194_ VGND net1933 net1691 sg13g2_o21ai_1
X_3068_ net1668 net112 net120 net1927 net96 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q
+ _1128_ VPWR VGND sg13g2_mux4_1
X_5709_ net1883 net1737 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_358 VPWR VGND sg13g2_fill_2
Xfanout1605 net1606 net1605 VPWR VGND sg13g2_buf_1
Xfanout1616 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 net1616 VPWR VGND sg13g2_buf_8
Xfanout1649 net1650 net1649 VPWR VGND sg13g2_buf_1
Xfanout1627 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 net1627 VPWR VGND
+ sg13g2_buf_8
Xfanout1638 net1639 net1638 VPWR VGND sg13g2_buf_1
XFILLER_68_104 VPWR VGND sg13g2_fill_1
XFILLER_78_70 VPWR VGND sg13g2_decap_8
XFILLER_78_81 VPWR VGND sg13g2_decap_4
X_4040_ _2043_ VPWR _2044_ VGND net62 net1679 sg13g2_o21ai_1
XFILLER_64_332 VPWR VGND sg13g2_fill_1
X_5991_ Tile_X0Y0_EE4END[11] net218 VPWR VGND sg13g2_buf_1
XFILLER_17_270 VPWR VGND sg13g2_fill_1
X_4942_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q VPWR _0485_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q _0483_ sg13g2_o21ai_1
X_4873_ net147 net1705 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q
+ _0420_ VPWR VGND sg13g2_mux2_1
X_3824_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q _1852_
+ _1853_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q sg13g2_a21oi_1
X_3755_ _1769_ VPWR _1785_ VGND _1784_ net1647 sg13g2_o21ai_1
X_2706_ _0778_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q _0784_
+ _0785_ VPWR VGND sg13g2_or3_1
X_3686_ _1721_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q net715
+ VPWR VGND sg13g2_nand2_1
Xoutput210 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 Tile_X0Y0_EE4BEG[14]
+ VPWR VGND sg13g2_buf_1
X_5425_ Tile_X0Y1_UserCLK net573 _0039_ _0022_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[1\]
+ VPWR VGND sg13g2_dfrbp_1
X_2637_ _0718_ VPWR _0719_ VGND net125 net1674 sg13g2_o21ai_1
Xoutput221 net221 Tile_X0Y0_FrameData_O[0] VPWR VGND sg13g2_buf_1
Xoutput243 net243 Tile_X0Y0_FrameData_O[2] VPWR VGND sg13g2_buf_1
Xoutput232 net232 Tile_X0Y0_FrameData_O[1] VPWR VGND sg13g2_buf_1
Xoutput254 net254 Tile_X0Y0_FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
Xoutput265 net265 Tile_X0Y0_FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
Xoutput276 net276 Tile_X0Y0_N1BEG[3] VPWR VGND sg13g2_buf_8
X_2568_ _0653_ VPWR _0654_ VGND net1682 net687 sg13g2_o21ai_1
X_5356_ net1992 net1839 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_2499_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q _0086_
+ _0588_ _0587_ sg13g2_a21oi_1
Xoutput298 net298 Tile_X0Y0_N4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput287 net287 Tile_X0Y0_N2BEGb[2] VPWR VGND sg13g2_buf_1
X_4307_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q net1936 net50
+ net167 net1551 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3
+ VPWR VGND sg13g2_mux4_1
X_5287_ net1981 net1732 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_212 VPWR VGND sg13g2_fill_2
X_4238_ net62 net1630 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q
+ _2199_ VPWR VGND sg13g2_mux2_1
X_4169_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q net1576 _2140_
+ VPWR VGND sg13g2_nor2_1
XFILLER_74_28 VPWR VGND sg13g2_fill_2
XFILLER_82_162 VPWR VGND sg13g2_decap_4
XFILLER_58_181 VPWR VGND sg13g2_fill_1
XFILLER_9_67 VPWR VGND sg13g2_fill_2
XFILLER_80_82 VPWR VGND sg13g2_decap_4
X_3540_ _1584_ VPWR _1585_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q
+ net1555 sg13g2_o21ai_1
X_3471_ net28 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q _1520_
+ VPWR VGND sg13g2_nor2_1
X_5210_ net1951 net1753 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_115_359 VPWR VGND sg13g2_fill_2
X_6190_ Tile_X0Y1_EE4END[9] net417 VPWR VGND sg13g2_buf_1
X_5141_ net1947 net1789 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_96_221 VPWR VGND sg13g2_decap_8
X_5072_ net1937 net1810 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_96_232 VPWR VGND sg13g2_fill_2
X_4023_ _2027_ _2020_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 VPWR VGND
+ sg13g2_nor2_2
XFILLER_56_129 VPWR VGND sg13g2_fill_1
Xfanout1980 Tile_X0Y0_FrameData[19] net1980 VPWR VGND sg13g2_buf_1
XFILLER_49_192 VPWR VGND sg13g2_decap_4
Xfanout1991 net1992 net1991 VPWR VGND sg13g2_buf_1
XFILLER_52_324 VPWR VGND sg13g2_fill_1
X_5974_ Tile_X0Y0_E6END[4] net197 VPWR VGND sg13g2_buf_1
X_4925_ _0469_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q _0178_
+ VPWR VGND sg13g2_nand2_1
X_4856_ _0403_ VPWR _0404_ VGND net1684 net69 sg13g2_o21ai_1
X_3807_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q VPWR _1836_ VGND
+ _0445_ _0456_ sg13g2_o21ai_1
X_4787_ net1584 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 net1692 _0338_
+ VPWR VGND sg13g2_mux2_1
X_3738_ _1769_ net1647 _0022_ VPWR VGND sg13g2_nand2_1
X_3669_ _1702_ _1704_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q
+ _1705_ VPWR VGND sg13g2_nand3_1
XFILLER_109_57 VPWR VGND sg13g2_fill_2
X_5408_ net1966 net1817 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_5339_ net1953 net1840 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_105_370 VPWR VGND sg13g2_fill_2
XFILLER_59_94 VPWR VGND sg13g2_decap_4
XFILLER_93_202 VPWR VGND sg13g2_fill_2
XFILLER_93_257 VPWR VGND sg13g2_fill_2
X_2971_ _1034_ _1033_ _1031_ VPWR VGND sg13g2_nand2_2
X_5690_ net1910 net1747 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_4710_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q _0262_
+ _0263_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q sg13g2_a21oi_1
X_4641_ net1657 net1563 _0198_ VPWR VGND sg13g2_nor2_1
X_4572_ VPWR _0129_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q VGND
+ sg13g2_inv_1
X_6311_ Tile_X0Y1_W6END[8] net534 VPWR VGND sg13g2_buf_1
X_3523_ _0143_ _1568_ _1569_ VPWR VGND sg13g2_and2_1
XFILLER_115_156 VPWR VGND sg13g2_decap_8
X_6242_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 net463 VPWR VGND sg13g2_buf_2
X_3454_ VGND VPWR net1645 _0136_ _1503_ net1650 sg13g2_a21oi_1
XFILLER_41_0 VPWR VGND sg13g2_decap_4
X_6173_ Tile_X0Y1_E6END[2] net394 VPWR VGND sg13g2_buf_1
X_3385_ _1426_ _1431_ _1437_ VPWR VGND sg13g2_nor2_1
X_5124_ net1973 net1785 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_5055_ net1964 net1809 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_4006_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q VPWR _2011_ VGND
+ _2009_ _2010_ sg13g2_o21ai_1
XFILLER_84_268 VPWR VGND sg13g2_fill_2
X_5957_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 net178 VPWR VGND sg13g2_buf_1
X_4908_ _0453_ VPWR _0454_ VGND net1933 net1677 sg13g2_o21ai_1
X_5888_ net1860 net1813 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_4839_ VGND VPWR _0386_ _0387_ net1539 net1685 sg13g2_a21oi_2
XFILLER_105_5 VPWR VGND sg13g2_fill_2
XFILLER_29_42 VPWR VGND sg13g2_fill_1
XFILLER_83_290 VPWR VGND sg13g2_fill_2
XFILLER_45_96 VPWR VGND sg13g2_fill_2
XFILLER_101_80 VPWR VGND sg13g2_decap_8
XFILLER_101_91 VPWR VGND sg13g2_fill_1
XFILLER_3_250 VPWR VGND sg13g2_fill_2
X_3170_ net1628 _1224_ _0702_ _1225_ VPWR VGND sg13g2_nand3_1
Xrebuffer29 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 net638 VPWR VGND
+ sg13g2_buf_2
X_5811_ net1895 net1836 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_5742_ net1884 net1726 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_2954_ _1017_ VPWR _1018_ VGND net24 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q
+ sg13g2_o21ai_1
X_2885_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q net1529 net1535
+ net1550 net1559 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q _0954_
+ VPWR VGND sg13g2_mux4_1
Xrebuffer119 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 net728 VPWR VGND
+ sg13g2_dlygate4sd1_1
Xrebuffer108 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 net717 VPWR VGND
+ sg13g2_dlygate4sd1_1
X_5673_ net1873 net1752 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_4624_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q net1598 net1611
+ net1603 net1633 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q _0181_
+ VPWR VGND sg13g2_mux4_1
X_4555_ VPWR _0112_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q VGND
+ sg13g2_inv_1
X_3506_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q VPWR _1553_ VGND
+ _0095_ net1669 sg13g2_o21ai_1
X_4486_ net1512 _1889_ _0043_ VPWR VGND sg13g2_nor2b_1
X_3437_ net1687 net1598 net1611 net1603 net1623 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q
+ _1488_ VPWR VGND sg13g2_mux4_1
X_6225_ net1887 net438 VPWR VGND sg13g2_buf_1
X_3368_ _1403_ _1395_ _1420_ VPWR VGND sg13g2_xor2_1
X_5107_ net1943 net1796 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_3299_ _1351_ _1350_ _1242_ VPWR VGND sg13g2_nand2b_1
X_6087_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 net299 VPWR VGND sg13g2_buf_1
X_5038_ net1995 net1852 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_25_176 VPWR VGND sg13g2_fill_1
XFILLER_40_157 VPWR VGND sg13g2_fill_1
XFILLER_31_76 VPWR VGND sg13g2_fill_2
XFILLER_103_2 VPWR VGND sg13g2_fill_1
XFILLER_0_220 VPWR VGND sg13g2_fill_1
Xinput110 Tile_X0Y1_EE4END[3] net110 VPWR VGND sg13g2_buf_1
Xinput121 Tile_X0Y1_N2END[6] net121 VPWR VGND sg13g2_buf_1
Xinput132 Tile_X0Y1_N4END[1] net132 VPWR VGND sg13g2_buf_1
Xinput154 Tile_X0Y1_W2END[3] net154 VPWR VGND sg13g2_buf_1
Xinput143 Tile_X0Y1_NN4END[4] net143 VPWR VGND sg13g2_buf_1
XFILLER_48_235 VPWR VGND sg13g2_fill_2
Xinput165 Tile_X0Y1_W2MID[6] net165 VPWR VGND sg13g2_buf_1
XFILLER_16_110 VPWR VGND sg13g2_fill_1
XFILLER_63_238 VPWR VGND sg13g2_decap_4
XFILLER_16_187 VPWR VGND sg13g2_fill_2
XFILLER_72_61 VPWR VGND sg13g2_decap_4
XFILLER_12_360 VPWR VGND sg13g2_fill_2
XFILLER_31_179 VPWR VGND sg13g2_decap_4
X_2670_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q _0750_
+ _0751_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q sg13g2_a21oi_1
XFILLER_117_218 VPWR VGND sg13g2_fill_2
XFILLER_8_375 VPWR VGND sg13g2_fill_2
X_4340_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q net1713 net1928
+ net147 net1559 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q _2272_
+ VPWR VGND sg13g2_mux4_1
X_4271_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q net1602 _0194_
+ net701 _0385_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0
+ VPWR VGND sg13g2_mux4_1
X_3222_ _1275_ VPWR _1276_ VGND _1272_ _1273_ sg13g2_o21ai_1
XFILLER_86_319 VPWR VGND sg13g2_fill_1
X_6010_ net1998 net222 VPWR VGND sg13g2_buf_1
X_3153_ _1208_ _1202_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q
+ _1209_ VPWR VGND sg13g2_nor3_2
XFILLER_39_246 VPWR VGND sg13g2_fill_1
X_3084_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q net142 net1927
+ net94 net1922 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q _1143_
+ VPWR VGND sg13g2_mux4_1
XFILLER_54_238 VPWR VGND sg13g2_fill_2
X_3986_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7
+ _1991_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q sg13g2_a21oi_1
X_5725_ net1918 net1737 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_2937_ _0106_ VPWR _1003_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q
+ _1002_ sg13g2_o21ai_1
X_5656_ net1906 net1758 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_2868_ VPWR _0938_ _0937_ VGND sg13g2_inv_1
X_4607_ VPWR _0164_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q VGND
+ sg13g2_inv_1
X_5587_ net1895 net1783 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_2799_ net1596 net1609 net1688 _0873_ VPWR VGND sg13g2_mux2_1
X_4538_ VPWR _0095_ net44 VGND sg13g2_inv_1
X_4469_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q
+ _2383_ VPWR VGND sg13g2_nor2b_1
Xfanout1809 net1811 net1809 VPWR VGND sg13g2_buf_1
X_6208_ net1861 net451 VPWR VGND sg13g2_buf_1
X_6139_ Tile_X0Y0_WW4END[6] net366 VPWR VGND sg13g2_buf_1
Xrebuffer9 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 net618 VPWR VGND sg13g2_buf_2
XFILLER_107_240 VPWR VGND sg13g2_fill_2
XFILLER_51_219 VPWR VGND sg13g2_decap_4
X_3840_ VPWR _1867_ _1866_ VGND sg13g2_inv_1
X_3771_ _1794_ VPWR _1801_ VGND _1799_ _1800_ sg13g2_o21ai_1
X_2722_ net50 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q
+ _0800_ VPWR VGND sg13g2_mux2_1
XFILLER_12_190 VPWR VGND sg13g2_fill_1
X_5510_ net1896 net1845 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_2653_ _0732_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q _0733_
+ _0734_ VPWR VGND sg13g2_a21o_1
X_5441_ Tile_X0Y1_UserCLK net557 _0055_ _0034_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[17\]
+ VPWR VGND sg13g2_dfrbp_1
X_2584_ _0668_ VPWR _0669_ VGND net1658 net1578 sg13g2_o21ai_1
Xoutput414 net414 Tile_X0Y1_EE4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput403 net403 Tile_X0Y1_E6BEG[7] VPWR VGND sg13g2_buf_1
Xoutput425 net425 Tile_X0Y1_FrameData_O[12] VPWR VGND sg13g2_buf_1
X_5372_ net1958 net1828 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_4323_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q net1577 net683
+ net1517 _1673_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2
+ VPWR VGND sg13g2_mux4_1
Xoutput469 net469 Tile_X0Y1_S2BEGb[3] VPWR VGND sg13g2_buf_1
Xoutput458 net458 Tile_X0Y1_S2BEG[0] VPWR VGND sg13g2_buf_1
Xoutput447 net447 Tile_X0Y1_FrameData_O[3] VPWR VGND sg13g2_buf_1
Xoutput436 net436 Tile_X0Y1_FrameData_O[22] VPWR VGND sg13g2_buf_1
X_4254_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q _1011_ _1483_
+ _0969_ net1576 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q _2213_
+ VPWR VGND sg13g2_mux4_1
X_3205_ _1259_ _0308_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q
+ _1260_ VPWR VGND sg13g2_mux2_1
X_4185_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q VPWR _2154_
+ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q _2153_ sg13g2_o21ai_1
X_3136_ _1193_ net1691 net1930 VPWR VGND sg13g2_nand2b_1
X_3067_ VGND VPWR _1122_ _1123_ _1127_ _1126_ sg13g2_a21oi_1
XFILLER_10_105 VPWR VGND sg13g2_fill_2
X_5708_ net1881 net1737 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_3969_ VGND VPWR _1975_ _1976_ _0034_ net1651 sg13g2_a21oi_2
X_5639_ net1919 net1769 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_88_38 VPWR VGND sg13g2_fill_2
Xfanout1606 net1607 net1606 VPWR VGND sg13g2_buf_1
Xfanout1617 net1617 net1618 VPWR VGND sg13g2_buf_16
Xfanout1628 _1148_ net1628 VPWR VGND sg13g2_buf_8
Xfanout1639 _0134_ net1639 VPWR VGND sg13g2_buf_1
XFILLER_37_20 VPWR VGND sg13g2_fill_1
XFILLER_58_352 VPWR VGND sg13g2_fill_1
XFILLER_64_355 VPWR VGND sg13g2_decap_4
X_5990_ Tile_X0Y0_EE4END[10] net217 VPWR VGND sg13g2_buf_1
X_4941_ net1936 net74 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q
+ _0484_ VPWR VGND sg13g2_mux2_1
X_4872_ _0418_ VPWR _0419_ VGND net1662 _0417_ sg13g2_o21ai_1
X_3823_ VGND VPWR net1678 net11 _1852_ _1851_ sg13g2_a21oi_1
X_3754_ VGND VPWR _1783_ _1784_ _0023_ net1643 sg13g2_a21oi_2
X_3685_ _1720_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q _1719_
+ VPWR VGND sg13g2_nand2_1
X_2705_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q _0780_
+ _0784_ _0783_ sg13g2_a21oi_1
Xoutput200 net200 Tile_X0Y0_E6BEG[5] VPWR VGND sg13g2_buf_1
X_5424_ Tile_X0Y1_UserCLK net574 _0038_ _0024_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[0\]
+ VPWR VGND sg13g2_dfrbp_1
X_2636_ _0718_ net1675 net137 VPWR VGND sg13g2_nand2b_1
Xoutput244 net244 Tile_X0Y0_FrameData_O[30] VPWR VGND sg13g2_buf_1
Xoutput222 net222 Tile_X0Y0_FrameData_O[10] VPWR VGND sg13g2_buf_1
Xoutput211 net211 Tile_X0Y0_EE4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput233 net233 Tile_X0Y0_FrameData_O[20] VPWR VGND sg13g2_buf_1
Xoutput255 net255 Tile_X0Y0_FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
Xoutput266 net266 Tile_X0Y0_FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
Xoutput277 net277 Tile_X0Y0_N2BEG[0] VPWR VGND sg13g2_buf_1
X_2567_ VGND VPWR net125 net1682 _0653_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q
+ sg13g2_a21oi_1
X_5355_ net1990 net1839 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_99_241 VPWR VGND sg13g2_fill_2
Xoutput299 net299 Tile_X0Y0_N4BEG[15] VPWR VGND sg13g2_buf_1
X_2498_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q net28 _0587_
+ VPWR VGND sg13g2_nor2_1
Xoutput288 net288 Tile_X0Y0_N2BEGb[3] VPWR VGND sg13g2_buf_1
X_4306_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q net38 net53
+ net1703 net1544 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2
+ VPWR VGND sg13g2_mux4_1
X_5286_ net1979 net1732 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_99_285 VPWR VGND sg13g2_decap_4
X_4237_ _2197_ VPWR _2198_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q
+ net681 sg13g2_o21ai_1
XFILLER_74_108 VPWR VGND sg13g2_fill_1
X_4168_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q _1482_
+ _2139_ _2138_ sg13g2_a21oi_1
XFILLER_55_322 VPWR VGND sg13g2_fill_2
X_3119_ _1175_ VPWR _1176_ VGND _1048_ _1051_ sg13g2_o21ai_1
X_4099_ VGND VPWR net1673 net1587 _2088_ _2087_ sg13g2_a21oi_1
XFILLER_82_196 VPWR VGND sg13g2_fill_1
XFILLER_99_26 VPWR VGND sg13g2_fill_1
XFILLER_0_26 VPWR VGND sg13g2_fill_1
XFILLER_61_314 VPWR VGND sg13g2_fill_1
XFILLER_73_196 VPWR VGND sg13g2_fill_2
XFILLER_9_46 VPWR VGND sg13g2_fill_1
X_3470_ _1518_ VPWR _1519_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q
+ _1516_ sg13g2_o21ai_1
X_5140_ net1945 net1789 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_5071_ net1997 net1810 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_96_244 VPWR VGND sg13g2_decap_4
Xfanout1970 Tile_X0Y0_FrameData[23] net1970 VPWR VGND sg13g2_buf_1
X_4022_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q
+ _2026_ _2022_ _2027_ _2025_ sg13g2_a221oi_1
Xfanout1981 net1982 net1981 VPWR VGND sg13g2_buf_1
Xfanout1992 Tile_X0Y0_FrameData[13] net1992 VPWR VGND sg13g2_buf_1
X_5973_ Tile_X0Y0_E6END[3] net196 VPWR VGND sg13g2_buf_1
X_4924_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q net1569
+ _0468_ _0467_ sg13g2_a21oi_1
X_4855_ _0403_ net1684 net1929 VPWR VGND sg13g2_nand2b_1
X_4786_ _0336_ VPWR _0337_ VGND net1692 net1631 sg13g2_o21ai_1
X_3806_ _1468_ VPWR _1835_ VGND _1832_ _1833_ sg13g2_o21ai_1
X_3737_ VGND VPWR _1765_ _1767_ _1764_ net1647 _1768_ _0020_ sg13g2_a221oi_1
XFILLER_118_143 VPWR VGND sg13g2_fill_1
XFILLER_109_25 VPWR VGND sg13g2_fill_1
X_3668_ _1703_ VPWR _1704_ VGND _0083_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q
+ sg13g2_o21ai_1
X_5407_ net1964 net1818 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_3599_ _1638_ VPWR _1639_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q
+ _0171_ sg13g2_o21ai_1
X_2619_ _0701_ net1642 Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[6\] VPWR VGND sg13g2_nand2b_1
X_5338_ net1951 net1840 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_5462__594 VPWR VGND net594 sg13g2_tiehi
X_5269_ net1947 net1740 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_18_44 VPWR VGND sg13g2_fill_1
XFILLER_55_141 VPWR VGND sg13g2_fill_1
XFILLER_11_222 VPWR VGND sg13g2_fill_1
XFILLER_119_0 VPWR VGND sg13g2_fill_1
XFILLER_109_165 VPWR VGND sg13g2_fill_2
XFILLER_46_130 VPWR VGND sg13g2_fill_1
XFILLER_61_100 VPWR VGND sg13g2_decap_4
X_2970_ _0933_ _1010_ _1030_ _1033_ VPWR VGND sg13g2_or3_1
X_4640_ _0197_ _0196_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q
+ VPWR VGND sg13g2_nand2b_1
X_6310_ Tile_X0Y1_W6END[7] net533 VPWR VGND sg13g2_buf_1
X_4571_ VPWR _0128_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q VGND
+ sg13g2_inv_1
X_3522_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q net1532 net1537
+ net1546 net1553 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q _1568_
+ VPWR VGND sg13g2_mux4_1
X_6241_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 net462 VPWR VGND sg13g2_buf_2
X_3453_ _1502_ net1638 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X
+ VPWR VGND sg13g2_nand2_1
X_5446__578 VPWR VGND net578 sg13g2_tiehi
X_6172_ net106 net393 VPWR VGND sg13g2_buf_1
XFILLER_103_319 VPWR VGND sg13g2_fill_1
X_5123_ net1972 net1785 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_34_0 VPWR VGND sg13g2_fill_1
X_3384_ _1436_ net682 _1435_ VPWR VGND sg13g2_nand2_2
X_5054_ net1961 net1809 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_4005_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q VPWR _2010_ VGND
+ _2001_ _2003_ sg13g2_o21ai_1
XFILLER_1_80 VPWR VGND sg13g2_fill_1
X_5956_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 net177 VPWR VGND sg13g2_buf_1
X_4907_ _0453_ net1677 net1930 VPWR VGND sg13g2_nand2b_1
X_5887_ net1859 net1812 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_4838_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q VPWR _0386_ VGND
+ net1684 _0175_ sg13g2_o21ai_1
X_4769_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q _0317_
+ _0320_ _0067_ sg13g2_a21oi_1
XFILLER_121_105 VPWR VGND sg13g2_fill_2
XFILLER_106_168 VPWR VGND sg13g2_decap_8
XFILLER_29_54 VPWR VGND sg13g2_decap_4
XFILLER_28_185 VPWR VGND sg13g2_fill_2
XFILLER_31_306 VPWR VGND sg13g2_fill_2
XFILLER_61_52 VPWR VGND sg13g2_decap_8
XFILLER_3_262 VPWR VGND sg13g2_fill_2
XFILLER_98_317 VPWR VGND sg13g2_fill_1
XFILLER_19_163 VPWR VGND sg13g2_fill_1
XFILLER_81_239 VPWR VGND sg13g2_fill_1
X_5810_ net1893 net1836 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_34_144 VPWR VGND sg13g2_fill_1
XFILLER_22_339 VPWR VGND sg13g2_fill_2
X_5741_ net1882 net1727 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_2953_ VGND VPWR _0062_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q
+ _1017_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q sg13g2_a21oi_1
X_2884_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q net1565 net1572
+ net1579 net1616 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q _0953_
+ VPWR VGND sg13g2_mux4_1
Xrebuffer109 _0416_ net718 VPWR VGND sg13g2_dlygate4sd1_1
X_5672_ net1871 net1752 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_4623_ net1535 _0180_ VPWR VGND sg13g2_inv_4
X_4554_ VPWR _0111_ net77 VGND sg13g2_inv_1
X_3505_ _1551_ VPWR _1552_ VGND _0416_ net1670 sg13g2_o21ai_1
X_4485_ net1512 _1886_ _0042_ VPWR VGND sg13g2_nor2_1
X_6224_ net1889 net437 VPWR VGND sg13g2_buf_1
X_3436_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q VPWR _1487_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q _1486_ sg13g2_o21ai_1
X_6155_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 net376 VPWR VGND sg13g2_buf_1
X_3367_ _1413_ _1418_ _1419_ VPWR VGND sg13g2_nor2_1
X_6086_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 net298 VPWR VGND sg13g2_buf_1
XFILLER_66_19 VPWR VGND sg13g2_fill_2
X_5106_ net1941 net1796 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_97_383 VPWR VGND sg13g2_fill_2
X_3298_ _1346_ _1349_ _1350_ VPWR VGND sg13g2_xor2_1
X_5037_ net1994 net1849 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_122_69 VPWR VGND sg13g2_fill_1
XFILLER_72_239 VPWR VGND sg13g2_fill_1
XFILLER_31_33 VPWR VGND sg13g2_fill_1
XFILLER_110_4 VPWR VGND sg13g2_fill_2
XFILLER_31_99 VPWR VGND sg13g2_fill_1
Xinput100 Tile_X0Y1_E2MID[1] net100 VPWR VGND sg13g2_buf_1
Xinput111 Tile_X0Y1_N1END[0] net111 VPWR VGND sg13g2_buf_1
Xinput133 Tile_X0Y1_N4END[2] net133 VPWR VGND sg13g2_buf_1
Xinput144 Tile_X0Y1_NN4END[5] net144 VPWR VGND sg13g2_buf_1
Xinput122 Tile_X0Y1_N2END[7] net122 VPWR VGND sg13g2_buf_1
Xinput155 Tile_X0Y1_W2END[4] net155 VPWR VGND sg13g2_buf_1
Xinput166 Tile_X0Y1_W2MID[7] net166 VPWR VGND sg13g2_buf_1
XFILLER_48_269 VPWR VGND sg13g2_fill_1
XFILLER_56_41 VPWR VGND sg13g2_decap_4
XFILLER_72_84 VPWR VGND sg13g2_fill_1
XFILLER_12_383 VPWR VGND sg13g2_fill_2
X_4270_ _2221_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 VGND _2227_
+ _2225_ sg13g2_o21ai_1
X_3221_ VGND VPWR _0129_ _1274_ _1275_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q
+ sg13g2_a21oi_1
XFILLER_98_158 VPWR VGND sg13g2_decap_4
X_3152_ VGND VPWR _1207_ _1208_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q
+ _1204_ sg13g2_a21oi_2
XFILLER_79_383 VPWR VGND sg13g2_fill_2
X_3083_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q _1140_
+ _1142_ _1141_ sg13g2_a21oi_1
X_3985_ VGND VPWR _1987_ _1989_ _1990_ _1986_ sg13g2_a21oi_1
X_5724_ net1916 net1737 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_2936_ net1661 net1710 net122 net1925 net98 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q
+ _1002_ VPWR VGND sg13g2_mux4_1
X_2867_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q net1599 net1612
+ net1605 net1625 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q _0937_
+ VPWR VGND sg13g2_mux4_1
X_5655_ net1905 net1761 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_4606_ VPWR _0163_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q
+ VGND sg13g2_inv_1
XFILLER_7_90 VPWR VGND sg13g2_fill_2
X_5586_ net1893 net1783 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_2798_ _0871_ VPWR _0872_ VGND net1688 net1621 sg13g2_o21ai_1
X_4537_ VPWR _0094_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q VGND
+ sg13g2_inv_1
XFILLER_89_103 VPWR VGND sg13g2_fill_2
X_4468_ _2378_ VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 VGND _2380_
+ _2382_ sg13g2_o21ai_1
X_6207_ net1863 net450 VPWR VGND sg13g2_buf_1
X_3419_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5
+ net43 net17 net78 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q _1471_
+ VPWR VGND sg13g2_mux4_1
XFILLER_89_169 VPWR VGND sg13g2_fill_1
X_4399_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q _1058_
+ _2323_ _2322_ sg13g2_a21oi_1
X_6138_ Tile_X0Y0_WW4END[5] net365 VPWR VGND sg13g2_buf_1
XFILLER_45_206 VPWR VGND sg13g2_fill_2
X_6069_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 net290 VPWR VGND sg13g2_buf_1
XFILLER_93_28 VPWR VGND sg13g2_fill_1
XFILLER_26_22 VPWR VGND sg13g2_fill_1
XFILLER_26_44 VPWR VGND sg13g2_fill_1
XFILLER_9_107 VPWR VGND sg13g2_fill_1
XFILLER_5_346 VPWR VGND sg13g2_fill_2
XFILLER_107_285 VPWR VGND sg13g2_fill_1
XFILLER_76_364 VPWR VGND sg13g2_fill_1
XFILLER_44_250 VPWR VGND sg13g2_decap_4
XFILLER_44_294 VPWR VGND sg13g2_fill_2
X_3770_ _0348_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q
+ _1800_ VPWR VGND sg13g2_a21o_1
X_2721_ _0792_ VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q
+ _0799_ sg13g2_o21ai_1
X_5440_ Tile_X0Y1_UserCLK net558 _0054_ _0032_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[16\]
+ VPWR VGND sg13g2_dfrbp_1
X_2652_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q VPWR _0733_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q _0731_ sg13g2_o21ai_1
Xoutput415 net415 Tile_X0Y1_EE4BEG[3] VPWR VGND sg13g2_buf_1
X_2583_ _0668_ net1658 net1617 VPWR VGND sg13g2_nand2b_1
Xoutput404 net404 Tile_X0Y1_E6BEG[8] VPWR VGND sg13g2_buf_1
Xoutput426 net426 Tile_X0Y1_FrameData_O[13] VPWR VGND sg13g2_buf_1
X_5371_ net1954 net1829 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput448 net448 Tile_X0Y1_FrameData_O[4] VPWR VGND sg13g2_buf_1
X_4322_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q net1573 net689
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 _0362_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 VPWR VGND sg13g2_mux4_1
Xoutput459 net459 Tile_X0Y1_S2BEG[1] VPWR VGND sg13g2_buf_1
Xoutput437 net437 Tile_X0Y1_FrameData_O[23] VPWR VGND sg13g2_buf_1
X_4253_ _2211_ VPWR _2212_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q
+ _2208_ sg13g2_o21ai_1
X_3204_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q net117 net93
+ net1935 net171 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q _1259_
+ VPWR VGND sg13g2_mux4_1
X_4184_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q net1588 net1523
+ net1519 net1540 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q _2153_
+ VPWR VGND sg13g2_mux4_1
X_3135_ _1191_ VPWR _1192_ VGND _0090_ net1691 sg13g2_o21ai_1
X_3066_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q VPWR _1126_ VGND
+ _1124_ _1125_ sg13g2_o21ai_1
XFILLER_103_27 VPWR VGND sg13g2_fill_1
X_3968_ net1651 _1974_ _1975_ VPWR VGND sg13g2_nor2_2
X_2919_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q _0985_
+ _0986_ _0102_ sg13g2_a21oi_1
X_5707_ net1879 net1735 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_3899_ VGND VPWR net11 net2005 _1913_ _1912_ sg13g2_a21oi_1
X_5638_ net1896 net1769 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_5569_ net1862 net1790 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
Xfanout1618 net1618 net1620 VPWR VGND sg13g2_buf_16
Xfanout1629 net1631 net1629 VPWR VGND sg13g2_buf_1
Xfanout1607 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 net1607 VPWR VGND
+ sg13g2_buf_8
XFILLER_33_209 VPWR VGND sg13g2_decap_4
XFILLER_110_203 VPWR VGND sg13g2_fill_2
XFILLER_76_161 VPWR VGND sg13g2_fill_1
XFILLER_17_250 VPWR VGND sg13g2_fill_2
X_4940_ _0482_ VPWR _0483_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q
+ net612 sg13g2_o21ai_1
XFILLER_32_220 VPWR VGND sg13g2_fill_1
X_4871_ VGND VPWR net1662 _0077_ _0418_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q
+ sg13g2_a21oi_1
X_3822_ net1678 net2001 _1851_ VPWR VGND sg13g2_nor2b_1
X_3753_ net1643 Tile_X0Y1_DSP_bot.C1 _1783_ VPWR VGND sg13g2_nor2_2
X_3684_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6
+ _1719_ _1718_ sg13g2_a21oi_1
X_2704_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q VPWR _0783_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q _0782_ sg13g2_o21ai_1
XFILLER_64_0 VPWR VGND sg13g2_fill_2
Xoutput201 net201 Tile_X0Y0_E6BEG[6] VPWR VGND sg13g2_buf_1
X_5423_ net1997 net1819 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_2635_ _0716_ VPWR _0717_ VGND net1 net1674 sg13g2_o21ai_1
Xoutput223 net223 Tile_X0Y0_FrameData_O[11] VPWR VGND sg13g2_buf_1
Xoutput234 net234 Tile_X0Y0_FrameData_O[21] VPWR VGND sg13g2_buf_1
X_5354_ net1987 net1839 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput212 net212 Tile_X0Y0_EE4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput267 net267 Tile_X0Y0_FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
Xoutput245 net245 Tile_X0Y0_FrameData_O[31] VPWR VGND sg13g2_buf_1
Xoutput256 net256 Tile_X0Y0_FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
X_4305_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q net1923 net41
+ net52 net1535 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1
+ VPWR VGND sg13g2_mux4_1
X_2566_ VGND VPWR _0651_ _0652_ _0650_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q
+ sg13g2_a21oi_2
Xoutput289 net289 Tile_X0Y0_N2BEGb[4] VPWR VGND sg13g2_buf_8
X_2497_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q _0585_ _0586_
+ VPWR VGND sg13g2_nor2b_1
Xoutput278 net278 Tile_X0Y0_N2BEG[1] VPWR VGND sg13g2_buf_1
X_5285_ net1975 net1731 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_4236_ VGND VPWR _0070_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q
+ _2197_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q sg13g2_a21oi_1
X_4167_ _0163_ VPWR _2138_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q
+ net1519 sg13g2_o21ai_1
XFILLER_67_150 VPWR VGND sg13g2_fill_1
XFILLER_67_194 VPWR VGND sg13g2_fill_2
X_3118_ _1174_ _1173_ _1175_ VPWR VGND sg13g2_and2_1
X_4098_ net1672 net1590 _2087_ VPWR VGND sg13g2_nor2_1
X_3049_ _1109_ _0930_ _1107_ VPWR VGND sg13g2_xnor2_1
XFILLER_48_31 VPWR VGND sg13g2_fill_2
XFILLER_65_109 VPWR VGND sg13g2_fill_2
XFILLER_61_348 VPWR VGND sg13g2_fill_2
XFILLER_96_212 VPWR VGND sg13g2_decap_4
X_5070_ net1995 net1810 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_4021_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q net26 net28 net54
+ net83 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q _2026_ VPWR VGND
+ sg13g2_mux4_1
Xfanout1960 Tile_X0Y0_FrameData[28] net1960 VPWR VGND sg13g2_buf_1
Xfanout1982 Tile_X0Y0_FrameData[18] net1982 VPWR VGND sg13g2_buf_1
Xfanout1971 Tile_X0Y0_FrameData[22] net1971 VPWR VGND sg13g2_buf_1
Xfanout1993 net1994 net1993 VPWR VGND sg13g2_buf_1
X_5972_ Tile_X0Y0_E6END[2] net193 VPWR VGND sg13g2_buf_1
X_4923_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q net1563 _0467_
+ VPWR VGND sg13g2_nor2_1
X_4854_ _0401_ VPWR _0402_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q
+ _0400_ sg13g2_o21ai_1
XFILLER_20_201 VPWR VGND sg13g2_fill_2
X_4785_ _0336_ net1692 net1590 VPWR VGND sg13g2_nand2_1
X_3805_ _1467_ _0235_ _1834_ VPWR VGND sg13g2_xor2_1
X_3736_ _1767_ net685 _1435_ VPWR VGND sg13g2_xnor2_1
X_3667_ VGND VPWR net104 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q
+ _1703_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q sg13g2_a21oi_1
X_5406_ net1961 net1820 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_3598_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q net1566
+ _1638_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q sg13g2_a21oi_1
X_2618_ _0527_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X
+ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q _0700_ sg13g2_o21ai_1
X_2549_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q net27 net35 net29
+ net1933 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q _0635_ VPWR
+ VGND sg13g2_mux4_1
X_5337_ net1999 net1721 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_87_212 VPWR VGND sg13g2_fill_2
X_5268_ net1945 net1740 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_4219_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q _2182_
+ _2184_ _2183_ sg13g2_a21oi_1
X_5199_ net1997 net1764 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_55_175 VPWR VGND sg13g2_fill_1
XFILLER_70_134 VPWR VGND sg13g2_fill_1
XFILLER_11_278 VPWR VGND sg13g2_fill_1
XFILLER_105_372 VPWR VGND sg13g2_fill_1
XFILLER_93_226 VPWR VGND sg13g2_fill_1
XFILLER_93_259 VPWR VGND sg13g2_fill_1
X_4570_ VPWR _0127_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q VGND
+ sg13g2_inv_1
X_3521_ VGND VPWR _0143_ _1566_ _1567_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q
+ sg13g2_a21oi_1
X_6240_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 net461 VPWR VGND sg13g2_buf_2
X_3452_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q _1500_ _1499_
+ _1483_ _1501_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X
+ VPWR VGND sg13g2_mux4_1
XFILLER_115_169 VPWR VGND sg13g2_fill_2
X_3383_ _1214_ net1548 _1427_ _1435_ VPWR VGND sg13g2_nor3_2
X_6171_ net105 net392 VPWR VGND sg13g2_buf_1
X_5122_ net1970 net1786 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_0 VPWR VGND sg13g2_fill_1
X_5053_ net1960 net1807 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_84_226 VPWR VGND sg13g2_decap_4
Xfanout1790 net1791 net1790 VPWR VGND sg13g2_buf_1
XFILLER_84_248 VPWR VGND sg13g2_fill_2
X_4004_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q _2005_
+ _2009_ _2008_ sg13g2_a21oi_1
XFILLER_25_359 VPWR VGND sg13g2_fill_2
X_5955_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 net176 VPWR VGND sg13g2_buf_8
X_4906_ VGND VPWR net35 net1677 _0452_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q
+ sg13g2_a21oi_1
X_5886_ net1856 net1812 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_4837_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q net137 net6 net72
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q
+ _0385_ VPWR VGND sg13g2_mux4_1
X_4768_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q net50
+ _0319_ _0318_ sg13g2_a21oi_1
X_3719_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q net120 net96
+ net59 net156 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q _1751_
+ VPWR VGND sg13g2_mux4_1
X_4699_ net85 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q
+ _0252_ VPWR VGND sg13g2_mux2_1
XFILLER_121_128 VPWR VGND sg13g2_fill_2
XFILLER_29_77 VPWR VGND sg13g2_fill_2
XFILLER_29_88 VPWR VGND sg13g2_fill_2
XFILLER_90_218 VPWR VGND sg13g2_decap_4
XFILLER_43_178 VPWR VGND sg13g2_decap_4
XFILLER_19_120 VPWR VGND sg13g2_fill_1
XFILLER_66_237 VPWR VGND sg13g2_fill_1
XFILLER_81_207 VPWR VGND sg13g2_fill_2
X_5740_ net1880 net1726 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_2952_ _1016_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q _1015_
+ VPWR VGND sg13g2_nand2_1
X_5671_ net1920 net1762 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_2883_ _0952_ _0941_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 VPWR VGND
+ sg13g2_nor2_2
X_4622_ VPWR _0179_ net1539 VGND sg13g2_inv_1
X_4553_ VPWR _0110_ net16 VGND sg13g2_inv_1
X_4484_ net1512 _1888_ _0041_ VPWR VGND sg13g2_nor2b_1
X_3504_ _1551_ net1670 _0682_ VPWR VGND sg13g2_nand2_1
X_3435_ net1635 net1586 net1687 _1486_ VPWR VGND sg13g2_mux2_1
X_6223_ net1891 net436 VPWR VGND sg13g2_buf_1
X_6154_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 net375 VPWR VGND sg13g2_buf_1
X_3366_ _1418_ _1416_ _1417_ VPWR VGND sg13g2_nand2_1
X_3297_ _1349_ _1299_ _1347_ VPWR VGND sg13g2_xnor2_1
X_5105_ net1939 net1795 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_6085_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 net297 VPWR VGND sg13g2_buf_1
X_5036_ net1992 net1849 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_15_24 VPWR VGND sg13g2_fill_1
X_5869_ net1882 net1813 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput101 Tile_X0Y1_E2MID[2] net101 VPWR VGND sg13g2_buf_1
Xinput123 Tile_X0Y1_N2MID[0] net123 VPWR VGND sg13g2_buf_1
Xinput145 Tile_X0Y1_NN4END[6] net145 VPWR VGND sg13g2_buf_1
Xinput134 Tile_X0Y1_N4END[3] net134 VPWR VGND sg13g2_buf_1
Xinput112 Tile_X0Y1_N1END[1] net112 VPWR VGND sg13g2_buf_1
XFILLER_48_215 VPWR VGND sg13g2_fill_2
Xinput167 Tile_X0Y1_W6END[0] net167 VPWR VGND sg13g2_buf_1
Xinput156 Tile_X0Y1_W2END[5] net156 VPWR VGND sg13g2_buf_1
XFILLER_48_237 VPWR VGND sg13g2_fill_1
XFILLER_56_97 VPWR VGND sg13g2_fill_2
XFILLER_112_70 VPWR VGND sg13g2_fill_1
XFILLER_16_189 VPWR VGND sg13g2_fill_1
X_3220_ net125 net101 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q
+ _1274_ VPWR VGND sg13g2_mux2_1
X_3151_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q VPWR _1207_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q _1206_ sg13g2_o21ai_1
XFILLER_94_310 VPWR VGND sg13g2_fill_2
X_3082_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q VPWR _1141_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q _1139_ sg13g2_o21ai_1
X_3984_ VGND VPWR _1977_ _1989_ _1978_ _1953_ sg13g2_a21oi_2
XFILLER_94_0 VPWR VGND sg13g2_fill_2
X_5723_ net1912 net1735 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_2935_ _1000_ _0997_ _1001_ VPWR VGND sg13g2_nor2b_1
X_5654_ net1903 net1761 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_2866_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q _0385_
+ _0936_ _0935_ sg13g2_a21oi_1
X_4605_ VPWR _0162_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q
+ VGND sg13g2_inv_1
XFILLER_108_209 VPWR VGND sg13g2_fill_2
X_5585_ net1891 net1783 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_2797_ _0871_ net1688 net1629 VPWR VGND sg13g2_nand2b_1
X_4536_ VPWR _0093_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q VGND
+ sg13g2_inv_1
XFILLER_117_48 VPWR VGND sg13g2_fill_1
X_4467_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q VPWR _2382_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q _2381_ sg13g2_o21ai_1
X_4398_ _0168_ VPWR _2322_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q
+ net1572 sg13g2_o21ai_1
X_6206_ net1865 net449 VPWR VGND sg13g2_buf_1
X_3418_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4
+ net77 net42 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q
+ _1470_ VPWR VGND sg13g2_mux4_1
X_3349_ _1400_ _1399_ _1401_ VPWR VGND sg13g2_nor2_2
X_6137_ Tile_X0Y0_WW4END[4] net358 VPWR VGND sg13g2_buf_1
XFILLER_97_170 VPWR VGND sg13g2_decap_8
X_6068_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 net289 VPWR VGND sg13g2_buf_8
XFILLER_85_354 VPWR VGND sg13g2_fill_1
X_5019_ net1953 net1853 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_91_379 VPWR VGND sg13g2_fill_2
X_2720_ _0798_ VPWR _0799_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q
+ _0793_ sg13g2_o21ai_1
X_2651_ net1582 net1619 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ _0732_ VPWR VGND sg13g2_mux2_1
Xoutput416 net416 Tile_X0Y1_EE4BEG[4] VPWR VGND sg13g2_buf_1
X_2582_ VGND VPWR net1658 net1569 _0667_ _0666_ sg13g2_a21oi_1
Xoutput405 net405 Tile_X0Y1_E6BEG[9] VPWR VGND sg13g2_buf_1
X_5370_ net1952 net1828 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_4321_ _2258_ VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 VGND _2253_
+ _2254_ sg13g2_o21ai_1
Xoutput449 net449 Tile_X0Y1_FrameData_O[5] VPWR VGND sg13g2_buf_1
Xoutput427 net427 Tile_X0Y1_FrameData_O[14] VPWR VGND sg13g2_buf_1
Xoutput438 net438 Tile_X0Y1_FrameData_O[24] VPWR VGND sg13g2_buf_1
X_4252_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q _2210_
+ _2211_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q sg13g2_a21oi_1
X_3203_ _1249_ VPWR _1258_ VGND _1246_ _1251_ sg13g2_o21ai_1
X_4183_ _2151_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q _2152_
+ VPWR VGND sg13g2_nor2b_1
X_3134_ VGND VPWR net37 net1691 _1191_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q
+ sg13g2_a21oi_1
XFILLER_27_207 VPWR VGND sg13g2_fill_1
X_3065_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q VPWR _1125_ VGND
+ net148 net1668 sg13g2_o21ai_1
XFILLER_50_276 VPWR VGND sg13g2_decap_8
X_3967_ VGND VPWR _1973_ _1974_ _0035_ net1645 sg13g2_a21oi_2
X_2918_ _0984_ VPWR _0985_ VGND net69 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q
+ sg13g2_o21ai_1
X_5706_ net1877 net1735 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_3898_ net2005 net2001 _1912_ VPWR VGND sg13g2_nor2b_1
X_2849_ net1667 net52 _0921_ VPWR VGND sg13g2_nor2b_1
X_5637_ net1874 net1769 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_5568_ net1860 net1790 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_4519_ VPWR _0076_ net82 VGND sg13g2_inv_1
XFILLER_104_201 VPWR VGND sg13g2_decap_8
X_5499_ net1913 net1848 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_5_8 VPWR VGND sg13g2_fill_2
Xfanout1619 net1620 net1619 VPWR VGND sg13g2_buf_1
Xfanout1608 _0768_ net1608 VPWR VGND sg13g2_buf_8
XFILLER_104_278 VPWR VGND sg13g2_decap_8
XFILLER_41_210 VPWR VGND sg13g2_fill_2
XFILLER_5_188 VPWR VGND sg13g2_fill_1
XFILLER_110_237 VPWR VGND sg13g2_decap_4
XFILLER_110_226 VPWR VGND sg13g2_fill_2
XFILLER_68_129 VPWR VGND sg13g2_fill_2
XFILLER_91_187 VPWR VGND sg13g2_fill_1
X_4870_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q net1629 net647
+ _0411_ _0385_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q _0417_
+ VPWR VGND sg13g2_mux4_1
X_3821_ _1849_ VPWR _1850_ VGND net1678 net622 sg13g2_o21ai_1
X_3752_ _1782_ VPWR Tile_X0Y1_DSP_bot.C1 VGND _1771_ _1773_ sg13g2_o21ai_1
X_3683_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q net161 _1718_
+ VPWR VGND sg13g2_nor2b_1
X_2703_ _0781_ VPWR _0782_ VGND net124 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q
+ sg13g2_o21ai_1
X_5422_ net1995 net1819 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_2634_ _0716_ net1674 net6 VPWR VGND sg13g2_nand2b_1
Xoutput224 net224 Tile_X0Y0_FrameData_O[12] VPWR VGND sg13g2_buf_1
Xoutput202 net202 Tile_X0Y0_E6BEG[7] VPWR VGND sg13g2_buf_1
X_5353_ net1986 net1841 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_2565_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q VPWR _0651_ VGND
+ _0649_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q sg13g2_o21ai_1
Xoutput235 net235 Tile_X0Y0_FrameData_O[22] VPWR VGND sg13g2_buf_1
Xoutput213 net213 Tile_X0Y0_EE4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput268 net268 Tile_X0Y0_FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
Xoutput246 net246 Tile_X0Y0_FrameData_O[3] VPWR VGND sg13g2_buf_1
Xoutput257 net257 Tile_X0Y0_FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
X_4304_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q net1921 net51
+ net1935 net1529 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0
+ VPWR VGND sg13g2_mux4_1
X_2496_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q net1516 net2003
+ net129 net10 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q _0585_
+ VPWR VGND sg13g2_mux4_1
Xoutput279 net279 Tile_X0Y0_N2BEG[2] VPWR VGND sg13g2_buf_1
X_5284_ net1973 net1731 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_99_265 VPWR VGND sg13g2_fill_2
X_4235_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 _2196_ VGND sg13g2_inv_1
X_4166_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q _2136_
+ _2137_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q sg13g2_a21oi_1
X_3117_ _1044_ _1046_ _1172_ _1174_ VPWR VGND sg13g2_or3_1
X_4097_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q _2085_ _2086_
+ VPWR VGND sg13g2_nor2_1
X_3048_ _1108_ _0807_ net1575 VPWR VGND sg13g2_nand2_1
XFILLER_70_327 VPWR VGND sg13g2_fill_2
XFILLER_23_298 VPWR VGND sg13g2_fill_2
X_4999_ _0539_ VPWR _0540_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q
+ _0538_ sg13g2_o21ai_1
XFILLER_58_162 VPWR VGND sg13g2_fill_2
XFILLER_104_71 VPWR VGND sg13g2_fill_1
XFILLER_61_327 VPWR VGND sg13g2_fill_1
XFILLER_120_92 VPWR VGND sg13g2_fill_2
XFILLER_50_7 VPWR VGND sg13g2_fill_2
X_4020_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q _2024_ _2025_
+ VPWR VGND sg13g2_nor2_1
Xfanout1961 net1962 net1961 VPWR VGND sg13g2_buf_1
Xfanout1950 Tile_X0Y0_FrameData[3] net1950 VPWR VGND sg13g2_buf_1
Xfanout1972 Tile_X0Y0_FrameData[22] net1972 VPWR VGND sg13g2_buf_1
Xfanout1983 net1984 net1983 VPWR VGND sg13g2_buf_1
Xfanout1994 Tile_X0Y0_FrameData[12] net1994 VPWR VGND sg13g2_buf_1
XFILLER_52_305 VPWR VGND sg13g2_fill_2
X_5971_ net19 net192 VPWR VGND sg13g2_buf_1
X_4922_ _0466_ _0465_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q
+ VPWR VGND sg13g2_nand2b_1
X_4853_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q _0399_
+ _0401_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q sg13g2_a21oi_1
XFILLER_20_246 VPWR VGND sg13g2_fill_1
X_4784_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q
+ _0334_ _0330_ _0335_ _0332_ sg13g2_a221oi_1
X_3804_ _0235_ _1467_ _1833_ VPWR VGND sg13g2_and2_1
X_3735_ _1766_ _1764_ _1765_ _0020_ net1647 VPWR VGND sg13g2_a22oi_1
X_5405_ net1960 net1820 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_3666_ _1701_ VPWR _1702_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q
+ _0594_ sg13g2_o21ai_1
X_3597_ VGND VPWR _0144_ _1636_ _1637_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q
+ sg13g2_a21oi_1
X_2617_ _0630_ _0698_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q
+ _0700_ VPWR VGND sg13g2_mux2_1
X_2548_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q _0633_
+ _0634_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q sg13g2_a21oi_1
X_5336_ net1977 net1721 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_5267_ net1943 net1740 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_2479_ _0569_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q _0568_
+ VPWR VGND sg13g2_nand2b_1
X_4218_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q VPWR _2183_
+ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q _2181_ sg13g2_o21ai_1
X_5198_ net1995 net1764 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_4149_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q net1539 _1470_
+ net623 _1020_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q _2123_
+ VPWR VGND sg13g2_mux4_1
XFILLER_55_132 VPWR VGND sg13g2_decap_8
XFILLER_70_102 VPWR VGND sg13g2_decap_4
XFILLER_70_168 VPWR VGND sg13g2_decap_8
XFILLER_109_101 VPWR VGND sg13g2_fill_1
XFILLER_109_167 VPWR VGND sg13g2_fill_1
XFILLER_59_86 VPWR VGND sg13g2_decap_4
XFILLER_46_187 VPWR VGND sg13g2_fill_2
X_3520_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q net111 net87
+ net115 net91 net1671 _1566_ VPWR VGND sg13g2_mux4_1
X_3451_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q net145 net48
+ net6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q
+ _1501_ VPWR VGND sg13g2_mux4_1
X_6170_ net104 net391 VPWR VGND sg13g2_buf_1
X_3382_ _1434_ _1213_ net1568 VPWR VGND sg13g2_nand2_2
XFILLER_69_224 VPWR VGND sg13g2_fill_1
X_5121_ net1967 net1787 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_111_365 VPWR VGND sg13g2_fill_2
X_5052_ net1958 net1807 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
Xfanout1791 net1792 net1791 VPWR VGND sg13g2_buf_1
Xfanout1780 net1784 net1780 VPWR VGND sg13g2_buf_1
X_4003_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q VPWR _2008_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q _2007_ sg13g2_o21ai_1
X_5954_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 net175 VPWR VGND sg13g2_buf_1
X_4905_ _0451_ net27 net1677 VPWR VGND sg13g2_nand2b_1
X_5885_ net1918 net1816 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_33_382 VPWR VGND sg13g2_fill_2
X_4836_ VPWR _0384_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 VGND sg13g2_inv_1
X_4767_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q net42 _0318_
+ VPWR VGND sg13g2_nor2b_1
X_3718_ _1750_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q _0362_
+ VPWR VGND sg13g2_nand2_1
X_4698_ _0251_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 VGND _0237_
+ _0243_ sg13g2_o21ai_1
XFILLER_106_115 VPWR VGND sg13g2_fill_2
X_3649_ _1685_ VPWR _1686_ VGND _0060_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q
+ sg13g2_o21ai_1
XFILLER_106_159 VPWR VGND sg13g2_fill_1
X_5319_ net1982 net1722 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_6299_ net161 net520 VPWR VGND sg13g2_buf_1
XFILLER_28_121 VPWR VGND sg13g2_decap_8
XFILLER_28_187 VPWR VGND sg13g2_fill_1
XFILLER_43_157 VPWR VGND sg13g2_decap_8
XFILLER_61_21 VPWR VGND sg13g2_fill_2
XFILLER_112_129 VPWR VGND sg13g2_decap_8
XFILLER_3_264 VPWR VGND sg13g2_fill_1
XFILLER_105_181 VPWR VGND sg13g2_fill_1
XFILLER_66_216 VPWR VGND sg13g2_fill_1
XFILLER_59_290 VPWR VGND sg13g2_fill_2
X_2951_ net72 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q
+ _1015_ VPWR VGND sg13g2_mux2_1
X_5670_ net1897 net1762 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_4621_ VPWR _0178_ net1616 VGND sg13g2_inv_1
XFILLER_30_341 VPWR VGND sg13g2_fill_2
X_5452__584 VPWR VGND net584 sg13g2_tiehi
X_2882_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q _0946_ _0951_
+ _0952_ VPWR VGND sg13g2_nor3_2
X_4552_ VPWR _0109_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q VGND
+ sg13g2_inv_1
X_4483_ net1512 _1883_ _0040_ VPWR VGND sg13g2_nor2b_1
X_3503_ _1543_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q _1550_
+ VPWR VGND sg13g2_nor2b_1
X_3434_ VGND VPWR net1687 net1539 _1485_ _1484_ sg13g2_a21oi_1
X_6222_ net1893 net435 VPWR VGND sg13g2_buf_1
X_6153_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 net374 VPWR VGND sg13g2_buf_1
X_3365_ net1568 _0807_ _1415_ _1417_ VPWR VGND sg13g2_a21o_1
X_3296_ _1348_ _1299_ _1347_ VPWR VGND sg13g2_nand2_1
X_5104_ net1937 net1795 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_6084_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 net296 VPWR VGND sg13g2_buf_1
X_5035_ net1989 net1852 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_5868_ net1880 net1813 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_5799_ net1919 net1716 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_4819_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q _0367_ _0365_
+ _0368_ VPWR VGND sg13g2_nand3_1
XFILLER_110_6 VPWR VGND sg13g2_fill_1
Xinput102 Tile_X0Y1_E2MID[3] net102 VPWR VGND sg13g2_buf_1
Xinput135 Tile_X0Y1_N4END[4] net135 VPWR VGND sg13g2_buf_1
Xinput124 Tile_X0Y1_N2MID[1] net124 VPWR VGND sg13g2_buf_1
Xinput113 Tile_X0Y1_N1END[2] net113 VPWR VGND sg13g2_buf_1
XFILLER_48_205 VPWR VGND sg13g2_decap_4
XFILLER_102_140 VPWR VGND sg13g2_fill_2
Xinput157 Tile_X0Y1_W2END[6] net157 VPWR VGND sg13g2_buf_1
Xinput146 Tile_X0Y1_NN4END[7] net146 VPWR VGND sg13g2_buf_1
Xinput168 Tile_X0Y1_W6END[1] net168 VPWR VGND sg13g2_buf_1
XFILLER_112_93 VPWR VGND sg13g2_fill_2
XFILLER_112_82 VPWR VGND sg13g2_decap_8
XFILLER_31_127 VPWR VGND sg13g2_fill_2
XFILLER_71_296 VPWR VGND sg13g2_fill_2
X_3150_ _1205_ VPWR _1206_ VGND net1706 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q
+ sg13g2_o21ai_1
X_3081_ net154 net168 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q
+ _1140_ VPWR VGND sg13g2_mux2_1
XFILLER_62_274 VPWR VGND sg13g2_decap_4
X_5722_ net1910 net1735 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_3983_ _1988_ _1987_ _1986_ VPWR VGND sg13g2_nand2b_1
X_2934_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q VPWR _1000_ VGND
+ _0998_ _0999_ sg13g2_o21ai_1
X_5653_ net1900 net1760 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_2865_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q _0934_ _0935_
+ VPWR VGND sg13g2_nor2b_1
X_5584_ net1888 net1783 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_4604_ VPWR _0161_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q
+ VGND sg13g2_inv_1
X_4535_ VPWR _0092_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q VGND
+ sg13g2_inv_1
X_2796_ VPWR _0870_ _0869_ VGND sg13g2_inv_1
XFILLER_117_16 VPWR VGND sg13g2_fill_2
X_4466_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q net1573 net1578
+ net1615 net1617 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q _2381_
+ VPWR VGND sg13g2_mux4_1
X_4397_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q _2320_ _2321_
+ VPWR VGND sg13g2_nor2_1
X_6205_ net1867 net448 VPWR VGND sg13g2_buf_1
X_3417_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q net128 net55
+ net9 net70 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q _1469_ VPWR
+ VGND sg13g2_mux4_1
X_3348_ _1400_ _1006_ net1568 VPWR VGND sg13g2_nand2_1
X_6067_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 net288 VPWR VGND sg13g2_buf_1
XFILLER_45_208 VPWR VGND sg13g2_fill_1
X_3279_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[0\] Tile_X0Y1_DSP_bot.B0 net1640 _1331_
+ VPWR VGND sg13g2_mux2_1
XFILLER_38_260 VPWR VGND sg13g2_fill_1
X_5018_ net1951 net1852 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_107_221 VPWR VGND sg13g2_fill_2
XFILLER_5_348 VPWR VGND sg13g2_fill_1
XFILLER_122_213 VPWR VGND sg13g2_fill_1
XFILLER_122_235 VPWR VGND sg13g2_fill_1
XFILLER_76_311 VPWR VGND sg13g2_fill_2
XFILLER_123_70 VPWR VGND sg13g2_fill_2
XFILLER_123_81 VPWR VGND sg13g2_fill_2
XFILLER_44_230 VPWR VGND sg13g2_fill_2
XFILLER_16_90 VPWR VGND sg13g2_fill_1
XFILLER_8_153 VPWR VGND sg13g2_fill_1
X_2650_ net1562 net1571 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ _0731_ VPWR VGND sg13g2_mux2_1
XFILLER_8_175 VPWR VGND sg13g2_fill_2
X_2581_ net1658 net1564 _0666_ VPWR VGND sg13g2_nor2_1
Xoutput406 net406 Tile_X0Y1_EE4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput417 net417 Tile_X0Y1_EE4BEG[5] VPWR VGND sg13g2_buf_1
X_4320_ _2258_ _2257_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q
+ VPWR VGND sg13g2_nand2b_1
Xoutput428 net428 Tile_X0Y1_FrameData_O[15] VPWR VGND sg13g2_buf_1
Xoutput439 net439 Tile_X0Y1_FrameData_O[25] VPWR VGND sg13g2_buf_1
X_4251_ VPWR _2210_ _2209_ VGND sg13g2_inv_1
XFILLER_113_279 VPWR VGND sg13g2_fill_1
X_3202_ _1256_ _1255_ _1257_ VPWR VGND sg13g2_nor2b_1
X_4182_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q _1011_ _1483_
+ _0969_ net1576 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q _2151_
+ VPWR VGND sg13g2_mux4_1
X_3133_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q _1189_
+ _1190_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q sg13g2_a21oi_1
X_3064_ net150 net1668 _1124_ VPWR VGND sg13g2_nor2b_1
XFILLER_82_336 VPWR VGND sg13g2_fill_2
X_5458__590 VPWR VGND net590 sg13g2_tiehi
X_3966_ net1644 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X
+ _1973_ VPWR VGND sg13g2_nor2_2
X_2917_ _0984_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q net1929
+ VPWR VGND sg13g2_nand2b_1
X_5705_ net1873 net1740 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_5636_ net1868 net1769 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_3897_ _1910_ VPWR _1911_ VGND _0597_ net2005 sg13g2_o21ai_1
X_2848_ VGND VPWR _0058_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q
+ _0920_ _0919_ sg13g2_a21oi_1
X_2779_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q VPWR _0854_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q _0852_ sg13g2_o21ai_1
X_5567_ net1858 net1792 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_5498_ net1911 net1848 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_4518_ VPWR _0075_ net21 VGND sg13g2_inv_1
X_4449_ _2364_ _2365_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 VPWR VGND sg13g2_mux2_1
Xfanout1609 net1609 net1614 VPWR VGND sg13g2_buf_16
XFILLER_58_366 VPWR VGND sg13g2_fill_1
X_6119_ net75 net340 VPWR VGND sg13g2_buf_1
XFILLER_53_22 VPWR VGND sg13g2_decap_4
XFILLER_53_99 VPWR VGND sg13g2_decap_8
XFILLER_5_123 VPWR VGND sg13g2_fill_1
XFILLER_78_63 VPWR VGND sg13g2_fill_2
XFILLER_78_85 VPWR VGND sg13g2_fill_1
XFILLER_94_95 VPWR VGND sg13g2_decap_4
XFILLER_17_252 VPWR VGND sg13g2_fill_1
X_3820_ VGND VPWR net1706 net1678 _1849_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q
+ sg13g2_a21oi_1
X_3751_ _1781_ VPWR _1782_ VGND _1774_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q
+ sg13g2_o21ai_1
X_2702_ _0781_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q net100
+ VPWR VGND sg13g2_nand2b_1
X_3682_ _1716_ VPWR _1717_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q
+ _1714_ sg13g2_o21ai_1
XFILLER_64_2 VPWR VGND sg13g2_fill_1
X_5421_ net1993 net1819 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_2633_ _0714_ VPWR _0715_ VGND net67 net1674 sg13g2_o21ai_1
Xoutput225 net225 Tile_X0Y0_FrameData_O[13] VPWR VGND sg13g2_buf_1
Xoutput203 net203 Tile_X0Y0_E6BEG[8] VPWR VGND sg13g2_buf_1
X_2564_ net1682 net1592 net1583 net1521 net699 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q
+ _0650_ VPWR VGND sg13g2_mux4_1
X_5352_ net1984 net1843 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_99_211 VPWR VGND sg13g2_decap_8
Xoutput214 net214 Tile_X0Y0_EE4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput258 net258 Tile_X0Y0_FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
Xoutput247 net247 Tile_X0Y0_FrameData_O[4] VPWR VGND sg13g2_buf_1
Xoutput236 net236 Tile_X0Y0_FrameData_O[23] VPWR VGND sg13g2_buf_1
X_4303_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q net1579 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2
+ _0596_ _0566_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3
+ VPWR VGND sg13g2_mux4_1
Xoutput269 net269 Tile_X0Y0_FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
X_2495_ _0583_ VPWR _0584_ VGND _0582_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q
+ sg13g2_o21ai_1
X_5283_ net1971 net1729 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_205 VPWR VGND sg13g2_decap_8
X_4234_ _2195_ VPWR _2196_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q
+ _2189_ sg13g2_o21ai_1
X_4165_ net26 net1634 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q
+ _2136_ VPWR VGND sg13g2_mux2_1
X_3116_ _1172_ VPWR _1173_ VGND _1046_ _1044_ sg13g2_o21ai_1
X_4096_ net1673 net1611 net1603 net1623 net1633 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q
+ _2085_ VPWR VGND sg13g2_mux4_1
X_3047_ _1107_ _0849_ _1103_ VPWR VGND sg13g2_nand2_1
XFILLER_82_166 VPWR VGND sg13g2_fill_1
X_4998_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q _0537_
+ _0539_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q sg13g2_a21oi_1
X_3949_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q VPWR _1958_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q _1956_ sg13g2_o21ai_1
XFILLER_23_58 VPWR VGND sg13g2_fill_2
X_5619_ net1895 net1772 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_61_339 VPWR VGND sg13g2_fill_1
XFILLER_80_75 VPWR VGND sg13g2_decap_8
XFILLER_80_86 VPWR VGND sg13g2_fill_2
XFILLER_108_360 VPWR VGND sg13g2_fill_2
XFILLER_89_73 VPWR VGND sg13g2_fill_2
XFILLER_123_374 VPWR VGND sg13g2_fill_2
Xfanout1951 Tile_X0Y0_FrameData[31] net1951 VPWR VGND sg13g2_buf_1
Xfanout1940 Tile_X0Y0_FrameData[8] net1940 VPWR VGND sg13g2_buf_1
Xfanout1973 net1974 net1973 VPWR VGND sg13g2_buf_1
Xfanout1962 Tile_X0Y0_FrameData[27] net1962 VPWR VGND sg13g2_buf_1
Xfanout1995 net1996 net1995 VPWR VGND sg13g2_buf_1
Xfanout1984 Tile_X0Y0_FrameData[17] net1984 VPWR VGND sg13g2_buf_1
X_5970_ net18 net191 VPWR VGND sg13g2_buf_1
X_4921_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q net1534 net1542
+ net1549 net1556 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q _0465_
+ VPWR VGND sg13g2_mux4_1
X_4852_ net1516 net1708 net1684 _0400_ VPWR VGND sg13g2_mux2_1
XFILLER_20_203 VPWR VGND sg13g2_fill_1
X_3803_ VGND VPWR _1477_ _1832_ _1831_ _1830_ sg13g2_a21oi_2
X_4783_ VPWR _0334_ _0333_ VGND sg13g2_inv_1
X_3734_ VGND VPWR net1643 _0154_ _1765_ net1647 sg13g2_a21oi_1
X_3665_ VGND VPWR net164 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q
+ _1701_ _0151_ sg13g2_a21oi_1
X_2616_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5
+ net43 net17 net78 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q _0699_
+ VPWR VGND sg13g2_mux4_1
X_5404_ net1958 net1818 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_3596_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q net114 net122
+ net90 net98 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q _1636_
+ VPWR VGND sg13g2_mux4_1
X_2547_ net2 net9 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q _0633_
+ VPWR VGND sg13g2_mux2_1
X_5335_ net1955 net1721 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_2478_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q net1565 net1572
+ net1579 net1618 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q _0568_
+ VPWR VGND sg13g2_mux4_1
X_5266_ net1941 net1740 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_87_214 VPWR VGND sg13g2_fill_1
X_4217_ net1576 _0835_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q
+ _2182_ VPWR VGND sg13g2_mux2_1
X_5197_ net1993 net1764 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_4148_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q net1527 net1933
+ net2004 net1594 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q _2122_
+ VPWR VGND sg13g2_mux4_1
XFILLER_28_336 VPWR VGND sg13g2_fill_2
X_4079_ _2075_ VPWR _2076_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q
+ _2074_ sg13g2_o21ai_1
XFILLER_43_328 VPWR VGND sg13g2_fill_2
XFILLER_59_21 VPWR VGND sg13g2_decap_4
XFILLER_78_225 VPWR VGND sg13g2_decap_4
XFILLER_59_98 VPWR VGND sg13g2_fill_1
XFILLER_115_82 VPWR VGND sg13g2_fill_2
XFILLER_115_149 VPWR VGND sg13g2_fill_2
X_3450_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2
+ net14 net1935 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q
+ _1500_ VPWR VGND sg13g2_mux4_1
XFILLER_41_4 VPWR VGND sg13g2_fill_2
X_3381_ _1430_ _1397_ _1433_ VPWR VGND sg13g2_xor2_1
X_5120_ net1966 net1787 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_5051_ net1954 net1807 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_69_269 VPWR VGND sg13g2_fill_1
X_4002_ VGND VPWR net1702 _0174_ _2007_ _2006_ sg13g2_a21oi_1
Xfanout1770 net1771 net1770 VPWR VGND sg13g2_buf_1
Xfanout1792 net1800 net1792 VPWR VGND sg13g2_buf_1
Xfanout1781 net1784 net1781 VPWR VGND sg13g2_buf_1
XFILLER_37_155 VPWR VGND sg13g2_decap_4
XFILLER_37_199 VPWR VGND sg13g2_fill_1
X_4904_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q
+ _0449_ _0446_ _0450_ _0447_ sg13g2_a221oi_1
X_5884_ net1916 net1816 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_4835_ _0270_ _0264_ _0383_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 VPWR
+ VGND sg13g2_a21o_2
X_4766_ net155 net167 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q
+ _0317_ VPWR VGND sg13g2_mux2_1
X_3717_ _1749_ _1748_ VPWR VGND sg13g2_inv_2
X_4697_ _0250_ VPWR _0251_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q
+ _0244_ sg13g2_o21ai_1
X_3648_ VGND VPWR net100 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q
+ _1685_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q sg13g2_a21oi_1
X_3579_ _1620_ net1648 _0008_ VPWR VGND sg13g2_nand2_1
X_5318_ net1980 net1722 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_6298_ net160 net519 VPWR VGND sg13g2_buf_1
X_5249_ net1968 net1742 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_29_79 VPWR VGND sg13g2_fill_1
XFILLER_28_100 VPWR VGND sg13g2_decap_8
XFILLER_28_133 VPWR VGND sg13g2_fill_2
XFILLER_16_339 VPWR VGND sg13g2_fill_2
XFILLER_45_56 VPWR VGND sg13g2_decap_4
XFILLER_24_372 VPWR VGND sg13g2_fill_1
XFILLER_117_0 VPWR VGND sg13g2_fill_2
X_2950_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q _1011_
+ _1014_ _1013_ sg13g2_a21oi_1
XFILLER_15_383 VPWR VGND sg13g2_fill_2
X_2881_ _0950_ _0948_ _0951_ VPWR VGND sg13g2_nor2b_1
XFILLER_89_4 VPWR VGND sg13g2_fill_1
X_4620_ VPWR _0177_ net1603 VGND sg13g2_inv_1
X_4551_ VPWR _0108_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q VGND
+ sg13g2_inv_1
X_4482_ net1512 _2057_ _0039_ VPWR VGND sg13g2_nor2_1
X_3502_ _1545_ _1548_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q
+ _1549_ VPWR VGND sg13g2_nand3_1
X_3433_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q VPWR _1484_ VGND
+ net1687 _0175_ sg13g2_o21ai_1
X_6221_ net1895 net434 VPWR VGND sg13g2_buf_1
X_6152_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 net364 VPWR VGND sg13g2_buf_8
XFILLER_106_18 VPWR VGND sg13g2_fill_2
X_3364_ _1416_ _1396_ _1414_ VPWR VGND sg13g2_nand2_2
X_5103_ net1997 net1797 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_6083_ Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A net295 VPWR VGND sg13g2_buf_1
X_3295_ net1511 _1104_ _1347_ VPWR VGND sg13g2_nor2_1
X_5034_ net1987 net1853 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_5867_ net1878 net1814 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_5798_ net1896 net1716 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_4818_ _0366_ VPWR _0367_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q
+ net1561 sg13g2_o21ai_1
X_4749_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q VPWR _0301_ VGND
+ net1666 net1579 sg13g2_o21ai_1
Xinput103 Tile_X0Y1_E2MID[4] net103 VPWR VGND sg13g2_buf_1
Xinput136 Tile_X0Y1_N4END[5] net136 VPWR VGND sg13g2_buf_1
Xinput125 Tile_X0Y1_N2MID[2] net125 VPWR VGND sg13g2_buf_8
Xinput114 Tile_X0Y1_N1END[3] net114 VPWR VGND sg13g2_buf_1
XFILLER_48_217 VPWR VGND sg13g2_fill_1
XFILLER_102_163 VPWR VGND sg13g2_fill_1
Xinput147 Tile_X0Y1_W1END[0] net147 VPWR VGND sg13g2_buf_1
Xinput158 Tile_X0Y1_W2END[7] net158 VPWR VGND sg13g2_buf_1
Xinput169 Tile_X0Y1_WW4END[0] net169 VPWR VGND sg13g2_buf_1
XFILLER_71_220 VPWR VGND sg13g2_decap_4
XFILLER_8_302 VPWR VGND sg13g2_fill_2
X_3080_ VGND VPWR net53 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q
+ _1139_ _1138_ sg13g2_a21oi_1
XFILLER_94_312 VPWR VGND sg13g2_fill_1
X_3982_ VGND VPWR _1987_ _1985_ _1932_ sg13g2_or2_1
X_2933_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q VPWR _0999_ VGND
+ net1661 net148 sg13g2_o21ai_1
X_5721_ net1909 net1739 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_94_2 VPWR VGND sg13g2_fill_1
X_5652_ net1899 net1760 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_2864_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q net125 net32
+ net6 net85 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q _0934_ VPWR
+ VGND sg13g2_mux4_1
X_5583_ net1886 net1783 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_2795_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5
+ net43 net17 net78 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q _0869_
+ VPWR VGND sg13g2_mux4_1
X_4603_ VPWR _0160_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[19\] VGND sg13g2_inv_1
X_4534_ VPWR _0091_ net27 VGND sg13g2_inv_1
X_4465_ _2379_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q _2380_
+ VPWR VGND sg13g2_nor2b_1
X_4396_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q net113 net1926
+ net149 net1544 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q _2320_
+ VPWR VGND sg13g2_mux4_1
X_6204_ net1869 net447 VPWR VGND sg13g2_buf_1
X_3416_ VGND VPWR _1468_ _0235_ _1467_ sg13g2_or2_1
X_6135_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 net347 VPWR VGND sg13g2_buf_1
X_3347_ VGND VPWR _1399_ _1373_ _1398_ sg13g2_or2_1
X_6066_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 net287 VPWR VGND sg13g2_buf_8
X_3278_ _1319_ VPWR Tile_X0Y1_DSP_bot.B0 VGND _1324_ _1330_ sg13g2_o21ai_1
X_5017_ _0557_ net1681 net1518 VPWR VGND sg13g2_nand2b_1
XFILLER_21_172 VPWR VGND sg13g2_fill_2
XFILLER_67_21 VPWR VGND sg13g2_fill_1
XFILLER_107_83 VPWR VGND sg13g2_decap_8
XFILLER_29_261 VPWR VGND sg13g2_fill_1
Xoutput407 net407 Tile_X0Y1_EE4BEG[10] VPWR VGND sg13g2_buf_1
X_2580_ _0665_ _0664_ _0089_ VPWR VGND sg13g2_nand2_2
Xoutput418 net418 Tile_X0Y1_EE4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput429 net429 Tile_X0Y1_FrameData_O[16] VPWR VGND sg13g2_buf_1
X_4250_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q net1605 net1635
+ net1625 net1594 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q _2209_
+ VPWR VGND sg13g2_mux4_1
XFILLER_4_371 VPWR VGND sg13g2_fill_2
X_3201_ _1227_ _1221_ _1256_ VPWR VGND sg13g2_xor2_1
X_4181_ _2149_ VPWR _2150_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q
+ _2146_ sg13g2_o21ai_1
X_3132_ VGND VPWR net11 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q
+ _1189_ _1188_ sg13g2_a21oi_1
X_3063_ VGND VPWR _0099_ net1668 _1123_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q
+ sg13g2_a21oi_1
XFILLER_94_186 VPWR VGND sg13g2_fill_2
X_3965_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q _1972_ _1971_
+ _1954_ _0647_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X
+ VPWR VGND sg13g2_mux4_1
X_2916_ VGND VPWR _0983_ _0982_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q
+ sg13g2_or2_1
X_5704_ net1871 net1740 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_3896_ VGND VPWR net1706 net2005 _1910_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q
+ sg13g2_a21oi_1
X_2847_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q VPWR _0919_ VGND
+ net153 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q sg13g2_o21ai_1
X_5635_ net1866 net1769 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_2778_ net1690 net1594 net1588 net1523 net1541 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q
+ _0853_ VPWR VGND sg13g2_mux4_1
X_5566_ net1856 net1792 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_308 VPWR VGND sg13g2_fill_2
X_5497_ net1909 net1850 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_4517_ VPWR _0074_ net126 VGND sg13g2_inv_1
X_4448_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q net1618 _1699_
+ _1759_ _0926_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q _2365_
+ VPWR VGND sg13g2_mux4_1
XFILLER_104_225 VPWR VGND sg13g2_decap_4
X_4379_ _2304_ _2305_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 VPWR VGND sg13g2_mux2_1
XFILLER_37_24 VPWR VGND sg13g2_decap_8
X_6118_ net74 net339 VPWR VGND sg13g2_buf_1
XFILLER_85_186 VPWR VGND sg13g2_fill_2
X_6049_ Tile_X0Y1_FrameStrobe[17] net261 VPWR VGND sg13g2_buf_1
XFILLER_26_220 VPWR VGND sg13g2_decap_4
XFILLER_26_242 VPWR VGND sg13g2_decap_4
XFILLER_78_42 VPWR VGND sg13g2_fill_2
XFILLER_110_228 VPWR VGND sg13g2_fill_1
XFILLER_1_374 VPWR VGND sg13g2_fill_2
XFILLER_49_301 VPWR VGND sg13g2_fill_2
X_3750_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q _1780_
+ _1781_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q sg13g2_a21oi_1
X_2701_ _0779_ VPWR _0780_ VGND net696 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q
+ sg13g2_o21ai_1
X_3681_ _1716_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q _1715_
+ VPWR VGND sg13g2_nand2b_1
X_5420_ net1991 net1819 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_2632_ _0714_ net1674 net81 VPWR VGND sg13g2_nand2b_1
Xoutput226 net226 Tile_X0Y0_FrameData_O[14] VPWR VGND sg13g2_buf_1
X_2563_ _0648_ _0649_ VPWR VGND sg13g2_inv_4
X_5351_ net1981 net1842 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput215 net215 Tile_X0Y0_EE4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput204 net204 Tile_X0Y0_E6BEG[9] VPWR VGND sg13g2_buf_1
Xoutput248 net248 Tile_X0Y0_FrameData_O[5] VPWR VGND sg13g2_buf_1
Xoutput237 net237 Tile_X0Y0_FrameData_O[24] VPWR VGND sg13g2_buf_1
Xoutput259 net259 Tile_X0Y0_FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
X_4302_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q net1572 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1
+ net1517 _1673_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2
+ VPWR VGND sg13g2_mux4_1
X_5282_ net1969 net1730 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_2494_ _0583_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q _0581_
+ VPWR VGND sg13g2_nand2b_1
X_4233_ _2194_ VPWR _2195_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q
+ _2191_ sg13g2_o21ai_1
XFILLER_99_267 VPWR VGND sg13g2_fill_1
XFILLER_99_289 VPWR VGND sg13g2_fill_1
X_4164_ _2134_ VPWR _2135_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q
+ net681 sg13g2_o21ai_1
X_3115_ _1172_ _1169_ _1170_ VPWR VGND sg13g2_xnor2_1
X_4095_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q net1621 net701
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 _0385_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 VPWR VGND sg13g2_mux4_1
X_3046_ _1106_ _1103_ _0899_ VPWR VGND sg13g2_nand2_2
X_4997_ net1708 net2003 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q
+ _0538_ VPWR VGND sg13g2_mux2_1
X_3948_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q net1634 net1524
+ net1594 net1519 net1700 _1957_ VPWR VGND sg13g2_mux4_1
X_3879_ _1896_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[10\] net1656 VPWR VGND sg13g2_nand2_1
X_5618_ net1893 net1772 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_5549_ net1882 net1793 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_48_23 VPWR VGND sg13g2_fill_2
XFILLER_58_131 VPWR VGND sg13g2_fill_1
XFILLER_73_123 VPWR VGND sg13g2_fill_2
XFILLER_100_294 VPWR VGND sg13g2_decap_8
X_5474__606 VPWR VGND net606 sg13g2_tiehi
XFILLER_14_223 VPWR VGND sg13g2_fill_1
XFILLER_120_61 VPWR VGND sg13g2_fill_1
Xfanout1930 net1931 net1930 VPWR VGND sg13g2_buf_1
Xfanout1941 net1942 net1941 VPWR VGND sg13g2_buf_1
XFILLER_96_248 VPWR VGND sg13g2_fill_1
Xfanout1952 Tile_X0Y0_FrameData[31] net1952 VPWR VGND sg13g2_buf_1
Xfanout1985 net1986 net1985 VPWR VGND sg13g2_buf_1
Xfanout1963 Tile_X0Y0_FrameData[26] net1963 VPWR VGND sg13g2_buf_1
Xfanout1974 Tile_X0Y0_FrameData[21] net1974 VPWR VGND sg13g2_buf_1
XFILLER_37_315 VPWR VGND sg13g2_fill_1
Xfanout1996 Tile_X0Y0_FrameData[11] net1996 VPWR VGND sg13g2_buf_1
XFILLER_37_359 VPWR VGND sg13g2_fill_2
XFILLER_52_307 VPWR VGND sg13g2_fill_1
X_4920_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q _0193_
+ _0464_ _0463_ sg13g2_a21oi_1
X_4851_ _0398_ VPWR _0399_ VGND net1684 net135 sg13g2_o21ai_1
X_3802_ _1831_ _1474_ _1476_ VPWR VGND sg13g2_xnor2_1
XFILLER_60_384 VPWR VGND sg13g2_fill_1
X_4782_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q net26 net30 net62
+ net1932 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q _0333_ VPWR
+ VGND sg13g2_mux4_1
X_3733_ _1764_ net1637 Tile_X0Y1_DSP_bot.C2 VPWR VGND sg13g2_nand2_2
XFILLER_20_259 VPWR VGND sg13g2_fill_2
X_3664_ _1700_ _1699_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_62_0 VPWR VGND sg13g2_decap_8
X_2615_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q _0697_ _0099_
+ _0098_ _0100_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q _0698_
+ VPWR VGND sg13g2_mux4_1
X_5403_ net1954 net1818 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_3595_ _1635_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q _1634_
+ VPWR VGND sg13g2_nand2_1
X_5334_ net1949 net1721 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_2546_ _0631_ VPWR _0632_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ net1527 sg13g2_o21ai_1
X_2477_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q net1529 net636
+ net1550 net1560 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q _0567_
+ VPWR VGND sg13g2_mux4_1
X_5265_ net1940 net1743 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_4216_ _2180_ VPWR _2181_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q
+ net1518 sg13g2_o21ai_1
X_5196_ net1991 net1764 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_28_304 VPWR VGND sg13g2_fill_1
X_4147_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 _2120_ _2121_ _2114_
+ _2116_ VPWR VGND sg13g2_a22oi_1
X_4078_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q _2072_
+ _2075_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q sg13g2_a21oi_1
X_3029_ _1089_ VPWR _1090_ VGND net109 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q
+ sg13g2_o21ai_1
XFILLER_61_104 VPWR VGND sg13g2_fill_1
XFILLER_91_31 VPWR VGND sg13g2_fill_1
XFILLER_91_42 VPWR VGND sg13g2_fill_2
XFILLER_42_384 VPWR VGND sg13g2_fill_1
X_3380_ _1432_ _1426_ _1431_ VPWR VGND sg13g2_nand2_1
X_5050_ net1952 net1807 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
Xfanout1760 net1761 net1760 VPWR VGND sg13g2_buf_1
X_4001_ net1701 net1633 _2006_ VPWR VGND sg13g2_nor2_1
Xfanout1771 Tile_X0Y1_FrameStrobe[4] net1771 VPWR VGND sg13g2_buf_1
Xfanout1793 net1800 net1793 VPWR VGND sg13g2_buf_1
Xfanout1782 net1783 net1782 VPWR VGND sg13g2_buf_1
XFILLER_92_251 VPWR VGND sg13g2_fill_1
XFILLER_92_273 VPWR VGND sg13g2_fill_1
X_4903_ VGND VPWR net9 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q
+ _0449_ _0448_ sg13g2_a21oi_1
X_5883_ net1914 net1816 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_33_384 VPWR VGND sg13g2_fill_1
X_4834_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q
+ _0382_ _0378_ _0383_ _0380_ sg13g2_a221oi_1
X_4765_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q net1711 net119
+ net95 net1923 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q _0316_
+ VPWR VGND sg13g2_mux4_1
X_3716_ _1748_ _1436_ _1438_ VPWR VGND sg13g2_xnor2_1
X_4696_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q _0249_ _0250_
+ VPWR VGND sg13g2_nor2_1
X_3647_ _1683_ VPWR _1684_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q
+ net696 sg13g2_o21ai_1
X_3578_ _1619_ _1618_ _1616_ VPWR VGND sg13g2_nand2b_1
X_5317_ net1976 net1722 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_114_150 VPWR VGND sg13g2_fill_1
X_2529_ _0615_ _0616_ VPWR VGND sg13g2_inv_4
X_6297_ net159 net518 VPWR VGND sg13g2_buf_1
XFILLER_29_47 VPWR VGND sg13g2_decap_8
XFILLER_29_58 VPWR VGND sg13g2_fill_2
X_5248_ net1966 net1742 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_5179_ net1953 net1764 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_181 VPWR VGND sg13g2_decap_4
XFILLER_61_45 VPWR VGND sg13g2_decap_8
XFILLER_101_96 VPWR VGND sg13g2_fill_1
XFILLER_59_292 VPWR VGND sg13g2_fill_1
X_2880_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q VPWR _0950_ VGND
+ _0113_ _0949_ sg13g2_o21ai_1
XFILLER_30_343 VPWR VGND sg13g2_fill_1
X_4550_ VPWR _0107_ net1660 VGND sg13g2_inv_1
X_4481_ net1512 _1884_ _0038_ VPWR VGND sg13g2_nor2_1
X_3501_ _1546_ _1547_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q
+ _1548_ VPWR VGND sg13g2_nand3_1
X_6220_ net1899 net432 VPWR VGND sg13g2_buf_1
X_3432_ VPWR _1483_ _1482_ VGND sg13g2_inv_1
X_3363_ net625 net1548 _1415_ VPWR VGND sg13g2_nor2_1
X_5102_ net1995 net1795 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_25_0 VPWR VGND sg13g2_fill_2
X_6082_ Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A net294 VPWR VGND sg13g2_buf_1
X_3294_ _1346_ _0807_ net1628 VPWR VGND sg13g2_nand2_1
X_5033_ net1985 net1854 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
Xfanout1590 _0174_ net1590 VPWR VGND sg13g2_buf_1
XFILLER_80_254 VPWR VGND sg13g2_fill_2
X_5866_ net1876 net1814 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_33_181 VPWR VGND sg13g2_decap_4
X_4817_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q net1573
+ _0366_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q sg13g2_a21oi_1
X_5797_ net1874 net1716 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_4748_ net1618 net1666 _0300_ VPWR VGND sg13g2_nor2b_1
X_4679_ net1636 VPWR _0233_ VGND net1638 _0027_ sg13g2_o21ai_1
Xinput104 Tile_X0Y1_E2MID[5] net104 VPWR VGND sg13g2_buf_1
Xinput115 Tile_X0Y1_N2END[0] net115 VPWR VGND sg13g2_buf_1
XFILLER_0_258 VPWR VGND sg13g2_fill_2
Xinput126 Tile_X0Y1_N2MID[3] net126 VPWR VGND sg13g2_buf_1
Xinput159 Tile_X0Y1_W2MID[0] net159 VPWR VGND sg13g2_buf_1
Xinput137 net137 Tile_X0Y1_N4END[6] VPWR VGND sg13g2_buf_16
Xinput148 Tile_X0Y1_W1END[1] net148 VPWR VGND sg13g2_buf_1
XFILLER_56_34 VPWR VGND sg13g2_decap_8
XFILLER_56_45 VPWR VGND sg13g2_fill_2
XFILLER_112_95 VPWR VGND sg13g2_fill_1
XFILLER_71_243 VPWR VGND sg13g2_fill_1
XFILLER_24_170 VPWR VGND sg13g2_fill_1
XFILLER_12_321 VPWR VGND sg13g2_fill_1
XFILLER_71_298 VPWR VGND sg13g2_fill_1
XFILLER_47_240 VPWR VGND sg13g2_fill_1
XFILLER_94_346 VPWR VGND sg13g2_fill_2
X_3981_ net700 _1985_ _1986_ VPWR VGND sg13g2_nor2b_1
X_5720_ net1906 net1739 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_2932_ net150 net1661 _0998_ VPWR VGND sg13g2_nor2b_1
XFILLER_15_181 VPWR VGND sg13g2_fill_1
X_5651_ net1894 net1759 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_2863_ _0850_ _0930_ _0933_ VPWR VGND sg13g2_nor2_1
X_5582_ net1884 net1782 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_2794_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q _0627_ _0110_
+ _0066_ _0867_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q _0868_
+ VPWR VGND sg13g2_mux4_1
X_4602_ VPWR _0159_ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[19\] VGND sg13g2_inv_1
X_4533_ VPWR _0090_ net29 VGND sg13g2_inv_1
XFILLER_117_18 VPWR VGND sg13g2_fill_1
XFILLER_7_380 VPWR VGND sg13g2_fill_1
X_4464_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q _0905_ _1130_
+ _1759_ _1699_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q _2379_
+ VPWR VGND sg13g2_mux4_1
X_6203_ net1875 net444 VPWR VGND sg13g2_buf_1
X_4395_ _2319_ _2316_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 VPWR VGND sg13g2_mux2_1
X_3415_ _1467_ _1466_ _1465_ VPWR VGND sg13g2_nand2_2
X_6134_ Tile_X0Y0_W6END[11] net357 VPWR VGND sg13g2_buf_1
X_3346_ _1398_ _1103_ net1628 VPWR VGND sg13g2_nand2_2
XFILLER_97_151 VPWR VGND sg13g2_fill_2
X_6065_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 net286 VPWR VGND sg13g2_buf_1
X_3277_ _0132_ VPWR _1330_ VGND _1326_ _1329_ sg13g2_o21ai_1
X_5016_ _0555_ VPWR _0556_ VGND net1680 net1590 sg13g2_o21ai_1
XFILLER_38_251 VPWR VGND sg13g2_fill_2
XFILLER_53_221 VPWR VGND sg13g2_decap_8
X_5849_ net1909 net1824 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_4 VPWR VGND sg13g2_fill_2
XFILLER_107_267 VPWR VGND sg13g2_fill_1
XFILLER_76_313 VPWR VGND sg13g2_fill_1
XFILLER_123_83 VPWR VGND sg13g2_fill_1
XFILLER_123_72 VPWR VGND sg13g2_fill_1
XFILLER_44_232 VPWR VGND sg13g2_fill_1
XFILLER_44_254 VPWR VGND sg13g2_fill_1
XFILLER_16_70 VPWR VGND sg13g2_fill_1
XFILLER_12_184 VPWR VGND sg13g2_fill_2
Xoutput408 net408 Tile_X0Y1_EE4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput419 net419 Tile_X0Y1_EE4BEG[7] VPWR VGND sg13g2_buf_1
X_3200_ _1254_ VPWR _1255_ VGND _1244_ _1245_ sg13g2_o21ai_1
X_4180_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q _2148_
+ _2149_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q sg13g2_a21oi_1
X_3131_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q net2001 _1188_
+ VPWR VGND sg13g2_nor2b_1
X_3062_ _1122_ _0615_ net1668 VPWR VGND sg13g2_nand2b_1
X_3964_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0
+ net73 net12 net727 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q
+ _1972_ VPWR VGND sg13g2_mux4_1
XFILLER_92_0 VPWR VGND sg13g2_fill_2
X_2915_ _0981_ VPWR _0982_ VGND _0059_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q
+ sg13g2_o21ai_1
X_5703_ net1920 net1750 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_3895_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q _1907_
+ _1909_ _1908_ sg13g2_a21oi_1
X_2846_ _0917_ VPWR _0918_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q
+ _0916_ sg13g2_o21ai_1
X_5634_ net1864 net1769 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_2777_ VPWR _0852_ _0851_ VGND sg13g2_inv_1
X_5565_ net1917 net1792 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_4516_ VPWR _0073_ net89 VGND sg13g2_inv_1
X_5496_ net1907 net1850 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_4447_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q net112 net148
+ _0616_ net1564 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q _2364_
+ VPWR VGND sg13g2_mux4_1
X_4378_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q net1620 _1699_
+ _1759_ _1210_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q _2305_
+ VPWR VGND sg13g2_mux4_1
X_6117_ net73 net338 VPWR VGND sg13g2_buf_1
X_3329_ _1381_ _1023_ net1568 VPWR VGND sg13g2_nand2_1
X_6048_ Tile_X0Y1_FrameStrobe[16] net260 VPWR VGND sg13g2_buf_1
XFILLER_73_338 VPWR VGND sg13g2_fill_2
XFILLER_41_224 VPWR VGND sg13g2_fill_2
XFILLER_78_65 VPWR VGND sg13g2_fill_1
XFILLER_94_20 VPWR VGND sg13g2_fill_2
XFILLER_76_198 VPWR VGND sg13g2_decap_8
XFILLER_32_246 VPWR VGND sg13g2_fill_1
X_2700_ _0779_ net160 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q
+ VPWR VGND sg13g2_nand2_1
X_3680_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q net133 net153
+ net60 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q
+ _1715_ VPWR VGND sg13g2_mux4_1
X_2631_ _0712_ VPWR _0713_ VGND net20 net1674 sg13g2_o21ai_1
X_2562_ net1682 net1596 net1602 net1621 net1630 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q
+ _0648_ VPWR VGND sg13g2_mux4_1
X_5350_ net1979 net1842 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput205 net205 Tile_X0Y0_EE4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput216 net216 Tile_X0Y0_EE4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput227 net227 Tile_X0Y0_FrameData_O[15] VPWR VGND sg13g2_buf_1
Xoutput249 net249 Tile_X0Y0_FrameData_O[6] VPWR VGND sg13g2_buf_1
Xoutput238 net238 Tile_X0Y0_FrameData_O[25] VPWR VGND sg13g2_buf_1
X_4301_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q net1565 net689
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 _0362_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 VPWR VGND sg13g2_mux4_1
X_5281_ net1967 net1729 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_2493_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q net1597 net1610
+ net649 net1623 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q _0582_
+ VPWR VGND sg13g2_mux4_1
X_4232_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q _2193_
+ _2194_ _0164_ sg13g2_a21oi_1
X_4163_ VGND VPWR _0061_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q
+ _2134_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q sg13g2_a21oi_1
XFILLER_67_121 VPWR VGND sg13g2_fill_1
X_3114_ _1171_ _1169_ _1170_ VPWR VGND sg13g2_nand2b_1
X_4094_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q net124 net1929
+ net135 net1522 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3
+ VPWR VGND sg13g2_mux4_1
X_3045_ VGND VPWR _1102_ _0898_ _1101_ _0123_ _1105_ _0897_ sg13g2_a221oi_1
X_4996_ _0536_ VPWR _0537_ VGND net8 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q
+ sg13g2_o21ai_1
X_3947_ VPWR _1956_ _1955_ VGND sg13g2_inv_1
XFILLER_109_307 VPWR VGND sg13g2_fill_1
X_3878_ _1895_ _1826_ _1827_ VPWR VGND sg13g2_xnor2_1
X_2829_ _0901_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3
+ VPWR VGND sg13g2_nand2_1
X_5617_ net1890 net1772 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_5548_ net1880 net1793 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_5479_ Tile_X0Y1_UserCLK net555 net709 _5479_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[19\]
+ VPWR VGND sg13g2_dfrbp_1
XFILLER_100_284 VPWR VGND sg13g2_fill_1
XFILLER_104_96 VPWR VGND sg13g2_decap_8
X_5448__580 VPWR VGND net580 sg13g2_tiehi
XFILLER_89_75 VPWR VGND sg13g2_fill_1
XFILLER_123_376 VPWR VGND sg13g2_fill_1
XFILLER_96_205 VPWR VGND sg13g2_fill_2
XFILLER_96_216 VPWR VGND sg13g2_fill_1
Xfanout1920 Tile_X0Y1_FrameData[0] net1920 VPWR VGND sg13g2_buf_1
Xfanout1942 Tile_X0Y0_FrameData[7] net1942 VPWR VGND sg13g2_buf_1
Xfanout1931 Tile_X0Y0_W1END[3] net1931 VPWR VGND sg13g2_buf_1
Xfanout1986 Tile_X0Y0_FrameData[16] net1986 VPWR VGND sg13g2_buf_1
Xfanout1964 Tile_X0Y0_FrameData[26] net1964 VPWR VGND sg13g2_buf_1
Xfanout1975 net1976 net1975 VPWR VGND sg13g2_buf_1
Xfanout1953 Tile_X0Y0_FrameData[30] net1953 VPWR VGND sg13g2_buf_1
Xfanout1997 Tile_X0Y0_FrameData[10] net1997 VPWR VGND sg13g2_buf_1
X_4850_ _0398_ net1684 net8 VPWR VGND sg13g2_nand2b_1
XFILLER_72_190 VPWR VGND sg13g2_fill_1
X_3801_ _1507_ VPWR _1830_ VGND _1829_ _1828_ sg13g2_o21ai_1
X_4781_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q _0331_
+ _0332_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q sg13g2_a21oi_1
X_3732_ Tile_X0Y1_DSP_bot.C2 _1763_ VPWR VGND sg13g2_inv_2
XFILLER_13_290 VPWR VGND sg13g2_fill_1
X_3663_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q net103 net163
+ net615 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q
+ _1699_ VPWR VGND sg13g2_mux4_1
X_2614_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 _0697_ VPWR VGND sg13g2_inv_8
X_5402_ net1952 net1818 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_3594_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q _0616_ _0723_
+ net1934 net1704 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q _1634_
+ VPWR VGND sg13g2_mux4_1
XFILLER_55_0 VPWR VGND sg13g2_fill_2
X_5333_ net1947 net1721 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_2545_ VGND VPWR _0083_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ _0631_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q sg13g2_a21oi_1
X_2476_ VPWR _0566_ net684 VGND sg13g2_inv_1
X_5264_ net1937 net1743 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_5195_ net1989 net1763 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_4215_ _2180_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q _1482_
+ VPWR VGND sg13g2_nand2_1
X_4146_ _2118_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q _2121_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_28_338 VPWR VGND sg13g2_fill_1
X_4077_ VGND VPWR net1693 net1602 _2074_ _2073_ sg13g2_a21oi_1
X_3028_ _1089_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q net52 VPWR
+ VGND sg13g2_nand2b_1
XFILLER_70_127 VPWR VGND sg13g2_decap_8
X_4979_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q VPWR _0520_ VGND
+ net82 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q sg13g2_o21ai_1
XFILLER_59_67 VPWR VGND sg13g2_fill_2
XFILLER_120_357 VPWR VGND sg13g2_fill_1
XFILLER_115_84 VPWR VGND sg13g2_fill_1
XFILLER_46_179 VPWR VGND sg13g2_fill_2
XFILLER_108_181 VPWR VGND sg13g2_fill_1
Xfanout1750 net1757 net1750 VPWR VGND sg13g2_buf_1
XFILLER_84_219 VPWR VGND sg13g2_decap_8
X_4000_ _2004_ VPWR _2005_ VGND net1702 net1586 sg13g2_o21ai_1
Xfanout1761 net1762 net1761 VPWR VGND sg13g2_buf_1
Xfanout1783 net1784 net1783 VPWR VGND sg13g2_buf_1
Xfanout1772 net1774 net1772 VPWR VGND sg13g2_buf_1
Xfanout1794 net1800 net1794 VPWR VGND sg13g2_buf_1
XFILLER_52_116 VPWR VGND sg13g2_fill_1
X_4902_ net1677 net2004 _0448_ VPWR VGND sg13g2_nor2b_1
X_5882_ net1911 net1815 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_4833_ VPWR _0382_ _0381_ VGND sg13g2_inv_1
X_4764_ _0310_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q _0314_
+ _0315_ VPWR VGND sg13g2_nand3_1
X_3715_ _0018_ net1648 _1746_ _1747_ VPWR VGND sg13g2_a21o_1
X_4695_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q _0245_
+ _0249_ _0248_ sg13g2_a21oi_1
X_3646_ VGND VPWR net160 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q
+ _1683_ _0150_ sg13g2_a21oi_1
X_3577_ _1617_ _1451_ _1618_ VPWR VGND sg13g2_xor2_1
X_5316_ net1974 net1722 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_6296_ net158 net517 VPWR VGND sg13g2_buf_1
X_2528_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q net1590 _0610_
+ _0613_ _0612_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q _0615_
+ VPWR VGND sg13g2_mux4_1
X_5247_ net1963 net1742 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_5178_ net1951 net1764 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_28_135 VPWR VGND sg13g2_fill_1
X_4129_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q _0598_ net1930
+ net2001 net1625 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q _2105_
+ VPWR VGND sg13g2_mux4_1
XFILLER_28_179 VPWR VGND sg13g2_fill_1
XFILLER_24_341 VPWR VGND sg13g2_fill_1
XFILLER_101_53 VPWR VGND sg13g2_fill_1
XFILLER_117_2 VPWR VGND sg13g2_fill_1
XFILLER_86_21 VPWR VGND sg13g2_fill_2
XFILLER_59_260 VPWR VGND sg13g2_fill_1
XFILLER_34_105 VPWR VGND sg13g2_fill_2
X_3500_ _1547_ net1670 net1616 VPWR VGND sg13g2_nand2_1
X_4480_ _2389_ VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q
+ _2393_ sg13g2_o21ai_1
X_3431_ _1482_ _1481_ _1479_ VPWR VGND sg13g2_nand2b_1
X_3362_ _0929_ net1568 _1414_ VPWR VGND sg13g2_and2_1
X_6150_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 net362 VPWR VGND sg13g2_buf_2
X_5101_ net1993 net1795 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_97_322 VPWR VGND sg13g2_fill_2
X_6081_ Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A net308 VPWR VGND sg13g2_buf_1
XFILLER_57_208 VPWR VGND sg13g2_fill_2
X_3293_ _1344_ _1342_ _1345_ VPWR VGND sg13g2_nor2_2
XFILLER_111_187 VPWR VGND sg13g2_fill_1
X_5032_ net1983 net1854 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
Xfanout1591 net1591 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 VPWR VGND
+ sg13g2_buf_16
XFILLER_18_0 VPWR VGND sg13g2_fill_1
Xfanout1580 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 net1580 VPWR VGND sg13g2_buf_8
X_5865_ net1872 net1814 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_4816_ _0364_ _0363_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q
+ _0365_ VPWR VGND sg13g2_nand3_1
XFILLER_119_221 VPWR VGND sg13g2_fill_1
X_5796_ net1868 net1716 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_4747_ VGND VPWR _0297_ _0298_ _0299_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q
+ sg13g2_a21oi_1
X_4678_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q _0231_ _0232_
+ _0213_ _0195_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X
+ VPWR VGND sg13g2_mux4_1
X_3629_ VGND VPWR Tile_X0Y1_DSP_bot.C8 _1666_ _1649_ sg13g2_or2_1
XFILLER_88_311 VPWR VGND sg13g2_fill_1
XFILLER_102_110 VPWR VGND sg13g2_decap_8
Xinput105 Tile_X0Y1_E2MID[6] net105 VPWR VGND sg13g2_buf_1
Xinput127 Tile_X0Y1_N2MID[4] net127 VPWR VGND sg13g2_buf_1
Xinput116 Tile_X0Y1_N2END[1] net116 VPWR VGND sg13g2_buf_1
X_6279_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 net491 VPWR VGND sg13g2_buf_8
Xinput149 Tile_X0Y1_W1END[2] net149 VPWR VGND sg13g2_buf_1
Xinput138 Tile_X0Y1_N4END[7] net138 VPWR VGND sg13g2_buf_1
XFILLER_112_63 VPWR VGND sg13g2_decap_8
XFILLER_72_34 VPWR VGND sg13g2_fill_1
XFILLER_122_0 VPWR VGND sg13g2_fill_2
XFILLER_62_222 VPWR VGND sg13g2_decap_8
XFILLER_62_233 VPWR VGND sg13g2_fill_2
XFILLER_46_90 VPWR VGND sg13g2_fill_2
X_3980_ _1985_ _1983_ _1984_ _0036_ net1649 VPWR VGND sg13g2_a22oi_1
X_2931_ _0996_ VPWR _0997_ VGND net1661 _0723_ sg13g2_o21ai_1
X_5650_ net1892 net1759 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_2862_ _0932_ _0849_ net714 VPWR VGND sg13g2_nand2_1
X_4601_ VPWR _0158_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q VGND
+ sg13g2_inv_1
X_5581_ net1882 net1782 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_2793_ VPWR _0867_ net615 VGND sg13g2_inv_1
X_4532_ VPWR _0089_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q VGND
+ sg13g2_inv_1
X_4463_ _2377_ VPWR _2378_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q
+ _2374_ sg13g2_o21ai_1
X_6202_ net1897 net433 VPWR VGND sg13g2_buf_1
X_3414_ _1179_ _1456_ _1464_ _1466_ VPWR VGND sg13g2_or3_1
X_4394_ _2317_ _2318_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q
+ _2319_ VPWR VGND sg13g2_mux2_1
X_6133_ Tile_X0Y0_W6END[10] net356 VPWR VGND sg13g2_buf_1
X_3345_ _1397_ net1628 _1213_ VPWR VGND sg13g2_nand2_1
X_6064_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 net285 VPWR VGND sg13g2_buf_1
X_3276_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q VPWR _1329_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q _1328_ sg13g2_o21ai_1
X_5015_ VGND VPWR net1680 net1583 _0555_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q
+ sg13g2_a21oi_1
XFILLER_13_108 VPWR VGND sg13g2_fill_1
X_5848_ net1907 net1824 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_5779_ net1894 net1714 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_174 VPWR VGND sg13g2_fill_1
XFILLER_115_290 VPWR VGND sg13g2_fill_2
XFILLER_29_296 VPWR VGND sg13g2_fill_2
Xoutput409 net409 Tile_X0Y1_EE4BEG[12] VPWR VGND sg13g2_buf_1
X_3130_ _1186_ VPWR _1187_ VGND net1691 net622 sg13g2_o21ai_1
X_3061_ _1120_ VPWR _1121_ VGND _1118_ _1119_ sg13g2_o21ai_1
XFILLER_82_306 VPWR VGND sg13g2_fill_1
XFILLER_94_166 VPWR VGND sg13g2_fill_2
XFILLER_94_188 VPWR VGND sg13g2_fill_1
XFILLER_50_203 VPWR VGND sg13g2_fill_1
X_3963_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q net611 net39
+ net13 net74 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q _1971_
+ VPWR VGND sg13g2_mux4_1
X_2914_ _0981_ net34 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q
+ VPWR VGND sg13g2_nand2_1
XFILLER_50_269 VPWR VGND sg13g2_decap_8
X_5702_ net1897 net1748 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_3894_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q VPWR _1908_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q _1906_ sg13g2_o21ai_1
X_2845_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q _0914_
+ _0917_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q sg13g2_a21oi_1
X_5633_ net1862 net1769 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_5564_ net1915 net1792 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_2776_ net1690 net1599 net1612 net1605 net1625 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q
+ _0851_ VPWR VGND sg13g2_mux4_1
X_4515_ VPWR _0072_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q VGND
+ sg13g2_inv_1
X_5495_ net1905 net1847 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_4446_ VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 _2363_ VGND sg13g2_inv_1
XFILLER_104_238 VPWR VGND sg13g2_fill_2
X_5465__597 VPWR VGND net597 sg13g2_tiehi
X_4377_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q net1712 net1927
+ _0616_ net1566 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q _2304_
+ VPWR VGND sg13g2_mux4_1
X_3328_ _1378_ _1377_ _1376_ _1380_ VPWR VGND sg13g2_a21o_1
X_6116_ net72 net337 VPWR VGND sg13g2_buf_1
X_6047_ Tile_X0Y1_FrameStrobe[15] net259 VPWR VGND sg13g2_buf_1
X_3259_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q net94 _1312_ VPWR
+ VGND sg13g2_nor2b_1
XFILLER_26_288 VPWR VGND sg13g2_fill_2
XFILLER_41_203 VPWR VGND sg13g2_fill_2
XFILLER_81_361 VPWR VGND sg13g2_fill_2
XFILLER_41_269 VPWR VGND sg13g2_fill_2
XFILLER_118_51 VPWR VGND sg13g2_fill_1
XFILLER_1_376 VPWR VGND sg13g2_fill_1
XFILLER_78_77 VPWR VGND sg13g2_fill_1
XFILLER_49_358 VPWR VGND sg13g2_fill_2
XFILLER_91_125 VPWR VGND sg13g2_fill_1
XFILLER_40_291 VPWR VGND sg13g2_fill_1
X_2630_ _0712_ net1674 net32 VPWR VGND sg13g2_nand2b_1
X_2561_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q net143 net65
+ net20 _0646_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q _0647_
+ VPWR VGND sg13g2_mux4_1
Xoutput206 net206 Tile_X0Y0_EE4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput217 net217 Tile_X0Y0_EE4BEG[6] VPWR VGND sg13g2_buf_1
X_2492_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q net1632 net1585
+ net1522 net1520 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q _0581_
+ VPWR VGND sg13g2_mux4_1
Xoutput228 net228 Tile_X0Y0_FrameData_O[16] VPWR VGND sg13g2_buf_1
Xoutput239 net239 Tile_X0Y0_FrameData_O[26] VPWR VGND sg13g2_buf_1
X_4300_ _2237_ VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q
+ _2246_ sg13g2_o21ai_1
X_5280_ net1965 net1730 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_4231_ _2192_ VPWR _2193_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q
+ _0868_ sg13g2_o21ai_1
X_4162_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 _2133_ VGND sg13g2_inv_1
X_4093_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q net1709 net138
+ net82 net1586 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2
+ VPWR VGND sg13g2_mux4_1
X_3113_ _1042_ _1040_ _1170_ VPWR VGND sg13g2_nor2_2
XFILLER_55_328 VPWR VGND sg13g2_fill_2
X_3044_ _1104_ _1103_ VPWR VGND sg13g2_inv_2
XFILLER_70_309 VPWR VGND sg13g2_fill_1
XFILLER_63_372 VPWR VGND sg13g2_fill_2
X_4995_ _0536_ _0059_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q
+ VPWR VGND sg13g2_nand2_1
X_3946_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q net1600 net1612
+ net1606 net1626 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q _1955_
+ VPWR VGND sg13g2_mux4_1
X_3877_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q net1558 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1
+ net1517 _1673_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2
+ VPWR VGND sg13g2_mux4_1
X_2828_ net1708 net103 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q
+ _0900_ VPWR VGND sg13g2_mux2_1
X_5616_ net1889 net1772 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_5547_ net1878 net1793 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_2759_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q net123 net30
+ net23 net65 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q _0835_
+ VPWR VGND sg13g2_mux4_1
X_5478_ Tile_X0Y1_UserCLK net554 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X
+ _0037_ _5478_/Q VPWR VGND sg13g2_dfrbp_1
X_4429_ _2345_ _2348_ _2349_ VPWR VGND sg13g2_nor2_1
XFILLER_48_25 VPWR VGND sg13g2_fill_1
XFILLER_100_230 VPWR VGND sg13g2_fill_2
XFILLER_46_339 VPWR VGND sg13g2_fill_2
XFILLER_73_125 VPWR VGND sg13g2_fill_1
XFILLER_64_24 VPWR VGND sg13g2_fill_1
XFILLER_14_203 VPWR VGND sg13g2_fill_2
XFILLER_80_12 VPWR VGND sg13g2_fill_1
XFILLER_13_50 VPWR VGND sg13g2_fill_1
XFILLER_96_228 VPWR VGND sg13g2_decap_4
Xfanout1932 net64 net1932 VPWR VGND sg13g2_buf_1
Xfanout1910 net1911 net1910 VPWR VGND sg13g2_buf_1
Xfanout1921 Tile_X0Y1_E6END[1] net1921 VPWR VGND sg13g2_buf_1
Xfanout1943 net1944 net1943 VPWR VGND sg13g2_buf_1
Xfanout1965 net1966 net1965 VPWR VGND sg13g2_buf_1
Xfanout1976 Tile_X0Y0_FrameData[20] net1976 VPWR VGND sg13g2_buf_1
Xfanout1954 Tile_X0Y0_FrameData[30] net1954 VPWR VGND sg13g2_buf_1
Xfanout1987 net1988 net1987 VPWR VGND sg13g2_buf_1
Xfanout1998 Tile_X0Y0_FrameData[10] net1998 VPWR VGND sg13g2_buf_1
XFILLER_45_383 VPWR VGND sg13g2_fill_2
X_4780_ net1 net4 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q _0331_
+ VPWR VGND sg13g2_mux2_1
X_3800_ _1829_ _1504_ _1506_ VPWR VGND sg13g2_xnor2_1
X_3731_ _1763_ _1762_ _1753_ VPWR VGND sg13g2_nand2_2
XFILLER_118_105 VPWR VGND sg13g2_fill_1
XFILLER_9_251 VPWR VGND sg13g2_fill_2
X_3662_ _1697_ VPWR _1698_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q
+ _1695_ sg13g2_o21ai_1
X_3593_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 _1632_ _1633_ _1625_
+ _1623_ VPWR VGND sg13g2_a22oi_1
X_2613_ VGND VPWR _0689_ _0697_ _0696_ _0693_ sg13g2_a21oi_2
X_5401_ net1999 net1827 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_2544_ _0630_ _0629_ VPWR VGND _0544_ sg13g2_nand2b_2
X_5332_ net1945 net1720 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_48_0 VPWR VGND sg13g2_fill_2
X_2475_ _0564_ VPWR _0565_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q
+ _0561_ sg13g2_o21ai_1
X_5263_ net1998 net1742 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_5194_ net1987 net1763 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_4214_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q _2178_
+ _2179_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q sg13g2_a21oi_1
X_4145_ _2120_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q _2119_
+ VPWR VGND sg13g2_nand2_1
X_4076_ net1693 net1609 _2073_ VPWR VGND sg13g2_nor2b_1
X_3027_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q _1086_
+ _1088_ _1087_ sg13g2_a21oi_1
XFILLER_63_191 VPWR VGND sg13g2_fill_1
XFILLER_34_38 VPWR VGND sg13g2_decap_8
XFILLER_51_375 VPWR VGND sg13g2_fill_2
X_4978_ net1511 net1515 _0519_ VPWR VGND sg13g2_nor2_1
X_3929_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q VPWR _1940_ VGND
+ _0099_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q sg13g2_o21ai_1
XFILLER_109_138 VPWR VGND sg13g2_decap_4
XFILLER_109_149 VPWR VGND sg13g2_fill_1
XFILLER_105_344 VPWR VGND sg13g2_fill_1
XFILLER_120_314 VPWR VGND sg13g2_fill_2
XFILLER_59_79 VPWR VGND sg13g2_decap_8
XFILLER_115_63 VPWR VGND sg13g2_fill_2
XFILLER_86_250 VPWR VGND sg13g2_decap_8
XFILLER_54_180 VPWR VGND sg13g2_fill_1
Xfanout1740 net1741 net1740 VPWR VGND sg13g2_buf_1
Xfanout1751 net1752 net1751 VPWR VGND sg13g2_buf_1
Xfanout1773 net1774 net1773 VPWR VGND sg13g2_buf_1
Xfanout1762 Tile_X0Y1_FrameStrobe[5] net1762 VPWR VGND sg13g2_buf_1
Xfanout1784 Tile_X0Y1_FrameStrobe[3] net1784 VPWR VGND sg13g2_buf_1
XFILLER_77_272 VPWR VGND sg13g2_fill_1
Xfanout1795 net1796 net1795 VPWR VGND sg13g2_buf_1
X_4901_ VGND VPWR net128 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q
+ _0447_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q sg13g2_a21oi_1
XFILLER_45_180 VPWR VGND sg13g2_fill_2
X_5881_ net1908 net1812 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_4832_ net1683 net21 net33 net68 net82 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q
+ _0381_ VPWR VGND sg13g2_mux4_1
X_4763_ _0313_ VPWR _0314_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q
+ _0311_ sg13g2_o21ai_1
X_3714_ VGND VPWR _1745_ _1746_ Tile_X0Y1_DSP_bot.C3 net1637 sg13g2_a21oi_2
X_4694_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q VPWR _0248_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q _0247_ sg13g2_o21ai_1
X_3645_ VGND VPWR _1681_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q
+ _1680_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q _1682_ _1679_
+ sg13g2_a221oi_1
X_3576_ _1343_ _1342_ _1617_ VPWR VGND sg13g2_xor2_1
X_5315_ net1971 net1723 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_6295_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 net516 VPWR VGND sg13g2_buf_2
X_2527_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q net723 net45
+ net19 net80 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q _0614_
+ VPWR VGND sg13g2_mux4_1
X_5246_ net1962 net1742 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_28_114 VPWR VGND sg13g2_decap_8
X_5177_ net1999 net1777 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_4128_ _2104_ _2103_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 VPWR VGND sg13g2_mux2_1
X_4059_ _2058_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[1\] net1652 VPWR VGND sg13g2_nand2_1
XFILLER_43_117 VPWR VGND sg13g2_fill_1
XFILLER_43_139 VPWR VGND sg13g2_fill_2
XFILLER_51_161 VPWR VGND sg13g2_decap_8
XFILLER_101_87 VPWR VGND sg13g2_decap_4
XFILLER_19_71 VPWR VGND sg13g2_fill_1
XFILLER_86_99 VPWR VGND sg13g2_fill_2
X_3430_ _1480_ VPWR _1481_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q
+ net616 sg13g2_o21ai_1
X_3361_ _1413_ _1373_ _1398_ VPWR VGND sg13g2_xnor2_1
X_6080_ Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A net307 VPWR VGND sg13g2_buf_1
X_5100_ net1991 net1795 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_3292_ _1343_ _1344_ VPWR VGND sg13g2_inv_4
X_5031_ net1982 net1854 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
Xfanout1570 net1571 net1570 VPWR VGND sg13g2_buf_1
Xfanout1581 net1582 net1581 VPWR VGND sg13g2_buf_1
Xfanout1592 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 net1592 VPWR VGND
+ sg13g2_buf_8
XFILLER_65_264 VPWR VGND sg13g2_fill_2
XFILLER_65_286 VPWR VGND sg13g2_fill_1
XFILLER_80_201 VPWR VGND sg13g2_decap_8
XFILLER_21_312 VPWR VGND sg13g2_fill_1
X_5864_ net1870 net1815 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_4815_ _0364_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q net1617
+ VPWR VGND sg13g2_nand2_2
X_5795_ net1866 net1716 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_4746_ _0298_ net1565 net1666 VPWR VGND sg13g2_nand2b_1
XFILLER_119_288 VPWR VGND sg13g2_fill_2
X_4677_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q net145 net5 net31
+ net66 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q _0232_ VPWR VGND
+ sg13g2_mux4_1
X_3628_ VGND VPWR _1665_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q
+ _1664_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q _1666_ _1663_
+ sg13g2_a221oi_1
X_3559_ _0138_ _1601_ _1602_ VPWR VGND sg13g2_nor2_1
Xinput117 Tile_X0Y1_N2END[2] net117 VPWR VGND sg13g2_buf_1
Xinput106 Tile_X0Y1_E2MID[7] net106 VPWR VGND sg13g2_buf_1
X_6278_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 net505 VPWR VGND sg13g2_buf_8
Xinput128 Tile_X0Y1_N2MID[5] net128 VPWR VGND sg13g2_buf_1
Xinput139 Tile_X0Y1_NN4END[0] net139 VPWR VGND sg13g2_buf_1
XFILLER_48_209 VPWR VGND sg13g2_fill_2
X_5229_ net1994 net1753 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_242 VPWR VGND sg13g2_decap_8
XFILLER_112_75 VPWR VGND sg13g2_decap_8
XFILLER_115_0 VPWR VGND sg13g2_fill_1
X_2930_ VGND VPWR _0081_ net1661 _0996_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q
+ sg13g2_a21oi_1
XFILLER_62_278 VPWR VGND sg13g2_fill_1
X_4600_ VPWR _0157_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q VGND
+ sg13g2_inv_1
X_2861_ _0931_ _0807_ _0899_ VPWR VGND sg13g2_nand2_1
X_2792_ _0866_ _0855_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 VPWR VGND
+ sg13g2_nor2_2
X_5580_ net1880 net1782 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_4531_ VPWR _0088_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q VGND
+ sg13g2_inv_1
X_4462_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q _2376_
+ _2377_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q sg13g2_a21oi_1
X_6201_ net1920 net422 VPWR VGND sg13g2_buf_1
X_3413_ _1464_ VPWR _1465_ VGND _1456_ _1179_ sg13g2_o21ai_1
X_4393_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q net1544 net1551
+ net1560 net1566 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q _2318_
+ VPWR VGND sg13g2_mux4_1
X_6132_ Tile_X0Y0_W6END[9] net355 VPWR VGND sg13g2_buf_1
XFILLER_30_0 VPWR VGND sg13g2_fill_2
X_3344_ net1548 _0808_ _1396_ VPWR VGND sg13g2_nor2_2
X_3275_ _1327_ VPWR _1328_ VGND net1706 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q
+ sg13g2_o21ai_1
X_5014_ _0554_ _0553_ _0108_ VPWR VGND sg13g2_nand2_2
XFILLER_38_253 VPWR VGND sg13g2_fill_1
XFILLER_21_131 VPWR VGND sg13g2_fill_2
X_5847_ net1904 net1826 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_5778_ net1892 net1714 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_4729_ _0281_ VPWR _0282_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q
+ _0279_ sg13g2_o21ai_1
XFILLER_107_214 VPWR VGND sg13g2_decap_8
XFILLER_107_64 VPWR VGND sg13g2_fill_2
XFILLER_88_164 VPWR VGND sg13g2_fill_2
XFILLER_91_307 VPWR VGND sg13g2_fill_2
XFILLER_44_223 VPWR VGND sg13g2_decap_8
X_3060_ _0127_ _1115_ _1120_ VPWR VGND sg13g2_nor2_2
X_3962_ _1970_ _1959_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 VPWR VGND
+ sg13g2_nor2_2
X_5701_ net1874 net1746 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_92_2 VPWR VGND sg13g2_fill_1
X_2913_ _0980_ _0102_ _0979_ VPWR VGND sg13g2_nand2_1
X_3893_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q net1634 net1523
+ net1593 net1519 net2005 _1907_ VPWR VGND sg13g2_mux4_1
X_2844_ VGND VPWR net1928 net1667 _0916_ _0915_ sg13g2_a21oi_1
X_5632_ net1860 net1769 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_5563_ net1912 net1791 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_4514_ VPWR _0071_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q VGND
+ sg13g2_inv_1
X_2775_ _0850_ _0807_ _0849_ VPWR VGND sg13g2_nand2_2
X_5494_ net1903 net1847 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_4445_ _2357_ VPWR _2363_ VGND _2359_ _2362_ sg13g2_o21ai_1
X_4376_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 _2299_ _2303_ _2297_
+ _2295_ VPWR VGND sg13g2_a22oi_1
X_3327_ _1379_ _1378_ _1376_ VPWR VGND sg13g2_nand2b_1
X_6115_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 net336 VPWR VGND sg13g2_buf_2
X_6046_ Tile_X0Y1_FrameStrobe[14] net258 VPWR VGND sg13g2_buf_1
X_3258_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q _0966_
+ _1311_ _1310_ sg13g2_a21oi_1
X_3189_ _1105_ _1213_ net1575 _1244_ VPWR VGND sg13g2_nand3_1
XFILLER_41_226 VPWR VGND sg13g2_fill_1
XFILLER_81_384 VPWR VGND sg13g2_fill_1
XFILLER_76_112 VPWR VGND sg13g2_fill_2
XFILLER_94_22 VPWR VGND sg13g2_fill_1
XFILLER_94_99 VPWR VGND sg13g2_fill_2
Xoutput207 net207 Tile_X0Y0_EE4BEG[11] VPWR VGND sg13g2_buf_1
X_2560_ _0646_ _0645_ VPWR VGND _0637_ sg13g2_nand2b_2
Xoutput229 net229 Tile_X0Y0_FrameData_O[17] VPWR VGND sg13g2_buf_1
X_2491_ VPWR _0580_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 VGND sg13g2_inv_1
XFILLER_99_204 VPWR VGND sg13g2_decap_8
Xoutput218 net218 Tile_X0Y0_EE4BEG[7] VPWR VGND sg13g2_buf_1
X_4230_ _2192_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q _1469_
+ VPWR VGND sg13g2_nand2_1
X_4161_ _2132_ VPWR _2133_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q
+ _2126_ sg13g2_o21ai_1
XFILLER_67_112 VPWR VGND sg13g2_decap_8
X_3112_ _1168_ _1164_ _1169_ VPWR VGND sg13g2_xor2_1
X_4092_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q net126 net137
+ net20 net1591 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1
+ VPWR VGND sg13g2_mux4_1
X_3043_ _1103_ _1101_ _1102_ VPWR VGND sg13g2_nand2_2
XFILLER_67_189 VPWR VGND sg13g2_fill_1
XFILLER_23_237 VPWR VGND sg13g2_fill_2
X_4994_ _0534_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q _0535_
+ VPWR VGND sg13g2_nor2b_1
X_3945_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q net124 net31
+ net25 net66 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q _1954_
+ VPWR VGND sg13g2_mux4_1
X_3876_ _1894_ VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 VGND net1654 _1893_
+ sg13g2_o21ai_1
X_5615_ net1886 net1772 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_2827_ VGND VPWR _0898_ _0899_ _0123_ _0897_ sg13g2_a21oi_2
XFILLER_117_353 VPWR VGND sg13g2_fill_2
X_5546_ net1877 net1793 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_2758_ VGND VPWR _0833_ _0834_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q
+ _0830_ sg13g2_a21oi_2
X_5477_ Tile_X0Y1_UserCLK net609 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X
+ _0035_ _5477_/Q VPWR VGND sg13g2_dfrbp_1
X_4428_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q VPWR _2348_ VGND
+ _2346_ _2347_ sg13g2_o21ai_1
X_2689_ _0766_ net1640 _0767_ _0768_ VPWR VGND sg13g2_a21o_1
X_4359_ _2288_ VPWR _2289_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q
+ _1278_ sg13g2_o21ai_1
XFILLER_100_220 VPWR VGND sg13g2_decap_8
XFILLER_100_242 VPWR VGND sg13g2_decap_4
X_6029_ net1958 net242 VPWR VGND sg13g2_buf_1
XFILLER_46_329 VPWR VGND sg13g2_fill_2
XFILLER_58_189 VPWR VGND sg13g2_fill_2
XFILLER_81_170 VPWR VGND sg13g2_fill_1
XFILLER_80_57 VPWR VGND sg13g2_fill_1
Xfanout1900 Tile_X0Y1_FrameData[18] net1900 VPWR VGND sg13g2_buf_1
XFILLER_96_207 VPWR VGND sg13g2_fill_1
Xfanout1933 net63 net1933 VPWR VGND sg13g2_buf_1
Xfanout1911 Tile_X0Y1_FrameData[13] net1911 VPWR VGND sg13g2_buf_1
Xfanout1922 Tile_X0Y1_E6END[1] net1922 VPWR VGND sg13g2_buf_1
Xfanout1966 Tile_X0Y0_FrameData[25] net1966 VPWR VGND sg13g2_buf_1
XFILLER_49_156 VPWR VGND sg13g2_fill_2
Xfanout1944 Tile_X0Y0_FrameData[6] net1944 VPWR VGND sg13g2_buf_1
Xfanout1977 net1978 net1977 VPWR VGND sg13g2_buf_1
Xfanout1955 net1956 net1955 VPWR VGND sg13g2_buf_1
Xfanout1999 Tile_X0Y0_FrameData[0] net1999 VPWR VGND sg13g2_buf_1
Xfanout1988 Tile_X0Y0_FrameData[15] net1988 VPWR VGND sg13g2_buf_1
XFILLER_64_148 VPWR VGND sg13g2_decap_8
XFILLER_45_362 VPWR VGND sg13g2_fill_1
X_3730_ _1761_ VPWR _1762_ VGND _1758_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q
+ sg13g2_o21ai_1
X_3661_ _1697_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q _1696_
+ VPWR VGND sg13g2_nand2b_1
X_3592_ VGND VPWR _1627_ _1630_ _1633_ _0149_ sg13g2_a21oi_1
X_2612_ _0695_ _0097_ _0696_ VPWR VGND sg13g2_nor2_2
X_5400_ net1977 net1827 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_2543_ _0628_ VPWR _0629_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q
+ _0627_ sg13g2_o21ai_1
X_5331_ net1944 net1720 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_2474_ _0564_ _0563_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q
+ VPWR VGND sg13g2_nand2_2
X_5262_ net1996 net1742 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_4213_ net62 net1631 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q
+ _2178_ VPWR VGND sg13g2_mux2_1
X_5193_ net1985 net1764 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_4144_ net1576 _0934_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q
+ _2119_ VPWR VGND sg13g2_mux2_1
XFILLER_18_18 VPWR VGND sg13g2_fill_1
X_4075_ net1621 net1629 net1693 _2072_ VPWR VGND sg13g2_mux2_1
X_3026_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q VPWR _1087_ VGND
+ net158 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q sg13g2_o21ai_1
XFILLER_36_384 VPWR VGND sg13g2_fill_1
X_4977_ VGND VPWR _0517_ _0518_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[7\] net1641 sg13g2_a21oi_2
X_3928_ _1938_ VPWR _1939_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q
+ _0697_ sg13g2_o21ai_1
X_3859_ _1884_ _1434_ net644 VPWR VGND sg13g2_xnor2_1
X_5529_ net1908 net1802 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_78_229 VPWR VGND sg13g2_fill_1
XFILLER_86_295 VPWR VGND sg13g2_fill_2
X_5439__559 VPWR VGND net559 sg13g2_tiehi
XFILLER_27_384 VPWR VGND sg13g2_fill_1
XFILLER_40_82 VPWR VGND sg13g2_decap_8
Xfanout1741 Tile_X0Y1_FrameStrobe[7] net1741 VPWR VGND sg13g2_buf_1
Xfanout1730 net1734 net1730 VPWR VGND sg13g2_buf_1
Xfanout1785 net1786 net1785 VPWR VGND sg13g2_buf_1
Xfanout1774 Tile_X0Y1_FrameStrobe[4] net1774 VPWR VGND sg13g2_buf_1
Xfanout1752 net1753 net1752 VPWR VGND sg13g2_buf_1
Xfanout1763 net1768 net1763 VPWR VGND sg13g2_buf_1
Xfanout1796 net1797 net1796 VPWR VGND sg13g2_buf_1
XFILLER_37_159 VPWR VGND sg13g2_fill_2
X_4900_ _0446_ net1527 net1677 VPWR VGND sg13g2_nand2b_1
X_5880_ net1906 net1812 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_4831_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q _0379_
+ _0380_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q sg13g2_a21oi_1
XFILLER_60_151 VPWR VGND sg13g2_fill_1
X_4762_ VGND VPWR _0067_ _0313_ _0312_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q
+ sg13g2_a21oi_2
X_3713_ net1636 VPWR _1745_ VGND net1637 _0019_ sg13g2_o21ai_1
X_4693_ VGND VPWR net33 net1676 _0247_ _0246_ sg13g2_a21oi_1
X_3644_ VGND VPWR net99 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q
+ _1681_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q sg13g2_a21oi_1
XFILLER_60_0 VPWR VGND sg13g2_fill_2
X_3575_ _0006_ net1651 _1615_ _1616_ VPWR VGND sg13g2_a21o_1
X_5314_ net1970 net1723 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_6294_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 net515 VPWR VGND sg13g2_buf_8
X_2526_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q _0435_ _0081_
+ _0080_ _0082_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q _0613_
+ VPWR VGND sg13g2_mux4_1
X_5245_ net1959 net1745 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_5176_ net1978 net1777 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_4127_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q net1516 net3
+ net1932 net1605 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q _2104_
+ VPWR VGND sg13g2_mux4_1
X_4058_ _2057_ _1805_ _1806_ VPWR VGND sg13g2_xnor2_1
XFILLER_45_27 VPWR VGND sg13g2_fill_2
X_3009_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 _1064_ _1071_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q
+ _1062_ VPWR VGND sg13g2_a22oi_1
XFILLER_61_26 VPWR VGND sg13g2_fill_2
XFILLER_61_59 VPWR VGND sg13g2_fill_2
XFILLER_3_236 VPWR VGND sg13g2_fill_1
Xoutput390 net390 Tile_X0Y1_E2BEGb[4] VPWR VGND sg13g2_buf_1
XFILLER_101_370 VPWR VGND sg13g2_fill_1
XFILLER_34_107 VPWR VGND sg13g2_fill_1
XFILLER_30_357 VPWR VGND sg13g2_fill_2
X_3360_ _1410_ _1411_ _1412_ VPWR VGND sg13g2_nor2b_1
XFILLER_111_134 VPWR VGND sg13g2_decap_8
XFILLER_32_4 VPWR VGND sg13g2_fill_2
X_3291_ _1343_ _1284_ _1291_ VPWR VGND sg13g2_xnor2_1
X_5030_ net1980 net1854 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
Xfanout1560 net719 net1560 VPWR VGND sg13g2_buf_1
Xfanout1593 net1594 net1593 VPWR VGND sg13g2_buf_1
Xfanout1571 _0173_ net1571 VPWR VGND sg13g2_buf_1
Xfanout1582 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 net1582 VPWR VGND sg13g2_buf_1
XFILLER_25_129 VPWR VGND sg13g2_fill_2
X_5863_ net1920 net1826 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_5794_ net1864 net1714 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_4814_ _0363_ net1578 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q
+ VPWR VGND sg13g2_nand2b_1
X_4745_ _0297_ net1666 net1572 VPWR VGND sg13g2_nand2_1
XFILLER_31_18 VPWR VGND sg13g2_fill_2
X_4676_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q net12 net73 net38
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q
+ _0231_ VPWR VGND sg13g2_mux4_1
X_3627_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4
+ _1665_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q sg13g2_a21oi_1
X_5429__569 VPWR VGND net569 sg13g2_tiehi
X_3558_ VGND VPWR net1705 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q
+ _1601_ _1600_ sg13g2_a21oi_1
X_2509_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q net1562 _0580_
+ _0595_ _0565_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q _0597_
+ VPWR VGND sg13g2_mux4_1
Xinput118 Tile_X0Y1_N2END[3] net118 VPWR VGND sg13g2_buf_1
Xinput107 Tile_X0Y1_EE4END[0] net107 VPWR VGND sg13g2_buf_1
X_3489_ _0004_ net1650 _1535_ _1536_ VPWR VGND sg13g2_a21o_1
X_6277_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 net504 VPWR VGND sg13g2_buf_1
Xinput129 Tile_X0Y1_N2MID[6] net129 VPWR VGND sg13g2_buf_1
X_5228_ net1992 net1751 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_5159_ net1982 net1778 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_112_32 VPWR VGND sg13g2_fill_1
XFILLER_71_213 VPWR VGND sg13g2_decap_8
XFILLER_71_224 VPWR VGND sg13g2_fill_2
XFILLER_122_2 VPWR VGND sg13g2_fill_1
XFILLER_108_0 VPWR VGND sg13g2_fill_2
XFILLER_46_92 VPWR VGND sg13g2_fill_1
X_2860_ _0930_ _0899_ net714 VPWR VGND sg13g2_nand2_1
X_2791_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q _0860_ _0865_
+ _0866_ VPWR VGND sg13g2_nor3_1
XFILLER_7_31 VPWR VGND sg13g2_fill_2
X_4530_ VPWR _0087_ net47 VGND sg13g2_inv_1
X_4461_ VPWR _2376_ _2375_ VGND sg13g2_inv_1
XFILLER_7_361 VPWR VGND sg13g2_fill_1
X_6200_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 net412 VPWR VGND sg13g2_buf_1
X_3412_ _1463_ _1457_ _1464_ VPWR VGND sg13g2_xor2_1
X_6131_ Tile_X0Y0_W6END[8] net354 VPWR VGND sg13g2_buf_1
X_4392_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q net89 net149
+ net1530 net1535 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q _2317_
+ VPWR VGND sg13g2_mux4_1
X_3343_ _1395_ _1379_ _1377_ VPWR VGND sg13g2_xnor2_1
X_3274_ _1327_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q net106
+ VPWR VGND sg13g2_nand2b_1
X_6062_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 net283 VPWR VGND sg13g2_buf_1
X_5013_ net1681 net1609 net1602 net1621 net1629 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q
+ _0553_ VPWR VGND sg13g2_mux4_1
XFILLER_53_235 VPWR VGND sg13g2_fill_1
XFILLER_42_17 VPWR VGND sg13g2_fill_2
X_5846_ net1902 net1832 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_5777_ net1891 net1718 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_2989_ _1052_ _1050_ _0772_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_198 VPWR VGND sg13g2_fill_1
X_4728_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q _0280_
+ _0281_ _0063_ sg13g2_a21oi_1
X_4659_ VGND VPWR net1699 net1539 _0215_ _0214_ sg13g2_a21oi_1
XFILLER_122_218 VPWR VGND sg13g2_fill_1
X_6329_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 net541 VPWR VGND sg13g2_buf_1
XFILLER_76_327 VPWR VGND sg13g2_fill_2
XFILLER_29_298 VPWR VGND sg13g2_fill_1
XFILLER_8_114 VPWR VGND sg13g2_fill_2
XFILLER_94_168 VPWR VGND sg13g2_fill_1
X_3961_ VGND VPWR _1969_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q
+ _1966_ _1961_ _1970_ _1964_ sg13g2_a221oi_1
X_2912_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q net1708 net135
+ net2003 net8 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q _0979_
+ VPWR VGND sg13g2_mux4_1
X_5700_ net1868 net1746 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_73_90 VPWR VGND sg13g2_fill_1
X_3892_ VPWR _1906_ _1905_ VGND sg13g2_inv_1
X_5631_ net1858 net1771 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_2843_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q net141 _0915_
+ VPWR VGND sg13g2_nor2b_1
X_5562_ net1910 net1791 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_2774_ _0849_ _0848_ VPWR VGND sg13g2_inv_8
X_4513_ VPWR _0070_ net26 VGND sg13g2_inv_1
X_5493_ net1901 net1846 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
Xhold136 _0024_ VPWR VGND net745 sg13g2_dlygate4sd3_1
X_4444_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q VPWR _2362_ VGND
+ _2360_ _2361_ sg13g2_o21ai_1
XFILLER_104_229 VPWR VGND sg13g2_fill_1
X_4375_ VPWR _2303_ _2302_ VGND sg13g2_inv_1
X_3326_ _1375_ VPWR _1378_ VGND net1608 _1104_ sg13g2_o21ai_1
X_6114_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 net335 VPWR VGND sg13g2_buf_1
X_6045_ Tile_X0Y1_FrameStrobe[13] net257 VPWR VGND sg13g2_buf_1
X_3257_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q VPWR _1310_ VGND
+ net171 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q sg13g2_o21ai_1
XFILLER_26_213 VPWR VGND sg13g2_decap_8
X_3188_ _1106_ _1242_ _1243_ VPWR VGND sg13g2_nor2_2
XFILLER_66_371 VPWR VGND sg13g2_fill_1
XFILLER_26_224 VPWR VGND sg13g2_fill_1
X_5829_ net1875 net1837 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_5_128 VPWR VGND sg13g2_fill_1
XFILLER_118_86 VPWR VGND sg13g2_fill_1
XFILLER_103_251 VPWR VGND sg13g2_decap_4
XFILLER_49_349 VPWR VGND sg13g2_fill_1
XFILLER_57_371 VPWR VGND sg13g2_fill_1
XFILLER_76_179 VPWR VGND sg13g2_fill_2
XFILLER_27_94 VPWR VGND sg13g2_fill_2
Xoutput208 net208 Tile_X0Y0_EE4BEG[12] VPWR VGND sg13g2_buf_1
X_2490_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 _0572_ _0579_ _0570_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q VPWR VGND sg13g2_a22oi_1
Xoutput219 net219 Tile_X0Y0_EE4BEG[8] VPWR VGND sg13g2_buf_1
X_4160_ _2131_ VPWR _2132_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q
+ _2128_ sg13g2_o21ai_1
X_3111_ _1168_ _1038_ _1166_ VPWR VGND sg13g2_xnor2_1
X_4091_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q net125 net136
+ net21 net1633 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0
+ VPWR VGND sg13g2_mux4_1
X_3042_ _1102_ Tile_X0Y1_DSP_bot.A1 net1641 VPWR VGND sg13g2_nand2b_1
XFILLER_67_168 VPWR VGND sg13g2_decap_4
XFILLER_63_352 VPWR VGND sg13g2_fill_2
XFILLER_63_374 VPWR VGND sg13g2_fill_1
X_4993_ VGND VPWR _0533_ _0534_ _0532_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q
+ sg13g2_a21oi_2
XFILLER_90_171 VPWR VGND sg13g2_fill_1
X_3944_ VGND VPWR _1948_ _1953_ _1951_ _1949_ sg13g2_a21oi_2
X_3875_ _1894_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[9\] net1654 VPWR VGND sg13g2_nand2_1
X_5614_ net1884 net1772 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_2826_ net1640 Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[6\] _0898_ VPWR VGND sg13g2_nor2_1
XFILLER_117_321 VPWR VGND sg13g2_fill_1
X_5545_ net1872 net1793 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_2757_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q VPWR _0833_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q _0832_ sg13g2_o21ai_1
X_2688_ net1640 Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[3\] _0767_ VPWR VGND sg13g2_nor2_1
X_5476_ Tile_X0Y1_UserCLK net608 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X
+ _0033_ _5476_/Q VPWR VGND sg13g2_dfrbp_1
X_4427_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q VPWR _2347_ VGND
+ _0169_ _1695_ sg13g2_o21ai_1
X_4358_ _2288_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q _1734_
+ VPWR VGND sg13g2_nand2_1
XFILLER_58_113 VPWR VGND sg13g2_fill_2
X_4289_ _2235_ VPWR _2236_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q
+ _2234_ sg13g2_o21ai_1
X_3309_ _1352_ _1351_ _1361_ VPWR VGND sg13g2_xor2_1
XFILLER_100_232 VPWR VGND sg13g2_fill_1
X_6028_ net1959 net241 VPWR VGND sg13g2_buf_1
XFILLER_73_116 VPWR VGND sg13g2_decap_8
XFILLER_54_363 VPWR VGND sg13g2_fill_2
XFILLER_64_48 VPWR VGND sg13g2_fill_2
XFILLER_14_205 VPWR VGND sg13g2_fill_1
Xfanout1912 net1913 net1912 VPWR VGND sg13g2_buf_1
Xfanout1901 Tile_X0Y1_FrameData[18] net1901 VPWR VGND sg13g2_buf_1
XFILLER_1_186 VPWR VGND sg13g2_fill_2
Xfanout1923 net1924 net1923 VPWR VGND sg13g2_buf_1
Xfanout1934 net45 net1934 VPWR VGND sg13g2_buf_1
Xfanout1967 net1968 net1967 VPWR VGND sg13g2_buf_1
Xfanout1945 Tile_X0Y0_FrameData[5] net1945 VPWR VGND sg13g2_buf_1
Xfanout1956 Tile_X0Y0_FrameData[2] net1956 VPWR VGND sg13g2_buf_1
Xfanout1989 net1990 net1989 VPWR VGND sg13g2_buf_1
Xfanout1978 Tile_X0Y0_FrameData[1] net1978 VPWR VGND sg13g2_buf_1
XFILLER_64_127 VPWR VGND sg13g2_decap_4
X_5455__587 VPWR VGND net587 sg13g2_tiehi
XFILLER_60_333 VPWR VGND sg13g2_fill_2
X_3660_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q net1922 net51
+ net172 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q
+ _1696_ VPWR VGND sg13g2_mux4_1
XFILLER_70_80 VPWR VGND sg13g2_fill_1
X_3591_ _1632_ _0148_ _1631_ VPWR VGND sg13g2_nand2_2
X_2611_ _0694_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q _0695_
+ VPWR VGND sg13g2_nor2_2
X_2542_ VGND VPWR net16 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q
+ _0628_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q sg13g2_a21oi_1
X_5330_ net1942 net1719 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_5261_ net1994 net1740 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_2473_ VGND VPWR _0562_ _0563_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q sg13g2_a21oi_2
X_4212_ _2176_ VPWR _2177_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q
+ net681 sg13g2_o21ai_1
X_5192_ net1983 net1767 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_4143_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q _1482_
+ _2118_ _2117_ sg13g2_a21oi_1
X_4074_ _0088_ VPWR _2071_ VGND _2069_ _2070_ sg13g2_o21ai_1
X_3025_ VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 _1086_ VGND sg13g2_inv_1
XFILLER_95_285 VPWR VGND sg13g2_fill_2
XFILLER_51_366 VPWR VGND sg13g2_fill_1
X_4976_ net1641 _0516_ _0517_ VPWR VGND sg13g2_nor2_2
X_3927_ VGND VPWR net17 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q
+ _1938_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q sg13g2_a21oi_1
X_3858_ _1883_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[2\] net1652 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ VPWR VGND sg13g2_mux2_1
X_3789_ _1731_ VPWR _1818_ VGND _1815_ _1816_ sg13g2_o21ai_1
X_2809_ net1688 net146 net2004 net7 net21 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q
+ _0883_ VPWR VGND sg13g2_mux4_1
X_5528_ net1906 net1802 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput550 net550 Tile_X0Y1_WW4BEG[6] VPWR VGND sg13g2_buf_1
X_5459_ Tile_X0Y1_UserCLK net591 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X
+ _5459_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[7\] VPWR VGND sg13g2_dfrbp_1
XFILLER_120_316 VPWR VGND sg13g2_fill_1
X_5478__554 VPWR VGND net554 sg13g2_tiehi
XFILLER_49_70 VPWR VGND sg13g2_fill_1
Xfanout1720 net1721 net1720 VPWR VGND sg13g2_buf_1
Xfanout1742 net1744 net1742 VPWR VGND sg13g2_buf_1
Xfanout1731 net1733 net1731 VPWR VGND sg13g2_buf_1
Xfanout1775 net1776 net1775 VPWR VGND sg13g2_buf_1
Xfanout1753 net1757 net1753 VPWR VGND sg13g2_buf_1
Xfanout1764 net1765 net1764 VPWR VGND sg13g2_buf_1
Xfanout1797 net1800 net1797 VPWR VGND sg13g2_buf_1
Xfanout1786 net1788 net1786 VPWR VGND sg13g2_buf_1
XFILLER_18_352 VPWR VGND sg13g2_fill_2
XFILLER_18_374 VPWR VGND sg13g2_fill_2
XFILLER_33_311 VPWR VGND sg13g2_fill_2
XFILLER_92_299 VPWR VGND sg13g2_fill_1
X_4830_ net138 net7 net1683 _0379_ VPWR VGND sg13g2_mux2_1
X_4761_ net1578 net1615 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q
+ _0312_ VPWR VGND sg13g2_mux2_1
X_3712_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q _1741_ _1742_
+ _1744_ _1743_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q Tile_X0Y1_DSP_bot.C3
+ VPWR VGND sg13g2_mux4_1
X_4692_ _0075_ net1676 _0246_ VPWR VGND sg13g2_nor2_1
X_3643_ _1680_ net1709 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q
+ VPWR VGND sg13g2_nand2b_1
X_5313_ net1968 net1723 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_3574_ VGND VPWR _1614_ _1615_ Tile_X0Y1_DSP_bot.C9 net1637 sg13g2_a21oi_2
XFILLER_53_0 VPWR VGND sg13g2_decap_4
X_6293_ net155 net514 VPWR VGND sg13g2_buf_1
X_2525_ VPWR _0612_ _0611_ VGND sg13g2_inv_1
X_5244_ net1957 net1745 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_5175_ net1956 net1777 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_4126_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q net1588 _0969_
+ _1011_ _1922_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q _2103_
+ VPWR VGND sg13g2_mux4_1
X_4057_ _2056_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[18\] net1655 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ VPWR VGND sg13g2_mux2_2
X_3008_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q _1070_ _1071_
+ VPWR VGND sg13g2_nor2_1
X_5438__560 VPWR VGND net560 sg13g2_tiehi
XFILLER_51_174 VPWR VGND sg13g2_decap_8
XFILLER_51_185 VPWR VGND sg13g2_fill_2
X_4959_ VGND VPWR _0062_ net1696 _0502_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q
+ sg13g2_a21oi_1
XFILLER_10_53 VPWR VGND sg13g2_fill_2
XFILLER_105_121 VPWR VGND sg13g2_fill_1
Xoutput380 net380 Tile_X0Y1_E2BEG[2] VPWR VGND sg13g2_buf_1
Xoutput391 net391 Tile_X0Y1_E2BEGb[5] VPWR VGND sg13g2_buf_1
XFILLER_19_138 VPWR VGND sg13g2_fill_2
XFILLER_27_171 VPWR VGND sg13g2_fill_2
X_3290_ _1341_ _1340_ _1339_ _1342_ VPWR VGND sg13g2_a21o_1
Xfanout1550 net1551 net1550 VPWR VGND sg13g2_buf_8
Xfanout1561 net1561 _0172_ VPWR VGND sg13g2_buf_16
Xfanout1572 net1573 net1572 VPWR VGND sg13g2_buf_1
Xfanout1583 net1583 net1584 VPWR VGND sg13g2_buf_16
Xfanout1594 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 net1594 VPWR VGND
+ sg13g2_buf_1
X_5470__602 VPWR VGND net602 sg13g2_tiehi
XFILLER_33_130 VPWR VGND sg13g2_fill_1
X_5862_ net1897 net1826 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_5793_ net1862 net1714 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_336 VPWR VGND sg13g2_fill_2
X_4813_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q net132 net59
+ net155 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q
+ _0362_ VPWR VGND sg13g2_mux4_1
X_4744_ VGND VPWR _0295_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q
+ _0294_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q _0296_ _0293_
+ sg13g2_a221oi_1
X_4675_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 net722 VGND sg13g2_inv_1
X_3626_ _1664_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q
+ VPWR VGND sg13g2_nand2b_1
X_3557_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q VPWR _1600_ VGND
+ _0095_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q sg13g2_o21ai_1
X_6276_ Tile_X0Y0_SS4END[15] net503 VPWR VGND sg13g2_buf_1
X_2508_ VPWR _0596_ net643 VGND sg13g2_inv_1
Xinput108 Tile_X0Y1_EE4END[1] net108 VPWR VGND sg13g2_buf_1
X_5227_ net1989 net1756 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_3488_ VGND VPWR net1638 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X
+ _1535_ _1534_ sg13g2_a21oi_1
Xinput119 Tile_X0Y1_N2END[4] net119 VPWR VGND sg13g2_buf_1
X_5158_ net1980 net1778 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_211 VPWR VGND sg13g2_fill_1
XFILLER_56_222 VPWR VGND sg13g2_fill_2
X_5089_ net1967 net1798 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_110_190 VPWR VGND sg13g2_decap_8
X_4109_ net1672 net2002 _2098_ VPWR VGND sg13g2_nor2b_1
XFILLER_16_108 VPWR VGND sg13g2_fill_2
XFILLER_97_23 VPWR VGND sg13g2_fill_2
XFILLER_97_56 VPWR VGND sg13g2_fill_2
XFILLER_79_347 VPWR VGND sg13g2_fill_1
XFILLER_47_288 VPWR VGND sg13g2_fill_1
XFILLER_62_214 VPWR VGND sg13g2_decap_4
XFILLER_62_247 VPWR VGND sg13g2_fill_2
XFILLER_62_269 VPWR VGND sg13g2_fill_2
X_2790_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q _0114_
+ _0864_ _0861_ _0865_ _0862_ sg13g2_a221oi_1
X_4460_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q net1543 net1551
+ net1558 net1564 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q _2375_
+ VPWR VGND sg13g2_mux4_1
X_4391_ _2315_ _2314_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q
+ _2316_ VPWR VGND sg13g2_mux2_1
X_3411_ _1462_ _1171_ _1463_ VPWR VGND sg13g2_xor2_1
X_6130_ Tile_X0Y0_W6END[7] net353 VPWR VGND sg13g2_buf_1
X_5428__570 VPWR VGND net570 sg13g2_tiehi
X_3342_ _1394_ _1392_ _1393_ VPWR VGND sg13g2_nand2b_1
X_6061_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 net282 VPWR VGND sg13g2_buf_1
X_3273_ VGND VPWR _0131_ _0347_ _1326_ _1325_ sg13g2_a21oi_1
X_5012_ _0550_ _0551_ _0552_ VPWR VGND sg13g2_nor2_2
XFILLER_97_177 VPWR VGND sg13g2_fill_2
XFILLER_16_0 VPWR VGND sg13g2_fill_2
XFILLER_53_203 VPWR VGND sg13g2_fill_1
X_5845_ net1901 net1832 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_5435__563 VPWR VGND net563 sg13g2_tiehi
XFILLER_21_133 VPWR VGND sg13g2_fill_1
X_5776_ net1889 net1717 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_2988_ _0772_ _1050_ _1051_ VPWR VGND sg13g2_nor2_1
X_4727_ net67 net1929 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q
+ _0280_ VPWR VGND sg13g2_mux2_1
X_4658_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q VPWR _0214_ VGND
+ net1699 _0175_ sg13g2_o21ai_1
Xinput90 Tile_X0Y1_E1END[3] net90 VPWR VGND sg13g2_buf_1
X_3609_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q VPWR _1648_ VGND
+ _1621_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q sg13g2_o21ai_1
X_4589_ VPWR _0146_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q VGND
+ sg13g2_inv_1
X_6328_ Tile_X0Y1_WW4END[15] net540 VPWR VGND sg13g2_buf_1
X_6259_ Tile_X0Y0_S4END[14] net486 VPWR VGND sg13g2_buf_1
X_5442__556 VPWR VGND net556 sg13g2_tiehi
XFILLER_91_309 VPWR VGND sg13g2_fill_1
XFILLER_120_0 VPWR VGND sg13g2_fill_2
XFILLER_113_208 VPWR VGND sg13g2_fill_2
XFILLER_67_317 VPWR VGND sg13g2_fill_2
XFILLER_67_328 VPWR VGND sg13g2_fill_1
XFILLER_67_339 VPWR VGND sg13g2_fill_1
XFILLER_94_125 VPWR VGND sg13g2_decap_8
XFILLER_75_350 VPWR VGND sg13g2_fill_1
X_3960_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q _1968_
+ _1969_ _0122_ sg13g2_a21oi_1
X_2911_ _0977_ VPWR _0978_ VGND _0976_ _0102_ sg13g2_o21ai_1
XFILLER_43_291 VPWR VGND sg13g2_fill_2
X_3891_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q net1599 net1612
+ net1605 net1625 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q _1905_
+ VPWR VGND sg13g2_mux4_1
X_5630_ net1856 net1771 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_2842_ net109 net1923 net1667 _0914_ VPWR VGND sg13g2_mux2_1
X_5561_ net1908 net1790 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_2773_ VGND VPWR _0847_ _0848_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q
+ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[7\] sg13g2_a21oi_2
X_5492_ net1899 net1845 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_4512_ VPWR _0069_ net1709 VGND sg13g2_inv_1
X_4443_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q VPWR _2361_ VGND
+ _0170_ _1147_ sg13g2_o21ai_1
X_4374_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q VPWR _2302_
+ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q _2301_ sg13g2_o21ai_1
X_3325_ net714 net1628 _1377_ VPWR VGND sg13g2_and2_1
X_6113_ net69 net334 VPWR VGND sg13g2_buf_1
X_6044_ net1818 net256 VPWR VGND sg13g2_buf_1
X_3256_ _1301_ VPWR _1309_ VGND _1298_ _1302_ sg13g2_o21ai_1
XFILLER_37_18 VPWR VGND sg13g2_fill_2
X_3187_ _1242_ net1575 _1213_ VPWR VGND sg13g2_nand2_1
XFILLER_41_217 VPWR VGND sg13g2_decap_8
X_5828_ net1869 net1837 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_5759_ net1858 net1725 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_5_118 VPWR VGND sg13g2_fill_1
XFILLER_72_331 VPWR VGND sg13g2_fill_2
Xoutput209 net209 Tile_X0Y0_EE4BEG[13] VPWR VGND sg13g2_buf_1
X_5425__573 VPWR VGND net573 sg13g2_tiehi
X_3110_ VGND VPWR _1167_ _1166_ _1038_ sg13g2_or2_1
X_4090_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q net1592 _0699_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 _0721_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 VPWR VGND sg13g2_mux4_1
X_3041_ _1101_ net1641 Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[1\] VPWR VGND sg13g2_nand2_1
X_4992_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q VPWR _0533_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q _0530_ sg13g2_o21ai_1
X_3943_ _1952_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[16\] net1656 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ VPWR VGND sg13g2_mux2_1
X_3874_ _1893_ _1824_ _1825_ VPWR VGND sg13g2_xnor2_1
X_5432__566 VPWR VGND net566 sg13g2_tiehi
X_5613_ net1882 net1772 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_2825_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X
+ _0897_ VGND sg13g2_inv_1
X_5544_ net1870 net1793 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_2756_ VGND VPWR net54 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q
+ _0832_ _0831_ sg13g2_a21oi_1
X_2687_ VPWR Tile_X0Y1_DSP_bot.B3 _0766_ VGND sg13g2_inv_1
X_5475_ Tile_X0Y1_UserCLK net607 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X
+ _0031_ _5475_/Q VPWR VGND sg13g2_dfrbp_1
X_4426_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q _1277_ _2346_
+ VPWR VGND sg13g2_nor2_1
X_4357_ _2286_ VPWR _2287_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q
+ net1573 sg13g2_o21ai_1
XFILLER_98_272 VPWR VGND sg13g2_fill_2
X_4288_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q _2233_
+ _2235_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q sg13g2_a21oi_1
X_3308_ _1360_ _1355_ _1359_ VPWR VGND sg13g2_xnor2_1
X_6027_ net1961 net240 VPWR VGND sg13g2_buf_1
XFILLER_58_158 VPWR VGND sg13g2_decap_4
X_3239_ VGND VPWR _1292_ _1291_ _1284_ sg13g2_or2_1
XFILLER_100_277 VPWR VGND sg13g2_decap_8
XFILLER_39_383 VPWR VGND sg13g2_fill_2
XFILLER_64_38 VPWR VGND sg13g2_fill_1
XFILLER_13_97 VPWR VGND sg13g2_fill_2
XFILLER_89_57 VPWR VGND sg13g2_fill_2
Xfanout1902 net1903 net1902 VPWR VGND sg13g2_buf_1
Xfanout1924 Tile_X0Y1_E6END[0] net1924 VPWR VGND sg13g2_buf_1
Xfanout1913 net1914 net1913 VPWR VGND sg13g2_buf_1
Xfanout1968 Tile_X0Y0_FrameData[24] net1968 VPWR VGND sg13g2_buf_1
Xfanout1935 net40 net1935 VPWR VGND sg13g2_buf_1
Xfanout1946 Tile_X0Y0_FrameData[5] net1946 VPWR VGND sg13g2_buf_1
Xfanout1957 Tile_X0Y0_FrameData[29] net1957 VPWR VGND sg13g2_buf_1
Xfanout1979 net1980 net1979 VPWR VGND sg13g2_buf_1
XFILLER_72_161 VPWR VGND sg13g2_decap_4
X_3590_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q net1532 net1536
+ net1546 net1553 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q _1631_
+ VPWR VGND sg13g2_mux4_1
X_2610_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q net1531 net1537
+ net1545 net1552 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q _0694_
+ VPWR VGND sg13g2_mux4_1
X_2541_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 _0627_ VPWR VGND sg13g2_inv_8
X_2472_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q net169 _0562_
+ VPWR VGND sg13g2_nor2b_1
X_5260_ net1992 net1740 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_4211_ VGND VPWR _0061_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q
+ _2176_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q sg13g2_a21oi_1
X_5191_ net1982 net1766 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_4142_ _0156_ VPWR _2117_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q
+ net1519 sg13g2_o21ai_1
X_4073_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q VPWR _2070_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q _2067_ sg13g2_o21ai_1
X_3024_ VGND VPWR _1082_ _1086_ _1085_ _0126_ sg13g2_a21oi_2
XFILLER_55_139 VPWR VGND sg13g2_fill_2
XFILLER_63_150 VPWR VGND sg13g2_fill_2
X_4975_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X
+ _0516_ VGND sg13g2_inv_1
X_3926_ _1936_ VPWR _1937_ VGND _0121_ _1934_ sg13g2_o21ai_1
X_3857_ _1883_ _1808_ _1807_ VPWR VGND sg13g2_xnor2_1
X_3788_ _1817_ _1728_ _1730_ VPWR VGND sg13g2_xnor2_1
X_2808_ _0881_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q _0882_
+ VPWR VGND sg13g2_nor2b_1
X_5527_ net1904 net1804 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_2739_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q VPWR _0816_ VGND
+ _0809_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q sg13g2_o21ai_1
Xoutput540 net540 Tile_X0Y1_WW4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput551 net551 Tile_X0Y1_WW4BEG[7] VPWR VGND sg13g2_buf_1
X_5458_ Tile_X0Y1_UserCLK net590 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X
+ _5458_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[6\] VPWR VGND sg13g2_dfrbp_1
X_4409_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q _2330_ _2331_
+ VPWR VGND sg13g2_nor2_1
X_5389_ net1993 net1831 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_75_59 VPWR VGND sg13g2_fill_2
XFILLER_61_109 VPWR VGND sg13g2_decap_4
XFILLER_10_231 VPWR VGND sg13g2_fill_1
XFILLER_6_246 VPWR VGND sg13g2_fill_2
XFILLER_6_279 VPWR VGND sg13g2_fill_2
XFILLER_108_163 VPWR VGND sg13g2_fill_1
XFILLER_123_166 VPWR VGND sg13g2_fill_2
Xfanout1710 net114 net1710 VPWR VGND sg13g2_buf_1
Xfanout1721 Tile_X0Y1_FrameStrobe[9] net1721 VPWR VGND sg13g2_buf_1
Xfanout1732 net1733 net1732 VPWR VGND sg13g2_buf_1
Xfanout1776 net1779 net1776 VPWR VGND sg13g2_buf_1
Xfanout1754 net1755 net1754 VPWR VGND sg13g2_buf_1
Xfanout1765 net1768 net1765 VPWR VGND sg13g2_buf_1
Xfanout1743 net1744 net1743 VPWR VGND sg13g2_buf_1
Xfanout1798 net1799 net1798 VPWR VGND sg13g2_buf_1
Xfanout1787 net1788 net1787 VPWR VGND sg13g2_buf_1
XFILLER_65_81 VPWR VGND sg13g2_decap_8
X_4760_ net1561 net1569 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q
+ _0311_ VPWR VGND sg13g2_mux2_1
X_3711_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q net141 net92
+ net1936 net152 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q _1744_
+ VPWR VGND sg13g2_mux4_1
XFILLER_81_91 VPWR VGND sg13g2_fill_2
X_4691_ net68 net84 net1676 _0245_ VPWR VGND sg13g2_mux2_1
X_3642_ _1678_ VPWR _1679_ VGND net159 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q
+ sg13g2_o21ai_1
XFILLER_60_2 VPWR VGND sg13g2_fill_1
X_5312_ net1966 net1723 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_3573_ net1636 VPWR _1614_ VGND net1637 _0007_ sg13g2_o21ai_1
X_6292_ net154 net513 VPWR VGND sg13g2_buf_1
XFILLER_46_0 VPWR VGND sg13g2_fill_2
X_2524_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q net136 net55
+ net69 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q
+ _0611_ VPWR VGND sg13g2_mux4_1
X_5243_ net1953 net1745 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_5174_ net1950 net1777 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_4125_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q net1596 _0699_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 _0721_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 VPWR VGND sg13g2_mux4_1
XFILLER_28_128 VPWR VGND sg13g2_fill_1
X_4056_ _2056_ _1989_ _1988_ VPWR VGND sg13g2_xnor2_1
X_3007_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q _1066_
+ _1070_ _1069_ sg13g2_a21oi_1
XFILLER_36_172 VPWR VGND sg13g2_decap_4
XFILLER_61_17 VPWR VGND sg13g2_decap_4
X_4958_ _0500_ VPWR _0501_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q
+ _0497_ sg13g2_o21ai_1
X_4889_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 _0435_ VPWR VGND sg13g2_inv_8
X_3909_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q net126 net7 net54
+ net68 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q _1922_ VPWR VGND
+ sg13g2_mux4_1
XFILLER_10_43 VPWR VGND sg13g2_fill_1
Xoutput370 net370 Tile_X0Y0_WW4BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_105_155 VPWR VGND sg13g2_fill_1
XFILLER_105_177 VPWR VGND sg13g2_decap_4
XFILLER_120_136 VPWR VGND sg13g2_fill_1
Xoutput381 net381 Tile_X0Y1_E2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput392 net392 Tile_X0Y1_E2BEGb[6] VPWR VGND sg13g2_buf_1
XFILLER_30_315 VPWR VGND sg13g2_fill_2
XFILLER_51_72 VPWR VGND sg13g2_fill_1
XFILLER_32_6 VPWR VGND sg13g2_fill_1
Xfanout1540 net1540 net1541 VPWR VGND sg13g2_buf_16
Xfanout1551 net1551 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 VPWR VGND sg13g2_buf_16
Xfanout1573 net1573 net1574 VPWR VGND sg13g2_buf_16
Xfanout1562 _0172_ net1562 VPWR VGND sg13g2_buf_1
Xfanout1584 net1584 net1589 VPWR VGND sg13g2_buf_16
XFILLER_80_215 VPWR VGND sg13g2_fill_1
X_5861_ net1875 net1823 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_4812_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 _0360_ _0361_ _0357_
+ _0350_ VPWR VGND sg13g2_a22oi_1
X_5792_ net1860 net1715 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_348 VPWR VGND sg13g2_fill_1
X_4743_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q _0180_
+ _0295_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q sg13g2_a21oi_1
XFILLER_119_214 VPWR VGND sg13g2_fill_1
X_4674_ _0221_ VPWR _0230_ VGND _0229_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q
+ sg13g2_o21ai_1
X_3625_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6
+ _1663_ _1662_ sg13g2_a21oi_1
X_3556_ _1598_ VPWR _1599_ VGND net718 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q
+ sg13g2_o21ai_1
X_6275_ Tile_X0Y0_SS4END[14] net502 VPWR VGND sg13g2_buf_1
X_2507_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q _0083_ _0084_
+ _0594_ _0085_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q _0595_
+ VPWR VGND sg13g2_mux4_1
Xinput109 Tile_X0Y1_EE4END[2] net109 VPWR VGND sg13g2_buf_1
X_5226_ net1987 net1756 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_3487_ _0135_ VPWR _1534_ VGND net1638 _0005_ sg13g2_o21ai_1
X_5157_ net1975 net1776 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_5088_ net1965 net1798 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_4108_ VGND VPWR net82 net1672 _2097_ _2096_ sg13g2_a21oi_1
X_4039_ _2043_ net1679 net1932 VPWR VGND sg13g2_nand2b_1
XFILLER_112_23 VPWR VGND sg13g2_decap_4
XFILLER_112_56 VPWR VGND sg13g2_decap_8
XFILLER_21_64 VPWR VGND sg13g2_fill_2
XFILLER_97_46 VPWR VGND sg13g2_fill_2
X_4390_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q net1574 net1580
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 net1618 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q
+ _2315_ VPWR VGND sg13g2_mux4_1
X_3410_ _1458_ _1460_ _1462_ VPWR VGND sg13g2_xor2_1
X_3341_ _1393_ _1366_ _1367_ VPWR VGND sg13g2_xnor2_1
X_3272_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q VPWR _1325_ VGND
+ net166 _0131_ sg13g2_o21ai_1
X_6060_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 net281 VPWR VGND sg13g2_buf_1
XFILLER_38_201 VPWR VGND sg13g2_decap_8
X_5011_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q VPWR _0551_ VGND
+ _0545_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q sg13g2_o21ai_1
X_5844_ net1899 net1824 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_42_19 VPWR VGND sg13g2_fill_1
X_5775_ net1887 net1716 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_2987_ _1050_ _1049_ _1048_ VPWR VGND sg13g2_nand2b_1
X_4726_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q net56
+ _0279_ _0278_ sg13g2_a21oi_1
X_4657_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q net611 net39
+ net13 net74 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q _0213_
+ VPWR VGND sg13g2_mux4_1
Xinput91 Tile_X0Y1_E2END[0] net91 VPWR VGND sg13g2_buf_1
X_3608_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6
+ _1647_ _1646_ sg13g2_a21oi_1
Xinput80 Tile_X0Y0_W2MID[7] net80 VPWR VGND sg13g2_buf_1
X_6327_ Tile_X0Y1_WW4END[14] net539 VPWR VGND sg13g2_buf_1
X_4588_ VPWR _0145_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q VGND
+ sg13g2_inv_1
XFILLER_107_12 VPWR VGND sg13g2_fill_2
XFILLER_107_23 VPWR VGND sg13g2_fill_2
X_3539_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q net1574
+ _1584_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q sg13g2_a21oi_1
X_6258_ Tile_X0Y0_S4END[13] net485 VPWR VGND sg13g2_buf_1
X_6189_ Tile_X0Y1_EE4END[8] net416 VPWR VGND sg13g2_buf_1
X_5209_ net2000 net1766 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_123_44 VPWR VGND sg13g2_fill_2
X_5477__609 VPWR VGND net609 sg13g2_tiehi
XFILLER_8_116 VPWR VGND sg13g2_fill_1
XFILLER_113_0 VPWR VGND sg13g2_fill_2
XFILLER_106_283 VPWR VGND sg13g2_fill_1
X_2910_ _0977_ _0102_ _0975_ VPWR VGND sg13g2_nand2b_1
X_3890_ _1904_ net1649 _0030_ VPWR VGND sg13g2_nand2_1
X_2841_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q _0912_ _0907_
+ _0913_ VPWR VGND sg13g2_nand3_1
X_5560_ net1906 net1790 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_2772_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q _0846_ _0847_
+ VPWR VGND sg13g2_nor2_2
X_5491_ net1894 net1848 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_4511_ VPWR _0068_ net41 VGND sg13g2_inv_1
X_4442_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q net1517 _2360_
+ VPWR VGND sg13g2_nor2_1
X_4373_ _2300_ VPWR _2301_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q
+ net1616 sg13g2_o21ai_1
X_3324_ net1608 _1104_ _1375_ _1376_ VPWR VGND sg13g2_nor3_2
X_6112_ net68 net333 VPWR VGND sg13g2_buf_1
X_3255_ VGND VPWR _1308_ net1548 _0703_ sg13g2_or2_1
X_6043_ net1830 net255 VPWR VGND sg13g2_buf_1
X_3186_ _1241_ _1234_ _1235_ VPWR VGND sg13g2_xnor2_1
X_5827_ net1867 net1836 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_5758_ net1856 net1725 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_4709_ net1622 net1630 net1683 _0262_ VPWR VGND sg13g2_mux2_1
XFILLER_118_11 VPWR VGND sg13g2_fill_2
X_5689_ net1908 net1749 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_76_159 VPWR VGND sg13g2_fill_2
XFILLER_27_96 VPWR VGND sg13g2_fill_1
XFILLER_72_354 VPWR VGND sg13g2_fill_2
XFILLER_32_218 VPWR VGND sg13g2_fill_2
XFILLER_25_292 VPWR VGND sg13g2_fill_1
XFILLER_99_218 VPWR VGND sg13g2_fill_1
XFILLER_67_148 VPWR VGND sg13g2_fill_2
X_3040_ Tile_X0Y1_DSP_bot.A1 _1099_ _1100_ _1094_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_48_362 VPWR VGND sg13g2_fill_1
XFILLER_48_384 VPWR VGND sg13g2_fill_1
XFILLER_63_354 VPWR VGND sg13g2_fill_1
X_4991_ _0531_ VPWR _0532_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q
+ net1521 sg13g2_o21ai_1
X_3942_ _1952_ _1950_ _1951_ VPWR VGND sg13g2_xnor2_1
X_3873_ _1892_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[7\] net1654 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ VPWR VGND sg13g2_mux2_1
X_5612_ net1880 net1772 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_2824_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q _0868_ _0870_
+ _0896_ _0894_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q _0897_
+ VPWR VGND sg13g2_mux4_1
X_5543_ net1919 net1801 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_76_0 VPWR VGND sg13g2_fill_2
XFILLER_117_312 VPWR VGND sg13g2_fill_1
X_2755_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q net135 _0831_
+ VPWR VGND sg13g2_nor2b_1
X_2686_ VGND VPWR _0765_ _0766_ _0756_ _0755_ sg13g2_a21oi_2
X_5474_ Tile_X0Y1_UserCLK net606 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X
+ _0029_ _5474_/Q VPWR VGND sg13g2_dfrbp_1
X_4425_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q _1058_
+ _2345_ _2344_ sg13g2_a21oi_1
X_4356_ _2286_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q _1058_
+ VPWR VGND sg13g2_nand2_1
X_3307_ _1357_ _1356_ _1359_ VPWR VGND sg13g2_xor2_1
X_4287_ _0180_ _0176_ net1664 _2234_ VPWR VGND sg13g2_mux2_1
X_6026_ net1963 net239 VPWR VGND sg13g2_buf_1
X_3238_ _1289_ _1288_ _1291_ VPWR VGND sg13g2_xor2_1
X_3169_ _1224_ _1150_ _1223_ VPWR VGND sg13g2_xnor2_1
XFILLER_54_354 VPWR VGND sg13g2_fill_2
XFILLER_66_192 VPWR VGND sg13g2_fill_1
XFILLER_108_378 VPWR VGND sg13g2_fill_2
Xfanout1925 net90 net1925 VPWR VGND sg13g2_buf_1
Xfanout1903 Tile_X0Y1_FrameData[17] net1903 VPWR VGND sg13g2_buf_1
Xfanout1914 Tile_X0Y1_FrameData[12] net1914 VPWR VGND sg13g2_buf_1
Xfanout1936 net39 net1936 VPWR VGND sg13g2_buf_1
Xfanout1947 Tile_X0Y0_FrameData[4] net1947 VPWR VGND sg13g2_buf_1
Xfanout1958 Tile_X0Y0_FrameData[29] net1958 VPWR VGND sg13g2_buf_1
Xfanout1969 Tile_X0Y0_FrameData[23] net1969 VPWR VGND sg13g2_buf_1
XFILLER_57_170 VPWR VGND sg13g2_fill_1
XFILLER_70_60 VPWR VGND sg13g2_fill_1
X_2540_ _0552_ _0626_ _0627_ VPWR VGND sg13g2_nor2b_2
X_2471_ net142 net53 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q _0561_
+ VPWR VGND sg13g2_mux2_1
X_4210_ _2173_ _2175_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 VPWR VGND
+ sg13g2_nor2_2
X_5190_ net1980 net1766 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_95_210 VPWR VGND sg13g2_fill_2
X_4141_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q _2115_
+ _2116_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q sg13g2_a21oi_1
X_4072_ VGND VPWR _0076_ net1694 _2069_ _2068_ sg13g2_a21oi_1
XFILLER_95_265 VPWR VGND sg13g2_fill_2
X_3023_ _1083_ _1084_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q
+ _1085_ VPWR VGND sg13g2_mux2_1
XFILLER_36_376 VPWR VGND sg13g2_fill_1
X_4974_ _0487_ _0515_ _0516_ VPWR VGND sg13g2_nor2_2
X_3925_ _1936_ _0121_ _1935_ VPWR VGND sg13g2_nand2b_1
X_3856_ _1882_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 VGND net1655
+ _1881_ sg13g2_o21ai_1
X_3787_ _1729_ _1730_ _1816_ VPWR VGND sg13g2_nor2_1
X_2807_ _0879_ _0880_ _0881_ VPWR VGND sg13g2_nor2_1
X_5526_ net1903 net1805 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_2738_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q _0813_
+ _0815_ _0814_ sg13g2_a21oi_1
X_5457_ Tile_X0Y1_UserCLK net589 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X
+ _5457_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[5\] VPWR VGND sg13g2_dfrbp_1
Xoutput530 net530 Tile_X0Y1_W6BEG[2] VPWR VGND sg13g2_buf_1
Xoutput541 net541 Tile_X0Y1_WW4BEG[12] VPWR VGND sg13g2_buf_1
X_4408_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q net1713 net1928
+ net147 net1559 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q _2330_
+ VPWR VGND sg13g2_mux4_1
Xoutput552 net552 Tile_X0Y1_WW4BEG[8] VPWR VGND sg13g2_buf_1
X_2669_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q net31 net47 net66
+ net82 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q _0750_ VPWR VGND
+ sg13g2_mux4_1
X_5388_ net1991 net1831 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_4339_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q _2269_ _2271_
+ _2268_ _2270_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A
+ VPWR VGND sg13g2_mux4_1
XFILLER_115_56 VPWR VGND sg13g2_decap_8
XFILLER_86_243 VPWR VGND sg13g2_decap_8
X_6009_ net1938 net252 VPWR VGND sg13g2_buf_1
XFILLER_27_343 VPWR VGND sg13g2_fill_2
XFILLER_24_42 VPWR VGND sg13g2_fill_1
XFILLER_6_225 VPWR VGND sg13g2_fill_2
XFILLER_40_41 VPWR VGND sg13g2_fill_1
XFILLER_108_153 VPWR VGND sg13g2_fill_2
XFILLER_6_0 VPWR VGND sg13g2_fill_2
Xfanout1700 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q net1700 VPWR
+ VGND sg13g2_buf_1
Xfanout1722 net1723 net1722 VPWR VGND sg13g2_buf_1
Xfanout1711 net113 net1711 VPWR VGND sg13g2_buf_1
Xfanout1733 net1734 net1733 VPWR VGND sg13g2_buf_1
X_5461__593 VPWR VGND net593 sg13g2_tiehi
Xfanout1744 Tile_X0Y1_FrameStrobe[7] net1744 VPWR VGND sg13g2_buf_1
Xfanout1755 net1756 net1755 VPWR VGND sg13g2_buf_1
Xfanout1766 net1767 net1766 VPWR VGND sg13g2_buf_1
Xfanout1799 net1800 net1799 VPWR VGND sg13g2_buf_1
Xfanout1788 Tile_X0Y1_FrameStrobe[3] net1788 VPWR VGND sg13g2_buf_1
Xfanout1777 net1779 net1777 VPWR VGND sg13g2_buf_1
XFILLER_18_376 VPWR VGND sg13g2_fill_1
XFILLER_33_313 VPWR VGND sg13g2_fill_1
XFILLER_33_335 VPWR VGND sg13g2_fill_1
X_3710_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q net110 net170
+ net50 _0323_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q _1743_
+ VPWR VGND sg13g2_mux4_1
XFILLER_60_198 VPWR VGND sg13g2_fill_2
X_4690_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q net126 net138
+ net2004 net7 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q _0244_
+ VPWR VGND sg13g2_mux4_1
X_3641_ _1678_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6
+ VPWR VGND sg13g2_nand2b_1
X_3572_ _1610_ _1613_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q
+ Tile_X0Y1_DSP_bot.C9 VPWR VGND sg13g2_mux2_1
X_2523_ _0610_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 VPWR VGND sg13g2_inv_2
X_5311_ net1963 net1719 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_6291_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 net512 VPWR VGND sg13g2_buf_2
X_5242_ net1951 net1745 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_39_0 VPWR VGND sg13g2_fill_2
X_5173_ net1948 net1777 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_4124_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q net1521 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1
+ net1576 _0647_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2
+ VPWR VGND sg13g2_mux4_1
XFILLER_28_107 VPWR VGND sg13g2_decap_8
Xinput1 Tile_X0Y0_E1END[0] net1 VPWR VGND sg13g2_buf_2
XFILLER_83_235 VPWR VGND sg13g2_decap_8
XFILLER_83_246 VPWR VGND sg13g2_fill_1
X_4055_ _2055_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[13\] net1655 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ VPWR VGND sg13g2_mux2_1
X_3006_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q VPWR _1069_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q _1068_ sg13g2_o21ai_1
X_4957_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q _0499_ _0500_
+ VPWR VGND sg13g2_nor2_1
X_4888_ _0424_ _0434_ _0435_ VPWR VGND sg13g2_nor2b_2
X_3908_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2
+ net75 net1935 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q
+ _1921_ VPWR VGND sg13g2_mux4_1
X_3839_ VGND VPWR net1649 _0028_ _1866_ _1865_ sg13g2_a21oi_1
X_5509_ net1874 net1845 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_10_55 VPWR VGND sg13g2_fill_1
XFILLER_10_77 VPWR VGND sg13g2_fill_2
X_5445__577 VPWR VGND net577 sg13g2_tiehi
Xoutput360 net360 Tile_X0Y0_WW4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput371 net371 Tile_X0Y0_WW4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput393 net393 Tile_X0Y1_E2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput382 net382 Tile_X0Y1_E2BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_86_37 VPWR VGND sg13g2_fill_2
XFILLER_27_173 VPWR VGND sg13g2_fill_1
XFILLER_35_96 VPWR VGND sg13g2_fill_1
Xfanout1530 net1530 net1533 VPWR VGND sg13g2_buf_16
Xfanout1541 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 net1541 VPWR VGND
+ sg13g2_buf_8
Xfanout1563 net1563 net1564 VPWR VGND sg13g2_buf_16
Xfanout1574 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 net1574 VPWR VGND sg13g2_buf_8
Xfanout1552 net1553 net1552 VPWR VGND sg13g2_buf_1
Xfanout1596 net1596 net1601 VPWR VGND sg13g2_buf_16
Xfanout1585 net1587 net1585 VPWR VGND sg13g2_buf_1
X_5860_ net1869 net1823 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_4811_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q _0358_
+ _0361_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q sg13g2_a21oi_1
X_5791_ net1859 net1717 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_338 VPWR VGND sg13g2_fill_1
X_4742_ VGND VPWR _0294_ net1529 net1666 sg13g2_or2_1
X_4673_ _0223_ VPWR _0229_ VGND _0225_ _0228_ sg13g2_o21ai_1
X_3624_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6
+ _1662_ VPWR VGND sg13g2_nor2b_1
X_3555_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q _1598_
+ net720 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q sg13g2_a21oi_2
X_6274_ Tile_X0Y0_SS4END[13] net501 VPWR VGND sg13g2_buf_1
X_2506_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 _0594_ VPWR VGND sg13g2_inv_8
X_3486_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X
+ _1532_ _1533_ _1514_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q
+ VPWR VGND sg13g2_a22oi_1
X_5225_ net1986 net1751 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_88_338 VPWR VGND sg13g2_fill_1
XFILLER_102_104 VPWR VGND sg13g2_fill_1
XFILLER_102_159 VPWR VGND sg13g2_decap_4
X_5156_ net1973 net1776 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_202 VPWR VGND sg13g2_decap_8
X_5087_ net1963 net1798 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_224 VPWR VGND sg13g2_fill_1
X_4107_ net1672 net66 _2096_ VPWR VGND sg13g2_nor2b_1
X_4038_ _2041_ VPWR _2042_ VGND _0070_ net1679 sg13g2_o21ai_1
X_5989_ Tile_X0Y0_EE4END[9] net216 VPWR VGND sg13g2_buf_1
XFILLER_12_338 VPWR VGND sg13g2_fill_1
XFILLER_20_371 VPWR VGND sg13g2_fill_2
XFILLER_97_25 VPWR VGND sg13g2_fill_1
Xoutput190 net190 Tile_X0Y0_E2BEGb[5] VPWR VGND sg13g2_buf_1
XFILLER_7_320 VPWR VGND sg13g2_fill_1
X_3340_ _1392_ _1388_ _1391_ VPWR VGND sg13g2_nand2_1
X_5010_ _0548_ _0549_ _0550_ VPWR VGND sg13g2_nor2_1
X_3271_ VGND VPWR _1323_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q
+ _0130_ _1320_ _1324_ _1322_ sg13g2_a221oi_1
XFILLER_16_2 VPWR VGND sg13g2_fill_1
X_5843_ net1895 net1824 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_61_293 VPWR VGND sg13g2_fill_1
XFILLER_21_179 VPWR VGND sg13g2_fill_2
X_5774_ net1885 net1716 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_2986_ _1035_ _1047_ _1031_ _1049_ VPWR VGND sg13g2_nand3_1
X_4725_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q net48 _0278_ VPWR
+ VGND sg13g2_nor2b_1
X_4656_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 _0206_ _0212_ _0204_
+ _0197_ VPWR VGND sg13g2_a22oi_1
X_4587_ VPWR _0144_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q VGND
+ sg13g2_inv_1
X_3607_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6
+ _1646_ VPWR VGND sg13g2_nor2b_1
Xinput70 Tile_X0Y0_W2END[5] net70 VPWR VGND sg13g2_buf_1
Xinput81 Tile_X0Y0_W6END[0] net81 VPWR VGND sg13g2_buf_8
Xinput92 Tile_X0Y1_E2END[1] net92 VPWR VGND sg13g2_buf_1
X_6326_ Tile_X0Y1_WW4END[13] net553 VPWR VGND sg13g2_buf_1
X_3538_ _1583_ _0140_ _1582_ VPWR VGND sg13g2_nand2_1
X_3469_ _1518_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q _1517_
+ VPWR VGND sg13g2_nand2b_1
X_6257_ Tile_X0Y0_S4END[12] net484 VPWR VGND sg13g2_buf_1
X_6188_ Tile_X0Y1_EE4END[7] net415 VPWR VGND sg13g2_buf_1
X_5208_ net1978 net1767 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_29_235 VPWR VGND sg13g2_decap_8
X_5139_ net1943 net1789 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_32_53 VPWR VGND sg13g2_fill_1
XFILLER_120_2 VPWR VGND sg13g2_fill_1
XFILLER_20_190 VPWR VGND sg13g2_fill_2
XFILLER_32_75 VPWR VGND sg13g2_decap_4
XFILLER_106_0 VPWR VGND sg13g2_fill_1
XFILLER_79_102 VPWR VGND sg13g2_fill_2
XFILLER_67_319 VPWR VGND sg13g2_fill_1
XFILLER_57_50 VPWR VGND sg13g2_fill_1
X_2840_ _0909_ _0911_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q
+ _0912_ VPWR VGND sg13g2_nand3_1
X_2771_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X
+ _0846_ VGND sg13g2_inv_1
X_4510_ VPWR _0067_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q VGND
+ sg13g2_inv_1
X_5490_ net1892 net1848 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_4441_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q _1780_
+ _2359_ _2358_ sg13g2_a21oi_1
X_4372_ _2300_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q _1780_
+ VPWR VGND sg13g2_nand2_1
X_6111_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 net332 VPWR VGND sg13g2_buf_1
X_3323_ VPWR _1375_ _1374_ VGND sg13g2_inv_1
X_3254_ _1305_ _1306_ _1307_ VPWR VGND sg13g2_nor2_1
X_6042_ net1844 net254 VPWR VGND sg13g2_buf_1
X_3185_ VPWR _1240_ _1239_ VGND sg13g2_inv_1
XFILLER_93_182 VPWR VGND sg13g2_fill_2
X_5826_ net1864 net1834 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_5757_ net1918 net1724 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_2969_ _1032_ _0770_ _0771_ VPWR VGND sg13g2_xnor2_1
X_4708_ _0260_ VPWR _0261_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q
+ net1596 sg13g2_o21ai_1
X_5688_ net1907 net1749 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_4639_ net1657 net1528 net1542 net1549 net1556 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q
+ _0196_ VPWR VGND sg13g2_mux4_1
X_6309_ Tile_X0Y1_W6END[6] net532 VPWR VGND sg13g2_buf_1
XFILLER_1_326 VPWR VGND sg13g2_fill_2
XFILLER_103_287 VPWR VGND sg13g2_decap_4
XFILLER_17_216 VPWR VGND sg13g2_fill_1
XFILLER_4_197 VPWR VGND sg13g2_fill_2
X_4990_ _0531_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q net1518
+ VPWR VGND sg13g2_nand2b_1
X_3941_ VGND VPWR _1927_ _1951_ _1900_ _1928_ sg13g2_a21oi_2
X_3872_ _1820_ _1821_ _1892_ VPWR VGND sg13g2_xor2_1
X_5611_ net1879 net1774 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_2823_ VPWR _0896_ _0895_ VGND sg13g2_inv_1
X_5542_ net1896 net1801 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_2754_ net1929 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q
+ _0830_ VPWR VGND sg13g2_mux2_1
XFILLER_69_0 VPWR VGND sg13g2_fill_2
X_2685_ _0762_ _0764_ _0765_ VPWR VGND sg13g2_nor2_1
X_5473_ Tile_X0Y1_UserCLK net605 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X
+ _0027_ _5473_/Q VPWR VGND sg13g2_dfrbp_1
X_4424_ net1570 _0169_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q
+ _2344_ VPWR VGND sg13g2_a21o_1
X_4355_ VGND VPWR _2284_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q
+ _2283_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q _2285_ _2282_
+ sg13g2_a221oi_1
X_3306_ _1358_ _1356_ _1357_ VPWR VGND sg13g2_nand2b_1
X_4286_ net1550 net1557 net1663 _2233_ VPWR VGND sg13g2_mux2_1
XFILLER_100_213 VPWR VGND sg13g2_decap_8
X_6025_ net1965 net238 VPWR VGND sg13g2_buf_1
X_3237_ _1290_ _1288_ _1289_ VPWR VGND sg13g2_nand2b_1
X_3168_ _1223_ _1006_ net1511 VPWR VGND sg13g2_nand2b_1
XFILLER_104_58 VPWR VGND sg13g2_fill_1
XFILLER_104_69 VPWR VGND sg13g2_fill_2
X_3099_ _1113_ _1155_ _1156_ VPWR VGND sg13g2_nor2b_1
X_5809_ net1891 net1836 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_13_99 VPWR VGND sg13g2_fill_1
XFILLER_89_59 VPWR VGND sg13g2_fill_1
Xfanout1904 Tile_X0Y1_FrameData[16] net1904 VPWR VGND sg13g2_buf_1
Xfanout1915 net1916 net1915 VPWR VGND sg13g2_buf_1
Xfanout1926 net89 net1926 VPWR VGND sg13g2_buf_1
XFILLER_49_138 VPWR VGND sg13g2_fill_1
Xfanout1959 Tile_X0Y0_FrameData[28] net1959 VPWR VGND sg13g2_buf_1
Xfanout1948 Tile_X0Y0_FrameData[4] net1948 VPWR VGND sg13g2_buf_1
Xfanout1937 net1938 net1937 VPWR VGND sg13g2_buf_1
XFILLER_54_40 VPWR VGND sg13g2_fill_1
XFILLER_62_7 VPWR VGND sg13g2_decap_4
X_2470_ VGND VPWR _0556_ _0559_ _0560_ _0109_ sg13g2_a21oi_1
XFILLER_114_349 VPWR VGND sg13g2_fill_2
X_4140_ net62 net1634 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q
+ _2115_ VPWR VGND sg13g2_mux2_1
X_4071_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q VPWR _2068_ VGND
+ net1693 net66 sg13g2_o21ai_1
X_3022_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q net1924 net153
+ net1935 net172 net1665 _1084_ VPWR VGND sg13g2_mux4_1
XFILLER_48_160 VPWR VGND sg13g2_decap_8
XFILLER_95_80 VPWR VGND sg13g2_fill_2
XFILLER_51_314 VPWR VGND sg13g2_fill_2
XFILLER_51_336 VPWR VGND sg13g2_fill_2
XFILLER_63_196 VPWR VGND sg13g2_fill_2
X_4973_ _0514_ _0512_ _0515_ VPWR VGND sg13g2_nor2_2
X_3924_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q net144 net35
+ net9 net70 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q _1935_ VPWR
+ VGND sg13g2_mux4_1
X_3855_ _1882_ net1655 Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[14\] VPWR VGND sg13g2_nand2_1
X_3786_ VGND VPWR _1740_ _1815_ _1813_ _1814_ sg13g2_a21oi_2
X_2806_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q VPWR _0880_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q _0877_ sg13g2_o21ai_1
X_5525_ net1900 net1805 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_2737_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q VPWR _0814_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q _0811_ sg13g2_o21ai_1
Xoutput520 net520 Tile_X0Y1_W2BEGb[2] VPWR VGND sg13g2_buf_1
X_5456_ Tile_X0Y1_UserCLK net588 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X
+ _5456_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[4\] VPWR VGND sg13g2_dfrbp_1
X_2668_ _0749_ _0748_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q
+ VPWR VGND sg13g2_nand2b_1
X_4407_ _2329_ _2328_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 VPWR VGND sg13g2_mux2_1
Xoutput553 net553 Tile_X0Y1_WW4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput542 net542 Tile_X0Y1_WW4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput531 net531 Tile_X0Y1_W6BEG[3] VPWR VGND sg13g2_buf_1
X_2599_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q _0095_
+ _0683_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q sg13g2_a21oi_1
X_5387_ net1990 net1829 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_4338_ net1581 _0905_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q
+ _2271_ VPWR VGND sg13g2_mux2_1
XFILLER_86_200 VPWR VGND sg13g2_fill_1
X_4269_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q VPWR _2227_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q _2226_ sg13g2_o21ai_1
XFILLER_75_17 VPWR VGND sg13g2_fill_2
XFILLER_27_300 VPWR VGND sg13g2_fill_1
XFILLER_46_119 VPWR VGND sg13g2_fill_1
X_6008_ net1940 net251 VPWR VGND sg13g2_buf_1
XFILLER_24_87 VPWR VGND sg13g2_fill_2
XFILLER_40_75 VPWR VGND sg13g2_decap_8
XFILLER_123_113 VPWR VGND sg13g2_fill_2
Xfanout1723 Tile_X0Y1_FrameStrobe[9] net1723 VPWR VGND sg13g2_buf_1
Xfanout1701 net1702 net1701 VPWR VGND sg13g2_buf_1
Xfanout1712 net112 net1712 VPWR VGND sg13g2_buf_1
XFILLER_77_222 VPWR VGND sg13g2_decap_8
Xfanout1734 Tile_X0Y1_FrameStrobe[8] net1734 VPWR VGND sg13g2_buf_1
Xfanout1745 Tile_X0Y1_FrameStrobe[7] net1745 VPWR VGND sg13g2_buf_1
Xfanout1756 net1757 net1756 VPWR VGND sg13g2_buf_1
Xfanout1767 net1768 net1767 VPWR VGND sg13g2_buf_1
Xfanout1778 net1779 net1778 VPWR VGND sg13g2_buf_1
Xfanout1789 Tile_X0Y1_FrameStrobe[3] net1789 VPWR VGND sg13g2_buf_1
XFILLER_92_269 VPWR VGND sg13g2_decap_4
X_3640_ _1677_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q _1676_
+ VPWR VGND sg13g2_nand2_1
X_3571_ _1613_ _1612_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q
+ _1611_ _1609_ VPWR VGND sg13g2_a22oi_1
XFILLER_114_102 VPWR VGND sg13g2_fill_1
X_6290_ net646 net511 VPWR VGND sg13g2_buf_1
X_2522_ VGND VPWR _0609_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 _0560_
+ _0554_ sg13g2_a21oi_2
X_5310_ net1962 net1719 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_5241_ net2000 net1755 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_5172_ net1946 net1777 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_4123_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q net1583 _0614_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 _0611_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 VPWR VGND sg13g2_mux4_1
Xinput2 Tile_X0Y0_E1END[1] net2 VPWR VGND sg13g2_buf_1
X_4054_ _2055_ _1834_ _1832_ VPWR VGND sg13g2_xnor2_1
X_3005_ VGND VPWR _0066_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q
+ _1068_ _1067_ sg13g2_a21oi_1
X_4956_ VGND VPWR _0059_ net1696 _0499_ _0498_ sg13g2_a21oi_1
X_4887_ _0428_ _0433_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q
+ _0434_ VPWR VGND sg13g2_nand3_1
X_3907_ _1920_ _1909_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 VPWR VGND
+ sg13g2_nor2_2
X_3838_ VGND VPWR net1638 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X
+ _1865_ _1864_ sg13g2_a21oi_1
X_5508_ net1869 net1845 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_3769_ VGND VPWR _1798_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q
+ _1797_ _1796_ _1799_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q
+ sg13g2_a221oi_1
X_5439_ Tile_X0Y1_UserCLK net559 _0053_ _0030_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[15\]
+ VPWR VGND sg13g2_dfrbp_1
Xoutput361 net361 Tile_X0Y0_WW4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput350 net350 Tile_X0Y0_W6BEG[2] VPWR VGND sg13g2_buf_1
Xoutput394 net394 Tile_X0Y1_E6BEG[0] VPWR VGND sg13g2_buf_1
Xoutput383 net383 Tile_X0Y1_E2BEG[5] VPWR VGND sg13g2_buf_1
Xoutput372 net372 Tile_X0Y0_WW4BEG[8] VPWR VGND sg13g2_buf_1
XFILLER_35_20 VPWR VGND sg13g2_fill_1
XFILLER_42_111 VPWR VGND sg13g2_decap_8
XFILLER_27_196 VPWR VGND sg13g2_decap_8
XFILLER_35_53 VPWR VGND sg13g2_fill_2
XFILLER_30_317 VPWR VGND sg13g2_fill_1
Xfanout1542 net1544 net1542 VPWR VGND sg13g2_buf_1
Xfanout1531 net1531 net1532 VPWR VGND sg13g2_buf_16
Xfanout1520 net1520 net726 VPWR VGND sg13g2_buf_16
Xfanout1553 net1554 net1553 VPWR VGND sg13g2_buf_1
Xfanout1564 net1564 net1567 VPWR VGND sg13g2_buf_16
Xfanout1575 _0973_ net1575 VPWR VGND sg13g2_buf_1
Xfanout1597 net1598 net1597 VPWR VGND sg13g2_buf_1
Xfanout1586 net1587 net1586 VPWR VGND sg13g2_buf_1
XFILLER_18_141 VPWR VGND sg13g2_fill_1
X_4810_ _0360_ _0359_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q
+ VPWR VGND sg13g2_nand2b_1
X_5790_ net1857 net1717 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_33_155 VPWR VGND sg13g2_decap_4
X_4741_ net1550 net1559 net1666 _0293_ VPWR VGND sg13g2_mux2_1
X_4672_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q VPWR _0228_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q _0227_ sg13g2_o21ai_1
X_3623_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 _1659_ _1661_ _1657_
+ _1651_ VPWR VGND sg13g2_a22oi_1
X_3554_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q _1595_ _1597_
+ _1594_ _1596_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7
+ VPWR VGND sg13g2_mux4_1
XFILLER_51_0 VPWR VGND sg13g2_fill_2
X_2505_ _0584_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q _0593_
+ _0594_ VPWR VGND sg13g2_a21o_2
X_6273_ Tile_X0Y0_SS4END[12] net500 VPWR VGND sg13g2_buf_1
X_3485_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q _0614_
+ _1533_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q sg13g2_a21oi_1
X_5224_ net1984 net1752 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_5155_ net1972 net1776 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_19 VPWR VGND sg13g2_fill_2
X_5086_ net1961 net1798 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_4106_ VGND VPWR net55 net1672 _2095_ _2094_ sg13g2_a21oi_1
X_4037_ VGND VPWR net30 net1679 _2041_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q
+ sg13g2_a21oi_1
XFILLER_112_47 VPWR VGND sg13g2_decap_4
X_5988_ Tile_X0Y0_EE4END[8] net215 VPWR VGND sg13g2_buf_1
X_4939_ _0482_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q net13 VPWR
+ VGND sg13g2_nand2b_1
XFILLER_21_66 VPWR VGND sg13g2_fill_1
Xoutput180 net180 Tile_X0Y0_E2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput191 net191 Tile_X0Y0_E2BEGb[6] VPWR VGND sg13g2_buf_1
XFILLER_62_239 VPWR VGND sg13g2_decap_4
XFILLER_30_147 VPWR VGND sg13g2_fill_2
XFILLER_7_310 VPWR VGND sg13g2_fill_1
XFILLER_116_219 VPWR VGND sg13g2_fill_1
X_3270_ net105 net624 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q
+ _1323_ VPWR VGND sg13g2_mux2_1
XFILLER_97_147 VPWR VGND sg13g2_decap_4
XFILLER_38_214 VPWR VGND sg13g2_fill_2
XFILLER_38_258 VPWR VGND sg13g2_fill_2
XFILLER_53_228 VPWR VGND sg13g2_decap_8
X_5842_ net1893 net1824 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_5773_ net1883 net1716 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_2985_ VGND VPWR _1047_ _1048_ _1035_ _1031_ sg13g2_a21oi_2
X_4724_ VGND VPWR _0274_ _0064_ _0276_ _0063_ _0277_ _0272_ sg13g2_a221oi_1
X_4655_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q _0211_ _0212_
+ VPWR VGND sg13g2_nor2_1
Xinput60 Tile_X0Y0_SS4END[6] net60 VPWR VGND sg13g2_buf_1
X_3606_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 _1644_ _1645_ _1637_ _1635_
+ VPWR VGND sg13g2_a22oi_1
X_4586_ VPWR _0143_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q VGND
+ sg13g2_inv_1
Xinput71 Tile_X0Y0_W2END[6] net71 VPWR VGND sg13g2_buf_1
Xinput82 Tile_X0Y0_W6END[1] net82 VPWR VGND sg13g2_buf_1
Xinput93 Tile_X0Y1_E2END[2] net93 VPWR VGND sg13g2_buf_1
X_6325_ Tile_X0Y1_WW4END[12] net552 VPWR VGND sg13g2_buf_1
X_3537_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q net1531 net1537
+ net1545 net1552 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q _1582_
+ VPWR VGND sg13g2_mux4_1
XFILLER_107_14 VPWR VGND sg13g2_fill_1
XFILLER_107_25 VPWR VGND sg13g2_fill_1
X_3468_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q net1632 net1585
+ net1525 net1520 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q _1517_
+ VPWR VGND sg13g2_mux4_1
X_6256_ Tile_X0Y0_S4END[11] net483 VPWR VGND sg13g2_buf_1
X_6187_ Tile_X0Y1_EE4END[6] net414 VPWR VGND sg13g2_buf_1
X_3399_ VGND VPWR _1370_ _1451_ _1450_ _1449_ sg13g2_a21oi_2
X_5207_ net1955 net1764 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_5138_ net1941 net1789 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_123_46 VPWR VGND sg13g2_fill_1
XFILLER_96_191 VPWR VGND sg13g2_fill_1
X_5069_ net1993 net1806 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_16_88 VPWR VGND sg13g2_fill_2
X_2770_ VGND VPWR _0837_ _0846_ _0845_ _0844_ sg13g2_a21oi_2
X_4440_ _0178_ _0170_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q
+ _2358_ VPWR VGND sg13g2_a21o_1
X_4371_ _2298_ VPWR _2299_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q
+ net1517 sg13g2_o21ai_1
X_6110_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 net331 VPWR VGND sg13g2_buf_1
X_3322_ net1511 _1214_ _1374_ VPWR VGND sg13g2_nor2_1
X_6041_ net1722 net272 VPWR VGND sg13g2_buf_1
X_3253_ _1306_ _1252_ _1253_ VPWR VGND sg13g2_xnor2_1
X_3184_ _1239_ _1234_ _1235_ _1237_ VPWR VGND sg13g2_and3_1
XFILLER_85_139 VPWR VGND sg13g2_fill_1
XFILLER_14_0 VPWR VGND sg13g2_fill_1
XFILLER_34_261 VPWR VGND sg13g2_fill_1
X_5825_ net1863 net1836 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_34_272 VPWR VGND sg13g2_fill_2
X_5756_ net1916 net1724 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_2968_ _1030_ VPWR _1031_ VGND _1010_ _0933_ sg13g2_o21ai_1
X_5687_ net1904 net1748 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_4707_ _0260_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q net1609
+ VPWR VGND sg13g2_nand2b_1
X_4638_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q net25 net84 net46
+ _0194_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q _0195_ VPWR
+ VGND sg13g2_mux4_1
X_2899_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2
+ net75 net14 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q
+ _0967_ VPWR VGND sg13g2_mux4_1
XFILLER_118_57 VPWR VGND sg13g2_fill_2
X_4569_ VPWR _0126_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q VGND
+ sg13g2_inv_1
X_6308_ Tile_X0Y1_W6END[5] net531 VPWR VGND sg13g2_buf_1
XFILLER_103_222 VPWR VGND sg13g2_decap_4
X_6239_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 net460 VPWR VGND sg13g2_buf_1
XFILLER_103_244 VPWR VGND sg13g2_decap_8
XFILLER_103_255 VPWR VGND sg13g2_fill_1
XFILLER_69_180 VPWR VGND sg13g2_fill_2
XFILLER_103_299 VPWR VGND sg13g2_fill_2
XFILLER_94_49 VPWR VGND sg13g2_fill_1
XFILLER_68_50 VPWR VGND sg13g2_decap_4
X_3940_ _1950_ _1949_ _1948_ VPWR VGND sg13g2_nand2b_1
X_3871_ _1891_ VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 VGND net1653 _1890_
+ sg13g2_o21ai_1
X_5610_ net1877 net1774 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_2822_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q net127 net8 net56
+ net69 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q _0895_ VPWR VGND
+ sg13g2_mux4_1
X_5541_ net1874 net1801 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_76_2 VPWR VGND sg13g2_fill_1
X_2753_ _0829_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 VGND _0816_
+ _0815_ sg13g2_o21ai_1
X_2684_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q VPWR _0764_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q _0763_ sg13g2_o21ai_1
X_5472_ Tile_X0Y1_UserCLK net604 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X
+ _0001_ _5472_/Q VPWR VGND sg13g2_dfrbp_1
X_4423_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q _2342_ _2343_
+ VPWR VGND sg13g2_nor2_1
X_4354_ VGND VPWR _0073_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q
+ _2284_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q sg13g2_a21oi_1
X_3305_ _1357_ _0702_ net1568 VPWR VGND sg13g2_nand2_1
XFILLER_98_264 VPWR VGND sg13g2_fill_2
X_6024_ net1967 net237 VPWR VGND sg13g2_buf_1
X_4285_ _2229_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q _2231_
+ _2232_ VPWR VGND sg13g2_a21o_1
X_3236_ _1232_ _1231_ _1289_ VPWR VGND sg13g2_xor2_1
XFILLER_39_375 VPWR VGND sg13g2_fill_2
X_3167_ _1222_ _1006_ net1608 VPWR VGND sg13g2_nand2b_1
XFILLER_66_172 VPWR VGND sg13g2_fill_2
X_3098_ _1155_ _1149_ _1153_ VPWR VGND sg13g2_xnor2_1
XFILLER_54_356 VPWR VGND sg13g2_fill_1
X_5808_ net1889 net1838 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_5739_ net1878 net1724 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_13_78 VPWR VGND sg13g2_fill_2
Xfanout1905 Tile_X0Y1_FrameData[16] net1905 VPWR VGND sg13g2_buf_1
Xfanout1916 Tile_X0Y1_FrameData[11] net1916 VPWR VGND sg13g2_buf_1
XFILLER_1_168 VPWR VGND sg13g2_fill_1
Xfanout1927 net88 net1927 VPWR VGND sg13g2_buf_1
Xfanout1949 net1950 net1949 VPWR VGND sg13g2_buf_1
Xfanout1938 Tile_X0Y0_FrameData[9] net1938 VPWR VGND sg13g2_buf_1
XFILLER_57_161 VPWR VGND sg13g2_decap_4
XFILLER_45_367 VPWR VGND sg13g2_fill_1
XFILLER_72_186 VPWR VGND sg13g2_decap_4
XFILLER_122_361 VPWR VGND sg13g2_fill_1
X_4070_ _2066_ VPWR _2067_ VGND net1694 net31 sg13g2_o21ai_1
X_3021_ net1665 net1713 net117 net133 net93 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q
+ _1083_ VPWR VGND sg13g2_mux4_1
XFILLER_95_267 VPWR VGND sg13g2_fill_1
X_4972_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q VPWR _0514_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q _0513_ sg13g2_o21ai_1
X_3923_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q net21 net47 net86
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q
+ _1934_ VPWR VGND sg13g2_mux4_1
X_3854_ _1881_ _1835_ _1880_ VPWR VGND sg13g2_xnor2_1
X_2805_ VGND VPWR net1688 net699 _0879_ _0878_ sg13g2_a21oi_1
XFILLER_81_0 VPWR VGND sg13g2_fill_2
X_3785_ _1739_ _1732_ _1814_ VPWR VGND sg13g2_xor2_1
X_5524_ net1898 net1805 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_2736_ _0812_ VPWR _0813_ VGND net1698 _0175_ sg13g2_o21ai_1
Xoutput510 net510 Tile_X0Y1_W2BEG[0] VPWR VGND sg13g2_buf_1
X_5455_ Tile_X0Y1_UserCLK net587 Tile_X0Y1_DSP_bot.B3 _5455_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[3\]
+ VPWR VGND sg13g2_dfrbp_1
X_2667_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q net144 net2002
+ net5 net21 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q _0748_ VPWR
+ VGND sg13g2_mux4_1
X_4406_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q net1710 net90
+ net1704 net1550 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q _2329_
+ VPWR VGND sg13g2_mux4_1
Xoutput521 net521 Tile_X0Y1_W2BEGb[3] VPWR VGND sg13g2_buf_1
Xoutput543 net543 Tile_X0Y1_WW4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput532 net532 Tile_X0Y1_W6BEG[4] VPWR VGND sg13g2_buf_1
X_5386_ net1988 net1829 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_2598_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q net1584 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1
+ net1576 _0647_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q _0682_
+ VPWR VGND sg13g2_mux4_1
X_4337_ _1130_ _1772_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q
+ _2270_ VPWR VGND sg13g2_mux2_1
XFILLER_86_223 VPWR VGND sg13g2_fill_2
X_4268_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q net1585 net1522
+ net1520 net1540 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q _2226_
+ VPWR VGND sg13g2_mux4_1
X_3219_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q VPWR _1273_ VGND
+ net161 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q sg13g2_o21ai_1
X_6007_ net1942 net250 VPWR VGND sg13g2_buf_1
X_4199_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q net1584 _0969_
+ _1011_ _1954_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q _2166_
+ VPWR VGND sg13g2_mux4_1
XFILLER_6_2 VPWR VGND sg13g2_fill_1
Xfanout1702 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q net1702 VPWR
+ VGND sg13g2_buf_1
Xfanout1724 net1726 net1724 VPWR VGND sg13g2_buf_1
Xfanout1713 net111 net1713 VPWR VGND sg13g2_buf_1
Xfanout1746 net1747 net1746 VPWR VGND sg13g2_buf_1
Xfanout1735 net1738 net1735 VPWR VGND sg13g2_buf_1
Xfanout1757 Tile_X0Y1_FrameStrobe[6] net1757 VPWR VGND sg13g2_buf_1
Xfanout1768 Tile_X0Y1_FrameStrobe[5] net1768 VPWR VGND sg13g2_buf_1
XFILLER_77_289 VPWR VGND sg13g2_fill_1
XFILLER_92_204 VPWR VGND sg13g2_fill_2
Xfanout1779 Tile_X0Y1_FrameStrobe[4] net1779 VPWR VGND sg13g2_buf_1
XFILLER_60_101 VPWR VGND sg13g2_decap_8
XFILLER_65_95 VPWR VGND sg13g2_decap_8
X_3570_ VGND VPWR _0137_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 _1612_
+ _1577_ sg13g2_a21oi_1
X_2521_ VGND VPWR _0608_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q
+ _0605_ _0600_ _0609_ _0603_ sg13g2_a221oi_1
XFILLER_53_4 VPWR VGND sg13g2_fill_1
X_5240_ net1978 net1755 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_102_309 VPWR VGND sg13g2_fill_1
XFILLER_39_2 VPWR VGND sg13g2_fill_1
X_5171_ net1944 net1777 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_122_191 VPWR VGND sg13g2_fill_1
X_4122_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q net1592 net701
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 _0385_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 VPWR VGND sg13g2_mux4_1
XFILLER_68_267 VPWR VGND sg13g2_fill_1
X_4053_ _2054_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 VGND net1655
+ _2053_ sg13g2_o21ai_1
X_3004_ net1924 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q _1067_
+ VPWR VGND sg13g2_nor2_1
Xinput3 Tile_X0Y0_E1END[2] net3 VPWR VGND sg13g2_buf_1
XFILLER_36_164 VPWR VGND sg13g2_decap_4
XFILLER_91_270 VPWR VGND sg13g2_decap_8
X_4955_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q VPWR _0498_ VGND
+ net6 net1695 sg13g2_o21ai_1
X_3906_ VGND VPWR _1919_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q
+ _1916_ _1914_ _1920_ _1911_ sg13g2_a221oi_1
X_4886_ _0432_ VPWR _0433_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q
+ _0430_ sg13g2_o21ai_1
X_3837_ net1636 VPWR _1864_ VGND net1639 _0029_ sg13g2_o21ai_1
X_3768_ VGND VPWR net105 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q
+ _1798_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q sg13g2_a21oi_1
X_5507_ net1866 net1846 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_2719_ _0794_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q _0797_
+ _0798_ VPWR VGND sg13g2_a21o_1
X_3699_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q net134 net53
+ net107 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q
+ _1733_ VPWR VGND sg13g2_mux4_1
XFILLER_10_79 VPWR VGND sg13g2_fill_1
Xoutput340 net340 Tile_X0Y0_W2BEGb[2] VPWR VGND sg13g2_buf_1
X_5438_ Tile_X0Y1_UserCLK net560 _0052_ _0028_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[14\]
+ VPWR VGND sg13g2_dfrbp_1
Xoutput362 net362 Tile_X0Y0_WW4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput351 net351 Tile_X0Y0_W6BEG[3] VPWR VGND sg13g2_buf_1
Xoutput384 net384 Tile_X0Y1_E2BEG[6] VPWR VGND sg13g2_buf_1
Xoutput395 net395 Tile_X0Y1_E6BEG[10] VPWR VGND sg13g2_buf_8
Xoutput373 net373 Tile_X0Y0_WW4BEG[9] VPWR VGND sg13g2_buf_1
X_5369_ net2000 net1844 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_86_39 VPWR VGND sg13g2_fill_1
XFILLER_111_117 VPWR VGND sg13g2_fill_2
Xfanout1532 net1532 net1533 VPWR VGND sg13g2_buf_16
Xfanout1521 net1521 net1526 VPWR VGND sg13g2_buf_16
Xfanout1565 net1567 net1565 VPWR VGND sg13g2_buf_1
Xfanout1554 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 net1554 VPWR VGND sg13g2_buf_1
Xfanout1543 net1543 net1544 VPWR VGND sg13g2_buf_16
XFILLER_76_83 VPWR VGND sg13g2_fill_1
Xfanout1576 _0681_ net1576 VPWR VGND sg13g2_buf_8
Xfanout1598 net1601 net1598 VPWR VGND sg13g2_buf_1
Xfanout1587 net1589 net1587 VPWR VGND sg13g2_buf_1
X_4740_ _0291_ VPWR _0292_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q
+ _0176_ sg13g2_o21ai_1
X_4671_ _0226_ VPWR _0227_ VGND _0070_ net1699 sg13g2_o21ai_1
X_3622_ VGND VPWR _0146_ _1660_ _1661_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q
+ sg13g2_a21oi_1
X_3553_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q net1533 net635
+ net1547 net1554 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q _1597_
+ VPWR VGND sg13g2_mux4_1
X_6272_ Tile_X0Y0_SS4END[11] net499 VPWR VGND sg13g2_buf_1
X_2504_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q _0586_ _0592_
+ _0593_ VPWR VGND sg13g2_nor3_1
XFILLER_44_0 VPWR VGND sg13g2_decap_8
X_3484_ _1531_ VPWR _1532_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q
+ _1515_ sg13g2_o21ai_1
X_5223_ net1981 net1754 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_102_117 VPWR VGND sg13g2_fill_2
X_5154_ net1970 net1776 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_4105_ _0075_ net1673 _2094_ VPWR VGND sg13g2_nor2_1
X_5085_ net1959 net1797 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_4036_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q _2039_ _2040_
+ VPWR VGND sg13g2_nor2_1
X_5987_ Tile_X0Y0_EE4END[7] net214 VPWR VGND sg13g2_buf_1
X_4938_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q _0464_ _0480_
+ _0481_ VPWR VGND sg13g2_nor3_1
X_5451__583 VPWR VGND net583 sg13g2_tiehi
X_4869_ _0416_ _0413_ _0415_ _0410_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q
+ VPWR VGND sg13g2_a22oi_1
Xoutput192 net192 Tile_X0Y0_E2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput181 net181 Tile_X0Y0_E2BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_62_207 VPWR VGND sg13g2_decap_8
XFILLER_62_229 VPWR VGND sg13g2_decap_4
XFILLER_102_81 VPWR VGND sg13g2_fill_2
XFILLER_70_295 VPWR VGND sg13g2_fill_1
XFILLER_62_85 VPWR VGND sg13g2_fill_1
XFILLER_7_344 VPWR VGND sg13g2_fill_2
XFILLER_93_376 VPWR VGND sg13g2_fill_1
X_5841_ net1891 net1821 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_5772_ net1880 net1718 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_61_284 VPWR VGND sg13g2_decap_4
X_2984_ _1045_ _0519_ _1047_ VPWR VGND sg13g2_xor2_1
X_4723_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q _0275_
+ _0276_ _0063_ sg13g2_a21oi_1
X_4654_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q _0208_
+ _0211_ _0210_ sg13g2_a21oi_1
Xinput61 Tile_X0Y0_SS4END[7] net61 VPWR VGND sg13g2_buf_1
Xinput50 Tile_X0Y0_S4END[4] net50 VPWR VGND sg13g2_buf_1
X_3605_ VGND VPWR _1639_ _1642_ _1645_ _0145_ sg13g2_a21oi_1
X_4585_ VPWR _0142_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q VGND
+ sg13g2_inv_1
Xinput72 Tile_X0Y0_W2END[7] net72 VPWR VGND sg13g2_buf_1
Xinput94 Tile_X0Y1_E2END[3] net94 VPWR VGND sg13g2_buf_1
X_6324_ Tile_X0Y1_WW4END[11] net551 VPWR VGND sg13g2_buf_1
X_3536_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q _1581_ _1580_
+ _1578_ _1579_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7
+ VPWR VGND sg13g2_mux4_1
Xinput83 Tile_X0Y0_WW4END[0] net83 VPWR VGND sg13g2_buf_1
XFILLER_115_253 VPWR VGND sg13g2_fill_2
X_6255_ Tile_X0Y0_S4END[10] net482 VPWR VGND sg13g2_buf_1
X_3467_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q net1597 net1610
+ net649 net1624 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q _1516_
+ VPWR VGND sg13g2_mux4_1
XFILLER_67_19 VPWR VGND sg13g2_fill_2
X_5206_ net1949 net1765 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_6186_ Tile_X0Y1_EE4END[5] net413 VPWR VGND sg13g2_buf_1
X_3398_ _1369_ _1368_ _1450_ VPWR VGND sg13g2_xor2_1
X_5137_ net1939 net1786 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_29_259 VPWR VGND sg13g2_fill_2
X_5068_ net1991 net1806 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_4019_ VGND VPWR net4 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q
+ _2024_ _2023_ sg13g2_a21oi_1
XFILLER_44_218 VPWR VGND sg13g2_fill_1
XFILLER_20_192 VPWR VGND sg13g2_fill_1
XFILLER_32_88 VPWR VGND sg13g2_fill_2
XFILLER_4_325 VPWR VGND sg13g2_fill_2
XFILLER_79_104 VPWR VGND sg13g2_fill_1
XFILLER_79_126 VPWR VGND sg13g2_decap_4
XFILLER_94_118 VPWR VGND sg13g2_decap_8
XFILLER_43_251 VPWR VGND sg13g2_fill_2
X_4370_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q _1316_
+ _2298_ _0167_ sg13g2_a21oi_1
X_3321_ _1373_ _1213_ net1608 VPWR VGND sg13g2_nand2b_1
XFILLER_112_267 VPWR VGND sg13g2_fill_1
X_3252_ _1305_ _1297_ _1304_ VPWR VGND sg13g2_nand2_1
X_6040_ net1731 net271 VPWR VGND sg13g2_buf_1
XFILLER_112_278 VPWR VGND sg13g2_fill_1
X_3183_ _1235_ _1234_ _1237_ _1238_ VPWR VGND sg13g2_a21o_1
XFILLER_93_184 VPWR VGND sg13g2_fill_1
X_5824_ net1861 net1836 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_5755_ net1913 net1727 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_2967_ _1029_ _1025_ _1030_ VPWR VGND sg13g2_xor2_1
X_2898_ _0966_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 VPWR VGND sg13g2_inv_4
X_5686_ net1902 net1748 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_4706_ _0256_ _0258_ _0259_ VPWR VGND sg13g2_nor2_1
X_4637_ VPWR _0194_ _0193_ VGND sg13g2_inv_1
XFILLER_1_306 VPWR VGND sg13g2_fill_2
X_4568_ VPWR _0125_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q VGND
+ sg13g2_inv_1
X_6307_ Tile_X0Y1_W6END[4] net530 VPWR VGND sg13g2_buf_1
X_3519_ _1564_ VPWR _1565_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q
+ _1561_ sg13g2_o21ai_1
X_4499_ net1513 _2056_ _0056_ VPWR VGND sg13g2_nor2b_1
X_6238_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 net459 VPWR VGND sg13g2_buf_1
X_6169_ net103 net390 VPWR VGND sg13g2_buf_1
XFILLER_27_22 VPWR VGND sg13g2_fill_2
XFILLER_84_151 VPWR VGND sg13g2_fill_1
XFILLER_68_95 VPWR VGND sg13g2_fill_2
XFILLER_63_313 VPWR VGND sg13g2_fill_2
XFILLER_75_195 VPWR VGND sg13g2_fill_1
X_3870_ _1891_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[6\] net1653 VPWR VGND sg13g2_nand2_1
XFILLER_31_265 VPWR VGND sg13g2_fill_2
X_2821_ _0892_ VPWR _0894_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q
+ _0893_ sg13g2_o21ai_1
XFILLER_83_4 VPWR VGND sg13g2_fill_2
X_5540_ net1868 net1801 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_2752_ _0822_ _0828_ _0829_ VPWR VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q
+ sg13g2_nand3b_1
XFILLER_117_326 VPWR VGND sg13g2_fill_1
X_5471_ Tile_X0Y1_UserCLK net603 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X
+ _0003_ _5471_/Q VPWR VGND sg13g2_dfrbp_1
X_4422_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q _0176_
+ _2342_ _2341_ sg13g2_a21oi_1
X_2683_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q net115 net38
+ net108 net151 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q _0763_
+ VPWR VGND sg13g2_mux4_1
XFILLER_69_2 VPWR VGND sg13g2_fill_1
X_4353_ VGND VPWR _2283_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q
+ net1711 sg13g2_or2_1
X_4284_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q VPWR _2231_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q _2230_ sg13g2_o21ai_1
X_3304_ _1348_ VPWR _1356_ VGND _1346_ _1349_ sg13g2_o21ai_1
X_3235_ _1288_ _1287_ _1257_ VPWR VGND sg13g2_nand2b_1
X_6023_ net1969 net236 VPWR VGND sg13g2_buf_1
XFILLER_39_365 VPWR VGND sg13g2_fill_1
X_3166_ _1221_ _1219_ _1220_ VPWR VGND sg13g2_xnor2_1
X_3097_ _1149_ _1153_ _1154_ VPWR VGND sg13g2_nor2b_1
XFILLER_22_232 VPWR VGND sg13g2_fill_2
X_5807_ net1887 net1835 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_3999_ _2004_ net1702 _0179_ VPWR VGND sg13g2_nand2_1
X_5738_ net1876 net1724 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_5669_ net1875 net1760 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
Xfanout1906 net1907 net1906 VPWR VGND sg13g2_buf_1
Xfanout1917 net1918 net1917 VPWR VGND sg13g2_buf_1
Xfanout1928 net87 net1928 VPWR VGND sg13g2_buf_1
Xfanout1939 net1940 net1939 VPWR VGND sg13g2_buf_1
XFILLER_45_313 VPWR VGND sg13g2_fill_1
XFILLER_54_86 VPWR VGND sg13g2_fill_2
X_3020_ _1075_ _1081_ _1082_ VPWR VGND sg13g2_nor2_1
XFILLER_63_132 VPWR VGND sg13g2_fill_2
XFILLER_63_187 VPWR VGND sg13g2_decap_4
X_4971_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q net1709 net4 net30
+ net86 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q _0513_ VPWR VGND
+ sg13g2_mux4_1
XFILLER_63_198 VPWR VGND sg13g2_fill_1
X_3922_ _1933_ net1649 _0032_ VPWR VGND sg13g2_nand2_1
X_3853_ _1880_ _1866_ _1878_ VPWR VGND sg13g2_xnor2_1
X_2804_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q VPWR _0878_ VGND
+ net1688 _0175_ sg13g2_o21ai_1
X_3784_ _1812_ VPWR _1813_ VGND _1747_ _1749_ sg13g2_o21ai_1
XFILLER_74_0 VPWR VGND sg13g2_fill_1
X_5523_ net1895 net1804 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_2735_ _0812_ net1698 net1518 VPWR VGND sg13g2_nand2_1
Xoutput511 net511 Tile_X0Y1_W2BEG[1] VPWR VGND sg13g2_buf_1
Xoutput500 net500 Tile_X0Y1_SS4BEG[4] VPWR VGND sg13g2_buf_1
X_5454_ Tile_X0Y1_UserCLK net586 Tile_X0Y1_DSP_bot.B2 _5454_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[2\]
+ VPWR VGND sg13g2_dfrbp_1
X_2666_ VGND VPWR _0103_ _0747_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q
+ _0746_ sg13g2_a21oi_2
XFILLER_105_318 VPWR VGND sg13g2_fill_1
X_4405_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q net1580 _0905_
+ _1130_ _1744_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q _2328_
+ VPWR VGND sg13g2_mux4_1
Xoutput522 net522 Tile_X0Y1_W2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput544 net544 Tile_X0Y1_WW4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput533 net533 Tile_X0Y1_W6BEG[5] VPWR VGND sg13g2_buf_1
X_5385_ net1985 net1828 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_4336_ net1710 net1925 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q
+ _2269_ VPWR VGND sg13g2_mux2_1
X_2597_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3
+ net15 net41 net76 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q _0681_
+ VPWR VGND sg13g2_mux4_1
XFILLER_113_384 VPWR VGND sg13g2_fill_1
XFILLER_113_373 VPWR VGND sg13g2_fill_2
X_4267_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q _2223_
+ _2225_ _2224_ sg13g2_a21oi_1
X_3218_ _1272_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q _1264_
+ _1271_ VPWR VGND sg13g2_and3_1
X_6006_ net1944 net249 VPWR VGND sg13g2_buf_1
X_4198_ _2159_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 VGND _2163_
+ _2165_ sg13g2_o21ai_1
XFILLER_39_184 VPWR VGND sg13g2_fill_2
XFILLER_54_110 VPWR VGND sg13g2_decap_8
X_3149_ _1205_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q net106
+ VPWR VGND sg13g2_nand2b_1
XFILLER_91_29 VPWR VGND sg13g2_fill_2
XFILLER_10_213 VPWR VGND sg13g2_fill_1
Xfanout1714 net1715 net1714 VPWR VGND sg13g2_buf_1
Xfanout1703 net168 net1703 VPWR VGND sg13g2_buf_1
XFILLER_104_362 VPWR VGND sg13g2_fill_2
Xfanout1758 net1762 net1758 VPWR VGND sg13g2_buf_1
Xfanout1736 net1738 net1736 VPWR VGND sg13g2_buf_1
Xfanout1725 net1726 net1725 VPWR VGND sg13g2_buf_1
XFILLER_49_75 VPWR VGND sg13g2_fill_2
XFILLER_49_86 VPWR VGND sg13g2_fill_2
Xfanout1747 net1757 net1747 VPWR VGND sg13g2_buf_1
Xfanout1769 net1771 net1769 VPWR VGND sg13g2_buf_1
XFILLER_65_52 VPWR VGND sg13g2_fill_1
XFILLER_65_74 VPWR VGND sg13g2_decap_8
X_2520_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q _0607_
+ _0608_ _0108_ sg13g2_a21oi_1
X_5170_ net1942 net1777 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_4121_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q net31 net46
+ net1929 net1622 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3
+ VPWR VGND sg13g2_mux4_1
XFILLER_110_365 VPWR VGND sg13g2_fill_2
X_4052_ _2054_ net1655 Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[19\] VPWR VGND sg13g2_nand2_1
X_3003_ _1065_ VPWR _1066_ VGND net155 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q
+ sg13g2_o21ai_1
XFILLER_36_110 VPWR VGND sg13g2_decap_8
Xinput4 Tile_X0Y0_E2END[0] net4 VPWR VGND sg13g2_buf_1
X_4954_ VGND VPWR net125 net1696 _0497_ _0496_ sg13g2_a21oi_1
XFILLER_51_168 VPWR VGND sg13g2_fill_2
X_3905_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q _1918_
+ _1919_ _0119_ sg13g2_a21oi_1
X_4885_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q _0431_
+ _0432_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q sg13g2_a21oi_1
X_3836_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X
+ _1861_ _1863_ _1843_ _1842_ VPWR VGND sg13g2_a22oi_1
X_3767_ _1797_ net1707 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q
+ VPWR VGND sg13g2_nand2b_1
X_5506_ net1864 net1848 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_2718_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q VPWR _0797_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q _0796_ sg13g2_o21ai_1
X_3698_ _1440_ _1439_ _1732_ VPWR VGND sg13g2_xor2_1
X_2649_ VGND VPWR _0729_ _0730_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q
+ _0725_ sg13g2_a21oi_2
Xoutput330 net330 Tile_X0Y0_W2BEG[0] VPWR VGND sg13g2_buf_1
Xoutput341 net341 Tile_X0Y0_W2BEGb[3] VPWR VGND sg13g2_buf_1
X_5437_ Tile_X0Y1_UserCLK net561 _0051_ _0026_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[13\]
+ VPWR VGND sg13g2_dfrbp_1
Xoutput352 net352 Tile_X0Y0_W6BEG[4] VPWR VGND sg13g2_buf_1
Xoutput385 net385 Tile_X0Y1_E2BEG[7] VPWR VGND sg13g2_buf_8
Xoutput374 net374 Tile_X0Y1_E1BEG[0] VPWR VGND sg13g2_buf_1
Xoutput396 net396 Tile_X0Y1_E6BEG[11] VPWR VGND sg13g2_buf_1
Xoutput363 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 Tile_X0Y0_WW4BEG[14]
+ VPWR VGND sg13g2_buf_1
X_5368_ net1978 net1844 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_4319_ _2256_ _2255_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q
+ _2257_ VPWR VGND sg13g2_mux2_1
X_5299_ net1943 net1727 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_321 VPWR VGND sg13g2_fill_2
XFILLER_82_271 VPWR VGND sg13g2_fill_1
Xfanout1522 net1525 net1522 VPWR VGND sg13g2_buf_1
Xfanout1533 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 net1533 VPWR VGND sg13g2_buf_8
Xfanout1511 _0462_ net1511 VPWR VGND sg13g2_buf_8
XFILLER_104_170 VPWR VGND sg13g2_fill_1
Xfanout1544 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 net1544 VPWR VGND sg13g2_buf_8
Xfanout1566 net1567 net1566 VPWR VGND sg13g2_buf_1
Xfanout1555 _0171_ net1555 VPWR VGND sg13g2_buf_8
Xfanout1599 net1600 net1599 VPWR VGND sg13g2_buf_1
Xfanout1588 net1589 net1588 VPWR VGND sg13g2_buf_1
Xfanout1577 net1577 net1578 VPWR VGND sg13g2_buf_16
XFILLER_80_208 VPWR VGND sg13g2_decap_8
XFILLER_73_282 VPWR VGND sg13g2_fill_2
XFILLER_14_382 VPWR VGND sg13g2_fill_2
X_4670_ _0226_ net28 net1699 VPWR VGND sg13g2_nand2_1
X_3621_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q net1710 net122
+ net1925 net98 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q _1660_
+ VPWR VGND sg13g2_mux4_1
X_3552_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q net1560 net1566
+ net1574 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q
+ _1596_ VPWR VGND sg13g2_mux4_1
X_2503_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q _0590_
+ _0592_ _0591_ sg13g2_a21oi_1
X_6271_ Tile_X0Y0_SS4END[10] net498 VPWR VGND sg13g2_buf_1
X_3483_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q _1530_
+ _1531_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q sg13g2_a21oi_1
X_5222_ net1979 net1754 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_5153_ net1967 net1778 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_37_0 VPWR VGND sg13g2_fill_1
X_4104_ VGND VPWR _2093_ _2092_ _2086_ sg13g2_or2_1
XFILLER_110_184 VPWR VGND sg13g2_fill_2
X_5084_ net1957 net1797 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_4035_ VGND VPWR net22 net1679 _2039_ _2038_ sg13g2_a21oi_1
XFILLER_112_27 VPWR VGND sg13g2_fill_1
X_5986_ Tile_X0Y0_EE4END[6] net213 VPWR VGND sg13g2_buf_1
X_4937_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q _0478_ _0479_
+ _0480_ VPWR VGND sg13g2_nor3_1
X_4868_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q _0414_ _0415_
+ VPWR VGND sg13g2_nor2_1
X_3819_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q _1846_
+ _1848_ _1847_ sg13g2_a21oi_1
X_4799_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q net1528 net1534
+ net1542 net1557 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q _0349_
+ VPWR VGND sg13g2_mux4_1
XFILLER_118_273 VPWR VGND sg13g2_fill_2
Xoutput182 net182 Tile_X0Y0_E2BEG[5] VPWR VGND sg13g2_buf_1
Xoutput193 net193 Tile_X0Y0_E6BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_47_238 VPWR VGND sg13g2_fill_2
XFILLER_47_249 VPWR VGND sg13g2_fill_1
XFILLER_102_71 VPWR VGND sg13g2_fill_1
XFILLER_62_53 VPWR VGND sg13g2_decap_8
XFILLER_62_64 VPWR VGND sg13g2_decap_4
XFILLER_30_149 VPWR VGND sg13g2_fill_1
XFILLER_109_240 VPWR VGND sg13g2_fill_2
XFILLER_7_48 VPWR VGND sg13g2_fill_2
XFILLER_7_378 VPWR VGND sg13g2_fill_2
XFILLER_97_127 VPWR VGND sg13g2_fill_2
XFILLER_38_216 VPWR VGND sg13g2_fill_1
X_5840_ net1889 net1821 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_5771_ net1879 net1717 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_2983_ net1511 net1515 _1045_ _1046_ VPWR VGND sg13g2_nor3_1
X_4722_ net1521 net1518 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q
+ _0275_ VPWR VGND sg13g2_mux2_1
Xinput40 Tile_X0Y0_S2MID[2] net40 VPWR VGND sg13g2_buf_1
X_4653_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q VPWR _0210_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q _0209_ sg13g2_o21ai_1
Xinput51 Tile_X0Y0_S4END[5] net51 VPWR VGND sg13g2_buf_1
X_3604_ _1644_ _0144_ _1643_ VPWR VGND sg13g2_nand2_2
X_4584_ VPWR _0141_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q VGND
+ sg13g2_inv_1
Xinput62 Tile_X0Y0_W1END[0] net62 VPWR VGND sg13g2_buf_1
Xinput73 Tile_X0Y0_W2MID[0] net73 VPWR VGND sg13g2_buf_1
Xinput95 Tile_X0Y1_E2END[4] net95 VPWR VGND sg13g2_buf_1
X_6323_ Tile_X0Y1_WW4END[10] net550 VPWR VGND sg13g2_buf_1
X_3535_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q net111 net1928
+ net115 net91 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q _1581_
+ VPWR VGND sg13g2_mux4_1
Xinput84 Tile_X0Y0_WW4END[1] net84 VPWR VGND sg13g2_buf_1
X_6254_ Tile_X0Y0_S4END[9] net481 VPWR VGND sg13g2_buf_1
X_3466_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 net18 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q
+ _1515_ VPWR VGND sg13g2_mux2_1
X_5205_ net1948 net1765 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_6185_ Tile_X0Y1_EE4END[4] net406 VPWR VGND sg13g2_buf_1
X_3397_ _1394_ VPWR _1449_ VGND _1446_ _1447_ sg13g2_o21ai_1
X_5136_ net1938 net1786 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_5067_ net1990 net1806 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_4018_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q VPWR _2023_ VGND
+ _0061_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q sg13g2_o21ai_1
XFILLER_16_68 VPWR VGND sg13g2_fill_2
X_5969_ net17 net190 VPWR VGND sg13g2_buf_1
XFILLER_113_92 VPWR VGND sg13g2_decap_8
XFILLER_43_274 VPWR VGND sg13g2_fill_2
X_3320_ _1007_ net1548 _1372_ VPWR VGND sg13g2_nor2_1
X_3251_ _1304_ _1303_ _1298_ VPWR VGND sg13g2_xnor2_1
X_3182_ _1236_ _1163_ _1237_ VPWR VGND sg13g2_and2_1
XFILLER_78_182 VPWR VGND sg13g2_fill_1
X_5823_ net1858 net1834 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_5754_ net1911 net1727 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_2966_ _1029_ _1027_ _0850_ VPWR VGND sg13g2_xnor2_1
X_5685_ net1900 net1746 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_2897_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q _0956_ _0965_
+ _0966_ VPWR VGND sg13g2_a21o_2
X_4705_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q VPWR _0258_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q _0257_ sg13g2_o21ai_1
X_4636_ _0184_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q _0192_
+ _0193_ VPWR VGND sg13g2_a21o_1
XFILLER_118_59 VPWR VGND sg13g2_fill_1
X_6306_ Tile_X0Y1_W6END[3] net529 VPWR VGND sg13g2_buf_1
X_4567_ VPWR _0124_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q VGND
+ sg13g2_inv_1
X_3518_ _0143_ _1563_ _1564_ VPWR VGND sg13g2_nor2_1
X_4498_ net1513 _1980_ _0055_ VPWR VGND sg13g2_nor2b_1
X_6237_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 net458 VPWR VGND sg13g2_buf_1
X_3449_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q net126 net7 net33
+ net84 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q _1499_ VPWR VGND
+ sg13g2_mux4_1
X_6168_ net102 net389 VPWR VGND sg13g2_buf_1
XFILLER_57_344 VPWR VGND sg13g2_fill_1
X_5119_ net1964 net1787 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_45 VPWR VGND sg13g2_fill_1
X_6099_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A net311 VPWR VGND sg13g2_buf_8
XFILLER_40_233 VPWR VGND sg13g2_fill_1
XFILLER_67_119 VPWR VGND sg13g2_fill_2
XFILLER_90_111 VPWR VGND sg13g2_fill_1
XFILLER_84_84 VPWR VGND sg13g2_fill_1
XFILLER_84_95 VPWR VGND sg13g2_decap_4
XFILLER_31_200 VPWR VGND sg13g2_fill_1
X_2820_ net144 net23 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q
+ _0893_ VPWR VGND sg13g2_mux2_1
X_2751_ _0827_ VPWR _0828_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q
+ _0824_ sg13g2_o21ai_1
X_2682_ _0758_ _0761_ _0762_ VPWR VGND sg13g2_nor2_1
X_5470_ Tile_X0Y1_UserCLK net602 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X
+ _0005_ _5470_/Q VPWR VGND sg13g2_dfrbp_1
X_4421_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q VPWR _2341_ VGND
+ net1705 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q sg13g2_o21ai_1
X_4352_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q _0176_
+ _2282_ _2281_ sg13g2_a21oi_1
X_4283_ net1561 net1570 net1663 _2230_ VPWR VGND sg13g2_mux2_1
X_3303_ VPWR _1355_ _1354_ VGND sg13g2_inv_1
X_6022_ net1972 net235 VPWR VGND sg13g2_buf_1
XFILLER_39_300 VPWR VGND sg13g2_fill_1
X_3234_ _1287_ _1286_ _1285_ VPWR VGND sg13g2_nand2b_1
XFILLER_98_266 VPWR VGND sg13g2_fill_1
XFILLER_39_322 VPWR VGND sg13g2_fill_1
XFILLER_39_377 VPWR VGND sg13g2_fill_1
X_3165_ _1109_ _1108_ _1220_ VPWR VGND sg13g2_xor2_1
XFILLER_66_174 VPWR VGND sg13g2_fill_1
X_3096_ _1152_ _0769_ _1153_ VPWR VGND sg13g2_xor2_1
X_3998_ _0158_ VPWR _2003_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q
+ _2002_ sg13g2_o21ai_1
X_5806_ net1885 net1838 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_5737_ net1872 net1724 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_2949_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q _1012_ _1013_
+ VPWR VGND sg13g2_nor2b_1
X_5668_ net1868 net1760 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_4619_ VPWR _0176_ net1544 VGND sg13g2_inv_1
X_5599_ net1858 net1781 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_1_115 VPWR VGND sg13g2_fill_2
Xfanout1907 Tile_X0Y1_FrameData[15] net1907 VPWR VGND sg13g2_buf_1
Xfanout1918 Tile_X0Y1_FrameData[10] net1918 VPWR VGND sg13g2_buf_1
Xfanout1929 net81 net1929 VPWR VGND sg13g2_buf_1
XFILLER_38_33 VPWR VGND sg13g2_decap_4
XFILLER_57_196 VPWR VGND sg13g2_fill_1
XFILLER_13_244 VPWR VGND sg13g2_fill_2
X_5473__605 VPWR VGND net605 sg13g2_tiehi
X_4970_ VGND VPWR _0511_ _0512_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q
+ _0508_ sg13g2_a21oi_2
X_3921_ VPWR _1932_ _1931_ VGND sg13g2_inv_1
X_3852_ _1878_ _1867_ _1879_ VPWR VGND sg13g2_nor2_2
X_2803_ _0876_ VPWR _0877_ VGND net1688 net1590 sg13g2_o21ai_1
X_3783_ _1812_ _1811_ _1810_ VPWR VGND sg13g2_nand2b_1
X_5522_ net1893 net1805 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_67_0 VPWR VGND sg13g2_fill_2
X_2734_ _0810_ VPWR _0811_ VGND net1697 net1592 sg13g2_o21ai_1
Xoutput501 net501 Tile_X0Y1_SS4BEG[5] VPWR VGND sg13g2_buf_1
X_5453_ Tile_X0Y1_UserCLK net585 Tile_X0Y1_DSP_bot.B1 _5453_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[1\]
+ VPWR VGND sg13g2_dfrbp_1
X_2665_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q net1592 net1583
+ net1521 net699 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q _0746_
+ VPWR VGND sg13g2_mux4_1
Xoutput512 net512 Tile_X0Y1_W2BEG[2] VPWR VGND sg13g2_buf_1
X_4404_ VGND VPWR _2326_ _2327_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0
+ _2321_ sg13g2_a21oi_1
Xoutput523 net523 Tile_X0Y1_W2BEGb[5] VPWR VGND sg13g2_buf_1
Xoutput545 net545 Tile_X0Y1_WW4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput534 net534 Tile_X0Y1_W6BEG[6] VPWR VGND sg13g2_buf_1
X_2596_ net633 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 VPWR VGND sg13g2_inv_16
X_5384_ net1983 net1828 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_4335_ _2267_ VPWR _2268_ VGND _0104_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q
+ sg13g2_o21ai_1
X_4266_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q VPWR _2224_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q _2222_ sg13g2_o21ai_1
XFILLER_86_225 VPWR VGND sg13g2_fill_1
X_3217_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 _1264_ _1271_ VPWR VGND
+ sg13g2_nand2_2
XFILLER_86_269 VPWR VGND sg13g2_fill_1
X_4197_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q VPWR _2165_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q _2164_ sg13g2_o21ai_1
X_6005_ net1946 net248 VPWR VGND sg13g2_buf_1
X_3148_ _1203_ VPWR _1204_ VGND _0347_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q
+ sg13g2_o21ai_1
X_3079_ _0068_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q _1138_
+ VPWR VGND sg13g2_nor2_1
XFILLER_50_383 VPWR VGND sg13g2_fill_2
XFILLER_40_89 VPWR VGND sg13g2_fill_1
Xfanout1715 net1718 net1715 VPWR VGND sg13g2_buf_1
Xfanout1704 net150 net1704 VPWR VGND sg13g2_buf_1
Xfanout1737 net1738 net1737 VPWR VGND sg13g2_buf_1
Xfanout1726 net1734 net1726 VPWR VGND sg13g2_buf_1
Xfanout1748 net1750 net1748 VPWR VGND sg13g2_buf_1
Xfanout1759 net1762 net1759 VPWR VGND sg13g2_buf_1
XFILLER_92_206 VPWR VGND sg13g2_fill_1
XFILLER_18_303 VPWR VGND sg13g2_fill_2
XFILLER_92_228 VPWR VGND sg13g2_fill_2
XFILLER_60_169 VPWR VGND sg13g2_fill_2
XFILLER_81_63 VPWR VGND sg13g2_fill_2
XFILLER_68_214 VPWR VGND sg13g2_decap_4
X_4120_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q net30 net82
+ net49 net648 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2
+ VPWR VGND sg13g2_mux4_1
X_4051_ _2052_ _1990_ _2053_ VPWR VGND sg13g2_xor2_1
X_3002_ _1065_ _0058_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q
+ VPWR VGND sg13g2_nand2_1
Xinput5 Tile_X0Y0_E2END[1] net5 VPWR VGND sg13g2_buf_1
X_4953_ net1696 net687 _0496_ VPWR VGND sg13g2_nor2_1
X_3904_ _1917_ VPWR _1918_ VGND net37 net2005 sg13g2_o21ai_1
X_4884_ net1546 net1553 net1662 _0431_ VPWR VGND sg13g2_mux2_1
X_3835_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q _1862_
+ _1863_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q sg13g2_a21oi_1
X_3766_ VGND VPWR _1795_ _1796_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 sg13g2_a21oi_2
X_5505_ net1862 net1849 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_2717_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q net52
+ _0796_ _0795_ sg13g2_a21oi_1
X_3697_ _1731_ _1729_ _1730_ VPWR VGND sg13g2_nand2_2
X_5436_ Tile_X0Y1_UserCLK net562 _0050_ _0000_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[12\]
+ VPWR VGND sg13g2_dfrbp_1
Xoutput320 net320 Tile_X0Y0_NN4BEG[5] VPWR VGND sg13g2_buf_1
X_2648_ VPWR _0729_ _0728_ VGND sg13g2_inv_1
Xoutput331 net331 Tile_X0Y0_W2BEG[1] VPWR VGND sg13g2_buf_1
Xoutput342 net342 Tile_X0Y0_W2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput353 net353 Tile_X0Y0_W6BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_120_119 VPWR VGND sg13g2_fill_2
Xoutput386 net386 Tile_X0Y1_E2BEGb[0] VPWR VGND sg13g2_buf_1
X_2579_ net1659 net1528 net1534 net1543 net1558 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q
+ _0664_ VPWR VGND sg13g2_mux4_1
Xoutput375 net375 Tile_X0Y1_E1BEG[1] VPWR VGND sg13g2_buf_1
X_5367_ net1955 net1841 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput364 net364 Tile_X0Y0_WW4BEG[15] VPWR VGND sg13g2_buf_8
XFILLER_113_182 VPWR VGND sg13g2_fill_1
Xoutput397 net397 Tile_X0Y1_E6BEG[1] VPWR VGND sg13g2_buf_1
X_4318_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q net140 net1925
+ net92 net1921 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q _2256_
+ VPWR VGND sg13g2_mux4_1
X_5298_ net1941 net1728 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_4249_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q net2002 net1931
+ net1599 net1612 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q _2208_
+ VPWR VGND sg13g2_mux4_1
XFILLER_35_45 VPWR VGND sg13g2_decap_4
XFILLER_35_78 VPWR VGND sg13g2_fill_2
Xfanout1512 net1514 net1512 VPWR VGND sg13g2_buf_8
Xfanout1523 net1524 net1523 VPWR VGND sg13g2_buf_1
Xfanout1534 net1535 net1534 VPWR VGND sg13g2_buf_8
Xfanout1556 net1556 net1557 VPWR VGND sg13g2_buf_16
Xfanout1545 net1546 net1545 VPWR VGND sg13g2_buf_1
Xfanout1578 net1578 net1580 VPWR VGND sg13g2_buf_16
Xfanout1567 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 net1567 VPWR VGND sg13g2_buf_8
Xfanout1589 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 net1589 VPWR VGND
+ sg13g2_buf_8
XFILLER_119_219 VPWR VGND sg13g2_fill_2
X_3620_ _1659_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q _1658_
+ VPWR VGND sg13g2_nand2_1
X_3551_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q net1713 net1928
+ net115 net91 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q _1595_
+ VPWR VGND sg13g2_mux4_1
X_2502_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q VPWR _0591_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q _0588_ sg13g2_o21ai_1
X_6270_ Tile_X0Y0_SS4END[9] net497 VPWR VGND sg13g2_buf_1
X_3482_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q net729
+ _1530_ _1529_ sg13g2_a21oi_1
X_5221_ net1976 net1753 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_5152_ net1965 net1778 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_4103_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q VPWR _2092_ VGND
+ _2090_ _2091_ sg13g2_o21ai_1
XFILLER_2_71 VPWR VGND sg13g2_fill_2
X_5083_ net1953 net1797 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_4034_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q VPWR _2038_ VGND
+ _0061_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q sg13g2_o21ai_1
XFILLER_2_93 VPWR VGND sg13g2_fill_1
XFILLER_49_280 VPWR VGND sg13g2_decap_8
X_5985_ Tile_X0Y0_EE4END[5] net212 VPWR VGND sg13g2_buf_1
X_4936_ net12 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q _0479_ VPWR
+ VGND sg13g2_nor2b_1
XFILLER_20_320 VPWR VGND sg13g2_fill_2
X_4867_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q net1629 _0414_
+ VPWR VGND sg13g2_nor2_1
X_3818_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q VPWR _1847_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q _1845_ sg13g2_o21ai_1
X_4798_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q net1706 net106
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 net166 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q
+ _0348_ VPWR VGND sg13g2_mux4_1
X_3749_ _1777_ VPWR _1780_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q
+ _1779_ sg13g2_o21ai_1
X_5419_ net1990 net1817 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput183 net183 Tile_X0Y0_E2BEG[6] VPWR VGND sg13g2_buf_1
Xoutput194 net194 Tile_X0Y0_E6BEG[10] VPWR VGND sg13g2_buf_1
X_5770_ net1877 net1717 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_61_264 VPWR VGND sg13g2_fill_1
X_2982_ _1045_ _1036_ _1043_ VPWR VGND sg13g2_xnor2_1
X_4721_ _0274_ _0273_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q
+ VPWR VGND sg13g2_nand2b_1
X_4652_ net1923 net1935 net1657 _0209_ VPWR VGND sg13g2_mux2_1
Xinput30 Tile_X0Y0_S2END[0] net30 VPWR VGND sg13g2_buf_1
X_3603_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q net1532 net1536
+ net1547 net1554 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q _1643_
+ VPWR VGND sg13g2_mux4_1
Xinput52 Tile_X0Y0_S4END[6] net52 VPWR VGND sg13g2_buf_1
Xinput41 Tile_X0Y0_S2MID[3] net41 VPWR VGND sg13g2_buf_1
X_4583_ VPWR _0140_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q VGND
+ sg13g2_inv_1
Xinput63 Tile_X0Y0_W1END[1] net63 VPWR VGND sg13g2_buf_1
Xinput96 Tile_X0Y1_E2END[5] net96 VPWR VGND sg13g2_buf_1
X_6322_ Tile_X0Y1_WW4END[9] net549 VPWR VGND sg13g2_buf_1
X_3534_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q net708 net147
+ net38 net1705 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q _1580_
+ VPWR VGND sg13g2_mux4_1
Xinput74 Tile_X0Y0_W2MID[1] net74 VPWR VGND sg13g2_buf_1
Xinput85 Tile_X0Y0_WW4END[2] net85 VPWR VGND sg13g2_buf_1
X_6253_ Tile_X0Y0_S4END[8] net474 VPWR VGND sg13g2_buf_1
X_3465_ _1513_ VPWR _1514_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q
+ _1512_ sg13g2_o21ai_1
X_5204_ net1946 net1765 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_6184_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 net396 VPWR VGND sg13g2_buf_1
X_3396_ _1448_ _1392_ _1393_ VPWR VGND sg13g2_xnor2_1
X_5135_ net1997 net1786 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_96_183 VPWR VGND sg13g2_decap_4
X_5066_ net1988 net1806 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_4017_ _2021_ VPWR _2022_ VGND net688 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q
+ sg13g2_o21ai_1
XFILLER_84_356 VPWR VGND sg13g2_fill_1
XFILLER_37_272 VPWR VGND sg13g2_fill_1
X_5968_ net16 net189 VPWR VGND sg13g2_buf_1
X_4919_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q VPWR _0463_ VGND
+ net38 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q sg13g2_o21ai_1
XFILLER_32_79 VPWR VGND sg13g2_fill_1
XFILLER_106_233 VPWR VGND sg13g2_decap_4
XFILLER_106_255 VPWR VGND sg13g2_decap_4
XFILLER_121_258 VPWR VGND sg13g2_fill_1
XFILLER_43_242 VPWR VGND sg13g2_fill_1
XFILLER_73_97 VPWR VGND sg13g2_fill_2
X_3250_ _1300_ _1247_ _1303_ VPWR VGND sg13g2_xor2_1
X_3181_ _1159_ _1162_ _1052_ _1236_ VPWR VGND sg13g2_nand3_1
XFILLER_19_250 VPWR VGND sg13g2_fill_2
XFILLER_34_242 VPWR VGND sg13g2_fill_2
X_5822_ net1856 net1836 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_34_286 VPWR VGND sg13g2_fill_1
X_5753_ net1909 net1728 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_97_0 VPWR VGND sg13g2_fill_2
X_2965_ VGND VPWR _1028_ _1026_ _0931_ sg13g2_or2_1
X_4704_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q net146 net36 net10
+ net71 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q _0257_ VPWR VGND
+ sg13g2_mux4_1
X_2896_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q _0958_ _0964_
+ _0965_ VPWR VGND sg13g2_nor3_1
X_5684_ net1898 net1746 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_4635_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q _0186_ _0191_
+ _0192_ VPWR VGND sg13g2_nor3_1
X_4566_ VPWR _0123_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q VGND
+ sg13g2_inv_1
X_6305_ Tile_X0Y1_W6END[2] net526 VPWR VGND sg13g2_buf_1
X_3517_ VGND VPWR net147 net1671 _1563_ _1562_ sg13g2_a21oi_1
XFILLER_1_308 VPWR VGND sg13g2_fill_1
X_4497_ net1514 _1952_ _0054_ VPWR VGND sg13g2_nor2b_1
X_3448_ VGND VPWR _0117_ _1498_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5
+ _1490_ sg13g2_a21oi_1
X_6167_ net101 net388 VPWR VGND sg13g2_buf_1
X_3379_ _1429_ VPWR _1431_ VGND _1397_ _1430_ sg13g2_o21ai_1
X_5118_ net1962 net1788 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_24 VPWR VGND sg13g2_fill_1
X_6098_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A net310 VPWR VGND sg13g2_buf_1
XFILLER_84_131 VPWR VGND sg13g2_fill_1
X_5049_ net1999 net1853 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_43_56 VPWR VGND sg13g2_decap_8
XFILLER_0_330 VPWR VGND sg13g2_fill_1
XFILLER_75_164 VPWR VGND sg13g2_fill_2
XFILLER_31_267 VPWR VGND sg13g2_fill_1
X_2750_ _0826_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q _0827_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_83_6 VPWR VGND sg13g2_fill_1
X_2681_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q VPWR _0761_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q _0760_ sg13g2_o21ai_1
X_4420_ _2339_ VPWR _2340_ VGND _0169_ _0682_ sg13g2_o21ai_1
X_4351_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q _0682_ _2281_
+ VPWR VGND sg13g2_nor2_1
X_4282_ net1579 net1617 net1663 _2229_ VPWR VGND sg13g2_mux2_1
X_3302_ _1024_ _1282_ _1354_ VPWR VGND sg13g2_nor2_1
XFILLER_98_256 VPWR VGND sg13g2_fill_2
X_6021_ net1973 net234 VPWR VGND sg13g2_buf_1
X_3233_ _1286_ _1255_ _1256_ VPWR VGND sg13g2_xnor2_1
XFILLER_12_0 VPWR VGND sg13g2_fill_2
XFILLER_39_356 VPWR VGND sg13g2_fill_1
X_3164_ _1216_ VPWR _1219_ VGND _1217_ _1218_ sg13g2_o21ai_1
X_3095_ net1511 _1024_ _1152_ VPWR VGND sg13g2_nor2_1
X_3997_ net1598 net1611 net1701 _2002_ VPWR VGND sg13g2_mux2_1
X_5805_ net1882 net1833 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_13_48 VPWR VGND sg13g2_fill_2
X_5736_ net1870 net1724 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_2948_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q net14 net75 net40
+ net705 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q _1012_ VPWR VGND
+ sg13g2_mux4_1
X_5667_ net1866 net1759 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_4618_ VPWR _0175_ net1525 VGND sg13g2_inv_1
X_2879_ net35 net1933 net1686 _0949_ VPWR VGND sg13g2_mux2_1
X_5598_ net1856 net1780 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_4549_ VPWR _0106_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q VGND
+ sg13g2_inv_1
Xfanout1908 net1909 net1908 VPWR VGND sg13g2_buf_1
Xfanout1919 Tile_X0Y1_FrameData[0] net1919 VPWR VGND sg13g2_buf_1
X_6219_ net1901 net431 VPWR VGND sg13g2_buf_1
XFILLER_54_88 VPWR VGND sg13g2_fill_1
XFILLER_13_267 VPWR VGND sg13g2_fill_2
XFILLER_0_182 VPWR VGND sg13g2_fill_1
XFILLER_48_153 VPWR VGND sg13g2_decap_8
XFILLER_63_134 VPWR VGND sg13g2_fill_1
X_3920_ _1931_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q VPWR VGND
+ _1903_ sg13g2_nand2b_2
X_3851_ _1878_ _1877_ _1876_ VPWR VGND sg13g2_nand2b_1
X_3782_ _1811_ _1747_ _1748_ VPWR VGND sg13g2_xnor2_1
X_2802_ _0876_ net1688 net1583 VPWR VGND sg13g2_nand2_1
X_5521_ net1890 net1805 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_2733_ _0810_ net1697 net1583 VPWR VGND sg13g2_nand2b_1
Xoutput502 net502 Tile_X0Y1_SS4BEG[6] VPWR VGND sg13g2_buf_1
X_5452_ Tile_X0Y1_UserCLK net584 Tile_X0Y1_DSP_bot.B0 _5452_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[0\]
+ VPWR VGND sg13g2_dfrbp_1
X_2664_ _0745_ _0744_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q
+ VPWR VGND sg13g2_nand2b_1
X_2595_ _0672_ VPWR _0680_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q
+ _0679_ sg13g2_o21ai_1
X_4403_ _2323_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q _2327_
+ VPWR VGND sg13g2_nor2b_1
Xoutput524 net524 Tile_X0Y1_W2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput513 net513 Tile_X0Y1_W2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput535 net535 Tile_X0Y1_W6BEG[7] VPWR VGND sg13g2_buf_1
X_5383_ net1981 net1828 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_113_320 VPWR VGND sg13g2_fill_1
Xoutput546 net546 Tile_X0Y1_WW4BEG[2] VPWR VGND sg13g2_buf_1
X_4334_ _2267_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q net1553
+ VPWR VGND sg13g2_nand2_1
XFILLER_113_353 VPWR VGND sg13g2_fill_2
X_4265_ _1470_ net623 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q
+ _2223_ VPWR VGND sg13g2_mux2_1
X_6004_ net1947 net247 VPWR VGND sg13g2_buf_1
XFILLER_39_131 VPWR VGND sg13g2_fill_1
X_3216_ _1271_ _1268_ _1270_ VPWR VGND sg13g2_nand2b_1
X_4196_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q net1588 net1524
+ net1519 net1540 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q _2164_
+ VPWR VGND sg13g2_mux4_1
X_3147_ _1203_ net166 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q
+ VPWR VGND sg13g2_nand2_1
X_3078_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q VPWR _1137_ VGND
+ _1136_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q sg13g2_o21ai_1
XFILLER_54_178 VPWR VGND sg13g2_fill_2
X_5719_ net1905 net1738 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
Xfanout1705 net149 net1705 VPWR VGND sg13g2_buf_1
Xfanout1716 net1718 net1716 VPWR VGND sg13g2_buf_1
XFILLER_49_88 VPWR VGND sg13g2_fill_1
Xfanout1749 net1757 net1749 VPWR VGND sg13g2_buf_1
Xfanout1727 net1728 net1727 VPWR VGND sg13g2_buf_1
Xfanout1738 net1741 net1738 VPWR VGND sg13g2_buf_1
XFILLER_60_115 VPWR VGND sg13g2_decap_4
X_4050_ _2052_ net700 _2051_ VPWR VGND sg13g2_xnor2_1
X_3001_ _1064_ _1063_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q
+ VPWR VGND sg13g2_nand2b_1
Xinput6 Tile_X0Y0_E2END[2] net6 VPWR VGND sg13g2_buf_8
X_4952_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q VPWR _0495_ VGND
+ _0494_ _0493_ sg13g2_o21ai_1
X_4883_ _0429_ VPWR _0430_ VGND net1662 net1531 sg13g2_o21ai_1
X_3903_ _1917_ net2005 net1930 VPWR VGND sg13g2_nand2b_1
X_3834_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q net724 net1934
+ net19 net80 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q _1862_
+ VPWR VGND sg13g2_mux4_1
X_3765_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q net165 _1795_
+ VPWR VGND sg13g2_nor2b_1
X_5504_ net1860 net1849 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_2716_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q net1935 _0795_
+ VPWR VGND sg13g2_nor2b_1
X_3696_ _1730_ _1441_ _1443_ VPWR VGND sg13g2_xnor2_1
Xoutput310 net310 Tile_X0Y0_NN4BEG[10] VPWR VGND sg13g2_buf_1
X_2647_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q _0727_ _0728_
+ VPWR VGND sg13g2_nor2_1
X_5435_ Tile_X0Y1_UserCLK net563 _0049_ _0002_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[11\]
+ VPWR VGND sg13g2_dfrbp_1
Xoutput321 net321 Tile_X0Y0_NN4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput332 net332 Tile_X0Y0_W2BEG[2] VPWR VGND sg13g2_buf_1
Xoutput343 net343 Tile_X0Y0_W2BEGb[5] VPWR VGND sg13g2_buf_1
Xoutput387 net387 Tile_X0Y1_E2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput376 net376 Tile_X0Y1_E1BEG[2] VPWR VGND sg13g2_buf_1
X_5366_ net1949 net1841 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput365 net365 Tile_X0Y0_WW4BEG[1] VPWR VGND sg13g2_buf_1
X_2578_ _0663_ _0652_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 VPWR VGND
+ sg13g2_nor2_2
Xoutput354 net354 Tile_X0Y0_W6BEG[6] VPWR VGND sg13g2_buf_1
Xoutput398 net398 Tile_X0Y1_E6BEG[2] VPWR VGND sg13g2_buf_1
X_4317_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q net1936 net51
+ net152 net1703 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q _2255_
+ VPWR VGND sg13g2_mux4_1
X_5297_ net1939 net1729 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_323 VPWR VGND sg13g2_fill_1
X_4248_ _2206_ _2207_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 VPWR VGND sg13g2_mux2_1
XFILLER_101_356 VPWR VGND sg13g2_fill_2
XFILLER_19_69 VPWR VGND sg13g2_fill_2
X_4179_ VPWR _2148_ _2147_ VGND sg13g2_inv_1
XFILLER_42_104 VPWR VGND sg13g2_decap_8
Xfanout1524 net1525 net1524 VPWR VGND sg13g2_buf_1
Xfanout1513 net1514 net1513 VPWR VGND sg13g2_buf_8
Xfanout1557 net1557 net1558 VPWR VGND sg13g2_buf_16
Xfanout1535 net637 net1535 VPWR VGND sg13g2_buf_8
Xfanout1546 net1547 net1546 VPWR VGND sg13g2_buf_1
XFILLER_104_194 VPWR VGND sg13g2_decap_8
Xfanout1579 net1580 net1579 VPWR VGND sg13g2_buf_1
Xfanout1568 _1331_ net1568 VPWR VGND sg13g2_buf_8
XFILLER_18_167 VPWR VGND sg13g2_fill_2
XFILLER_33_148 VPWR VGND sg13g2_decap_8
XFILLER_33_159 VPWR VGND sg13g2_fill_1
XFILLER_25_90 VPWR VGND sg13g2_fill_1
XFILLER_14_384 VPWR VGND sg13g2_fill_1
X_3550_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q net703 _0682_
+ net58 net169 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q _1594_
+ VPWR VGND sg13g2_mux4_1
X_2501_ _0589_ VPWR _0590_ VGND net62 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q
+ sg13g2_o21ai_1
X_5220_ net1974 net1753 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_3481_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q net79 _1529_
+ VPWR VGND sg13g2_nor2b_1
X_5151_ net1964 net1778 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_5082_ net1951 net1797 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_4102_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q VPWR _2091_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q _2088_ sg13g2_o21ai_1
X_4033_ _2036_ VPWR _2037_ VGND net1679 net687 sg13g2_o21ai_1
XFILLER_110_197 VPWR VGND sg13g2_fill_2
XFILLER_112_18 VPWR VGND sg13g2_fill_1
X_5984_ Tile_X0Y0_EE4END[4] net205 VPWR VGND sg13g2_buf_1
X_4935_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0
+ _0478_ VPWR VGND sg13g2_nor2_1
XFILLER_32_181 VPWR VGND sg13g2_decap_8
X_4866_ _0413_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q _0412_
+ VPWR VGND sg13g2_nand2_1
X_3817_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q net1634 net1523
+ net1593 net1540 net1678 _1846_ VPWR VGND sg13g2_mux4_1
X_4797_ _0347_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 VPWR VGND sg13g2_inv_4
XFILLER_118_220 VPWR VGND sg13g2_fill_2
X_3748_ _1778_ VPWR _1779_ VGND _0074_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q
+ sg13g2_o21ai_1
XFILLER_118_275 VPWR VGND sg13g2_fill_1
X_3679_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q net118 net94
+ net58 net154 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q _1714_
+ VPWR VGND sg13g2_mux4_1
X_5418_ net1988 net1817 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput195 net195 Tile_X0Y0_E6BEG[11] VPWR VGND sg13g2_buf_1
X_5349_ net1976 net1842 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput173 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 Tile_X0Y0_E1BEG[0]
+ VPWR VGND sg13g2_buf_1
Xoutput184 net184 Tile_X0Y0_E2BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_101_175 VPWR VGND sg13g2_fill_2
XFILLER_15_104 VPWR VGND sg13g2_fill_2
XFILLER_15_137 VPWR VGND sg13g2_fill_2
XFILLER_109_253 VPWR VGND sg13g2_decap_8
XFILLER_109_297 VPWR VGND sg13g2_fill_1
Xfanout2000 Tile_X0Y0_FrameData[0] net2000 VPWR VGND sg13g2_buf_1
XFILLER_97_129 VPWR VGND sg13g2_fill_1
X_2981_ _1043_ _1036_ _1044_ VPWR VGND sg13g2_and2_1
XFILLER_99_4 VPWR VGND sg13g2_fill_1
X_4720_ net1592 net1583 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q
+ _0273_ VPWR VGND sg13g2_mux2_1
X_4651_ _0207_ VPWR _0208_ VGND net1657 net153 sg13g2_o21ai_1
Xinput31 Tile_X0Y0_S2END[1] net31 VPWR VGND sg13g2_buf_1
X_3602_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q _1641_
+ _1642_ _0144_ sg13g2_a21oi_1
Xinput20 Tile_X0Y0_E6END[0] net20 VPWR VGND sg13g2_buf_2
Xinput53 Tile_X0Y0_S4END[7] net53 VPWR VGND sg13g2_buf_1
Xinput42 Tile_X0Y0_S2MID[4] net42 VPWR VGND sg13g2_buf_1
X_4582_ VPWR _0139_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q VGND
+ sg13g2_inv_1
Xinput64 Tile_X0Y0_W1END[2] net64 VPWR VGND sg13g2_buf_1
Xinput97 Tile_X0Y1_E2END[6] net97 VPWR VGND sg13g2_buf_1
X_6321_ Tile_X0Y1_WW4END[8] net548 VPWR VGND sg13g2_buf_1
XFILLER_6_380 VPWR VGND sg13g2_fill_1
X_3533_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q net1558 net1564
+ net1574 net1619 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q _1579_
+ VPWR VGND sg13g2_mux4_1
Xinput75 Tile_X0Y0_W2MID[2] net75 VPWR VGND sg13g2_buf_1
Xinput86 Tile_X0Y0_WW4END[3] net86 VPWR VGND sg13g2_buf_1
XFILLER_115_234 VPWR VGND sg13g2_fill_2
X_6252_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 net473 VPWR VGND sg13g2_buf_1
X_3464_ _1513_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q _1511_
+ VPWR VGND sg13g2_nand2_1
X_6183_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 net395 VPWR VGND sg13g2_buf_8
X_5203_ net1943 net1763 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_3395_ _1392_ _1393_ _1447_ VPWR VGND sg13g2_nor2b_1
XFILLER_69_343 VPWR VGND sg13g2_fill_2
X_5134_ net1995 net1786 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_5065_ net1986 net1809 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_4016_ VGND VPWR net1709 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q
+ _2021_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q sg13g2_a21oi_1
X_5967_ net15 net188 VPWR VGND sg13g2_buf_1
X_4918_ _0461_ VPWR _0462_ VGND _0123_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[4\] sg13g2_o21ai_1
XFILLER_32_36 VPWR VGND sg13g2_fill_2
X_4849_ _0396_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q _0397_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_106_278 VPWR VGND sg13g2_fill_2
XFILLER_87_173 VPWR VGND sg13g2_fill_2
XFILLER_98_73 VPWR VGND sg13g2_fill_2
X_3180_ _1235_ _1160_ _1161_ VPWR VGND sg13g2_xnor2_1
X_5821_ net1917 net1834 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_5752_ net1907 net1728 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_2964_ _1027_ _1006_ _0899_ VPWR VGND sg13g2_nand2_2
X_4703_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q _0252_
+ _0256_ _0255_ sg13g2_a21oi_1
X_2895_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q _0962_
+ _0964_ _0963_ sg13g2_a21oi_1
X_5683_ net1894 net1749 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_4634_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q _0189_
+ _0191_ _0190_ sg13g2_a21oi_1
X_4565_ VPWR _0122_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q VGND
+ sg13g2_inv_1
X_3516_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q VPWR _1562_ VGND
+ _0077_ net1671 sg13g2_o21ai_1
X_6304_ net166 net525 VPWR VGND sg13g2_buf_1
X_4496_ net1513 _1930_ _0053_ VPWR VGND sg13g2_nor2b_1
X_3447_ VGND VPWR _0116_ _1491_ _1498_ _1497_ sg13g2_a21oi_1
X_6235_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 net456 VPWR VGND sg13g2_buf_1
XFILLER_103_226 VPWR VGND sg13g2_fill_1
X_3378_ _1430_ _1428_ _1414_ VPWR VGND sg13g2_xnor2_1
X_6166_ net100 net387 VPWR VGND sg13g2_buf_1
X_5117_ net1960 net1785 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_6097_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A net324 VPWR VGND sg13g2_buf_8
X_5048_ net1977 net1853 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_72_316 VPWR VGND sg13g2_fill_2
XFILLER_25_232 VPWR VGND sg13g2_fill_2
XFILLER_4_136 VPWR VGND sg13g2_fill_1
XFILLER_108_50 VPWR VGND sg13g2_fill_2
X_5464__596 VPWR VGND net596 sg13g2_tiehi
XFILLER_16_232 VPWR VGND sg13g2_fill_2
XFILLER_16_298 VPWR VGND sg13g2_fill_2
XFILLER_16_287 VPWR VGND sg13g2_fill_2
X_2680_ VGND VPWR net58 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q
+ _0760_ _0759_ sg13g2_a21oi_1
X_4350_ _2280_ _2279_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q
+ Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A VPWR VGND sg13g2_mux2_1
X_3301_ _1351_ _1352_ _1353_ VPWR VGND sg13g2_nor2_1
X_4281_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q net1557 net693
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 _0308_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 VPWR VGND sg13g2_mux4_1
X_6020_ net1975 net233 VPWR VGND sg13g2_buf_1
X_3232_ _1285_ _1258_ _1283_ VPWR VGND sg13g2_xnor2_1
X_3163_ _1218_ _1105_ _1215_ VPWR VGND sg13g2_xnor2_1
X_3094_ VPWR _1151_ _1150_ VGND sg13g2_inv_1
XFILLER_81_124 VPWR VGND sg13g2_decap_4
X_5804_ net1880 net1833 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_3996_ VGND VPWR net1701 net1623 _2001_ _2000_ sg13g2_a21oi_1
X_5735_ net1920 net1739 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_2947_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3
+ net15 net41 net76 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q _1011_
+ VPWR VGND sg13g2_mux4_1
X_5666_ net1864 net1759 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_4617_ VPWR _0174_ net1591 VGND sg13g2_inv_1
X_2878_ _0947_ VPWR _0948_ VGND _0091_ net1686 sg13g2_o21ai_1
X_5597_ net1917 net1781 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_4548_ VPWR _0105_ net148 VGND sg13g2_inv_1
X_4479_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q _2392_
+ _2393_ _2391_ sg13g2_a21oi_1
Xfanout1909 Tile_X0Y1_FrameData[14] net1909 VPWR VGND sg13g2_buf_1
X_6218_ net1903 net430 VPWR VGND sg13g2_buf_1
XFILLER_38_24 VPWR VGND sg13g2_fill_1
X_6149_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 net361 VPWR VGND sg13g2_buf_1
XFILLER_48_198 VPWR VGND sg13g2_decap_8
XFILLER_63_146 VPWR VGND sg13g2_decap_4
X_3850_ _1868_ _1875_ _1465_ _1877_ VPWR VGND sg13g2_nand3_1
X_3781_ _1768_ _1809_ _1810_ VPWR VGND sg13g2_nor2_2
X_2801_ _0874_ VPWR _0875_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q
+ _0873_ sg13g2_o21ai_1
X_5520_ net1888 net1805 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_2732_ net1697 net1596 net1609 net1621 net1629 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q
+ _0809_ VPWR VGND sg13g2_mux4_1
XFILLER_117_148 VPWR VGND sg13g2_fill_2
X_2663_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q net1609 net1602
+ net1621 net1629 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q _0744_
+ VPWR VGND sg13g2_mux4_1
X_5451_ Tile_X0Y1_UserCLK net583 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X
+ _5451_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[7\] VPWR VGND sg13g2_dfrbp_1
X_4402_ _2326_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q _2325_
+ VPWR VGND sg13g2_nand2_1
X_2594_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q _0674_ _0676_
+ _0678_ _0677_ _0089_ _0679_ VPWR VGND sg13g2_mux4_1
Xoutput525 net525 Tile_X0Y1_W2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput514 net514 Tile_X0Y1_W2BEG[4] VPWR VGND sg13g2_buf_1
Xoutput503 net503 Tile_X0Y1_SS4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput536 net536 Tile_X0Y1_W6BEG[8] VPWR VGND sg13g2_buf_1
X_5382_ net1979 net1828 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_4333_ VGND VPWR _2265_ _2266_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A _2260_ sg13g2_a21oi_1
Xoutput547 net547 Tile_X0Y1_WW4BEG[3] VPWR VGND sg13g2_buf_1
X_4264_ _0630_ _0868_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q
+ _2222_ VPWR VGND sg13g2_mux2_1
X_6003_ net1950 net246 VPWR VGND sg13g2_buf_1
X_3215_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q VPWR _1270_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q _1269_ sg13g2_o21ai_1
X_4195_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q _2161_
+ _2163_ _2162_ sg13g2_a21oi_1
X_3146_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q _1199_ _1201_
+ _1202_ VPWR VGND sg13g2_nor3_1
X_3077_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q net1529 net1535
+ net1550 net1559 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q _1136_
+ VPWR VGND sg13g2_mux4_1
X_5718_ net1903 net1738 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_3979_ VGND VPWR net1644 _0155_ _1984_ net1651 sg13g2_a21oi_1
XFILLER_108_115 VPWR VGND sg13g2_fill_1
X_5649_ net1890 net1758 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_159 VPWR VGND sg13g2_decap_4
Xfanout1706 net130 net1706 VPWR VGND sg13g2_buf_1
Xfanout1717 net1718 net1717 VPWR VGND sg13g2_buf_1
Xfanout1728 net1734 net1728 VPWR VGND sg13g2_buf_1
Xfanout1739 net1741 net1739 VPWR VGND sg13g2_buf_1
XFILLER_18_305 VPWR VGND sg13g2_fill_1
XFILLER_65_88 VPWR VGND sg13g2_decap_8
XFILLER_81_43 VPWR VGND sg13g2_fill_2
XFILLER_81_65 VPWR VGND sg13g2_fill_1
XFILLER_81_87 VPWR VGND sg13g2_decap_4
X_3000_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q net1711 net119
+ net131 net95 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q _1063_
+ VPWR VGND sg13g2_mux4_1
Xinput7 Tile_X0Y0_E2END[3] net7 VPWR VGND sg13g2_buf_1
XFILLER_36_124 VPWR VGND sg13g2_fill_2
X_4951_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q VPWR _0494_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q _0491_ sg13g2_o21ai_1
X_4882_ _0429_ net1662 _0180_ VPWR VGND sg13g2_nand2_1
X_3902_ _1915_ VPWR _1916_ VGND _0091_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q
+ sg13g2_o21ai_1
X_3833_ _1861_ _1860_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q
+ VPWR VGND sg13g2_nand2b_1
X_3764_ _1791_ _1793_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q
+ _1794_ VPWR VGND sg13g2_nand3_1
X_2715_ net153 net167 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q
+ _0794_ VPWR VGND sg13g2_mux2_1
X_3695_ _1728_ _1729_ VPWR VGND sg13g2_inv_4
X_5503_ net1859 net1849 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput300 net300 Tile_X0Y0_N4BEG[1] VPWR VGND sg13g2_buf_1
X_2646_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q _0726_ _0727_
+ VPWR VGND sg13g2_nor2_1
X_5434_ Tile_X0Y1_UserCLK net564 _0048_ _0004_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[10\]
+ VPWR VGND sg13g2_dfrbp_1
Xoutput322 net322 Tile_X0Y0_NN4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput311 net311 Tile_X0Y0_NN4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput333 net333 Tile_X0Y0_W2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput344 net344 Tile_X0Y0_W2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput377 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 Tile_X0Y1_E1BEG[3]
+ VPWR VGND sg13g2_buf_1
X_5365_ net1947 net1841 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput366 net366 Tile_X0Y0_WW4BEG[2] VPWR VGND sg13g2_buf_1
X_2577_ VGND VPWR _0662_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q
+ _0659_ _0654_ _0663_ _0657_ sg13g2_a221oi_1
Xoutput355 net355 Tile_X0Y0_W6BEG[7] VPWR VGND sg13g2_buf_1
Xoutput399 net399 Tile_X0Y1_E6BEG[3] VPWR VGND sg13g2_buf_1
Xoutput388 net388 Tile_X0Y1_E2BEGb[2] VPWR VGND sg13g2_buf_1
X_4316_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q VPWR _2254_ VGND
+ _2248_ _2251_ sg13g2_o21ai_1
X_5296_ net1937 net1729 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_4247_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q net1539 _1470_
+ net623 _0525_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q _2207_
+ VPWR VGND sg13g2_mux4_1
XFILLER_59_238 VPWR VGND sg13g2_fill_2
XFILLER_101_368 VPWR VGND sg13g2_fill_2
XFILLER_101_379 VPWR VGND sg13g2_fill_2
X_4178_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q net1606 net1634
+ net1626 net1593 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q _2147_
+ VPWR VGND sg13g2_mux4_1
XFILLER_67_293 VPWR VGND sg13g2_fill_2
X_3129_ VGND VPWR net130 net1691 _1186_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q
+ sg13g2_a21oi_1
Xfanout1514 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr net1514 VPWR VGND sg13g2_buf_8
Xfanout1547 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 net1547 VPWR VGND sg13g2_buf_1
Xfanout1536 net635 net1536 VPWR VGND sg13g2_buf_8
Xfanout1525 net1526 net1525 VPWR VGND sg13g2_buf_1
Xfanout1569 net1571 net1569 VPWR VGND sg13g2_buf_1
Xfanout1558 net1558 net721 VPWR VGND sg13g2_buf_16
XFILLER_26_190 VPWR VGND sg13g2_fill_2
X_2500_ _0589_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q net1932
+ VPWR VGND sg13g2_nand2b_1
X_3480_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 _1527_ _1528_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q
+ _1519_ VPWR VGND sg13g2_a22oi_1
X_5150_ net1961 net1778 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_96_300 VPWR VGND sg13g2_fill_2
X_5081_ net1999 net1810 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_4101_ VGND VPWR net1673 _0179_ _2090_ _2089_ sg13g2_a21oi_1
X_4032_ VGND VPWR net1709 net1679 _2036_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q
+ sg13g2_a21oi_1
X_5983_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 net195 VPWR VGND sg13g2_buf_1
X_4934_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 _0475_ _0477_ _0466_
+ _0473_ VPWR VGND sg13g2_a22oi_1
XFILLER_20_322 VPWR VGND sg13g2_fill_1
X_4865_ VPWR _0412_ _0411_ VGND sg13g2_inv_1
X_3816_ VPWR _1845_ _1844_ VGND sg13g2_inv_1
X_4796_ _0335_ _0346_ _0347_ VPWR VGND sg13g2_nor2b_2
X_3747_ _1778_ net102 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q
+ VPWR VGND sg13g2_nand2_1
X_3678_ _1713_ net1647 _0014_ VPWR VGND sg13g2_nand2_1
X_5417_ net1986 net1819 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_2629_ _0101_ _0710_ _0711_ VPWR VGND sg13g2_nor2_1
X_5348_ net1974 net1843 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput174 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 Tile_X0Y0_E1BEG[1]
+ VPWR VGND sg13g2_buf_1
Xoutput185 net185 Tile_X0Y0_E2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput196 net196 Tile_X0Y0_E6BEG[1] VPWR VGND sg13g2_buf_1
X_5279_ net1963 net1732 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_198 VPWR VGND sg13g2_decap_8
XFILLER_70_211 VPWR VGND sg13g2_decap_8
XFILLER_15_127 VPWR VGND sg13g2_fill_2
XFILLER_11_71 VPWR VGND sg13g2_fill_1
Xfanout2001 net2002 net2001 VPWR VGND sg13g2_buf_1
XFILLER_87_53 VPWR VGND sg13g2_fill_2
XFILLER_38_208 VPWR VGND sg13g2_fill_2
XFILLER_61_211 VPWR VGND sg13g2_decap_4
X_2980_ _1043_ _1037_ _1041_ VPWR VGND sg13g2_xnor2_1
X_4650_ _0207_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q _0058_
+ VPWR VGND sg13g2_nand2_1
X_3601_ _1640_ VPWR _1641_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q
+ net1582 sg13g2_o21ai_1
Xinput10 Tile_X0Y0_E2END[6] net10 VPWR VGND sg13g2_buf_1
Xinput21 Tile_X0Y0_E6END[1] net21 VPWR VGND sg13g2_buf_1
Xinput54 Tile_X0Y0_SS4END[0] net54 VPWR VGND sg13g2_buf_1
Xinput32 net32 Tile_X0Y0_S2END[2] VPWR VGND sg13g2_buf_16
Xinput43 Tile_X0Y0_S2MID[5] net43 VPWR VGND sg13g2_buf_1
X_6320_ Tile_X0Y1_WW4END[7] net547 VPWR VGND sg13g2_buf_1
X_4581_ VPWR _0138_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q VGND
+ sg13g2_inv_1
Xinput98 Tile_X0Y1_E2END[7] net98 VPWR VGND sg13g2_buf_1
Xinput87 Tile_X0Y1_E1END[0] net87 VPWR VGND sg13g2_buf_1
X_3532_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q net1532 net1536
+ net1546 net1553 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q _1578_
+ VPWR VGND sg13g2_mux4_1
Xinput76 Tile_X0Y0_W2MID[3] net76 VPWR VGND sg13g2_buf_1
Xinput65 Tile_X0Y0_W2END[0] net65 VPWR VGND sg13g2_buf_1
X_6251_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 net472 VPWR VGND sg13g2_buf_1
X_3463_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q net130 net24
+ net37 net72 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q _1512_
+ VPWR VGND sg13g2_mux4_1
X_6182_ Tile_X0Y1_E6END[11] net405 VPWR VGND sg13g2_buf_1
X_5202_ net1941 net1763 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_5133_ net1993 net1785 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_35_0 VPWR VGND sg13g2_fill_2
X_3394_ VGND VPWR _1412_ _1446_ _1445_ _1444_ sg13g2_a21oi_2
XFILLER_69_366 VPWR VGND sg13g2_fill_2
X_5064_ net1984 net1809 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_4015_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q _2018_
+ _2020_ _2019_ sg13g2_a21oi_1
X_5966_ net14 net187 VPWR VGND sg13g2_buf_1
X_4917_ _0461_ net1640 _0460_ VPWR VGND sg13g2_nand2_2
X_4848_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q _0393_ _0395_
+ _0396_ VPWR VGND sg13g2_nor3_1
XFILLER_32_26 VPWR VGND sg13g2_fill_1
X_4779_ _0329_ VPWR _0330_ VGND net1692 _0327_ sg13g2_o21ai_1
XFILLER_113_40 VPWR VGND sg13g2_fill_2
XFILLER_113_84 VPWR VGND sg13g2_decap_4
XFILLER_73_55 VPWR VGND sg13g2_decap_4
XFILLER_73_77 VPWR VGND sg13g2_fill_2
XFILLER_73_88 VPWR VGND sg13g2_fill_2
X_5469__601 VPWR VGND net601 sg13g2_tiehi
XFILLER_22_70 VPWR VGND sg13g2_fill_1
XFILLER_7_189 VPWR VGND sg13g2_fill_1
XFILLER_78_141 VPWR VGND sg13g2_fill_1
XFILLER_34_222 VPWR VGND sg13g2_fill_2
X_5820_ net1915 net1834 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_5751_ net1905 net1725 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_2963_ _1026_ _0849_ _1006_ VPWR VGND sg13g2_nand2_1
X_4702_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q VPWR _0255_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q _0254_ sg13g2_o21ai_1
X_2894_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q VPWR _0963_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q _0960_ sg13g2_o21ai_1
X_5682_ net1892 net1749 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_4633_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q VPWR _0190_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q _0187_ sg13g2_o21ai_1
X_4564_ VPWR _0121_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q VGND
+ sg13g2_inv_1
X_3515_ _1560_ VPWR _1561_ VGND net1671 _0416_ sg13g2_o21ai_1
X_6303_ net165 net524 VPWR VGND sg13g2_buf_1
X_6234_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 net455 VPWR VGND sg13g2_buf_8
X_4495_ net1513 _1881_ _0052_ VPWR VGND sg13g2_nor2_1
X_3446_ _1493_ _1496_ _1497_ VPWR VGND sg13g2_nor2_1
X_6165_ net99 net386 VPWR VGND sg13g2_buf_1
X_3377_ _1429_ _1414_ _1428_ VPWR VGND sg13g2_nand2_1
X_5116_ net1958 net1785 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_6096_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A net323 VPWR VGND sg13g2_buf_1
XFILLER_57_369 VPWR VGND sg13g2_fill_2
X_5047_ net1955 net1851 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_25_222 VPWR VGND sg13g2_fill_2
XFILLER_4_104 VPWR VGND sg13g2_fill_1
XFILLER_108_40 VPWR VGND sg13g2_fill_1
XFILLER_108_95 VPWR VGND sg13g2_fill_2
XFILLER_48_336 VPWR VGND sg13g2_fill_2
XFILLER_84_21 VPWR VGND sg13g2_fill_1
XFILLER_75_166 VPWR VGND sg13g2_fill_1
XFILLER_16_255 VPWR VGND sg13g2_fill_1
X_3300_ _1352_ _1297_ _1304_ VPWR VGND sg13g2_xnor2_1
X_4280_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 _2228_ VPWR VGND sg13g2_inv_2
X_3231_ _1284_ _1258_ _1283_ VPWR VGND sg13g2_nand2_2
XFILLER_98_258 VPWR VGND sg13g2_fill_1
X_3162_ _1217_ net714 net1575 VPWR VGND sg13g2_nand2_1
XFILLER_66_111 VPWR VGND sg13g2_fill_2
XFILLER_66_166 VPWR VGND sg13g2_fill_1
X_3093_ net1608 _1024_ _1150_ VPWR VGND sg13g2_nor2_1
XFILLER_81_114 VPWR VGND sg13g2_decap_4
XFILLER_22_225 VPWR VGND sg13g2_decap_8
X_5803_ net1878 net1833 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_3995_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q VPWR _2000_ VGND
+ net1702 _0177_ sg13g2_o21ai_1
X_5734_ net1897 net1739 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_2946_ _1009_ _1008_ _1010_ VPWR VGND sg13g2_nor2_2
X_5665_ net1863 net1761 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_2877_ VGND VPWR net29 net1686 _0947_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q
+ sg13g2_a21oi_1
X_4616_ VPWR _0173_ net1572 VGND sg13g2_inv_1
X_5596_ net1915 net1780 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_4547_ VPWR _0104_ net1704 VGND sg13g2_inv_1
X_4478_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q net159 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 net614 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q
+ _2392_ VPWR VGND sg13g2_mux4_1
X_6217_ net1905 net429 VPWR VGND sg13g2_buf_1
X_3429_ VGND VPWR net15 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q
+ _1480_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q sg13g2_a21oi_1
X_6148_ Tile_X0Y0_WW4END[15] net360 VPWR VGND sg13g2_buf_1
X_6079_ Tile_X0Y1_N4END[15] net306 VPWR VGND sg13g2_buf_1
XFILLER_70_34 VPWR VGND sg13g2_fill_1
XFILLER_70_78 VPWR VGND sg13g2_fill_2
XFILLER_107_330 VPWR VGND sg13g2_fill_2
XFILLER_119_94 VPWR VGND sg13g2_fill_2
XFILLER_28_80 VPWR VGND sg13g2_fill_2
X_3780_ _1807_ _1808_ _1809_ VPWR VGND sg13g2_nor2b_1
X_2800_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q _0872_
+ _0874_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q sg13g2_a21oi_1
X_2731_ _0808_ _0807_ VPWR VGND sg13g2_inv_8
X_5450_ Tile_X0Y1_UserCLK net582 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X
+ _5450_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[6\] VPWR VGND sg13g2_dfrbp_1
X_4401_ _2324_ VPWR _2325_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q
+ _1278_ sg13g2_o21ai_1
X_2662_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q VPWR _0743_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q net159 sg13g2_o21ai_1
X_5381_ net1975 net1827 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_2593_ net119 net131 net1658 _0678_ VPWR VGND sg13g2_mux2_1
Xoutput515 net515 Tile_X0Y1_W2BEG[5] VPWR VGND sg13g2_buf_1
Xoutput504 net504 Tile_X0Y1_SS4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput526 net526 Tile_X0Y1_W6BEG[0] VPWR VGND sg13g2_buf_1
X_4332_ _2262_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q _2266_
+ VPWR VGND sg13g2_nor2b_1
Xoutput537 net537 Tile_X0Y1_W6BEG[9] VPWR VGND sg13g2_buf_1
Xoutput548 net548 Tile_X0Y1_WW4BEG[4] VPWR VGND sg13g2_buf_1
X_4263_ _2220_ VPWR _2221_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q
+ _2217_ sg13g2_o21ai_1
X_3214_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q net1533 net635
+ net1547 net1554 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q _1269_
+ VPWR VGND sg13g2_mux4_1
X_6002_ net1956 net243 VPWR VGND sg13g2_buf_1
X_4194_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q VPWR _2162_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q _2160_ sg13g2_o21ai_1
XFILLER_39_166 VPWR VGND sg13g2_fill_1
X_3145_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q net633
+ _1201_ _1200_ sg13g2_a21oi_1
X_3076_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q _1132_
+ _1135_ _1134_ sg13g2_a21oi_1
XFILLER_39_199 VPWR VGND sg13g2_decap_4
X_3978_ _1983_ net1638 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X
+ VPWR VGND sg13g2_nand2_1
X_5717_ net1901 net1737 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_2929_ _0994_ VPWR _0995_ VGND _0992_ _0993_ sg13g2_o21ai_1
X_5648_ net1888 net1758 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_5579_ net1879 net1782 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_104_300 VPWR VGND sg13g2_fill_2
XFILLER_116_193 VPWR VGND sg13g2_fill_1
Xfanout1707 net129 net1707 VPWR VGND sg13g2_buf_1
XFILLER_49_68 VPWR VGND sg13g2_fill_2
Xfanout1718 Tile_X0Y1_FrameStrobe[9] net1718 VPWR VGND sg13g2_buf_1
Xfanout1729 net1734 net1729 VPWR VGND sg13g2_buf_1
XFILLER_45_136 VPWR VGND sg13g2_fill_2
XFILLER_26_383 VPWR VGND sg13g2_fill_2
XFILLER_110_325 VPWR VGND sg13g2_fill_2
Xinput8 Tile_X0Y0_E2END[4] net8 VPWR VGND sg13g2_buf_1
XFILLER_76_272 VPWR VGND sg13g2_fill_2
XFILLER_36_136 VPWR VGND sg13g2_fill_2
XFILLER_91_231 VPWR VGND sg13g2_fill_1
XFILLER_17_361 VPWR VGND sg13g2_fill_1
X_4950_ VGND VPWR net1695 _0179_ _0493_ _0492_ sg13g2_a21oi_1
X_4881_ _0427_ VPWR _0428_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q
+ _0425_ sg13g2_o21ai_1
X_3901_ VGND VPWR net29 net2005 _1915_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q
+ sg13g2_a21oi_1
X_3832_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6
+ net18 net44 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q
+ _1860_ VPWR VGND sg13g2_mux4_1
X_3763_ _1793_ _1792_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q
+ VPWR VGND sg13g2_nand2b_1
X_5502_ net1857 net1849 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_2714_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q net1713 net117
+ net93 net1923 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q _0793_
+ VPWR VGND sg13g2_mux4_1
X_3694_ _1713_ VPWR _1728_ VGND _1727_ net1647 sg13g2_o21ai_1
XFILLER_65_0 VPWR VGND sg13g2_fill_2
Xoutput301 net301 Tile_X0Y0_N4BEG[2] VPWR VGND sg13g2_buf_1
X_5433_ Tile_X0Y1_UserCLK net565 _0047_ _0006_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[9\]
+ VPWR VGND sg13g2_dfrbp_1
X_2645_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q net1712 net120
+ net88 net96 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q _0726_
+ VPWR VGND sg13g2_mux4_1
Xoutput323 net323 Tile_X0Y0_NN4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput312 net312 Tile_X0Y0_NN4BEG[12] VPWR VGND sg13g2_buf_1
X_5364_ net1945 net1841 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput334 net334 Tile_X0Y0_W2BEG[4] VPWR VGND sg13g2_buf_1
Xoutput378 net378 Tile_X0Y1_E2BEG[0] VPWR VGND sg13g2_buf_1
X_4315_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q _2252_ _2253_
+ VPWR VGND sg13g2_nor2_1
Xoutput345 net345 Tile_X0Y0_W2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput367 net367 Tile_X0Y0_WW4BEG[3] VPWR VGND sg13g2_buf_1
X_2576_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q _0661_
+ _0662_ _0094_ sg13g2_a21oi_1
Xoutput356 net356 Tile_X0Y0_W6BEG[8] VPWR VGND sg13g2_buf_1
XFILLER_99_331 VPWR VGND sg13g2_fill_2
Xoutput389 net389 Tile_X0Y1_E2BEGb[3] VPWR VGND sg13g2_buf_1
X_5295_ net1997 net1733 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_99_375 VPWR VGND sg13g2_fill_2
X_4246_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q _0376_ net63
+ net27 net1591 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q _2206_
+ VPWR VGND sg13g2_mux4_1
X_4177_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q net2001 net1930
+ net1599 net1613 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q _2146_
+ VPWR VGND sg13g2_mux4_1
X_3128_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q _1183_
+ _1185_ _1184_ sg13g2_a21oi_1
XFILLER_27_114 VPWR VGND sg13g2_fill_1
XFILLER_82_253 VPWR VGND sg13g2_fill_1
X_3059_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q VPWR _1119_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q _1116_ sg13g2_o21ai_1
XFILLER_35_59 VPWR VGND sg13g2_fill_2
XFILLER_50_172 VPWR VGND sg13g2_decap_8
XFILLER_2_213 VPWR VGND sg13g2_fill_1
XFILLER_4_4 VPWR VGND sg13g2_fill_2
Xfanout1515 _0518_ net1515 VPWR VGND sg13g2_buf_8
Xfanout1537 net1537 net635 VPWR VGND sg13g2_buf_16
Xfanout1548 _1282_ net1548 VPWR VGND sg13g2_buf_8
Xfanout1526 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 net1526 VPWR VGND
+ sg13g2_buf_8
Xfanout1559 net1560 net1559 VPWR VGND sg13g2_buf_8
XFILLER_58_250 VPWR VGND sg13g2_fill_1
XFILLER_18_169 VPWR VGND sg13g2_fill_1
XFILLER_33_128 VPWR VGND sg13g2_fill_2
X_5080_ net1977 net1810 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_4100_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q VPWR _2089_ VGND
+ net1673 net1522 sg13g2_o21ai_1
X_4031_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q _2033_
+ _2035_ _2034_ sg13g2_a21oi_1
XFILLER_56_209 VPWR VGND sg13g2_fill_2
XFILLER_49_294 VPWR VGND sg13g2_decap_8
XFILLER_64_242 VPWR VGND sg13g2_fill_1
XFILLER_64_253 VPWR VGND sg13g2_fill_2
X_5982_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 net194 VPWR VGND sg13g2_buf_1
X_4933_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q _0476_
+ _0477_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q sg13g2_a21oi_1
X_4864_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q net611 net1936
+ net13 net74 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q _0411_
+ VPWR VGND sg13g2_mux4_1
X_3815_ net1678 net1600 net1612 net1605 net1625 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q
+ _1844_ VPWR VGND sg13g2_mux4_1
X_4795_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q _0345_ _0340_
+ _0346_ VPWR VGND sg13g2_nand3_1
XFILLER_118_222 VPWR VGND sg13g2_fill_1
X_3746_ _1777_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q _1776_
+ VPWR VGND sg13g2_nand2_1
X_3677_ _1710_ _1711_ _1712_ VPWR VGND sg13g2_nor2_1
X_5416_ net1984 net1819 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_2628_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q _0708_
+ _0710_ _0709_ sg13g2_a21oi_1
X_2559_ _0645_ _0642_ _0644_ VPWR VGND sg13g2_nand2b_1
X_5347_ net1971 net1842 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput175 net175 Tile_X0Y0_E1BEG[2] VPWR VGND sg13g2_buf_1
Xoutput186 net186 Tile_X0Y0_E2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput197 net197 Tile_X0Y0_E6BEG[2] VPWR VGND sg13g2_buf_1
X_5278_ net1961 net1732 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_4229_ _2190_ VPWR _2191_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q
+ net1526 sg13g2_o21ai_1
XFILLER_101_177 VPWR VGND sg13g2_fill_1
XFILLER_46_36 VPWR VGND sg13g2_fill_2
XFILLER_102_64 VPWR VGND sg13g2_decap_8
XFILLER_109_211 VPWR VGND sg13g2_decap_8
XFILLER_11_50 VPWR VGND sg13g2_fill_2
Xfanout2002 Tile_X0Y0_E1END[3] net2002 VPWR VGND sg13g2_buf_1
XFILLER_46_264 VPWR VGND sg13g2_fill_1
XFILLER_14_150 VPWR VGND sg13g2_fill_2
X_3600_ _1640_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q net1620
+ VPWR VGND sg13g2_nand2b_1
X_4580_ VPWR _0137_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q VGND
+ sg13g2_inv_1
Xinput22 Tile_X0Y0_EE4END[0] net22 VPWR VGND sg13g2_buf_1
Xinput11 Tile_X0Y0_E2END[7] net11 VPWR VGND sg13g2_buf_1
Xinput55 Tile_X0Y0_SS4END[1] net55 VPWR VGND sg13g2_buf_1
Xinput33 Tile_X0Y0_S2END[3] net33 VPWR VGND sg13g2_buf_1
Xinput44 Tile_X0Y0_S2MID[6] net44 VPWR VGND sg13g2_buf_1
X_3531_ VGND VPWR _1565_ _1567_ _1577_ _1576_ sg13g2_a21oi_1
Xinput88 Tile_X0Y1_E1END[1] net88 VPWR VGND sg13g2_buf_1
Xinput66 Tile_X0Y0_W2END[1] net66 VPWR VGND sg13g2_buf_1
Xinput77 Tile_X0Y0_W2MID[4] net77 VPWR VGND sg13g2_buf_1
Xinput99 Tile_X0Y1_E2MID[0] net99 VPWR VGND sg13g2_buf_1
X_6250_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 net471 VPWR VGND sg13g2_buf_1
X_3462_ VPWR _1511_ _1510_ VGND sg13g2_inv_1
X_6181_ Tile_X0Y1_E6END[10] net404 VPWR VGND sg13g2_buf_1
X_3393_ _1445_ _1410_ _1411_ VPWR VGND sg13g2_xnor2_1
X_5201_ net1940 net1766 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_5132_ net1991 net1785 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_69_345 VPWR VGND sg13g2_fill_1
XFILLER_84_304 VPWR VGND sg13g2_fill_2
X_5063_ net1982 net1809 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_4014_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q VPWR _2019_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q _2017_ sg13g2_o21ai_1
Xfanout1890 net1891 net1890 VPWR VGND sg13g2_buf_1
X_5965_ net13 net186 VPWR VGND sg13g2_buf_1
X_4916_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X
+ net707 VGND sg13g2_inv_1
X_4847_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q _0394_ _0395_
+ VPWR VGND sg13g2_nor2_1
XFILLER_32_38 VPWR VGND sg13g2_fill_1
XFILLER_20_175 VPWR VGND sg13g2_fill_1
X_4778_ VGND VPWR _0069_ net1692 _0329_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ sg13g2_a21oi_1
X_3729_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q _1760_
+ _1761_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q sg13g2_a21oi_1
XFILLER_121_239 VPWR VGND sg13g2_fill_2
XFILLER_75_348 VPWR VGND sg13g2_fill_2
XFILLER_90_318 VPWR VGND sg13g2_fill_1
XFILLER_98_86 VPWR VGND sg13g2_fill_2
XFILLER_34_201 VPWR VGND sg13g2_decap_8
X_5750_ net1903 net1725 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_2962_ _1025_ net1575 _1023_ VPWR VGND sg13g2_nand2_1
X_5681_ net1890 net1749 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_4701_ VGND VPWR net57 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q
+ _0254_ _0253_ sg13g2_a21oi_1
X_2893_ _0961_ VPWR _0962_ VGND net154 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q
+ sg13g2_o21ai_1
X_4632_ _0188_ VPWR _0189_ VGND net69 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q
+ sg13g2_o21ai_1
X_4563_ VPWR _0120_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q VGND
+ sg13g2_inv_1
X_6302_ net164 net523 VPWR VGND sg13g2_buf_1
X_3514_ _1560_ net1671 _0682_ VPWR VGND sg13g2_nand2_1
X_4494_ net1514 _2055_ _0051_ VPWR VGND sg13g2_nor2b_1
X_3445_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q VPWR _1496_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q _1495_ sg13g2_o21ai_1
X_6233_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 net454 VPWR VGND sg13g2_buf_8
X_6164_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 net385 VPWR VGND sg13g2_buf_8
X_3376_ _1104_ net1548 _1428_ VPWR VGND sg13g2_nor2_2
X_5115_ net1954 net1788 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_6095_ Tile_X0Y1_NN4END[15] net322 VPWR VGND sg13g2_buf_1
X_5046_ net1949 net1851 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_72_318 VPWR VGND sg13g2_fill_1
X_5879_ net1904 net1812 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_52 VPWR VGND sg13g2_fill_1
XFILLER_75_123 VPWR VGND sg13g2_fill_2
XFILLER_75_145 VPWR VGND sg13g2_fill_2
XFILLER_84_99 VPWR VGND sg13g2_fill_2
XFILLER_16_289 VPWR VGND sg13g2_fill_1
XFILLER_71_384 VPWR VGND sg13g2_fill_1
X_3230_ _1282_ net1515 _1283_ VPWR VGND sg13g2_nor2_2
X_3161_ _1216_ _1105_ _1215_ VPWR VGND sg13g2_nand2_1
X_3092_ _1149_ _1148_ _0518_ VPWR VGND sg13g2_nand2b_1
X_5802_ net1876 net1833 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_3994_ VGND VPWR _1998_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q
+ _1995_ _0158_ _1999_ _1993_ sg13g2_a221oi_1
XFILLER_13_18 VPWR VGND sg13g2_fill_1
X_5733_ net1875 net1737 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_2945_ _1009_ _0931_ _0932_ VPWR VGND sg13g2_xnor2_1
X_5664_ net1861 net1761 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_2876_ VGND VPWR _0945_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q
+ _0944_ _0113_ _0946_ _0943_ sg13g2_a221oi_1
X_4615_ _0172_ net1563 VPWR VGND sg13g2_inv_8
X_5595_ net1912 net1781 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_4546_ VPWR _0103_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q VGND
+ sg13g2_inv_1
X_4477_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q _2390_ _2391_
+ VPWR VGND sg13g2_nor2b_1
X_6216_ net1907 net428 VPWR VGND sg13g2_buf_1
X_3428_ VGND VPWR net76 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q
+ _1479_ _1478_ sg13g2_a21oi_1
X_6147_ Tile_X0Y0_WW4END[14] net359 VPWR VGND sg13g2_buf_1
X_3359_ _1411_ _1389_ _1390_ VPWR VGND sg13g2_xnor2_1
X_6078_ Tile_X0Y1_N4END[14] net305 VPWR VGND sg13g2_buf_1
X_5029_ net1976 net1851 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_54_36 VPWR VGND sg13g2_decap_4
XFILLER_70_24 VPWR VGND sg13g2_fill_2
XFILLER_21_281 VPWR VGND sg13g2_fill_1
XFILLER_107_353 VPWR VGND sg13g2_fill_2
XFILLER_95_21 VPWR VGND sg13g2_fill_1
XFILLER_95_229 VPWR VGND sg13g2_decap_8
XFILLER_36_318 VPWR VGND sg13g2_fill_2
XFILLER_44_384 VPWR VGND sg13g2_fill_1
X_2730_ Tile_X0Y1_DSP_bot.A3 Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[3\] net1641 _0807_
+ VPWR VGND sg13g2_mux2_2
X_2661_ _0124_ _0730_ _0740_ _0742_ VPWR VGND sg13g2_nor3_1
X_4400_ _2324_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q _1674_
+ VPWR VGND sg13g2_nand2_1
X_5380_ net1973 net1827 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_2592_ net1926 net95 net1659 _0677_ VPWR VGND sg13g2_mux2_1
Xoutput527 net527 Tile_X0Y1_W6BEG[10] VPWR VGND sg13g2_buf_1
Xoutput516 net516 Tile_X0Y1_W2BEG[6] VPWR VGND sg13g2_buf_1
Xoutput505 net505 Tile_X0Y1_SS4BEG[9] VPWR VGND sg13g2_buf_8
X_4331_ _2264_ VPWR _2265_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q
+ _1277_ sg13g2_o21ai_1
Xoutput538 net538 Tile_X0Y1_WW4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput549 net549 Tile_X0Y1_WW4BEG[5] VPWR VGND sg13g2_buf_1
X_4262_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q _2219_
+ _2220_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q sg13g2_a21oi_1
X_3213_ _1266_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q _1267_
+ _1268_ VPWR VGND sg13g2_a21o_1
X_6001_ net1978 net232 VPWR VGND sg13g2_buf_1
X_4193_ _1470_ net623 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q
+ _2161_ VPWR VGND sg13g2_mux2_1
X_3144_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q VPWR _1200_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q net165 sg13g2_o21ai_1
X_3075_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q VPWR _1134_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q _1133_ sg13g2_o21ai_1
XFILLER_50_310 VPWR VGND sg13g2_fill_2
X_5454__586 VPWR VGND net586 sg13g2_tiehi
X_3977_ _1982_ _1981_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X VPWR
+ VGND sg13g2_mux2_1
X_5716_ net1899 net1737 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_2928_ _0106_ _0989_ _0994_ VPWR VGND sg13g2_nor2_2
X_5647_ net1887 net1761 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_2859_ _0928_ _0929_ VPWR VGND sg13g2_inv_4
X_5578_ net1876 net1782 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_4529_ VPWR _0086_ net36 VGND sg13g2_inv_1
XFILLER_77_229 VPWR VGND sg13g2_fill_1
Xfanout1719 net1720 net1719 VPWR VGND sg13g2_buf_1
Xfanout1708 net127 net1708 VPWR VGND sg13g2_buf_1
XFILLER_105_75 VPWR VGND sg13g2_decap_4
XFILLER_81_45 VPWR VGND sg13g2_fill_1
XFILLER_5_255 VPWR VGND sg13g2_fill_2
XFILLER_30_60 VPWR VGND sg13g2_decap_4
XFILLER_107_161 VPWR VGND sg13g2_fill_2
XFILLER_36_126 VPWR VGND sg13g2_fill_1
Xinput9 Tile_X0Y0_E2END[5] net9 VPWR VGND sg13g2_buf_1
X_4880_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q _0426_
+ _0427_ _0078_ sg13g2_a21oi_1
X_3900_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q _1913_
+ _1914_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q sg13g2_a21oi_1
X_3831_ _1848_ _1859_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 VPWR VGND
+ sg13g2_nor2_2
XFILLER_32_343 VPWR VGND sg13g2_fill_2
X_3762_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q net122 net109
+ net1934 net158 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q _1792_
+ VPWR VGND sg13g2_mux4_1
X_5501_ net1917 net1846 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_3693_ VGND VPWR _1726_ _1727_ _0015_ net1643 sg13g2_a21oi_2
X_2713_ _0791_ VPWR _0792_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q
+ _0786_ sg13g2_o21ai_1
X_5432_ Tile_X0Y1_UserCLK net566 _0046_ _0008_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[8\]
+ VPWR VGND sg13g2_dfrbp_1
X_2644_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q net645 _0724_
+ _0099_ _0105_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q _0725_
+ VPWR VGND sg13g2_mux4_1
Xoutput313 net313 Tile_X0Y0_NN4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput302 net302 Tile_X0Y0_N4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput324 net324 Tile_X0Y0_NN4BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_58_0 VPWR VGND sg13g2_decap_4
Xoutput335 net335 Tile_X0Y0_W2BEG[5] VPWR VGND sg13g2_buf_1
X_2575_ _0660_ VPWR _0661_ VGND net67 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q
+ sg13g2_o21ai_1
X_5363_ net1943 net1843 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_4314_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q net1534 net1542
+ net1549 net1557 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q _2252_
+ VPWR VGND sg13g2_mux4_1
Xoutput368 net368 Tile_X0Y0_WW4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput346 net346 Tile_X0Y0_W6BEG[0] VPWR VGND sg13g2_buf_1
Xoutput357 net357 Tile_X0Y0_W6BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_99_354 VPWR VGND sg13g2_fill_1
Xoutput379 net379 Tile_X0Y1_E2BEG[1] VPWR VGND sg13g2_buf_1
X_5294_ net1995 net1733 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_4245_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 _2202_ _2205_ _2198_
+ _2200_ VPWR VGND sg13g2_a22oi_1
X_4176_ _2144_ _2145_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 VPWR VGND sg13g2_mux2_1
X_3127_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q VPWR _1184_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q _1182_ sg13g2_o21ai_1
XFILLER_42_118 VPWR VGND sg13g2_fill_2
X_3058_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q _0178_
+ _1118_ _1117_ sg13g2_a21oi_1
Xfanout1516 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 net1516 VPWR VGND
+ sg13g2_buf_8
Xfanout1527 _0376_ net1527 VPWR VGND sg13g2_buf_1
XFILLER_104_175 VPWR VGND sg13g2_decap_8
Xfanout1549 net1549 net1551 VPWR VGND sg13g2_buf_16
XFILLER_41_81 VPWR VGND sg13g2_fill_2
X_4030_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q VPWR _2034_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q _2032_ sg13g2_o21ai_1
XFILLER_110_178 VPWR VGND sg13g2_fill_1
X_5981_ Tile_X0Y0_E6END[11] net204 VPWR VGND sg13g2_buf_1
X_4932_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q net1921 net152
+ net59 net1703 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q _0476_
+ VPWR VGND sg13g2_mux4_1
XFILLER_32_162 VPWR VGND sg13g2_fill_2
X_4863_ net647 _0385_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q
+ _0410_ VPWR VGND sg13g2_mux2_1
XFILLER_20_357 VPWR VGND sg13g2_fill_1
X_4794_ _0344_ VPWR _0345_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ _0342_ sg13g2_o21ai_1
X_3814_ _1840_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q _1843_
+ VPWR VGND sg13g2_nor2b_1
X_3745_ _1775_ VPWR _1776_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 sg13g2_o21ai_1
X_3676_ _1711_ _1444_ _1445_ VPWR VGND sg13g2_xnor2_1
X_5415_ net1982 net1817 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_2627_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q VPWR _0709_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q _0706_ sg13g2_o21ai_1
X_2558_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q VPWR _0644_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q _0643_ sg13g2_o21ai_1
X_5346_ net1969 net1842 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput176 net176 Tile_X0Y0_E1BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_99_140 VPWR VGND sg13g2_decap_8
X_2489_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q _0578_ _0579_
+ VPWR VGND sg13g2_nor2_1
X_5277_ net1960 net1732 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_99_184 VPWR VGND sg13g2_fill_2
Xoutput187 net187 Tile_X0Y0_E2BEGb[2] VPWR VGND sg13g2_buf_1
Xoutput198 net198 Tile_X0Y0_E6BEG[3] VPWR VGND sg13g2_buf_1
X_4228_ _2190_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q _0630_
+ VPWR VGND sg13g2_nand2_1
XFILLER_87_368 VPWR VGND sg13g2_fill_1
X_4159_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q _2130_
+ _2131_ _0161_ sg13g2_a21oi_1
Xfanout2003 net3 net2003 VPWR VGND sg13g2_buf_1
XFILLER_87_55 VPWR VGND sg13g2_fill_1
XFILLER_61_202 VPWR VGND sg13g2_fill_2
Xinput12 Tile_X0Y0_E2MID[0] net12 VPWR VGND sg13g2_buf_1
Xinput34 Tile_X0Y0_S2END[4] net34 VPWR VGND sg13g2_buf_1
Xinput45 Tile_X0Y0_S2MID[7] net45 VPWR VGND sg13g2_buf_1
X_3530_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q VPWR _1576_ VGND
+ _1569_ _1575_ sg13g2_o21ai_1
Xinput23 Tile_X0Y0_EE4END[1] net23 VPWR VGND sg13g2_buf_1
Xinput56 Tile_X0Y0_SS4END[2] net56 VPWR VGND sg13g2_buf_1
Xinput89 Tile_X0Y1_E1END[2] net89 VPWR VGND sg13g2_buf_1
Xinput67 Tile_X0Y0_W2END[2] net67 VPWR VGND sg13g2_buf_8
Xinput78 Tile_X0Y0_W2MID[5] net78 VPWR VGND sg13g2_buf_1
X_3461_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q net138 net7 net68
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q
+ _1510_ VPWR VGND sg13g2_mux4_1
X_6180_ Tile_X0Y1_E6END[9] net403 VPWR VGND sg13g2_buf_1
X_3392_ _1425_ VPWR _1444_ VGND _1441_ _1442_ sg13g2_o21ai_1
X_5200_ net1937 net1766 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_123_281 VPWR VGND sg13g2_fill_2
X_5131_ net1989 net1785 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_35_2 VPWR VGND sg13g2_fill_1
X_5062_ net1980 net1809 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_69_368 VPWR VGND sg13g2_fill_1
XFILLER_96_132 VPWR VGND sg13g2_fill_2
X_4013_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q net1632 net1586
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 net1539 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q
+ _2018_ VPWR VGND sg13g2_mux4_1
XFILLER_96_176 VPWR VGND sg13g2_decap_8
Xfanout1891 Tile_X0Y1_FrameData[22] net1891 VPWR VGND sg13g2_buf_1
Xfanout1880 net1881 net1880 VPWR VGND sg13g2_buf_1
X_5964_ net12 net185 VPWR VGND sg13g2_buf_1
X_5895_ net1920 net1816 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_4915_ VGND VPWR _0259_ _0460_ _0440_ _0459_ sg13g2_a21oi_2
X_4846_ net1597 net1611 net1685 _0394_ VPWR VGND sg13g2_mux2_1
X_4777_ _0326_ VPWR _0328_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q
+ _0292_ sg13g2_o21ai_1
X_3728_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q net128 net104
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 net164 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q
+ _1760_ VPWR VGND sg13g2_mux4_1
X_3659_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q net140 net96
+ net43 net156 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q _1695_
+ VPWR VGND sg13g2_mux4_1
XFILLER_106_226 VPWR VGND sg13g2_decap_8
XFILLER_106_237 VPWR VGND sg13g2_fill_1
XFILLER_106_259 VPWR VGND sg13g2_fill_2
X_5329_ net1940 net1720 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_43_235 VPWR VGND sg13g2_decap_8
XFILLER_98_21 VPWR VGND sg13g2_fill_2
XFILLER_34_224 VPWR VGND sg13g2_fill_1
X_2961_ VPWR _1024_ _1023_ VGND sg13g2_inv_1
X_5680_ net1888 net1749 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_4700_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q net7 _0253_ VPWR
+ VGND sg13g2_nor2b_1
X_2892_ _0961_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q net170
+ VPWR VGND sg13g2_nand2b_1
X_4631_ _0188_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q net1929
+ VPWR VGND sg13g2_nand2b_1
X_4562_ VPWR _0119_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q VGND
+ sg13g2_inv_1
X_6301_ net163 net522 VPWR VGND sg13g2_buf_1
X_3513_ VPWR _1559_ net717 VGND sg13g2_inv_1
X_4493_ net1513 _1898_ _0050_ VPWR VGND sg13g2_nor2_1
X_3444_ _1494_ VPWR _1495_ VGND _0070_ net1687 sg13g2_o21ai_1
X_6232_ net1871 net446 VPWR VGND sg13g2_buf_1
X_6163_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 net384 VPWR VGND sg13g2_buf_1
X_3375_ _1427_ _1103_ net1568 VPWR VGND sg13g2_nand2_2
X_5114_ net1952 net1786 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_6094_ Tile_X0Y1_NN4END[14] net321 VPWR VGND sg13g2_buf_1
X_5045_ net1947 net1851 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_39 VPWR VGND sg13g2_fill_2
XFILLER_65_371 VPWR VGND sg13g2_fill_1
X_5878_ net1902 net1812 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_4829_ _0377_ VPWR _0378_ VGND net1683 net1527 sg13g2_o21ai_1
XFILLER_102_251 VPWR VGND sg13g2_decap_8
XFILLER_56_382 VPWR VGND sg13g2_fill_2
X_3160_ _0848_ _1214_ _1215_ VPWR VGND sg13g2_nor2_1
X_3091_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[2\] Tile_X0Y1_DSP_bot.B2 net1640 _1148_
+ VPWR VGND sg13g2_mux2_1
XFILLER_66_113 VPWR VGND sg13g2_fill_1
XFILLER_54_308 VPWR VGND sg13g2_fill_1
X_5801_ net1872 net1833 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_5732_ net1869 net1737 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_3993_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q _1997_
+ _1998_ _0158_ sg13g2_a21oi_1
X_2944_ _1008_ _0973_ _1006_ VPWR VGND sg13g2_nand2_2
XFILLER_88_0 VPWR VGND sg13g2_fill_2
X_2875_ VGND VPWR net9 net1686 _0945_ _0113_ sg13g2_a21oi_1
X_5663_ net1859 net1762 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_5594_ net1910 net1781 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_4614_ VPWR _0171_ net1558 VGND sg13g2_inv_1
X_4545_ VPWR _0102_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q VGND
+ sg13g2_inv_1
X_4476_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q net1707 net99
+ net105 net642 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q _2390_
+ VPWR VGND sg13g2_mux4_1
X_6215_ net1909 net427 VPWR VGND sg13g2_buf_1
X_3427_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q VPWR _1478_ VGND
+ _0068_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q sg13g2_o21ai_1
X_6146_ Tile_X0Y0_WW4END[13] net373 VPWR VGND sg13g2_buf_1
X_3358_ _1406_ _1409_ _1410_ VPWR VGND sg13g2_nor2_2
XFILLER_97_282 VPWR VGND sg13g2_fill_2
X_6077_ Tile_X0Y1_N4END[13] net304 VPWR VGND sg13g2_buf_1
XFILLER_57_168 VPWR VGND sg13g2_fill_2
X_3289_ _1341_ _1337_ _1338_ VPWR VGND sg13g2_xnor2_1
X_5028_ net1974 net1851 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_65_190 VPWR VGND sg13g2_fill_2
XFILLER_13_205 VPWR VGND sg13g2_fill_1
XFILLER_70_58 VPWR VGND sg13g2_fill_2
XFILLER_107_310 VPWR VGND sg13g2_fill_1
XFILLER_119_96 VPWR VGND sg13g2_fill_1
XFILLER_0_164 VPWR VGND sg13g2_fill_1
XFILLER_48_146 VPWR VGND sg13g2_decap_8
XFILLER_95_99 VPWR VGND sg13g2_fill_1
XFILLER_28_82 VPWR VGND sg13g2_fill_1
XFILLER_63_127 VPWR VGND sg13g2_fill_1
XFILLER_8_253 VPWR VGND sg13g2_fill_2
X_2660_ VGND VPWR _0741_ _0740_ _0730_ sg13g2_or2_1
Xoutput506 net506 Tile_X0Y1_W1BEG[0] VPWR VGND sg13g2_buf_1
X_2591_ VGND VPWR _0058_ net1658 _0676_ _0675_ sg13g2_a21oi_1
Xoutput517 net517 Tile_X0Y1_W2BEG[7] VPWR VGND sg13g2_buf_1
X_4330_ _0166_ _2263_ _2264_ VPWR VGND sg13g2_nor2_1
Xoutput539 net539 Tile_X0Y1_WW4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput528 net528 Tile_X0Y1_W6BEG[11] VPWR VGND sg13g2_buf_1
X_4261_ VPWR _2219_ _2218_ VGND sg13g2_inv_1
X_3212_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q VPWR _1267_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q _1265_ sg13g2_o21ai_1
X_6000_ net2000 net221 VPWR VGND sg13g2_buf_1
XFILLER_79_271 VPWR VGND sg13g2_fill_2
X_4192_ _0630_ _0868_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q
+ _2160_ VPWR VGND sg13g2_mux2_1
X_3143_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q _1197_ _1198_
+ _1199_ VPWR VGND sg13g2_nor3_1
X_3074_ net1561 net1570 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q
+ _1133_ VPWR VGND sg13g2_mux2_1
XFILLER_50_322 VPWR VGND sg13g2_fill_2
XFILLER_50_366 VPWR VGND sg13g2_fill_1
X_3976_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q
+ _1982_ VPWR VGND sg13g2_mux4_1
X_5715_ net1894 net1736 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_2927_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q VPWR _0993_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q _0990_ sg13g2_o21ai_1
XFILLER_40_17 VPWR VGND sg13g2_fill_2
X_5646_ net1885 net1761 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_2858_ _0927_ VPWR _0928_ VGND Tile_X0Y1_DSP_bot.A2 net1641 sg13g2_o21ai_1
X_2789_ _0863_ VPWR _0864_ VGND net1933 net1690 sg13g2_o21ai_1
X_5577_ net1872 net1782 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_4528_ VPWR _0085_ net164 VGND sg13g2_inv_1
X_4459_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q net1926 net1705
+ net1528 net1535 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q _2374_
+ VPWR VGND sg13g2_mux4_1
Xfanout1709 net123 net1709 VPWR VGND sg13g2_buf_1
X_6129_ Tile_X0Y0_W6END[6] net352 VPWR VGND sg13g2_buf_1
XFILLER_65_36 VPWR VGND sg13g2_fill_1
XFILLER_45_138 VPWR VGND sg13g2_fill_1
XFILLER_60_108 VPWR VGND sg13g2_decap_8
XFILLER_60_119 VPWR VGND sg13g2_fill_2
XFILLER_36_138 VPWR VGND sg13g2_fill_1
XFILLER_91_277 VPWR VGND sg13g2_fill_1
X_3830_ VGND VPWR _1858_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q
+ _1855_ _1850_ _1859_ _1853_ sg13g2_a221oi_1
X_3761_ _1791_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q _1790_
+ VPWR VGND sg13g2_nand2_1
X_5500_ net1915 net1845 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_2712_ _0790_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q _0791_
+ VPWR VGND sg13g2_nor2b_1
X_3692_ net1643 Tile_X0Y1_DSP_bot.C5 _1726_ VPWR VGND sg13g2_nor2_2
X_5431_ Tile_X0Y1_UserCLK net567 _0045_ _0010_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[7\]
+ VPWR VGND sg13g2_dfrbp_1
X_2643_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q _0175_ _0384_
+ _0698_ _0722_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q _0724_
+ VPWR VGND sg13g2_mux4_1
Xoutput325 net325 Tile_X0Y0_UserCLKo VPWR VGND sg13g2_buf_1
Xoutput303 net303 Tile_X0Y0_N4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput314 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 Tile_X0Y0_NN4BEG[14]
+ VPWR VGND sg13g2_buf_1
X_2574_ _0660_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q net86 VPWR
+ VGND sg13g2_nand2b_1
X_5362_ net1942 net1843 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_4313_ _2251_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q _2250_
+ VPWR VGND sg13g2_nand2_1
Xoutput336 net336 Tile_X0Y0_W2BEG[6] VPWR VGND sg13g2_buf_1
Xoutput358 net358 Tile_X0Y0_WW4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput369 net369 Tile_X0Y0_WW4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput347 net347 Tile_X0Y0_W6BEG[10] VPWR VGND sg13g2_buf_1
XFILLER_99_333 VPWR VGND sg13g2_fill_1
X_5293_ net1994 net1732 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_338 VPWR VGND sg13g2_fill_2
X_4244_ _2204_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q _2205_
+ VPWR VGND sg13g2_nor2b_1
X_4175_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q net1540 _1470_
+ net623 _0974_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q _2145_
+ VPWR VGND sg13g2_mux4_1
XFILLER_67_241 VPWR VGND sg13g2_fill_1
X_3126_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q net1634 net1523
+ net1593 net1540 net1691 _1183_ VPWR VGND sg13g2_mux4_1
X_3057_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q VPWR _1117_ VGND
+ net1668 net1582 sg13g2_o21ai_1
X_3959_ _1967_ VPWR _1968_ VGND net37 net1700 sg13g2_o21ai_1
X_5629_ net1917 net1771 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_4_6 VPWR VGND sg13g2_fill_1
XFILLER_104_110 VPWR VGND sg13g2_fill_2
Xfanout1539 net1539 net1540 VPWR VGND sg13g2_buf_16
Xfanout1517 _1724_ net1517 VPWR VGND sg13g2_buf_1
Xfanout1528 net1530 net1528 VPWR VGND sg13g2_buf_8
XFILLER_104_187 VPWR VGND sg13g2_decap_8
XFILLER_18_105 VPWR VGND sg13g2_fill_1
XFILLER_73_222 VPWR VGND sg13g2_decap_8
XFILLER_73_233 VPWR VGND sg13g2_fill_1
Xrebuffer90 net1541 net699 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_25_50 VPWR VGND sg13g2_fill_2
XFILLER_44_7 VPWR VGND sg13g2_fill_1
X_5980_ Tile_X0Y0_E6END[10] net203 VPWR VGND sg13g2_buf_1
X_4931_ _0475_ _0474_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q
+ VPWR VGND sg13g2_nand2b_1
X_4862_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 _0409_ _0402_ _0397_ _0391_
+ VPWR VGND sg13g2_a22oi_1
XFILLER_32_174 VPWR VGND sg13g2_decap_8
X_3813_ _1842_ _1841_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q
+ VPWR VGND sg13g2_nand2b_1
X_4793_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q _0343_
+ _0344_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q sg13g2_a21oi_1
X_3744_ _1775_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q net162
+ VPWR VGND sg13g2_nand2b_1
XFILLER_70_0 VPWR VGND sg13g2_fill_1
X_3675_ VPWR _1710_ _1709_ VGND sg13g2_inv_1
X_2626_ _0707_ VPWR _0708_ VGND net1675 net1522 sg13g2_o21ai_1
X_5414_ net1980 net1817 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_2557_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q net1599 net1613
+ net1606 net1626 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q _0643_
+ VPWR VGND sg13g2_mux4_1
X_5345_ net1968 net1840 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput177 net177 Tile_X0Y0_E2BEG[0] VPWR VGND sg13g2_buf_1
Xoutput199 net199 Tile_X0Y0_E6BEG[4] VPWR VGND sg13g2_buf_1
X_5276_ net1957 net1733 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_2488_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q _0574_
+ _0578_ _0577_ sg13g2_a21oi_1
Xoutput188 net188 Tile_X0Y0_E2BEGb[3] VPWR VGND sg13g2_buf_1
X_4227_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q _0598_ net1931
+ net29 net1622 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q _2189_
+ VPWR VGND sg13g2_mux4_1
XFILLER_101_157 VPWR VGND sg13g2_fill_1
XFILLER_46_38 VPWR VGND sg13g2_fill_1
X_4158_ _2129_ VPWR _2130_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q
+ _0868_ sg13g2_o21ai_1
X_3109_ _1166_ _0702_ _0899_ VPWR VGND sg13g2_nand2_2
X_4089_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q net1633 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1
+ net694 _0647_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2
+ VPWR VGND sg13g2_mux4_1
XFILLER_70_225 VPWR VGND sg13g2_fill_2
XFILLER_102_77 VPWR VGND sg13g2_decap_4
XFILLER_109_246 VPWR VGND sg13g2_decap_8
Xfanout2004 net2 net2004 VPWR VGND sg13g2_buf_1
XFILLER_78_358 VPWR VGND sg13g2_fill_1
XFILLER_14_152 VPWR VGND sg13g2_fill_1
Xinput13 Tile_X0Y0_E2MID[1] net13 VPWR VGND sg13g2_buf_1
Xinput46 Tile_X0Y0_S4END[0] net46 VPWR VGND sg13g2_buf_1
Xinput35 Tile_X0Y0_S2END[5] net35 VPWR VGND sg13g2_buf_1
Xinput24 Tile_X0Y0_EE4END[2] net24 VPWR VGND sg13g2_buf_1
Xinput57 Tile_X0Y0_SS4END[3] net57 VPWR VGND sg13g2_buf_1
Xinput79 Tile_X0Y0_W2MID[6] net79 VPWR VGND sg13g2_buf_1
Xinput68 Tile_X0Y0_W2END[3] net68 VPWR VGND sg13g2_buf_1
X_3460_ _1453_ _1508_ _1509_ VPWR VGND sg13g2_nor2b_2
X_3391_ _1443_ _1423_ _1424_ VPWR VGND sg13g2_xnor2_1
X_5130_ net1987 net1786 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_5061_ net1975 net1808 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_4012_ VPWR _2017_ _2016_ VGND sg13g2_inv_1
Xfanout1870 Tile_X0Y1_FrameData[31] net1870 VPWR VGND sg13g2_buf_1
XFILLER_84_328 VPWR VGND sg13g2_fill_2
Xfanout1881 Tile_X0Y1_FrameData[27] net1881 VPWR VGND sg13g2_buf_1
Xfanout1892 net1893 net1892 VPWR VGND sg13g2_buf_1
XFILLER_77_380 VPWR VGND sg13g2_fill_1
X_5963_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 net184 VPWR VGND sg13g2_buf_8
X_4914_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q _0458_ _0459_
+ VPWR VGND sg13g2_nor2_1
X_5894_ net1897 net1816 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_4845_ VGND VPWR net1685 net1633 _0393_ _0392_ sg13g2_a21oi_1
X_4776_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q net1543 _0289_
+ net710 _0308_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q _0327_
+ VPWR VGND sg13g2_mux4_1
X_3727_ _1758_ _1759_ VPWR VGND sg13g2_inv_4
X_3658_ _1694_ _1693_ _1692_ VPWR VGND sg13g2_nand2b_1
X_3589_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q _1629_
+ _1630_ _0148_ sg13g2_a21oi_1
X_2609_ _0691_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q _0692_
+ _0693_ VPWR VGND sg13g2_a21o_1
XFILLER_87_111 VPWR VGND sg13g2_fill_2
X_5328_ net1938 net1719 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_114_282 VPWR VGND sg13g2_fill_2
XFILLER_57_48 VPWR VGND sg13g2_fill_2
X_5259_ net1989 net1745 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_118_0 VPWR VGND sg13g2_fill_2
XFILLER_0_0 VPWR VGND sg13g2_fill_1
XFILLER_78_122 VPWR VGND sg13g2_decap_4
X_5476__608 VPWR VGND net608 sg13g2_tiehi
XFILLER_19_299 VPWR VGND sg13g2_fill_1
XFILLER_74_383 VPWR VGND sg13g2_fill_2
X_2960_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[5\] net1642 _1023_ VPWR VGND sg13g2_mux2_2
X_2891_ VGND VPWR _0068_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q
+ _0960_ _0959_ sg13g2_a21oi_1
X_4630_ net34 net46 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q _0187_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_75 VPWR VGND sg13g2_fill_1
X_4561_ VPWR _0118_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q VGND
+ sg13g2_inv_1
X_6300_ net162 net521 VPWR VGND sg13g2_buf_1
X_3512_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 _1558_ _1556_ _1550_
+ _1549_ VPWR VGND sg13g2_a22oi_1
X_4492_ net1513 _1897_ _0049_ VPWR VGND sg13g2_nor2b_1
X_3443_ _1494_ net28 net1687 VPWR VGND sg13g2_nand2_1
XFILLER_6_192 VPWR VGND sg13g2_fill_2
X_6231_ net1873 net445 VPWR VGND sg13g2_buf_1
X_6162_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 net383 VPWR VGND sg13g2_buf_1
X_3374_ _1418_ _1413_ _1426_ VPWR VGND sg13g2_xor2_1
X_5113_ net1999 net1796 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_6093_ Tile_X0Y1_NN4END[13] net320 VPWR VGND sg13g2_buf_1
XFILLER_111_296 VPWR VGND sg13g2_fill_2
X_5044_ net1945 net1851 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_5877_ net1900 net1813 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_4828_ VGND VPWR _0074_ net1683 _0377_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q
+ sg13g2_a21oi_1
X_4759_ _0310_ _0067_ _0309_ VPWR VGND sg13g2_nand2b_1
XFILLER_75_125 VPWR VGND sg13g2_fill_1
X_3090_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q _1130_ _1131_
+ _1147_ _1146_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q Tile_X0Y1_DSP_bot.B2
+ VPWR VGND sg13g2_mux4_1
XFILLER_81_128 VPWR VGND sg13g2_fill_1
X_5800_ net1870 net1833 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_3992_ VGND VPWR net62 net1701 _1997_ _1996_ sg13g2_a21oi_1
X_5731_ net1866 net1735 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_2943_ VPWR _1007_ _1006_ VGND sg13g2_inv_1
X_5662_ net1857 net1762 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_2874_ _0944_ net2004 net1686 VPWR VGND sg13g2_nand2b_1
X_5593_ net1908 net1781 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_4613_ VPWR _0170_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q VGND
+ sg13g2_inv_1
X_4544_ VPWR _0101_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q VGND
+ sg13g2_inv_1
X_6214_ net1911 net426 VPWR VGND sg13g2_buf_1
X_4475_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q VPWR _2389_ VGND
+ _2385_ _2388_ sg13g2_o21ai_1
X_3426_ VGND VPWR _1473_ _1476_ _1472_ _0000_ _1477_ net1650 sg13g2_a221oi_1
X_3357_ _1407_ _1408_ _1409_ VPWR VGND sg13g2_nor2b_1
X_6145_ Tile_X0Y0_WW4END[12] net372 VPWR VGND sg13g2_buf_1
X_6076_ Tile_X0Y1_N4END[12] net303 VPWR VGND sg13g2_buf_1
XFILLER_57_103 VPWR VGND sg13g2_fill_1
X_3288_ _1332_ _1309_ _1334_ _1340_ VPWR VGND sg13g2_a21o_1
X_5027_ net1971 net1852 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_72_139 VPWR VGND sg13g2_fill_1
XFILLER_53_364 VPWR VGND sg13g2_fill_2
XFILLER_80_194 VPWR VGND sg13g2_decap_8
XFILLER_119_75 VPWR VGND sg13g2_fill_2
XFILLER_122_303 VPWR VGND sg13g2_fill_2
XFILLER_88_261 VPWR VGND sg13g2_decap_4
XFILLER_88_283 VPWR VGND sg13g2_fill_2
XFILLER_63_139 VPWR VGND sg13g2_decap_4
XFILLER_60_70 VPWR VGND sg13g2_fill_1
X_2590_ net155 net1658 _0675_ VPWR VGND sg13g2_nor2_1
Xoutput507 net507 Tile_X0Y1_W1BEG[1] VPWR VGND sg13g2_buf_1
Xoutput518 net518 Tile_X0Y1_W2BEGb[0] VPWR VGND sg13g2_buf_1
XFILLER_5_10 VPWR VGND sg13g2_fill_1
Xoutput529 net529 Tile_X0Y1_W6BEG[1] VPWR VGND sg13g2_buf_1
X_4260_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q net649 net1632
+ net1624 net1591 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q _2218_
+ VPWR VGND sg13g2_mux4_1
X_3211_ net1582 net1619 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q
+ _1266_ VPWR VGND sg13g2_mux2_1
X_4191_ _2158_ VPWR _2159_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q
+ _2155_ sg13g2_o21ai_1
X_3142_ net1707 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q _1198_
+ VPWR VGND sg13g2_nor2_1
X_3073_ net1579 net1616 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q
+ _1132_ VPWR VGND sg13g2_mux2_1
XFILLER_54_117 VPWR VGND sg13g2_fill_2
X_3975_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 _0646_ net727 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q
+ _1981_ VPWR VGND sg13g2_mux4_1
X_5714_ net1892 net1735 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_2926_ VGND VPWR net1661 _0178_ _0992_ _0991_ sg13g2_a21oi_1
X_5645_ net1883 net1760 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_2857_ _0927_ net1641 Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[2\] VPWR VGND sg13g2_nand2b_1
X_2788_ _0863_ net1690 net1930 VPWR VGND sg13g2_nand2b_1
X_5576_ net1870 net1782 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_4527_ VPWR _0084_ net104 VGND sg13g2_inv_1
X_4458_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q _2366_ _2367_
+ _2373_ _2372_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0
+ VPWR VGND sg13g2_mux4_1
X_3409_ _1461_ _1458_ _1460_ VPWR VGND sg13g2_nand2b_1
X_6128_ Tile_X0Y0_W6END[5] net351 VPWR VGND sg13g2_buf_1
X_4389_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q _0905_ _1130_
+ _1759_ _1699_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q _2314_
+ VPWR VGND sg13g2_mux4_1
XFILLER_85_231 VPWR VGND sg13g2_fill_1
X_6059_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 net280 VPWR VGND sg13g2_buf_1
XFILLER_14_41 VPWR VGND sg13g2_fill_1
XFILLER_100_0 VPWR VGND sg13g2_fill_2
XFILLER_122_166 VPWR VGND sg13g2_fill_1
XFILLER_36_117 VPWR VGND sg13g2_decap_8
XFILLER_32_345 VPWR VGND sg13g2_fill_1
XFILLER_32_356 VPWR VGND sg13g2_fill_2
X_3760_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q net134 net94
+ net154 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q
+ _1790_ VPWR VGND sg13g2_mux4_1
X_2711_ VGND VPWR _0789_ _0790_ _0788_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q
+ sg13g2_a21oi_2
X_3691_ VGND VPWR _1725_ Tile_X0Y1_DSP_bot.C5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q
+ _1717_ sg13g2_a21oi_2
X_5430_ Tile_X0Y1_UserCLK net568 _0044_ _0012_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[6\]
+ VPWR VGND sg13g2_dfrbp_1
X_2642_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q net1521 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2
+ _0699_ _0721_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q _0723_
+ VPWR VGND sg13g2_mux4_1
Xoutput315 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 Tile_X0Y0_NN4BEG[15]
+ VPWR VGND sg13g2_buf_1
Xoutput304 net304 Tile_X0Y0_N4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput326 net326 Tile_X0Y0_W1BEG[0] VPWR VGND sg13g2_buf_1
X_5361_ net1939 net1841 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_2573_ _0658_ VPWR _0659_ VGND _0059_ net1682 sg13g2_o21ai_1
X_4312_ _2249_ VPWR _2250_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q
+ net1564 sg13g2_o21ai_1
Xoutput337 net337 Tile_X0Y0_W2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput359 net359 Tile_X0Y0_WW4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput348 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 Tile_X0Y0_W6BEG[11]
+ VPWR VGND sg13g2_buf_1
X_5292_ net1992 net1731 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_99_323 VPWR VGND sg13g2_decap_4
X_4243_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q _0896_
+ _2204_ _2203_ sg13g2_a21oi_1
X_4174_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q net1527 net27
+ net2004 net1593 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q _2144_
+ VPWR VGND sg13g2_mux4_1
X_5460__592 VPWR VGND net592 sg13g2_tiehi
X_3125_ VPWR _1182_ _1181_ VGND sg13g2_inv_1
X_3056_ net1562 net1571 net1668 _1116_ VPWR VGND sg13g2_mux2_1
X_3958_ _1967_ net1700 net1930 VPWR VGND sg13g2_nand2b_1
X_2909_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q net1591 net1585
+ net1522 net1520 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q _0976_
+ VPWR VGND sg13g2_mux4_1
X_3889_ _1902_ _1876_ _1874_ _1903_ VPWR VGND sg13g2_nor3_2
X_5628_ net1915 net1771 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_5559_ net1904 net1794 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_104_144 VPWR VGND sg13g2_fill_1
Xfanout1529 net1529 net1530 VPWR VGND sg13g2_buf_16
Xfanout1518 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 net1518 VPWR VGND
+ sg13g2_buf_8
XFILLER_104_166 VPWR VGND sg13g2_decap_4
XFILLER_18_139 VPWR VGND sg13g2_fill_2
XFILLER_18_117 VPWR VGND sg13g2_fill_1
Xrebuffer80 _0348_ net689 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer91 _1931_ net700 VPWR VGND sg13g2_buf_8
X_5437__561 VPWR VGND net561 sg13g2_tiehi
X_5444__576 VPWR VGND net576 sg13g2_tiehi
XFILLER_66_80 VPWR VGND sg13g2_decap_4
X_4930_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q net116 net132
+ net1925 net92 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q _0474_
+ VPWR VGND sg13g2_mux4_1
X_4861_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q _0408_ _0409_
+ VPWR VGND sg13g2_nor2_1
X_3812_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q net1706 net37
+ net11 net83 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q _1841_
+ VPWR VGND sg13g2_mux4_1
X_4792_ net1607 net1622 net1692 _0343_ VPWR VGND sg13g2_mux2_1
X_3743_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q net125 net101
+ net715 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q
+ _1774_ VPWR VGND sg13g2_mux4_1
X_3674_ _1709_ _1707_ _1708_ _0012_ net1648 VPWR VGND sg13g2_a22oi_1
XFILLER_63_0 VPWR VGND sg13g2_fill_2
X_2625_ _0707_ net1675 net1520 VPWR VGND sg13g2_nand2b_1
X_5413_ net1975 net1817 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_5344_ net1966 net1839 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_2556_ _0641_ VPWR _0642_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q
+ _0639_ sg13g2_o21ai_1
X_2487_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q VPWR _0577_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q _0576_ sg13g2_o21ai_1
XFILLER_99_164 VPWR VGND sg13g2_fill_2
XFILLER_99_186 VPWR VGND sg13g2_fill_1
Xoutput189 net189 Tile_X0Y0_E2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput178 net178 Tile_X0Y0_E2BEG[1] VPWR VGND sg13g2_buf_1
X_5275_ net1953 net1733 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_4226_ _2188_ _2187_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 VPWR VGND sg13g2_mux2_1
X_4157_ _2129_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q _1512_
+ VPWR VGND sg13g2_nand2_1
X_3108_ _0703_ _0848_ _1165_ VPWR VGND sg13g2_nor2_1
X_4088_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q net1622 _0614_
+ _2084_ _0611_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1
+ VPWR VGND sg13g2_mux4_1
X_3039_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q _1091_
+ _1100_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q sg13g2_a21oi_1
XFILLER_70_204 VPWR VGND sg13g2_decap_8
XFILLER_23_175 VPWR VGND sg13g2_fill_2
XFILLER_11_326 VPWR VGND sg13g2_fill_1
Xfanout2005 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q net2005 VPWR
+ VGND sg13g2_buf_1
XFILLER_87_13 VPWR VGND sg13g2_fill_1
XFILLER_87_35 VPWR VGND sg13g2_fill_2
XFILLER_61_204 VPWR VGND sg13g2_fill_1
XFILLER_61_215 VPWR VGND sg13g2_fill_1
XFILLER_61_237 VPWR VGND sg13g2_fill_2
Xinput36 Tile_X0Y0_S2END[6] net36 VPWR VGND sg13g2_buf_1
Xinput25 Tile_X0Y0_EE4END[3] net25 VPWR VGND sg13g2_buf_1
Xinput14 Tile_X0Y0_E2MID[2] net14 VPWR VGND sg13g2_buf_1
Xinput58 Tile_X0Y0_SS4END[4] net58 VPWR VGND sg13g2_buf_1
Xinput47 Tile_X0Y0_S4END[1] net47 VPWR VGND sg13g2_buf_1
Xinput69 Tile_X0Y0_W2END[4] net69 VPWR VGND sg13g2_buf_1
X_3390_ _1424_ _1423_ _1442_ VPWR VGND sg13g2_nor2b_1
XFILLER_123_283 VPWR VGND sg13g2_fill_1
X_5060_ net1973 net1808 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_4011_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q net1598 net1610
+ net649 net1623 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q _2016_
+ VPWR VGND sg13g2_mux4_1
Xfanout1860 Tile_X0Y1_FrameData[7] net1860 VPWR VGND sg13g2_buf_1
Xfanout1882 Tile_X0Y1_FrameData[26] net1882 VPWR VGND sg13g2_buf_1
Xfanout1871 Tile_X0Y1_FrameData[31] net1871 VPWR VGND sg13g2_buf_1
Xfanout1893 Tile_X0Y1_FrameData[21] net1893 VPWR VGND sg13g2_buf_1
X_5962_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 net183 VPWR VGND sg13g2_buf_1
XFILLER_52_259 VPWR VGND sg13g2_fill_1
X_4913_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q _0457_ _0458_
+ VPWR VGND sg13g2_nor2_1
X_5893_ net1875 net1814 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_4844_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q VPWR _0392_ VGND
+ net1685 _0177_ sg13g2_o21ai_1
XFILLER_32_19 VPWR VGND sg13g2_fill_2
XFILLER_60_270 VPWR VGND sg13g2_fill_2
X_4775_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q _0308_ _0325_
+ _0326_ VPWR VGND sg13g2_a21o_1
X_3726_ _1758_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q _1757_
+ _1756_ _1754_ VPWR VGND sg13g2_a22oi_1
X_3657_ _1693_ _1446_ _1448_ VPWR VGND sg13g2_xnor2_1
X_3588_ _1628_ VPWR _1629_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q
+ net1581 sg13g2_o21ai_1
X_2608_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q VPWR _0692_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q _0690_ sg13g2_o21ai_1
X_5427__571 VPWR VGND net571 sg13g2_tiehi
X_2539_ _0625_ VPWR _0626_ VGND _0618_ _0622_ sg13g2_o21ai_1
X_5327_ net1998 net1719 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_5258_ net1987 net1745 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_5189_ net1976 net1763 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_4209_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q _2174_ _2175_
+ VPWR VGND sg13g2_nor2_1
XFILLER_113_99 VPWR VGND sg13g2_decap_4
XFILLER_73_59 VPWR VGND sg13g2_fill_1
X_5434__564 VPWR VGND net564 sg13g2_tiehi
XFILLER_11_145 VPWR VGND sg13g2_fill_2
XFILLER_98_23 VPWR VGND sg13g2_fill_1
XFILLER_98_45 VPWR VGND sg13g2_fill_2
X_5441__557 VPWR VGND net557 sg13g2_tiehi
XFILLER_66_329 VPWR VGND sg13g2_fill_2
XFILLER_74_340 VPWR VGND sg13g2_fill_2
X_2890_ net1922 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q _0959_
+ VPWR VGND sg13g2_nor2_1
X_4560_ VPWR _0117_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q VGND
+ sg13g2_inv_1
X_3511_ VGND VPWR _0142_ _1557_ _1558_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q
+ sg13g2_a21oi_1
X_4491_ net1513 _1895_ _0048_ VPWR VGND sg13g2_nor2_1
X_3442_ VGND VPWR net64 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q
+ _1493_ _1492_ sg13g2_a21oi_1
X_6230_ net1877 net443 VPWR VGND sg13g2_buf_1
X_6161_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 net382 VPWR VGND sg13g2_buf_1
X_3373_ _1425_ _1424_ _1423_ VPWR VGND sg13g2_nand2b_1
X_5112_ net1977 net1796 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_6092_ Tile_X0Y1_NN4END[12] net319 VPWR VGND sg13g2_buf_1
X_5043_ net1943 net1851 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
Xfanout1690 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q net1690 VPWR
+ VGND sg13g2_buf_1
XFILLER_25_215 VPWR VGND sg13g2_fill_2
X_5876_ net1898 net1812 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_4827_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q net1549 net689
+ _0375_ _0362_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q _0376_
+ VPWR VGND sg13g2_mux4_1
X_4758_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q net1528 net1534
+ net1543 net1556 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q _0309_
+ VPWR VGND sg13g2_mux4_1
X_3709_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q net124 net100
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 net160 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q
+ _1742_ VPWR VGND sg13g2_mux4_1
X_4689_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q VPWR _0243_ VGND
+ _0241_ _0242_ sg13g2_o21ai_1
XFILLER_75_104 VPWR VGND sg13g2_fill_2
XFILLER_84_36 VPWR VGND sg13g2_fill_2
XFILLER_56_384 VPWR VGND sg13g2_fill_1
XFILLER_58_70 VPWR VGND sg13g2_fill_2
XFILLER_66_159 VPWR VGND sg13g2_fill_2
XFILLER_81_118 VPWR VGND sg13g2_fill_2
X_3991_ net1701 net30 _1996_ VPWR VGND sg13g2_nor2b_1
X_5730_ net1864 net1735 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_2942_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[4\] net1642 _1006_ VPWR VGND sg13g2_mux2_2
X_5661_ net1917 net1760 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_2873_ _0942_ VPWR _0943_ VGND _0376_ net1686 sg13g2_o21ai_1
X_4612_ VPWR _0169_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q VGND
+ sg13g2_inv_1
X_5592_ net1906 net1781 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_4543_ VPWR _0100_ net78 VGND sg13g2_inv_1
X_4474_ VGND VPWR _1559_ _2383_ _2388_ _2387_ sg13g2_a21oi_1
X_6213_ net1914 net425 VPWR VGND sg13g2_buf_1
X_3425_ _1476_ _1475_ _1456_ VPWR VGND sg13g2_nand2b_1
X_6144_ Tile_X0Y0_WW4END[11] net371 VPWR VGND sg13g2_buf_1
X_3356_ _1404_ _1405_ _1408_ VPWR VGND sg13g2_xor2_1
X_6075_ Tile_X0Y1_N4END[11] net302 VPWR VGND sg13g2_buf_1
X_5424__574 VPWR VGND net574 sg13g2_tiehi
X_3287_ _1337_ _1338_ _1339_ VPWR VGND sg13g2_nor2b_1
X_5026_ net1969 net1852 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_5859_ net1867 net1821 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_5431__567 VPWR VGND net567 sg13g2_tiehi
XFILLER_119_194 VPWR VGND sg13g2_fill_2
XFILLER_79_25 VPWR VGND sg13g2_fill_2
XFILLER_122_359 VPWR VGND sg13g2_fill_2
XFILLER_29_340 VPWR VGND sg13g2_fill_2
XFILLER_8_255 VPWR VGND sg13g2_fill_1
Xoutput508 net508 Tile_X0Y1_W1BEG[2] VPWR VGND sg13g2_buf_1
Xoutput519 net519 Tile_X0Y1_W2BEGb[1] VPWR VGND sg13g2_buf_1
X_3210_ net1562 net1571 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q
+ _1265_ VPWR VGND sg13g2_mux2_1
XFILLER_69_80 VPWR VGND sg13g2_decap_8
XFILLER_69_91 VPWR VGND sg13g2_fill_1
X_4190_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q _2157_
+ _2158_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q sg13g2_a21oi_1
X_3141_ net624 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q _1197_
+ VPWR VGND sg13g2_nor2b_1
X_3072_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q net128 net104
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 net164 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q
+ _1131_ VPWR VGND sg13g2_mux4_1
XFILLER_62_151 VPWR VGND sg13g2_fill_1
XFILLER_62_195 VPWR VGND sg13g2_decap_4
X_3974_ _1980_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[17\] net1655 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ VPWR VGND sg13g2_mux2_1
XFILLER_93_0 VPWR VGND sg13g2_fill_2
X_5713_ net1890 net1736 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_2925_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q VPWR _0991_ VGND
+ net1661 net1581 sg13g2_o21ai_1
X_2856_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q _0905_ _0926_
+ _0596_ _0925_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q Tile_X0Y1_DSP_bot.A2
+ VPWR VGND sg13g2_mux4_1
X_5644_ net1881 net1760 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_40_19 VPWR VGND sg13g2_fill_1
X_2787_ VGND VPWR net35 net1690 _0862_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q
+ sg13g2_a21oi_1
X_5575_ net1919 net1790 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_4526_ VPWR _0083_ net128 VGND sg13g2_inv_1
X_4457_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q net1573 net1577
+ net1615 net1617 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q _2373_
+ VPWR VGND sg13g2_mux4_1
X_3408_ _1460_ _1165_ _1459_ VPWR VGND sg13g2_xnor2_1
XFILLER_104_348 VPWR VGND sg13g2_fill_1
X_6127_ Tile_X0Y0_W6END[4] net350 VPWR VGND sg13g2_buf_1
X_4388_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q _2306_ _2307_
+ _2313_ _2312_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0
+ VPWR VGND sg13g2_mux4_1
X_3339_ _1391_ _1390_ _1389_ VPWR VGND sg13g2_nand2b_1
XFILLER_45_107 VPWR VGND sg13g2_fill_1
X_6058_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 net279 VPWR VGND sg13g2_buf_1
XFILLER_45_129 VPWR VGND sg13g2_decap_8
X_5009_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q VPWR _0549_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q _0546_ sg13g2_o21ai_1
XFILLER_41_357 VPWR VGND sg13g2_fill_2
XFILLER_5_269 VPWR VGND sg13g2_fill_1
XFILLER_122_189 VPWR VGND sg13g2_fill_2
XFILLER_39_61 VPWR VGND sg13g2_fill_2
XFILLER_29_181 VPWR VGND sg13g2_decap_8
XFILLER_44_151 VPWR VGND sg13g2_decap_4
X_2710_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q VPWR _0789_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q _0787_ sg13g2_o21ai_1
X_3690_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q
+ _1724_ _1720_ _1725_ _1723_ sg13g2_a221oi_1
X_2641_ _0722_ _0721_ VPWR VGND sg13g2_inv_2
Xoutput316 net316 Tile_X0Y0_NN4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput305 net305 Tile_X0Y0_N4BEG[6] VPWR VGND sg13g2_buf_1
X_5360_ net1937 net1841 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_2572_ VGND VPWR net32 net1682 _0658_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q
+ sg13g2_a21oi_1
X_4311_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q net1569
+ _2249_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q sg13g2_a21oi_1
Xoutput327 net327 Tile_X0Y0_W1BEG[1] VPWR VGND sg13g2_buf_1
Xoutput338 net338 Tile_X0Y0_W2BEGb[0] VPWR VGND sg13g2_buf_1
X_5291_ net1990 net1730 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput349 net349 Tile_X0Y0_W6BEG[1] VPWR VGND sg13g2_buf_1
X_4242_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q VPWR _2203_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q net694 sg13g2_o21ai_1
X_4173_ VGND VPWR _2143_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 _2137_
+ _2135_ sg13g2_a21oi_2
X_3124_ net1691 net1599 net1612 net1605 net1625 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q
+ _1181_ VPWR VGND sg13g2_mux4_1
X_3055_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q _1114_ _1115_
+ VPWR VGND sg13g2_nor2_2
X_3957_ _1965_ VPWR _1966_ VGND _0091_ net1700 sg13g2_o21ai_1
X_2908_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q net1597 net1610
+ net649 net1632 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q _0975_
+ VPWR VGND sg13g2_mux4_1
X_3888_ _1870_ _1901_ _1902_ VPWR VGND sg13g2_and2_1
X_5627_ net1912 net1770 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_2839_ _0911_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q _0910_
+ VPWR VGND sg13g2_nand2_1
X_5558_ net1902 net1794 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_4509_ VPWR _0066_ net42 VGND sg13g2_inv_1
XFILLER_104_112 VPWR VGND sg13g2_fill_1
X_5489_ net1890 net1848 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
Xfanout1519 net1520 net1519 VPWR VGND sg13g2_buf_2
XFILLER_58_276 VPWR VGND sg13g2_decap_8
Xrebuffer81 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 net690 VPWR VGND
+ sg13g2_dlygate4sd1_1
XFILLER_25_52 VPWR VGND sg13g2_fill_1
XFILLER_14_335 VPWR VGND sg13g2_fill_1
Xrebuffer92 _0411_ net701 VPWR VGND sg13g2_buf_8
XFILLER_110_104 VPWR VGND sg13g2_fill_1
XFILLER_2_12 VPWR VGND sg13g2_fill_2
XFILLER_110_159 VPWR VGND sg13g2_fill_1
XFILLER_49_287 VPWR VGND sg13g2_decap_8
X_4860_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q _0404_
+ _0408_ _0407_ sg13g2_a21oi_1
X_3811_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q _1837_
+ _1840_ _1839_ sg13g2_a21oi_1
X_4791_ _0341_ VPWR _0342_ VGND net1692 net1601 sg13g2_o21ai_1
X_3742_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q VPWR _1773_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q _1772_ sg13g2_o21ai_1
X_3673_ VGND VPWR net1643 _0152_ _1708_ net1648 sg13g2_a21oi_1
X_2624_ net690 net1587 net1674 _0706_ VPWR VGND sg13g2_mux2_1
X_5412_ net1973 net1817 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_0 VPWR VGND sg13g2_decap_8
X_5343_ net1963 net1839 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_2555_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q _0640_
+ _0641_ _0092_ sg13g2_a21oi_1
XFILLER_99_154 VPWR VGND sg13g2_decap_4
X_2486_ _0575_ VPWR _0576_ VGND _0068_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q
+ sg13g2_o21ai_1
XFILLER_87_327 VPWR VGND sg13g2_fill_1
Xoutput179 net179 Tile_X0Y0_E2BEG[2] VPWR VGND sg13g2_buf_1
X_5274_ net1951 net1733 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_4225_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2
+ net28 net1932 net1607 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q
+ _2188_ VPWR VGND sg13g2_mux4_1
X_4156_ _2127_ VPWR _2128_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q
+ net1524 sg13g2_o21ai_1
X_3107_ _1164_ net1575 net1515 VPWR VGND sg13g2_nand2b_1
X_4087_ _2083_ VPWR _2084_ VGND _2065_ _2071_ sg13g2_o21ai_1
X_3038_ _1097_ VPWR _1099_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q
+ _1098_ sg13g2_o21ai_1
XFILLER_70_227 VPWR VGND sg13g2_fill_1
XFILLER_102_46 VPWR VGND sg13g2_fill_2
X_4989_ net1592 net1584 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q
+ _0530_ VPWR VGND sg13g2_mux2_1
XFILLER_11_21 VPWR VGND sg13g2_fill_1
XFILLER_11_43 VPWR VGND sg13g2_fill_2
X_5467__599 VPWR VGND net599 sg13g2_tiehi
XFILLER_93_319 VPWR VGND sg13g2_fill_2
XFILLER_100_192 VPWR VGND sg13g2_decap_4
Xinput37 Tile_X0Y0_S2END[7] net37 VPWR VGND sg13g2_buf_1
Xinput26 Tile_X0Y0_S1END[0] net26 VPWR VGND sg13g2_buf_1
Xinput15 Tile_X0Y0_E2MID[3] net15 VPWR VGND sg13g2_buf_1
Xinput59 Tile_X0Y0_SS4END[5] net59 VPWR VGND sg13g2_buf_1
Xinput48 Tile_X0Y0_S4END[2] net48 VPWR VGND sg13g2_buf_1
X_4010_ _1992_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q _2014_
+ _2015_ VPWR VGND sg13g2_nand3_1
Xfanout1861 Tile_X0Y1_FrameData[7] net1861 VPWR VGND sg13g2_buf_1
Xfanout1850 Tile_X0Y1_FrameStrobe[0] net1850 VPWR VGND sg13g2_buf_1
Xfanout1883 Tile_X0Y1_FrameData[26] net1883 VPWR VGND sg13g2_buf_1
Xfanout1894 net1895 net1894 VPWR VGND sg13g2_buf_1
XFILLER_37_224 VPWR VGND sg13g2_decap_4
Xfanout1872 Tile_X0Y1_FrameData[30] net1872 VPWR VGND sg13g2_buf_1
X_5961_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 net182 VPWR VGND sg13g2_buf_1
X_4912_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q net18 net79 net44
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q
+ _0457_ VPWR VGND sg13g2_mux4_1
X_5892_ net1869 net1814 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_4843_ VGND VPWR _0391_ _0387_ _0390_ sg13g2_or2_1
XFILLER_20_135 VPWR VGND sg13g2_fill_2
X_4774_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q VPWR _0325_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q _0324_ sg13g2_o21ai_1
X_3725_ net163 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q
+ _1757_ VPWR VGND sg13g2_mux2_1
X_3656_ _1672_ VPWR _1692_ VGND _1691_ _1690_ sg13g2_o21ai_1
X_3587_ _1628_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q net1619
+ VPWR VGND sg13g2_nand2b_1
X_2607_ net1581 net1619 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ _0691_ VPWR VGND sg13g2_mux2_1
X_2538_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q _0624_ _0625_
+ VPWR VGND sg13g2_nor2_1
X_5326_ net1996 net1719 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_114_273 VPWR VGND sg13g2_fill_1
X_5257_ net1985 net1744 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_2469_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q _0558_
+ _0559_ _0108_ sg13g2_a21oi_1
X_4208_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q _0598_ net1931
+ net2001 net1622 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q _2174_
+ VPWR VGND sg13g2_mux4_1
XFILLER_68_382 VPWR VGND sg13g2_fill_2
X_5188_ net1974 net1763 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_4139_ _2113_ VPWR _2114_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q
+ net681 sg13g2_o21ai_1
XFILLER_43_216 VPWR VGND sg13g2_fill_2
XFILLER_118_2 VPWR VGND sg13g2_fill_1
XFILLER_22_97 VPWR VGND sg13g2_fill_1
XFILLER_3_345 VPWR VGND sg13g2_fill_2
XFILLER_93_105 VPWR VGND sg13g2_fill_1
X_3510_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q net1711 net1926
+ net121 net97 net1669 _1557_ VPWR VGND sg13g2_mux4_1
X_4490_ net1514 _1893_ _0047_ VPWR VGND sg13g2_nor2_1
X_3441_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q VPWR _1492_ VGND
+ _0086_ net1687 sg13g2_o21ai_1
XFILLER_6_194 VPWR VGND sg13g2_fill_1
X_6160_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 net381 VPWR VGND sg13g2_buf_1
X_3372_ _1424_ _1407_ _1408_ VPWR VGND sg13g2_xnor2_1
X_5111_ net1955 net1796 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_6091_ Tile_X0Y1_NN4END[11] net318 VPWR VGND sg13g2_buf_1
X_5042_ net1941 net1851 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
Xfanout1691 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q net1691 VPWR
+ VGND sg13g2_buf_1
Xfanout1680 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q net1680 VPWR
+ VGND sg13g2_buf_1
XFILLER_84_149 VPWR VGND sg13g2_fill_2
X_5875_ net1894 net1812 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_4826_ _0375_ _0372_ _0374_ _0370_ _0368_ VPWR VGND sg13g2_a22oi_1
X_4757_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q net133 net93
+ net158 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q
+ _0308_ VPWR VGND sg13g2_mux4_1
X_3708_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q net99 net159
+ net642 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q
+ _1741_ VPWR VGND sg13g2_mux4_1
X_4688_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q VPWR _0242_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q _0239_ sg13g2_o21ai_1
X_3639_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q _1673_
+ _1676_ _1675_ sg13g2_a21oi_1
X_5309_ net1959 net1719 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_6289_ net151 net510 VPWR VGND sg13g2_buf_1
XFILLER_102_265 VPWR VGND sg13g2_fill_2
XFILLER_33_30 VPWR VGND sg13g2_fill_1
XFILLER_33_63 VPWR VGND sg13g2_fill_1
XFILLER_33_74 VPWR VGND sg13g2_fill_2
XFILLER_123_0 VPWR VGND sg13g2_fill_2
XFILLER_74_171 VPWR VGND sg13g2_fill_2
X_3990_ _1994_ VPWR _1995_ VGND _0070_ net1701 sg13g2_o21ai_1
X_2941_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q _1004_ _1005_
+ _0974_ _0721_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X
+ VPWR VGND sg13g2_mux4_1
X_5660_ net1915 net1761 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_30_230 VPWR VGND sg13g2_decap_8
X_4611_ VPWR _0168_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q
+ VGND sg13g2_inv_1
X_2872_ _0942_ _0083_ net1686 VPWR VGND sg13g2_nand2_1
X_5591_ net1904 net1783 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_4542_ VPWR _0099_ net43 VGND sg13g2_inv_1
XFILLER_116_324 VPWR VGND sg13g2_fill_2
X_4473_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q VPWR _2387_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q _2386_ sg13g2_o21ai_1
X_6212_ net1916 net424 VPWR VGND sg13g2_buf_1
X_3424_ _1238_ _1455_ _1180_ _1475_ VPWR VGND sg13g2_a21o_1
X_6143_ Tile_X0Y0_WW4END[10] net370 VPWR VGND sg13g2_buf_1
X_3355_ VGND VPWR _1401_ _1407_ _1402_ _1396_ sg13g2_a21oi_2
X_6074_ Tile_X0Y1_N4END[10] net301 VPWR VGND sg13g2_buf_1
X_3286_ _1338_ _1285_ _1286_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_330 VPWR VGND sg13g2_fill_1
X_5025_ net1968 net1854 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_54_29 VPWR VGND sg13g2_decap_8
XFILLER_53_366 VPWR VGND sg13g2_fill_1
XFILLER_110_24 VPWR VGND sg13g2_fill_2
XFILLER_110_68 VPWR VGND sg13g2_fill_2
X_5858_ net1865 net1821 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_4809_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q net119 net95
+ net1926 net1923 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q _0359_
+ VPWR VGND sg13g2_mux4_1
X_5789_ net1918 net1717 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_48_105 VPWR VGND sg13g2_fill_2
XFILLER_28_41 VPWR VGND sg13g2_fill_1
XFILLER_48_127 VPWR VGND sg13g2_fill_2
XFILLER_71_174 VPWR VGND sg13g2_fill_1
XFILLER_44_73 VPWR VGND sg13g2_fill_1
Xoutput509 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 Tile_X0Y1_W1BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_60_94 VPWR VGND sg13g2_decap_8
X_3140_ _1196_ _1185_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 VPWR VGND
+ sg13g2_nor2_2
XFILLER_10_4 VPWR VGND sg13g2_fill_2
X_3071_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q net1708 net103
+ net615 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q
+ _1130_ VPWR VGND sg13g2_mux4_1
XFILLER_94_255 VPWR VGND sg13g2_fill_2
XFILLER_35_333 VPWR VGND sg13g2_fill_2
X_5712_ net1888 net1736 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_3973_ _1980_ _1953_ _1979_ VPWR VGND sg13g2_xnor2_1
X_2924_ net1555 net1562 net1661 _0990_ VPWR VGND sg13g2_mux2_1
X_5643_ net1878 net1759 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_2855_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q net119 net42 net107
+ net155 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q _0926_ VPWR VGND
+ sg13g2_mux4_1
X_5574_ net1896 net1790 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_2786_ _0861_ net27 net1690 VPWR VGND sg13g2_nand2b_1
X_4525_ VPWR _0082_ net80 VGND sg13g2_inv_1
X_4456_ _2372_ _2371_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q
+ _2369_ _2368_ VPWR VGND sg13g2_a22oi_1
X_4387_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q net1572 net1579
+ net1615 net1618 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q _2313_
+ VPWR VGND sg13g2_mux4_1
X_3407_ net1515 _0899_ _1459_ VPWR VGND sg13g2_nor2b_1
X_6126_ Tile_X0Y0_W6END[3] net349 VPWR VGND sg13g2_buf_1
X_3338_ _1390_ _1386_ _1387_ VPWR VGND sg13g2_xnor2_1
XFILLER_112_382 VPWR VGND sg13g2_fill_2
XFILLER_85_222 VPWR VGND sg13g2_decap_8
X_3269_ VPWR _1322_ _1321_ VGND sg13g2_inv_1
X_6057_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 net278 VPWR VGND sg13g2_buf_1
XFILLER_26_322 VPWR VGND sg13g2_fill_2
X_5008_ VGND VPWR net1660 _0178_ _0548_ _0547_ sg13g2_a21oi_1
XFILLER_30_53 VPWR VGND sg13g2_decap_8
XFILLER_100_2 VPWR VGND sg13g2_fill_1
XFILLER_44_141 VPWR VGND sg13g2_fill_1
XFILLER_32_358 VPWR VGND sg13g2_fill_1
X_2640_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q net146 net83 net49
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q
+ _0721_ VPWR VGND sg13g2_mux4_1
Xoutput306 net306 Tile_X0Y0_N4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput317 net317 Tile_X0Y0_NN4BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_58_4 VPWR VGND sg13g2_fill_1
X_2571_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q _0656_
+ _0657_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q sg13g2_a21oi_1
X_4310_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q _0178_
+ _2248_ _2247_ sg13g2_a21oi_1
Xoutput328 net328 Tile_X0Y0_W1BEG[2] VPWR VGND sg13g2_buf_1
Xoutput339 net339 Tile_X0Y0_W2BEGb[1] VPWR VGND sg13g2_buf_1
X_5290_ net1988 net1730 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_4241_ _1482_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q _2201_
+ _2202_ VPWR VGND sg13g2_a21o_1
X_4172_ _2139_ _2142_ _2143_ VPWR VGND sg13g2_nor2_1
X_3123_ _1180_ _1178_ _1163_ VPWR VGND sg13g2_xnor2_1
X_3054_ net1668 net1531 net1536 net1545 net1552 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q
+ _1114_ VPWR VGND sg13g2_mux4_1
X_3956_ VGND VPWR net29 net1700 _1965_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q
+ sg13g2_a21oi_1
X_2907_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q net1707 net10
+ net57 net71 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q _0974_ VPWR
+ VGND sg13g2_mux4_1
X_5626_ net1910 net1770 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_3887_ _1901_ _1166_ _1872_ VPWR VGND sg13g2_nand2b_1
X_2838_ net1577 net1617 net1667 _0910_ VPWR VGND sg13g2_mux2_1
X_5557_ net1900 net1794 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_2769_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q _0412_
+ _0845_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q sg13g2_a21oi_1
X_4508_ VPWR _0065_ net113 VGND sg13g2_inv_1
X_5488_ net1888 net1848 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_218 VPWR VGND sg13g2_fill_1
X_4439_ _2356_ VPWR _2357_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q
+ _2353_ sg13g2_o21ai_1
X_6109_ net65 net330 VPWR VGND sg13g2_buf_1
XFILLER_100_352 VPWR VGND sg13g2_fill_1
Xrebuffer60 _0565_ net669 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer82 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 net691 VPWR VGND
+ sg13g2_dlygate4sd1_1
XFILLER_41_155 VPWR VGND sg13g2_fill_1
XFILLER_41_177 VPWR VGND sg13g2_fill_2
XFILLER_41_52 VPWR VGND sg13g2_fill_1
XFILLER_41_74 VPWR VGND sg13g2_decap_8
XFILLER_96_306 VPWR VGND sg13g2_decap_8
XFILLER_49_200 VPWR VGND sg13g2_fill_1
XFILLER_66_60 VPWR VGND sg13g2_fill_2
XFILLER_17_196 VPWR VGND sg13g2_fill_2
X_4790_ _0341_ net1692 net1614 VPWR VGND sg13g2_nand2b_1
X_3810_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q VPWR _1839_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q _1838_ sg13g2_o21ai_1
X_3741_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q net118 net94
+ net41 net170 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q _1772_
+ VPWR VGND sg13g2_mux4_1
XFILLER_32_188 VPWR VGND sg13g2_fill_1
XFILLER_13_380 VPWR VGND sg13g2_fill_1
X_3672_ _1707_ net1637 Tile_X0Y1_DSP_bot.C6 VPWR VGND sg13g2_nand2_1
X_5411_ net1972 net1818 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_63_2 VPWR VGND sg13g2_fill_1
X_2623_ _0705_ _0704_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q
+ VPWR VGND sg13g2_nand2b_1
X_2554_ net1524 net1520 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ _0640_ VPWR VGND sg13g2_mux2_1
X_5342_ net1962 net1842 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_99_133 VPWR VGND sg13g2_decap_8
X_2485_ _0575_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q net53 VPWR
+ VGND sg13g2_nand2_1
X_5273_ net2000 net1742 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_99_166 VPWR VGND sg13g2_fill_1
X_4224_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q net1584 _0969_
+ _1011_ _1935_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q _2187_
+ VPWR VGND sg13g2_mux4_1
X_4155_ _2127_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q _0630_
+ VPWR VGND sg13g2_nand2_1
X_3106_ _1162_ _1159_ _1052_ _1163_ VPWR VGND sg13g2_a21o_1
X_4086_ _2076_ _2082_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q
+ _2083_ VPWR VGND sg13g2_nand3_1
X_3037_ net101 net715 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q
+ _1098_ VPWR VGND sg13g2_mux2_1
XFILLER_23_177 VPWR VGND sg13g2_fill_1
X_4988_ _0529_ _0528_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q
+ VPWR VGND sg13g2_nand2b_1
X_3939_ _1949_ _1931_ _1947_ VPWR VGND sg13g2_nand2_2
X_5609_ net1873 net1774 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_46_269 VPWR VGND sg13g2_fill_1
XFILLER_54_280 VPWR VGND sg13g2_decap_8
XFILLER_52_40 VPWR VGND sg13g2_fill_1
Xinput27 Tile_X0Y0_S1END[1] net27 VPWR VGND sg13g2_buf_1
X_5450__582 VPWR VGND net582 sg13g2_tiehi
Xinput16 Tile_X0Y0_E2MID[4] net16 VPWR VGND sg13g2_buf_1
Xinput49 Tile_X0Y0_S4END[3] net49 VPWR VGND sg13g2_buf_1
Xinput38 Tile_X0Y0_S2MID[0] net38 VPWR VGND sg13g2_buf_1
XFILLER_6_365 VPWR VGND sg13g2_fill_1
Xfanout1840 net1841 net1840 VPWR VGND sg13g2_buf_1
Xfanout1851 net1853 net1851 VPWR VGND sg13g2_buf_1
Xfanout1862 Tile_X0Y1_FrameData[6] net1862 VPWR VGND sg13g2_buf_1
Xfanout1884 Tile_X0Y1_FrameData[25] net1884 VPWR VGND sg13g2_buf_1
Xfanout1873 Tile_X0Y1_FrameData[30] net1873 VPWR VGND sg13g2_buf_1
XFILLER_77_361 VPWR VGND sg13g2_fill_2
Xfanout1895 Tile_X0Y1_FrameData[20] net1895 VPWR VGND sg13g2_buf_1
XFILLER_52_206 VPWR VGND sg13g2_fill_1
X_5960_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 net181 VPWR VGND sg13g2_buf_1
X_5891_ net1867 net1819 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_4911_ _0445_ _0456_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 VPWR VGND
+ sg13g2_nor2_1
X_4842_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q VPWR _0390_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q _0389_ sg13g2_o21ai_1
X_4773_ net713 _0324_ VPWR VGND sg13g2_inv_4
X_3724_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q _1755_ _1756_
+ VPWR VGND sg13g2_nor2_1
X_3655_ net1636 VPWR _1691_ VGND net1639 _0011_ sg13g2_o21ai_1
X_2606_ net1555 net1571 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ _0690_ VPWR VGND sg13g2_mux2_1
XFILLER_106_219 VPWR VGND sg13g2_decap_8
X_3586_ _1626_ VPWR _1627_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q
+ net1555 sg13g2_o21ai_1
X_2537_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q _0623_ _0624_
+ VPWR VGND sg13g2_nor2_1
X_5325_ net1993 net1722 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_2468_ _0557_ VPWR _0558_ VGND net1680 net1521 sg13g2_o21ai_1
X_5256_ net1983 net1744 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_4207_ VGND VPWR _2172_ _2173_ _2169_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q
+ sg13g2_a21oi_2
XFILLER_68_372 VPWR VGND sg13g2_fill_2
X_5187_ net1971 net1763 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_4138_ VGND VPWR _0061_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q
+ _2113_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q sg13g2_a21oi_1
X_4069_ _2066_ net1694 _0087_ VPWR VGND sg13g2_nand2_1
XFILLER_11_147 VPWR VGND sg13g2_fill_1
XFILLER_11_169 VPWR VGND sg13g2_fill_2
XFILLER_22_54 VPWR VGND sg13g2_fill_2
XFILLER_98_47 VPWR VGND sg13g2_fill_1
XFILLER_86_180 VPWR VGND sg13g2_fill_2
XFILLER_6_140 VPWR VGND sg13g2_fill_1
XFILLER_6_151 VPWR VGND sg13g2_fill_1
X_3440_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q net1516 net2003
+ net1707 net10 net1687 _1491_ VPWR VGND sg13g2_mux4_1
X_3371_ VGND VPWR _1419_ _1420_ _1423_ _1422_ sg13g2_a21oi_1
X_6090_ Tile_X0Y1_NN4END[10] net317 VPWR VGND sg13g2_buf_1
X_5110_ net1949 net1796 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_69_147 VPWR VGND sg13g2_fill_1
X_5041_ net1939 net1854 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
Xfanout1670 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q net1670 VPWR
+ VGND sg13g2_buf_1
Xfanout1681 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q net1681 VPWR
+ VGND sg13g2_buf_1
Xfanout1692 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q net1692 VPWR
+ VGND sg13g2_buf_1
XFILLER_25_217 VPWR VGND sg13g2_fill_1
XFILLER_92_161 VPWR VGND sg13g2_fill_2
X_5874_ net1892 net1813 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_4825_ VGND VPWR _0071_ _0373_ _0374_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q
+ sg13g2_a21oi_1
X_4756_ _0307_ VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 VGND _0303_
+ _0296_ sg13g2_o21ai_1
X_3707_ _1732_ _1739_ _1740_ VPWR VGND sg13g2_nor2_1
X_4687_ VGND VPWR net1676 _0179_ _0241_ _0240_ sg13g2_a21oi_1
X_3638_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q _1674_ _1675_
+ VPWR VGND sg13g2_nor2b_1
X_3569_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7
+ _1611_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q sg13g2_a21oi_1
X_5308_ net1957 net1719 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_5239_ net1956 net1754 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_320 VPWR VGND sg13g2_fill_1
XFILLER_56_353 VPWR VGND sg13g2_fill_2
XFILLER_71_378 VPWR VGND sg13g2_fill_1
XFILLER_24_283 VPWR VGND sg13g2_fill_1
XFILLER_116_0 VPWR VGND sg13g2_fill_1
XFILLER_62_356 VPWR VGND sg13g2_fill_2
X_2940_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7
+ net45 net19 net80 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q _1005_
+ VPWR VGND sg13g2_mux4_1
X_2871_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q _0939_
+ _0941_ _0940_ sg13g2_a21oi_1
X_4610_ VPWR _0167_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q
+ VGND sg13g2_inv_1
XFILLER_30_275 VPWR VGND sg13g2_fill_2
X_5590_ net1902 net1783 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_4541_ VPWR _0098_ net17 VGND sg13g2_inv_1
X_4472_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q net712 _2386_
+ VPWR VGND sg13g2_nor2_1
X_6211_ net1918 net423 VPWR VGND sg13g2_buf_1
X_3423_ _1474_ _1472_ _1473_ net1650 _0000_ VPWR VGND sg13g2_a22oi_1
X_6142_ Tile_X0Y0_WW4END[9] net369 VPWR VGND sg13g2_buf_1
XFILLER_31_0 VPWR VGND sg13g2_fill_1
X_3354_ _1404_ _1405_ _1406_ VPWR VGND sg13g2_nor2_1
XFILLER_97_231 VPWR VGND sg13g2_fill_1
X_6073_ Tile_X0Y1_N4END[9] net300 VPWR VGND sg13g2_buf_1
X_3285_ VGND VPWR _1335_ _1336_ _1337_ _1307_ sg13g2_a21oi_1
X_5024_ net1965 net1854 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_65_183 VPWR VGND sg13g2_decap_8
XFILLER_110_36 VPWR VGND sg13g2_fill_2
X_5857_ net1863 net1821 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_70_18 VPWR VGND sg13g2_fill_2
X_4808_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q net42 net50 net155
+ net171 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q _0358_ VPWR
+ VGND sg13g2_mux4_1
X_5788_ net1916 net1715 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_4739_ _0291_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q _0289_
+ VPWR VGND sg13g2_nand2_1
XFILLER_119_196 VPWR VGND sg13g2_fill_1
XFILLER_79_27 VPWR VGND sg13g2_fill_1
XFILLER_29_353 VPWR VGND sg13g2_fill_1
XFILLER_71_131 VPWR VGND sg13g2_fill_1
XFILLER_8_235 VPWR VGND sg13g2_fill_1
X_3070_ _1121_ VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 VGND _1127_
+ _1129_ sg13g2_o21ai_1
X_5711_ net1886 net1739 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_3972_ _1977_ _1978_ _1979_ VPWR VGND sg13g2_nor2b_1
XFILLER_93_2 VPWR VGND sg13g2_fill_1
X_2923_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q _0988_ _0989_
+ VPWR VGND sg13g2_nor2_2
X_5642_ net1876 net1758 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_2854_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q net132 net1703
+ net1921 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q
+ _0925_ VPWR VGND sg13g2_mux4_1
X_2785_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q
+ _0859_ _0856_ _0860_ _0857_ sg13g2_a221oi_1
X_5573_ net1874 net1791 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_4524_ VPWR _0081_ net1934 VGND sg13g2_inv_1
XFILLER_116_188 VPWR VGND sg13g2_fill_1
X_4455_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q net1517
+ _2371_ _2370_ sg13g2_a21oi_1
X_4386_ _2312_ _2311_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q
+ _2309_ _2308_ VPWR VGND sg13g2_a22oi_1
X_3406_ _1167_ VPWR _1458_ VGND _1164_ _1168_ sg13g2_o21ai_1
X_6125_ Tile_X0Y0_W6END[2] net346 VPWR VGND sg13g2_buf_1
X_3337_ VGND VPWR _1380_ _1382_ _1389_ _1384_ sg13g2_a21oi_1
X_3268_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q VPWR _1321_ VGND
+ net165 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q sg13g2_o21ai_1
X_6056_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 net277 VPWR VGND sg13g2_buf_1
XFILLER_38_172 VPWR VGND sg13g2_decap_8
X_5007_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q VPWR _0547_ VGND
+ net1660 net1581 sg13g2_o21ai_1
X_3199_ _1254_ _1252_ _1253_ VPWR VGND sg13g2_nand2_1
XFILLER_53_120 VPWR VGND sg13g2_fill_2
XFILLER_41_304 VPWR VGND sg13g2_fill_1
XFILLER_39_63 VPWR VGND sg13g2_fill_1
XFILLER_76_212 VPWR VGND sg13g2_decap_4
XFILLER_39_85 VPWR VGND sg13g2_fill_2
XFILLER_29_172 VPWR VGND sg13g2_fill_1
XFILLER_29_194 VPWR VGND sg13g2_fill_2
XFILLER_55_40 VPWR VGND sg13g2_decap_4
XFILLER_71_61 VPWR VGND sg13g2_fill_1
Xoutput307 net307 Tile_X0Y0_N4BEG[8] VPWR VGND sg13g2_buf_1
X_2570_ VGND VPWR net6 net1682 _0656_ _0655_ sg13g2_a21oi_1
Xoutput318 net318 Tile_X0Y0_NN4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput329 net329 Tile_X0Y0_W1BEG[3] VPWR VGND sg13g2_buf_1
X_4240_ _0165_ VPWR _2201_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q
+ net1518 sg13g2_o21ai_1
X_4171_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q VPWR _2142_
+ VGND _2140_ _2141_ sg13g2_o21ai_1
X_3122_ _1163_ _1178_ _1179_ VPWR VGND sg13g2_nor2b_1
X_3053_ _1113_ _1111_ _1112_ VPWR VGND sg13g2_xnor2_1
X_3955_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q _1963_
+ _1964_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q sg13g2_a21oi_1
X_2906_ _0972_ VPWR _0973_ VGND _0971_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q
+ sg13g2_o21ai_1
X_5625_ net1908 net1770 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_3886_ VGND VPWR _1879_ _1900_ _1880_ _1835_ sg13g2_a21oi_2
X_2837_ _0908_ VPWR _0909_ VGND net1667 net1563 sg13g2_o21ai_1
X_5556_ net1898 net1794 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_2768_ _0840_ _0838_ _0843_ _0844_ VPWR VGND sg13g2_a21o_1
X_2699_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q _0777_ _0774_
+ _0778_ VPWR VGND sg13g2_nor3_2
X_5487_ net1886 net1849 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_4507_ VPWR _0064_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q VGND
+ sg13g2_inv_1
XFILLER_104_103 VPWR VGND sg13g2_decap_8
X_4438_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q _2355_ _2356_
+ VPWR VGND sg13g2_nor2_1
X_4369_ VGND VPWR _0167_ _2296_ _2297_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q
+ sg13g2_a21oi_1
XFILLER_76_28 VPWR VGND sg13g2_fill_2
X_6108_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 net329 VPWR VGND sg13g2_buf_1
XFILLER_100_342 VPWR VGND sg13g2_fill_2
XFILLER_73_215 VPWR VGND sg13g2_decap_8
X_6039_ net1743 net270 VPWR VGND sg13g2_buf_1
Xrebuffer72 _0327_ net681 VPWR VGND sg13g2_buf_8
Xrebuffer94 _0417_ net703 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer83 _0289_ net692 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_49_223 VPWR VGND sg13g2_fill_2
XFILLER_49_245 VPWR VGND sg13g2_fill_1
X_3740_ _1770_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q _1771_
+ VPWR VGND sg13g2_nor2b_1
X_3671_ Tile_X0Y1_DSP_bot.C6 _1700_ _1706_ _1698_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q
+ VPWR VGND sg13g2_a22oi_1
X_5410_ net1970 net1818 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_2622_ net1675 net1598 net1603 net1623 net1633 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q
+ _0704_ VPWR VGND sg13g2_mux4_1
X_2553_ _0638_ VPWR _0639_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ net1593 sg13g2_o21ai_1
X_5341_ net1959 net1842 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_2484_ _0573_ VPWR _0574_ VGND net154 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q
+ sg13g2_o21ai_1
X_5272_ net1977 net1742 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_4223_ _2185_ _2186_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 VPWR VGND sg13g2_mux2_1
X_4154_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q _0598_ net2001
+ net29 net1626 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q _2126_
+ VPWR VGND sg13g2_mux4_1
X_3105_ _1162_ _1160_ _1161_ VPWR VGND sg13g2_nand2b_1
X_4085_ _2078_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q _2081_
+ _2082_ VPWR VGND sg13g2_a21o_1
XFILLER_95_384 VPWR VGND sg13g2_fill_1
X_3036_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q _1097_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q _1096_ sg13g2_a21oi_2
XFILLER_70_218 VPWR VGND sg13g2_decap_8
X_4987_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q net1596 net1609
+ net1602 net1630 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q _0528_
+ VPWR VGND sg13g2_mux4_1
X_3938_ _1931_ _1947_ _1948_ VPWR VGND sg13g2_nor2_2
X_3869_ _1890_ _1818_ _1819_ VPWR VGND sg13g2_xnor2_1
X_5608_ net1871 net1774 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_117_261 VPWR VGND sg13g2_fill_1
X_5539_ net1866 net1801 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_78_329 VPWR VGND sg13g2_fill_1
XFILLER_100_161 VPWR VGND sg13g2_decap_4
XFILLER_52_74 VPWR VGND sg13g2_fill_2
Xinput28 Tile_X0Y0_S1END[2] net28 VPWR VGND sg13g2_buf_1
XFILLER_52_96 VPWR VGND sg13g2_fill_2
Xinput17 Tile_X0Y0_E2MID[5] net17 VPWR VGND sg13g2_buf_1
Xinput39 Tile_X0Y0_S2MID[1] net39 VPWR VGND sg13g2_buf_1
XFILLER_6_344 VPWR VGND sg13g2_fill_2
XFILLER_108_283 VPWR VGND sg13g2_fill_2
XFILLER_69_329 VPWR VGND sg13g2_fill_1
XFILLER_96_104 VPWR VGND sg13g2_decap_4
XFILLER_96_115 VPWR VGND sg13g2_fill_2
Xfanout1841 net1844 net1841 VPWR VGND sg13g2_buf_1
Xfanout1852 net1853 net1852 VPWR VGND sg13g2_buf_1
Xfanout1830 net1831 net1830 VPWR VGND sg13g2_buf_1
Xfanout1874 Tile_X0Y1_FrameData[2] net1874 VPWR VGND sg13g2_buf_1
Xfanout1863 Tile_X0Y1_FrameData[6] net1863 VPWR VGND sg13g2_buf_1
Xfanout1885 Tile_X0Y1_FrameData[25] net1885 VPWR VGND sg13g2_buf_1
XFILLER_77_351 VPWR VGND sg13g2_fill_2
Xfanout1896 Tile_X0Y1_FrameData[1] net1896 VPWR VGND sg13g2_buf_1
X_4910_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q _0450_ _0455_
+ _0456_ VPWR VGND sg13g2_nor3_1
X_5890_ net1865 net1816 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_4841_ _0388_ VPWR _0389_ VGND net1684 net1590 sg13g2_o21ai_1
XFILLER_20_137 VPWR VGND sg13g2_fill_1
X_4772_ _0315_ VPWR _0323_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q
+ _0322_ sg13g2_o21ai_1
X_3723_ net1708 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q _1755_
+ VPWR VGND sg13g2_nor2_1
X_3654_ net1646 _1689_ _1690_ VPWR VGND sg13g2_nor2_1
X_2605_ VGND VPWR _0688_ _0689_ _0684_ _0686_ sg13g2_a21oi_2
X_3585_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q net1567
+ _1626_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q sg13g2_a21oi_1
X_2536_ net1660 net1712 net120 net1927 net96 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q
+ _0623_ VPWR VGND sg13g2_mux4_1
X_5324_ net1991 net1722 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_5255_ net1981 net1743 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_4206_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q VPWR _2172_
+ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q _2171_ sg13g2_o21ai_1
XFILLER_68_362 VPWR VGND sg13g2_fill_2
X_5186_ net1969 net1763 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_28_215 VPWR VGND sg13g2_fill_1
XFILLER_68_384 VPWR VGND sg13g2_fill_1
X_4137_ _2106_ _2112_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 VPWR VGND
+ sg13g2_nor2_1
X_4068_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q
+ _2064_ _2061_ _2065_ _2062_ sg13g2_a221oi_1
X_3019_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q VPWR _1081_ VGND
+ _1077_ _1080_ sg13g2_o21ai_1
XFILLER_51_273 VPWR VGND sg13g2_decap_4
XFILLER_3_303 VPWR VGND sg13g2_fill_2
XFILLER_3_347 VPWR VGND sg13g2_fill_1
Xoutput490 net490 Tile_X0Y1_SS4BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_78_159 VPWR VGND sg13g2_fill_2
XFILLER_47_52 VPWR VGND sg13g2_fill_2
XFILLER_27_292 VPWR VGND sg13g2_fill_2
X_3370_ _0807_ net1568 _1415_ _1420_ _1422_ VPWR VGND sg13g2_and4_1
X_5040_ net1938 net1855 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
Xfanout1660 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q net1660 VPWR
+ VGND sg13g2_buf_1
Xfanout1671 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q net1671 VPWR
+ VGND sg13g2_buf_1
Xfanout1693 net1694 net1693 VPWR VGND sg13g2_buf_1
Xfanout1682 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q net1682 VPWR
+ VGND sg13g2_buf_1
X_5457__589 VPWR VGND net589 sg13g2_tiehi
XFILLER_92_195 VPWR VGND sg13g2_decap_4
X_5873_ net1891 net1814 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_4824_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q net1710 net92
+ net116 net1921 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q _0373_
+ VPWR VGND sg13g2_mux4_1
X_4755_ _0307_ _0306_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q
+ VPWR VGND sg13g2_nand2b_1
X_3706_ _0016_ net1648 _1738_ _1739_ VPWR VGND sg13g2_a21o_1
X_4686_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q VPWR _0240_ VGND
+ net1676 net1525 sg13g2_o21ai_1
X_3637_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q net116 net110
+ net1936 net152 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q _1674_
+ VPWR VGND sg13g2_mux4_1
X_3568_ _0137_ net725 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q
+ _1610_ VPWR VGND sg13g2_mux4_1
X_5307_ net1953 net1721 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_2519_ _0606_ VPWR _0607_ VGND net66 net1681 sg13g2_o21ai_1
X_6287_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 net508 VPWR VGND sg13g2_buf_1
X_3499_ _1546_ net1581 net1669 VPWR VGND sg13g2_nand2b_1
X_5238_ net1950 net1754 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_310 VPWR VGND sg13g2_fill_2
X_5169_ net1940 net1775 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_68_192 VPWR VGND sg13g2_fill_1
XFILLER_83_151 VPWR VGND sg13g2_fill_1
XFILLER_33_76 VPWR VGND sg13g2_fill_1
XFILLER_123_2 VPWR VGND sg13g2_fill_1
XFILLER_109_0 VPWR VGND sg13g2_fill_2
XFILLER_3_199 VPWR VGND sg13g2_fill_1
XFILLER_59_181 VPWR VGND sg13g2_decap_8
XFILLER_47_365 VPWR VGND sg13g2_fill_2
XFILLER_59_192 VPWR VGND sg13g2_fill_1
XFILLER_74_162 VPWR VGND sg13g2_fill_1
XFILLER_74_173 VPWR VGND sg13g2_fill_1
XFILLER_15_240 VPWR VGND sg13g2_fill_1
X_2870_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q VPWR _0940_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q _0938_ sg13g2_o21ai_1
X_4540_ VPWR _0097_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q VGND
+ sg13g2_inv_1
X_4471_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q _2384_ _2385_
+ VPWR VGND sg13g2_nor2b_1
X_6210_ net1857 net453 VPWR VGND sg13g2_buf_1
X_3422_ VGND VPWR _0133_ net1645 _1473_ net1650 sg13g2_a21oi_1
X_6141_ Tile_X0Y0_WW4END[8] net368 VPWR VGND sg13g2_buf_1
X_3353_ _1405_ _1371_ _1385_ VPWR VGND sg13g2_xnor2_1
X_6072_ Tile_X0Y1_N4END[8] net293 VPWR VGND sg13g2_buf_1
X_3284_ _1306_ _1305_ _1336_ VPWR VGND sg13g2_xor2_1
X_5023_ net1963 net1855 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_65_162 VPWR VGND sg13g2_decap_8
X_5856_ net1861 net1821 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_243 VPWR VGND sg13g2_decap_4
X_4807_ _0356_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q _0357_
+ VPWR VGND sg13g2_nor2b_1
X_2999_ _1061_ VPWR _1062_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q
+ _1059_ sg13g2_o21ai_1
X_5787_ net1912 net1714 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_4738_ VPWR _0290_ net692 VGND sg13g2_inv_1
X_4669_ VGND VPWR net64 net1699 _0225_ _0224_ sg13g2_a21oi_1
XFILLER_88_254 VPWR VGND sg13g2_decap_8
XFILLER_88_265 VPWR VGND sg13g2_fill_1
XFILLER_44_335 VPWR VGND sg13g2_fill_2
XFILLER_71_165 VPWR VGND sg13g2_fill_1
XFILLER_44_64 VPWR VGND sg13g2_fill_2
XFILLER_60_63 VPWR VGND sg13g2_decap_8
XFILLER_39_129 VPWR VGND sg13g2_fill_2
XFILLER_47_195 VPWR VGND sg13g2_fill_2
X_3971_ _1978_ _1932_ _1976_ VPWR VGND sg13g2_nand2_2
XFILLER_50_349 VPWR VGND sg13g2_fill_1
X_2922_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q net1531 net1537
+ net1545 net1552 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q _0988_
+ VPWR VGND sg13g2_mux4_1
X_5710_ net1884 net1739 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_5641_ net1872 net1758 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_2853_ _0913_ VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q
+ _0924_ sg13g2_o21ai_1
X_2784_ VGND VPWR net9 net1690 _0859_ _0858_ sg13g2_a21oi_1
X_5572_ net1868 net1791 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_4523_ VPWR _0080_ net19 VGND sg13g2_inv_1
XFILLER_116_134 VPWR VGND sg13g2_fill_1
X_4454_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q _1780_ _2370_
+ VPWR VGND sg13g2_nor2_1
X_4385_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q net1517
+ _2311_ _2310_ sg13g2_a21oi_1
X_3405_ _1457_ _1173_ _1176_ VPWR VGND sg13g2_nand2_1
X_3336_ _1388_ _1387_ _1386_ VPWR VGND sg13g2_nand2b_1
X_6124_ net80 net345 VPWR VGND sg13g2_buf_1
XFILLER_112_384 VPWR VGND sg13g2_fill_1
X_6055_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 net276 VPWR VGND sg13g2_buf_8
X_5006_ net1561 net1571 net1660 _0546_ VPWR VGND sg13g2_mux2_1
X_3267_ _0626_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q _1320_
+ VPWR VGND _0552_ sg13g2_nand3b_1
X_3198_ _1253_ _1243_ _1245_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_324 VPWR VGND sg13g2_fill_1
X_5472__604 VPWR VGND net604 sg13g2_tiehi
X_5839_ net1887 net1821 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_29_162 VPWR VGND sg13g2_fill_2
XFILLER_44_121 VPWR VGND sg13g2_decap_4
XFILLER_17_379 VPWR VGND sg13g2_fill_2
XFILLER_44_165 VPWR VGND sg13g2_fill_1
Xoutput308 net308 Tile_X0Y0_N4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput319 net319 Tile_X0Y0_NN4BEG[4] VPWR VGND sg13g2_buf_1
X_4170_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q VPWR _2141_
+ VGND _0162_ _0257_ sg13g2_o21ai_1
X_3121_ _1177_ _1176_ _1178_ VPWR VGND sg13g2_and2_1
XFILLER_96_81 VPWR VGND sg13g2_fill_1
X_3052_ _1009_ _1008_ _1112_ VPWR VGND sg13g2_xor2_1
XFILLER_82_249 VPWR VGND sg13g2_decap_4
XFILLER_35_198 VPWR VGND sg13g2_fill_2
XFILLER_90_260 VPWR VGND sg13g2_decap_8
XFILLER_90_271 VPWR VGND sg13g2_fill_2
X_3954_ VGND VPWR net11 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q
+ _1963_ _1962_ sg13g2_a21oi_1
XFILLER_91_0 VPWR VGND sg13g2_fill_1
XFILLER_50_179 VPWR VGND sg13g2_decap_8
X_2905_ _0972_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[5\]
+ VPWR VGND sg13g2_nand2_1
X_3885_ _1899_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 VGND _1898_
+ net1656 sg13g2_o21ai_1
X_5624_ net1906 net1770 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_2836_ VGND VPWR net1667 net1569 _0908_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q
+ sg13g2_a21oi_1
X_5555_ net1894 net1794 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_2767_ _0843_ _0842_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q
+ VPWR VGND sg13g2_nand2b_1
X_2698_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q _0775_ _0776_
+ _0777_ VPWR VGND sg13g2_nor3_1
X_5486_ net1884 net1849 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_4506_ VPWR _0063_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q VGND
+ sg13g2_inv_1
X_4437_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q net1555
+ _2355_ _2354_ sg13g2_a21oi_1
XFILLER_104_137 VPWR VGND sg13g2_decap_8
X_4368_ net1713 net1928 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q
+ _2296_ VPWR VGND sg13g2_mux2_1
X_6107_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 net328 VPWR VGND sg13g2_buf_1
X_4299_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q _2241_ _2245_
+ _2239_ _2243_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q _2246_
+ VPWR VGND sg13g2_mux4_1
X_3319_ _1371_ _1242_ _1350_ VPWR VGND sg13g2_xnor2_1
X_6038_ net1755 net269 VPWR VGND sg13g2_buf_1
Xrebuffer73 _1433_ net682 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer40 net649 net648 VPWR VGND sg13g2_buf_16
Xrebuffer84 _0289_ net693 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer95 _1801_ net704 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_41_113 VPWR VGND sg13g2_fill_2
Xrebuffer130 net740 net739 VPWR VGND sg13g2_buf_2
XFILLER_41_87 VPWR VGND sg13g2_fill_1
XFILLER_103_170 VPWR VGND sg13g2_fill_2
XFILLER_66_51 VPWR VGND sg13g2_fill_1
XFILLER_66_62 VPWR VGND sg13g2_fill_1
XFILLER_57_290 VPWR VGND sg13g2_decap_4
XFILLER_17_198 VPWR VGND sg13g2_fill_1
X_3670_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q _1705_ _1706_
+ VPWR VGND sg13g2_nor2b_1
X_2621_ _0701_ VPWR _0703_ VGND net1642 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X
+ sg13g2_o21ai_1
X_2552_ _0638_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q net1588
+ VPWR VGND sg13g2_nand2b_1
X_5340_ net1957 net1842 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_5271_ net1955 net1744 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_99_113 VPWR VGND sg13g2_fill_1
X_2483_ _0573_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q net168
+ VPWR VGND sg13g2_nand2b_1
X_4222_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q net699 _1470_
+ net623 _0513_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q _2186_
+ VPWR VGND sg13g2_mux4_1
XFILLER_101_118 VPWR VGND sg13g2_fill_1
X_4153_ _2125_ _2124_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 VPWR VGND sg13g2_mux2_1
X_3104_ _1158_ _1157_ _1161_ VPWR VGND sg13g2_xor2_1
X_4084_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q VPWR _2081_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q _2080_ sg13g2_o21ai_1
X_3035_ VGND VPWR _1095_ _1096_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 sg13g2_a21oi_2
X_4986_ _0524_ _0521_ _0526_ _0527_ VPWR VGND sg13g2_a21o_1
X_3937_ _1933_ VPWR _1947_ VGND _1946_ net1649 sg13g2_o21ai_1
XFILLER_109_218 VPWR VGND sg13g2_fill_1
X_3868_ _1889_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[5\] net1652 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ VPWR VGND sg13g2_mux2_1
X_5607_ net1919 net1781 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_2819_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q
+ _0891_ _0892_ VPWR VGND sg13g2_a21o_1
X_3799_ VGND VPWR _1538_ _1828_ _1826_ _1827_ sg13g2_a21oi_2
X_5538_ net1864 net1801 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_5469_ Tile_X0Y1_UserCLK net601 Tile_X0Y1_DSP_bot.C9 _0007_ _5469_/Q VPWR VGND sg13g2_dfrbp_1
XFILLER_86_330 VPWR VGND sg13g2_fill_1
XFILLER_46_249 VPWR VGND sg13g2_fill_2
XFILLER_36_54 VPWR VGND sg13g2_fill_1
XFILLER_52_20 VPWR VGND sg13g2_decap_8
Xinput18 Tile_X0Y0_E2MID[6] net18 VPWR VGND sg13g2_buf_1
Xinput29 Tile_X0Y0_S1END[3] net29 VPWR VGND sg13g2_buf_1
XFILLER_6_378 VPWR VGND sg13g2_fill_2
XFILLER_69_319 VPWR VGND sg13g2_fill_2
Xfanout1820 Tile_X0Y1_FrameStrobe[12] net1820 VPWR VGND sg13g2_buf_1
Xfanout1831 net1832 net1831 VPWR VGND sg13g2_buf_1
Xfanout1842 net1843 net1842 VPWR VGND sg13g2_buf_1
Xfanout1875 Tile_X0Y1_FrameData[2] net1875 VPWR VGND sg13g2_buf_1
Xfanout1864 Tile_X0Y1_FrameData[5] net1864 VPWR VGND sg13g2_buf_1
Xfanout1853 net1855 net1853 VPWR VGND sg13g2_buf_1
Xfanout1897 Tile_X0Y1_FrameData[1] net1897 VPWR VGND sg13g2_buf_1
Xfanout1886 Tile_X0Y1_FrameData[24] net1886 VPWR VGND sg13g2_buf_1
XFILLER_45_260 VPWR VGND sg13g2_decap_4
X_4840_ _0388_ net1684 net1585 VPWR VGND sg13g2_nand2_1
X_4771_ _0321_ VPWR _0322_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q
+ _0316_ sg13g2_o21ai_1
X_3722_ _1754_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q _0867_
+ VPWR VGND sg13g2_nand2_1
XFILLER_9_183 VPWR VGND sg13g2_fill_2
X_3653_ VPWR Tile_X0Y1_DSP_bot.C7 _1689_ VGND sg13g2_inv_1
X_2604_ _0097_ VPWR _0688_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q
+ _0687_ sg13g2_o21ai_1
X_3584_ VGND VPWR _0148_ _1624_ _1625_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q
+ sg13g2_a21oi_1
XFILLER_54_0 VPWR VGND sg13g2_decap_8
X_5323_ net1989 net1722 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_2535_ VPWR _0622_ _0621_ VGND sg13g2_inv_1
X_5254_ net1979 net1743 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_4205_ _2170_ VPWR _2171_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q
+ net1526 sg13g2_o21ai_1
X_5185_ net1967 net1766 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_4136_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q _2108_
+ _2112_ _2111_ sg13g2_a21oi_1
X_4067_ VGND VPWR _0075_ net1694 _2064_ _2063_ sg13g2_a21oi_1
X_3018_ _1080_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q _1079_
+ VPWR VGND sg13g2_nand2_1
X_4969_ _0511_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q _0510_
+ VPWR VGND sg13g2_nand2_1
XFILLER_22_56 VPWR VGND sg13g2_fill_1
Xoutput480 net480 Tile_X0Y1_S4BEG[15] VPWR VGND sg13g2_buf_1
XFILLER_105_254 VPWR VGND sg13g2_fill_1
Xoutput491 net491 Tile_X0Y1_SS4BEG[10] VPWR VGND sg13g2_buf_8
XFILLER_19_205 VPWR VGND sg13g2_fill_2
XFILLER_47_86 VPWR VGND sg13g2_fill_2
XFILLER_42_241 VPWR VGND sg13g2_decap_8
XFILLER_8_25 VPWR VGND sg13g2_fill_2
XFILLER_6_186 VPWR VGND sg13g2_fill_2
XFILLER_111_235 VPWR VGND sg13g2_fill_2
XFILLER_26_4 VPWR VGND sg13g2_fill_1
Xfanout1650 net1651 net1650 VPWR VGND sg13g2_buf_1
Xfanout1661 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q net1661 VPWR
+ VGND sg13g2_buf_1
Xfanout1694 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q net1694 VPWR
+ VGND sg13g2_buf_1
XFILLER_77_182 VPWR VGND sg13g2_fill_2
Xfanout1683 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q net1683 VPWR
+ VGND sg13g2_buf_1
Xfanout1672 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q net1672 VPWR
+ VGND sg13g2_buf_1
XFILLER_65_355 VPWR VGND sg13g2_fill_2
XFILLER_92_141 VPWR VGND sg13g2_fill_2
XFILLER_92_163 VPWR VGND sg13g2_fill_1
X_5872_ net1889 net1814 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_4823_ _0372_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q _0371_
+ VPWR VGND sg13g2_nand2_1
X_4754_ _0305_ _0304_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q
+ _0306_ VPWR VGND sg13g2_mux2_1
X_3705_ VGND VPWR net1637 Tile_X0Y1_DSP_bot.C4 _1738_ _1737_ sg13g2_a21oi_1
X_4685_ VGND VPWR net1676 net1585 _0239_ _0238_ sg13g2_a21oi_1
X_3636_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q net139 net151
+ net1923 _0741_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q _1673_
+ VPWR VGND sg13g2_mux4_1
X_3567_ _1609_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 _0137_ VPWR VGND
+ sg13g2_nand2_2
X_6286_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 net507 VPWR VGND sg13g2_buf_8
XFILLER_0_307 VPWR VGND sg13g2_fill_2
X_5306_ net1951 net1721 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_2518_ _0606_ _0076_ net1681 VPWR VGND sg13g2_nand2_1
X_3498_ _1544_ VPWR _1545_ VGND net1669 net1555 sg13g2_o21ai_1
X_5237_ net1947 net1751 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_68_160 VPWR VGND sg13g2_fill_1
X_5168_ net1938 net1775 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_5099_ net1989 net1795 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_4119_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q net20 net48
+ net33 net1609 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1
+ VPWR VGND sg13g2_mux4_1
XFILLER_71_369 VPWR VGND sg13g2_fill_2
XFILLER_3_156 VPWR VGND sg13g2_fill_1
XFILLER_58_63 VPWR VGND sg13g2_fill_2
XFILLER_47_344 VPWR VGND sg13g2_fill_2
XFILLER_62_358 VPWR VGND sg13g2_fill_1
XFILLER_30_244 VPWR VGND sg13g2_fill_2
X_4470_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3
+ net617 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q _2384_ VPWR VGND sg13g2_mux4_1
X_3421_ _1472_ net1638 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X
+ VPWR VGND sg13g2_nand2_1
X_6140_ Tile_X0Y0_WW4END[7] net367 VPWR VGND sg13g2_buf_1
X_3352_ _1404_ _1395_ _1403_ VPWR VGND sg13g2_nand2_2
X_6071_ net725 net292 VPWR VGND sg13g2_buf_1
X_3283_ _1333_ _1308_ _1335_ VPWR VGND sg13g2_xor2_1
XFILLER_97_255 VPWR VGND sg13g2_decap_8
X_5022_ net1962 net1855 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_97_288 VPWR VGND sg13g2_fill_2
XFILLER_97_299 VPWR VGND sg13g2_fill_2
XFILLER_17_0 VPWR VGND sg13g2_fill_2
XFILLER_110_38 VPWR VGND sg13g2_fill_1
X_5855_ net1858 net1823 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_4806_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q _0354_
+ _0356_ _0355_ sg13g2_a21oi_1
XFILLER_119_110 VPWR VGND sg13g2_fill_1
X_2998_ _1061_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q _1060_
+ VPWR VGND sg13g2_nand2b_1
X_5786_ net1910 net1714 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_4737_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q net124 net100
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 net160 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q
+ _0289_ VPWR VGND sg13g2_mux4_1
X_4668_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q VPWR _0224_ VGND
+ _0086_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q sg13g2_o21ai_1
X_3619_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q _0723_ net148
+ net1934 net1704 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q _1658_
+ VPWR VGND sg13g2_mux4_1
XFILLER_102_8 VPWR VGND sg13g2_fill_1
X_4599_ VPWR _0156_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q VGND
+ sg13g2_inv_1
XFILLER_115_371 VPWR VGND sg13g2_fill_2
X_6269_ Tile_X0Y0_SS4END[8] net490 VPWR VGND sg13g2_buf_1
XFILLER_121_0 VPWR VGND sg13g2_fill_2
XFILLER_69_73 VPWR VGND sg13g2_decap_8
XFILLER_94_203 VPWR VGND sg13g2_fill_2
XFILLER_47_152 VPWR VGND sg13g2_fill_2
X_3970_ _1976_ _1932_ _1977_ VPWR VGND sg13g2_nor2_2
X_2921_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 _0980_ _0987_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q
+ _0978_ VPWR VGND sg13g2_a22oi_1
X_5640_ net1870 net1758 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_2852_ _0918_ VPWR _0924_ VGND _0920_ _0923_ sg13g2_o21ai_1
X_2783_ net1690 net2004 _0858_ VPWR VGND sg13g2_nor2b_1
X_5571_ net1866 net1790 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_4522_ VPWR _0079_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q VGND
+ sg13g2_inv_1
X_4453_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q _1277_
+ _2369_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q sg13g2_a21oi_1
X_3404_ _1456_ _1455_ _1238_ _1180_ VPWR VGND sg13g2_and3_1
XFILLER_104_319 VPWR VGND sg13g2_fill_1
X_4384_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q _1780_ _2310_
+ VPWR VGND sg13g2_nor2_1
X_3335_ _1387_ _1360_ _1361_ VPWR VGND sg13g2_xnor2_1
X_6123_ net79 net344 VPWR VGND sg13g2_buf_1
X_3266_ _1318_ VPWR _1319_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q
+ _1315_ sg13g2_o21ai_1
X_5005_ net1660 net1532 net1536 net1545 net1552 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q
+ _0545_ VPWR VGND sg13g2_mux4_1
X_3197_ _1252_ _1246_ _1250_ VPWR VGND sg13g2_xnor2_1
XFILLER_41_317 VPWR VGND sg13g2_fill_2
X_5838_ net1885 net1821 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_5769_ net1873 net1717 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_5_207 VPWR VGND sg13g2_fill_1
XFILLER_29_196 VPWR VGND sg13g2_fill_1
XFILLER_44_111 VPWR VGND sg13g2_fill_2
XFILLER_40_361 VPWR VGND sg13g2_fill_1
Xoutput309 net309 Tile_X0Y0_NN4BEG[0] VPWR VGND sg13g2_buf_1
X_3120_ _1048_ _1051_ _1175_ _1177_ VPWR VGND sg13g2_or3_1
X_3051_ _1110_ VPWR _1111_ VGND _0932_ _1106_ sg13g2_o21ai_1
X_3953_ net1700 net2001 _1962_ VPWR VGND sg13g2_nor2b_1
X_2904_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X
+ _0971_ VGND sg13g2_inv_1
X_3884_ _1899_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[12\] net1656 VPWR VGND sg13g2_nand2_1
X_2835_ VGND VPWR _0907_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q
+ _0906_ sg13g2_or2_1
X_5623_ net1904 net1773 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_84_0 VPWR VGND sg13g2_fill_2
X_5554_ net1892 net1794 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_2766_ _0841_ VPWR _0842_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 sg13g2_o21ai_1
X_5485_ net1883 net1845 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_2697_ net1709 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q _0776_
+ VPWR VGND sg13g2_nor2_1
X_4505_ VPWR _0062_ net48 VGND sg13g2_inv_1
X_4436_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q VPWR _2354_ VGND
+ net147 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q sg13g2_o21ai_1
XFILLER_116_48 VPWR VGND sg13g2_fill_2
X_4367_ _2294_ VPWR _2295_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q
+ net703 sg13g2_o21ai_1
X_6106_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 net327 VPWR VGND sg13g2_buf_1
X_3318_ _1368_ _1369_ _1370_ VPWR VGND sg13g2_nor2_1
X_4298_ VGND VPWR net1936 net1663 _2245_ _2244_ sg13g2_a21oi_1
X_3249_ _1247_ _1300_ _1302_ VPWR VGND sg13g2_nor2_1
X_6037_ net1767 net268 VPWR VGND sg13g2_buf_1
Xrebuffer30 net638 net639 VPWR VGND sg13g2_buf_1
Xrebuffer74 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 net683 VPWR VGND
+ sg13g2_dlygate4sd1_1
Xrebuffer85 _0681_ net694 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer96 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 net705 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer120 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 net729 VPWR VGND
+ sg13g2_dlygate4sd1_1
Xrebuffer131 net741 net740 VPWR VGND sg13g2_buf_2
XFILLER_1_221 VPWR VGND sg13g2_fill_2
XFILLER_9_343 VPWR VGND sg13g2_fill_1
X_2620_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[6\] net1642 _0702_ VPWR VGND sg13g2_mux2_2
X_2551_ VGND VPWR _0632_ _0634_ _0637_ _0636_ sg13g2_a21oi_1
X_2482_ _0572_ _0571_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q
+ VPWR VGND sg13g2_nand2b_1
X_5270_ net1949 net1744 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_4221_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q net1527 net1933
+ net2004 net691 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q _2185_
+ VPWR VGND sg13g2_mux4_1
XFILLER_99_147 VPWR VGND sg13g2_decap_8
XFILLER_99_158 VPWR VGND sg13g2_fill_2
X_4152_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q net1516 net28
+ net3 net1606 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q _2125_
+ VPWR VGND sg13g2_mux4_1
X_3103_ _1152_ _0769_ _1154_ _1160_ VPWR VGND sg13g2_a21o_1
X_4083_ VGND VPWR net1693 net1584 _2080_ _2079_ sg13g2_a21oi_1
X_3034_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q net161 _1095_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_63_294 VPWR VGND sg13g2_fill_2
X_4985_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q VPWR _0526_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q _0525_ sg13g2_o21ai_1
X_3936_ VGND VPWR net1644 _0033_ _1946_ _1945_ sg13g2_a21oi_1
X_3867_ _1889_ _1815_ _1817_ VPWR VGND sg13g2_xnor2_1
X_5606_ net1896 net1780 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_2818_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q VPWR _0891_ VGND
+ _0087_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q sg13g2_o21ai_1
X_3798_ _1827_ _1536_ _1509_ VPWR VGND sg13g2_xnor2_1
XFILLER_117_252 VPWR VGND sg13g2_fill_2
X_5537_ net1862 net1801 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_2749_ VGND VPWR _0076_ net1698 _0826_ _0825_ sg13g2_a21oi_1
XFILLER_11_69 VPWR VGND sg13g2_fill_2
X_5468_ Tile_X0Y1_UserCLK net600 Tile_X0Y1_DSP_bot.C8 _0009_ _5468_/Q VPWR VGND sg13g2_dfrbp_1
XFILLER_78_309 VPWR VGND sg13g2_fill_2
X_4419_ VGND VPWR _0065_ _0169_ _2339_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q
+ sg13g2_a21oi_1
X_5399_ net1956 net1827 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_36_11 VPWR VGND sg13g2_decap_4
XFILLER_52_76 VPWR VGND sg13g2_fill_1
XFILLER_52_98 VPWR VGND sg13g2_fill_1
Xinput19 Tile_X0Y0_E2MID[7] net19 VPWR VGND sg13g2_buf_1
XFILLER_10_375 VPWR VGND sg13g2_fill_2
XFILLER_108_285 VPWR VGND sg13g2_fill_1
XFILLER_96_117 VPWR VGND sg13g2_fill_1
Xfanout1821 net1823 net1821 VPWR VGND sg13g2_buf_1
Xfanout1832 Tile_X0Y1_FrameStrobe[11] net1832 VPWR VGND sg13g2_buf_1
Xfanout1810 net1811 net1810 VPWR VGND sg13g2_buf_1
Xfanout1843 net1844 net1843 VPWR VGND sg13g2_buf_1
Xfanout1865 Tile_X0Y1_FrameData[5] net1865 VPWR VGND sg13g2_buf_1
Xfanout1876 Tile_X0Y1_FrameData[29] net1876 VPWR VGND sg13g2_buf_1
Xfanout1854 net1855 net1854 VPWR VGND sg13g2_buf_1
Xfanout1898 Tile_X0Y1_FrameData[19] net1898 VPWR VGND sg13g2_buf_1
XFILLER_37_217 VPWR VGND sg13g2_decap_8
XFILLER_37_228 VPWR VGND sg13g2_fill_1
Xfanout1887 Tile_X0Y1_FrameData[24] net1887 VPWR VGND sg13g2_buf_1
XFILLER_20_117 VPWR VGND sg13g2_fill_1
X_4770_ _0320_ VPWR _0321_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q
+ _0319_ sg13g2_o21ai_1
X_3721_ _1750_ _1752_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q
+ _1753_ VPWR VGND sg13g2_nand3_1
X_3652_ _1677_ VPWR _1689_ VGND _1688_ _1682_ sg13g2_o21ai_1
X_3583_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q net114 net122
+ net1925 net98 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q _1624_
+ VPWR VGND sg13g2_mux4_1
X_2603_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q net1711 net1926
+ net121 net97 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q _0687_
+ VPWR VGND sg13g2_mux4_1
X_5322_ net1988 net1723 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_2534_ _0620_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q _0621_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_114_233 VPWR VGND sg13g2_fill_2
XFILLER_47_0 VPWR VGND sg13g2_fill_1
X_5253_ net1976 net1741 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_68_320 VPWR VGND sg13g2_fill_1
X_4204_ _2170_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q _0630_
+ VPWR VGND sg13g2_nand2_2
X_5184_ net1965 net1767 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_68_364 VPWR VGND sg13g2_fill_1
X_4135_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q VPWR _2111_
+ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q _2110_ sg13g2_o21ai_1
XFILLER_113_27 VPWR VGND sg13g2_decap_4
X_4066_ net1694 net5 _2063_ VPWR VGND sg13g2_nor2_1
X_3017_ _1078_ VPWR _1079_ VGND net1665 net1565 sg13g2_o21ai_1
X_4968_ _0509_ VPWR _0510_ VGND net135 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q
+ sg13g2_o21ai_1
X_4899_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q _0443_
+ _0445_ _0444_ sg13g2_a21oi_1
XFILLER_11_139 VPWR VGND sg13g2_fill_2
X_3919_ _1930_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[15\] net1655 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ VPWR VGND sg13g2_mux2_2
XFILLER_3_305 VPWR VGND sg13g2_fill_1
Xoutput470 net470 Tile_X0Y1_S2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput492 net492 Tile_X0Y1_SS4BEG[11] VPWR VGND sg13g2_buf_8
Xoutput481 net481 Tile_X0Y1_S4BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_78_139 VPWR VGND sg13g2_fill_2
XFILLER_59_342 VPWR VGND sg13g2_fill_1
XFILLER_47_54 VPWR VGND sg13g2_fill_1
XFILLER_63_42 VPWR VGND sg13g2_decap_8
XFILLER_63_86 VPWR VGND sg13g2_fill_2
XFILLER_8_48 VPWR VGND sg13g2_fill_2
XFILLER_2_360 VPWR VGND sg13g2_fill_1
Xfanout1651 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q net1651 VPWR
+ VGND sg13g2_buf_1
Xfanout1640 _0123_ net1640 VPWR VGND sg13g2_buf_1
Xfanout1684 net1685 net1684 VPWR VGND sg13g2_buf_1
Xfanout1662 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q net1662 VPWR
+ VGND sg13g2_buf_1
XFILLER_77_150 VPWR VGND sg13g2_fill_2
Xfanout1673 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q net1673 VPWR
+ VGND sg13g2_buf_1
Xfanout1695 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q net1695 VPWR
+ VGND sg13g2_buf_1
X_5871_ net1887 net1814 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_4822_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q net1936 net51
+ net152 net1703 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q _0371_
+ VPWR VGND sg13g2_mux4_1
X_4753_ net1666 net1712 net118 net134 net94 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q
+ _0305_ VPWR VGND sg13g2_mux4_1
X_3704_ net1636 VPWR _1737_ VGND net1639 _0017_ sg13g2_o21ai_1
X_4684_ net1676 net1590 _0238_ VPWR VGND sg13g2_nor2_1
X_3635_ _1672_ net1651 _0010_ VPWR VGND sg13g2_nand2_1
X_3566_ VGND VPWR _1604_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 _1608_
+ _1607_ sg13g2_a21oi_2
X_6285_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 net506 VPWR VGND sg13g2_buf_1
X_3497_ VGND VPWR net1669 net1574 _1544_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q
+ sg13g2_a21oi_1
X_2517_ _0604_ VPWR _0605_ VGND _0075_ net1680 sg13g2_o21ai_1
X_5305_ net1999 net1729 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_5236_ net1945 net1751 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_102_258 VPWR VGND sg13g2_decap_8
XFILLER_84_19 VPWR VGND sg13g2_fill_2
X_5167_ net1997 net1775 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_5098_ net1987 net1795 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_4118_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q net21 net47
+ net32 net1596 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0
+ VPWR VGND sg13g2_mux4_1
X_4049_ _2050_ VPWR _2051_ VGND net1636 _0160_ sg13g2_o21ai_1
XFILLER_71_326 VPWR VGND sg13g2_fill_2
XFILLER_33_67 VPWR VGND sg13g2_decap_8
XFILLER_58_31 VPWR VGND sg13g2_fill_1
XFILLER_59_150 VPWR VGND sg13g2_fill_1
XFILLER_47_367 VPWR VGND sg13g2_fill_1
XFILLER_62_315 VPWR VGND sg13g2_fill_1
XFILLER_90_40 VPWR VGND sg13g2_fill_2
X_3420_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q _1470_ _1471_
+ _1469_ _0611_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X
+ VPWR VGND sg13g2_mux4_1
X_3351_ _1402_ _1396_ _1403_ VPWR VGND sg13g2_xor2_1
X_5463__595 VPWR VGND net595 sg13g2_tiehi
X_3282_ _1308_ _1333_ _1334_ VPWR VGND sg13g2_nor2_1
X_6070_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 net291 VPWR VGND sg13g2_buf_1
XFILLER_57_109 VPWR VGND sg13g2_fill_1
X_5021_ net1959 net1853 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_97_278 VPWR VGND sg13g2_decap_4
XFILLER_80_156 VPWR VGND sg13g2_fill_2
X_5854_ net1856 net1822 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_4805_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q VPWR _0355_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q _0352_ sg13g2_o21ai_1
X_2997_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q net1563 net1573
+ net1578 net1615 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q _1060_
+ VPWR VGND sg13g2_mux4_1
X_5785_ net1908 net1715 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_4736_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 _0288_ VPWR VGND sg13g2_inv_2
X_4667_ _0223_ _0222_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q
+ VPWR VGND sg13g2_nand2b_1
X_3618_ VGND VPWR _1653_ _1656_ _1657_ _0147_ sg13g2_a21oi_1
X_4598_ VPWR _0155_ _0037_ VGND sg13g2_inv_1
X_3549_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 _1591_ _1593_ _1589_
+ _1583_ VPWR VGND sg13g2_a22oi_1
X_6268_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 net480 VPWR VGND sg13g2_buf_1
X_6199_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 net411 VPWR VGND sg13g2_buf_1
X_5219_ net1971 net1751 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_44_337 VPWR VGND sg13g2_fill_1
XFILLER_44_33 VPWR VGND sg13g2_fill_2
XFILLER_44_44 VPWR VGND sg13g2_fill_2
XFILLER_52_370 VPWR VGND sg13g2_fill_1
XFILLER_114_0 VPWR VGND sg13g2_fill_2
X_5447__579 VPWR VGND net579 sg13g2_tiehi
XFILLER_94_215 VPWR VGND sg13g2_fill_2
XFILLER_47_164 VPWR VGND sg13g2_decap_4
XFILLER_85_95 VPWR VGND sg13g2_fill_2
XFILLER_62_156 VPWR VGND sg13g2_decap_8
X_2920_ VGND VPWR _0983_ _0986_ _0987_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q
+ sg13g2_a21oi_1
XFILLER_62_189 VPWR VGND sg13g2_fill_2
X_2851_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q VPWR _0923_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q _0922_ sg13g2_o21ai_1
X_2782_ VGND VPWR net128 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q
+ _0857_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q sg13g2_a21oi_1
X_5570_ net1864 net1790 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_4521_ VPWR _0078_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q VGND
+ sg13g2_inv_1
X_4452_ VGND VPWR _2368_ _1058_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q
+ sg13g2_or2_1
X_3403_ _1239_ _1293_ _1453_ _1455_ VPWR VGND sg13g2_or3_1
X_4383_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q _1277_
+ _2309_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q sg13g2_a21oi_1
X_3334_ _1386_ _1371_ _1385_ VPWR VGND sg13g2_nand2_2
X_6122_ net78 net343 VPWR VGND sg13g2_buf_1
X_3265_ VPWR _1318_ _1317_ VGND sg13g2_inv_1
X_6053_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 net274 VPWR VGND sg13g2_buf_1
X_5004_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3
+ _0544_ _0543_ sg13g2_a21oi_1
XFILLER_38_131 VPWR VGND sg13g2_fill_1
X_3196_ VPWR _1251_ _1250_ VGND sg13g2_inv_1
X_5837_ net1883 net1825 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_5768_ net1871 net1717 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_4719_ VPWR _0272_ _0271_ VGND sg13g2_inv_1
X_5699_ net1866 net1748 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_3050_ VGND VPWR _1110_ _1109_ _1108_ sg13g2_or2_1
XFILLER_35_101 VPWR VGND sg13g2_decap_8
X_3952_ _1960_ VPWR _1961_ VGND net1700 net620 sg13g2_o21ai_1
XFILLER_50_126 VPWR VGND sg13g2_fill_2
X_3883_ _1898_ _1830_ _1831_ VPWR VGND sg13g2_xnor2_1
X_2903_ _0970_ _0936_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q
+ _0971_ VPWR VGND sg13g2_mux2_1
X_2834_ net1667 net1528 net1542 net1549 net1556 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q
+ _0906_ VPWR VGND sg13g2_mux4_1
X_5622_ net1902 net1773 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_5553_ net1890 net1794 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_77_0 VPWR VGND sg13g2_fill_2
X_2765_ VGND VPWR _0077_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q
+ _0841_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q sg13g2_a21oi_1
X_4504_ VPWR _0061_ net1 VGND sg13g2_inv_1
X_5484_ net1881 net1845 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_2696_ net99 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q _0775_ VPWR
+ VGND sg13g2_nor2b_1
X_4435_ _2352_ VPWR _2353_ VGND net1713 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q
+ sg13g2_o21ai_1
X_4366_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q net1555
+ _2294_ _0167_ sg13g2_a21oi_1
X_3317_ _1369_ _1340_ _1341_ VPWR VGND sg13g2_xnor2_1
X_6105_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 net326 VPWR VGND sg13g2_buf_1
XFILLER_100_301 VPWR VGND sg13g2_decap_4
X_4297_ net1663 net1921 _2244_ VPWR VGND sg13g2_nor2b_1
X_3248_ _1301_ _1248_ _1299_ VPWR VGND sg13g2_nand2_1
X_6036_ net1779 net267 VPWR VGND sg13g2_buf_1
X_3179_ _1230_ _1229_ _1233_ _1234_ VPWR VGND sg13g2_a21o_1
XFILLER_73_229 VPWR VGND sg13g2_decap_4
Xrebuffer97 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 net706 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer75 _0565_ net684 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer86 _0288_ net695 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer110 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 net719 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_41_45 VPWR VGND sg13g2_fill_2
Xrebuffer121 net731 net730 VPWR VGND sg13g2_buf_2
Xrebuffer132 net742 net741 VPWR VGND sg13g2_buf_2
XFILLER_103_172 VPWR VGND sg13g2_fill_1
XFILLER_32_104 VPWR VGND sg13g2_decap_4
XFILLER_32_126 VPWR VGND sg13g2_fill_2
XFILLER_72_295 VPWR VGND sg13g2_fill_2
X_2550_ _0093_ VPWR _0636_ VGND _0092_ _0635_ sg13g2_o21ai_1
X_2481_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q net1712 net118
+ net94 net1922 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q _0571_
+ VPWR VGND sg13g2_mux4_1
X_4220_ VGND VPWR _2184_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 _2179_
+ _2177_ sg13g2_a21oi_2
XFILLER_95_321 VPWR VGND sg13g2_fill_1
X_4151_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q net1588 _0969_
+ _1011_ _1841_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q _2124_
+ VPWR VGND sg13g2_mux4_1
X_3102_ _1159_ _1157_ _1158_ VPWR VGND sg13g2_nand2b_1
X_4082_ net1693 net1590 _2079_ VPWR VGND sg13g2_nor2_1
X_3033_ _1092_ VPWR _1094_ VGND _1088_ _1093_ sg13g2_o21ai_1
X_4984_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q net1708 net34
+ net22 net69 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q _0525_ VPWR
+ VGND sg13g2_mux4_1
X_3935_ net1644 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X
+ _1945_ VPWR VGND sg13g2_nor2_1
X_5605_ net1874 net1781 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_3866_ _1888_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[3\] net1652 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ VPWR VGND sg13g2_mux2_2
X_3797_ _1619_ VPWR _1826_ VGND _1825_ _1824_ sg13g2_o21ai_1
X_2817_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 _0884_ _0890_ _0875_
+ _0882_ VPWR VGND sg13g2_a22oi_1
XFILLER_117_220 VPWR VGND sg13g2_fill_1
X_5536_ net1860 net1801 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_2748_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q VPWR _0825_ VGND
+ net68 net1697 sg13g2_o21ai_1
X_5467_ Tile_X0Y1_UserCLK net599 Tile_X0Y1_DSP_bot.C7 _0011_ _5467_/Q VPWR VGND sg13g2_dfrbp_1
X_4418_ _2338_ _2337_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 VPWR VGND sg13g2_mux2_1
X_2679_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q net131 _0759_
+ VPWR VGND sg13g2_nor2b_1
X_5398_ net1950 net1830 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_4349_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q net1712 net148
+ net1927 net1566 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q _2280_
+ VPWR VGND sg13g2_mux4_1
X_6019_ net1979 net231 VPWR VGND sg13g2_buf_1
XFILLER_54_240 VPWR VGND sg13g2_fill_1
XFILLER_54_262 VPWR VGND sg13g2_fill_2
XFILLER_54_273 VPWR VGND sg13g2_decap_8
XFILLER_10_354 VPWR VGND sg13g2_fill_2
XFILLER_7_0 VPWR VGND sg13g2_fill_2
Xfanout1800 Tile_X0Y1_FrameStrobe[2] net1800 VPWR VGND sg13g2_buf_1
Xfanout1811 Tile_X0Y1_FrameStrobe[1] net1811 VPWR VGND sg13g2_buf_1
Xfanout1822 net1823 net1822 VPWR VGND sg13g2_buf_1
Xfanout1833 net1835 net1833 VPWR VGND sg13g2_buf_1
XFILLER_77_41 VPWR VGND sg13g2_fill_1
XFILLER_77_52 VPWR VGND sg13g2_fill_2
XFILLER_77_332 VPWR VGND sg13g2_fill_2
Xfanout1866 net1867 net1866 VPWR VGND sg13g2_buf_1
Xfanout1855 Tile_X0Y1_FrameStrobe[0] net1855 VPWR VGND sg13g2_buf_1
Xfanout1844 Tile_X0Y1_FrameStrobe[10] net1844 VPWR VGND sg13g2_buf_1
Xfanout1888 net1889 net1888 VPWR VGND sg13g2_buf_1
Xfanout1899 Tile_X0Y1_FrameData[19] net1899 VPWR VGND sg13g2_buf_1
Xfanout1877 Tile_X0Y1_FrameData[29] net1877 VPWR VGND sg13g2_buf_1
XFILLER_93_95 VPWR VGND sg13g2_decap_4
X_3720_ _1752_ _1751_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q
+ VPWR VGND sg13g2_nand2b_1
X_3651_ _1688_ _1687_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q
+ VPWR VGND sg13g2_nand2b_1
X_3582_ _1623_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q _1622_
+ VPWR VGND sg13g2_nand2_1
X_2602_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q _0685_
+ _0686_ _0096_ sg13g2_a21oi_1
X_5321_ net1985 net1723 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_2533_ VGND VPWR _0104_ net1660 _0620_ _0619_ sg13g2_a21oi_1
X_5252_ net1974 net1741 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_4203_ _2168_ VPWR _2169_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q
+ _0868_ sg13g2_o21ai_1
X_5183_ net1964 net1766 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_4134_ _2109_ VPWR _2110_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q
+ net1523 sg13g2_o21ai_1
X_4065_ VGND VPWR _0060_ net1694 _2062_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q
+ sg13g2_a21oi_1
X_3016_ VGND VPWR net1665 net1570 _1078_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q
+ sg13g2_a21oi_1
XFILLER_51_254 VPWR VGND sg13g2_fill_2
X_4967_ VGND VPWR _0059_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q
+ _0509_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q sg13g2_a21oi_1
X_4898_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q VPWR _0444_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q _0442_ sg13g2_o21ai_1
X_3918_ _1930_ _1929_ _1900_ VPWR VGND sg13g2_xnor2_1
X_3849_ VGND VPWR _1875_ _1876_ _1868_ _1465_ sg13g2_a21oi_2
X_5519_ net1886 net1804 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput471 net471 Tile_X0Y1_S2BEGb[5] VPWR VGND sg13g2_buf_1
Xoutput460 net460 Tile_X0Y1_S2BEG[2] VPWR VGND sg13g2_buf_1
Xoutput493 net493 Tile_X0Y1_SS4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput482 net482 Tile_X0Y1_S4BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_19_207 VPWR VGND sg13g2_fill_1
XFILLER_47_88 VPWR VGND sg13g2_fill_1
XFILLER_103_50 VPWR VGND sg13g2_fill_2
XFILLER_6_122 VPWR VGND sg13g2_fill_1
XFILLER_6_199 VPWR VGND sg13g2_fill_1
XFILLER_88_40 VPWR VGND sg13g2_fill_1
XFILLER_111_237 VPWR VGND sg13g2_fill_1
Xfanout1641 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q net1641 VPWR
+ VGND sg13g2_buf_1
Xfanout1630 net1630 net1631 VPWR VGND sg13g2_buf_16
Xfanout1685 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q net1685 VPWR
+ VGND sg13g2_buf_1
Xfanout1663 net1664 net1663 VPWR VGND sg13g2_buf_1
Xfanout1652 net1653 net1652 VPWR VGND sg13g2_buf_1
Xfanout1674 net1675 net1674 VPWR VGND sg13g2_buf_1
XFILLER_65_357 VPWR VGND sg13g2_fill_1
Xfanout1696 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q net1696 VPWR
+ VGND sg13g2_buf_1
XFILLER_92_143 VPWR VGND sg13g2_fill_1
X_5870_ net1884 net1813 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_4821_ VGND VPWR _0071_ _0369_ _0370_ _0072_ sg13g2_a21oi_1
X_4752_ net1666 net1921 net41 net154 net1703 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q
+ _0304_ VPWR VGND sg13g2_mux4_1
X_5468__600 VPWR VGND net600 sg13g2_tiehi
X_3703_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q _1735_ _1736_
+ _1734_ _1733_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q Tile_X0Y1_DSP_bot.C4
+ VPWR VGND sg13g2_mux4_1
X_4683_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q _0236_ _0237_
+ VPWR VGND sg13g2_nor2_1
X_3634_ _1669_ _1670_ _1671_ VPWR VGND sg13g2_nor2b_1
X_3565_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q _1605_
+ _1608_ _0139_ sg13g2_a21oi_1
X_6284_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 net496 VPWR VGND sg13g2_buf_1
X_3496_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q
+ _1542_ _1539_ _1543_ _1540_ sg13g2_a221oi_1
X_2516_ VGND VPWR net31 net1681 _0604_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q
+ sg13g2_a21oi_1
X_5304_ net1977 net1729 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_5235_ net1943 net1751 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_5166_ net1996 net1775 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_5097_ net1986 net1798 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_4117_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q net1583 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2
+ _0699_ _0721_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3
+ VPWR VGND sg13g2_mux4_1
X_4048_ _2049_ VPWR _2050_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X
+ net1644 sg13g2_o21ai_1
XFILLER_24_243 VPWR VGND sg13g2_decap_8
X_5999_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 net211 VPWR VGND sg13g2_buf_8
Xoutput290 net290 Tile_X0Y0_N2BEGb[5] VPWR VGND sg13g2_buf_1
XFILLER_101_270 VPWR VGND sg13g2_fill_1
XFILLER_47_379 VPWR VGND sg13g2_fill_1
XFILLER_62_305 VPWR VGND sg13g2_fill_2
XFILLER_74_143 VPWR VGND sg13g2_fill_2
XFILLER_15_298 VPWR VGND sg13g2_fill_1
XFILLER_90_63 VPWR VGND sg13g2_fill_1
X_3350_ _1400_ _1399_ _1402_ VPWR VGND sg13g2_xor2_1
XFILLER_97_224 VPWR VGND sg13g2_fill_2
X_3281_ _1333_ _1309_ _1332_ VPWR VGND sg13g2_xnor2_1
X_5020_ net1957 net1853 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_38_357 VPWR VGND sg13g2_fill_2
XFILLER_65_176 VPWR VGND sg13g2_decap_8
X_5853_ net1917 net1822 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_213 VPWR VGND sg13g2_fill_2
X_5784_ net1906 net1715 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_4804_ _0353_ VPWR _0354_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q
+ net1578 sg13g2_o21ai_1
X_2996_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q net1530 net1534
+ net1543 net1556 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q _1059_
+ VPWR VGND sg13g2_mux4_1
X_4735_ VGND VPWR _0277_ _0288_ _0287_ _0282_ sg13g2_a21oi_2
X_4666_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q net1516 net2003
+ net1707 net10 net1699 _0222_ VPWR VGND sg13g2_mux4_1
X_4597_ VPWR _0154_ _0021_ VGND sg13g2_inv_1
X_3617_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q _1655_
+ _1656_ _0146_ sg13g2_a21oi_1
X_3548_ VGND VPWR _0140_ _1592_ _1593_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q
+ sg13g2_a21oi_1
X_3479_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q _1525_ _1528_
+ VPWR VGND sg13g2_nor2_1
X_6267_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 net479 VPWR VGND sg13g2_buf_1
X_6198_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 net410 VPWR VGND sg13g2_buf_1
X_5218_ net1969 net1751 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_5149_ net1960 net1776 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_176 VPWR VGND sg13g2_fill_2
XFILLER_100_73 VPWR VGND sg13g2_fill_1
XFILLER_100_95 VPWR VGND sg13g2_decap_8
XFILLER_20_290 VPWR VGND sg13g2_fill_1
XFILLER_79_202 VPWR VGND sg13g2_fill_2
XFILLER_47_176 VPWR VGND sg13g2_fill_2
X_2850_ VGND VPWR net1667 net60 _0922_ _0921_ sg13g2_a21oi_1
X_2781_ _0856_ net1527 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q
+ VPWR VGND sg13g2_nand2b_1
X_4520_ VPWR _0077_ net38 VGND sg13g2_inv_1
X_4451_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q net1542 net1549
+ net1556 net1563 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q _2367_
+ VPWR VGND sg13g2_mux4_1
X_3402_ _1453_ _1293_ _1454_ VPWR VGND sg13g2_nor2_2
X_4382_ VGND VPWR _2308_ _1058_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q
+ sg13g2_or2_1
X_6121_ net77 net342 VPWR VGND sg13g2_buf_1
X_3333_ _1385_ _1372_ _1383_ VPWR VGND sg13g2_xnor2_1
XFILLER_22_0 VPWR VGND sg13g2_fill_2
X_3264_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q VPWR _1317_ VGND
+ _1311_ _1314_ sg13g2_o21ai_1
X_6052_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 net273 VPWR VGND sg13g2_buf_1
X_5003_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q VPWR _0543_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q _0111_ sg13g2_o21ai_1
X_3195_ _1250_ _1222_ _1248_ VPWR VGND sg13g2_xnor2_1
XFILLER_41_319 VPWR VGND sg13g2_fill_1
X_5836_ net1881 net1824 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_5767_ net1919 net1725 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_2979_ _1037_ _1041_ _1042_ VPWR VGND sg13g2_nor2b_1
X_5698_ net1865 net1748 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_4718_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q net1596 net1602
+ net1621 net1629 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q _0271_
+ VPWR VGND sg13g2_mux4_1
X_4649_ _0206_ _0205_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q
+ VPWR VGND sg13g2_nand2b_1
X_6319_ Tile_X0Y1_WW4END[6] net546 VPWR VGND sg13g2_buf_1
XFILLER_76_205 VPWR VGND sg13g2_decap_8
XFILLER_103_376 VPWR VGND sg13g2_fill_1
XFILLER_29_121 VPWR VGND sg13g2_fill_1
XFILLER_55_44 VPWR VGND sg13g2_fill_1
XFILLER_25_382 VPWR VGND sg13g2_fill_2
X_3951_ VGND VPWR net1706 net1700 _1960_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q
+ sg13g2_a21oi_1
X_2902_ VGND VPWR _0968_ _0970_ _0969_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q
+ sg13g2_a21oi_2
XFILLER_31_352 VPWR VGND sg13g2_fill_2
X_3882_ _1897_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[11\] net1656 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ VPWR VGND sg13g2_mux2_1
X_2833_ VPWR _0905_ _0904_ VGND sg13g2_inv_1
XFILLER_31_363 VPWR VGND sg13g2_fill_1
X_5621_ net1900 net1773 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_5552_ net1888 net1794 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_2764_ _0839_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q _0840_
+ VPWR VGND sg13g2_nor2b_1
X_4503_ VPWR _0060_ net124 VGND sg13g2_inv_1
X_5483_ net1878 net1847 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_2695_ VGND VPWR _0773_ _0774_ net712 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q
+ sg13g2_a21oi_2
X_4434_ _2352_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q net718
+ VPWR VGND sg13g2_nand2_1
X_4365_ _2292_ _2293_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 VPWR VGND sg13g2_mux2_1
XFILLER_104_129 VPWR VGND sg13g2_fill_2
XFILLER_112_140 VPWR VGND sg13g2_fill_2
X_6104_ Tile_X0Y1_UserCLK net325 VPWR VGND sg13g2_buf_1
X_3316_ VGND VPWR _1366_ _1367_ _1368_ _1365_ sg13g2_a21oi_1
X_6035_ net1787 net266 VPWR VGND sg13g2_buf_1
X_4296_ VGND VPWR net1703 net1663 _2243_ _2242_ sg13g2_a21oi_1
XFILLER_100_324 VPWR VGND sg13g2_fill_1
X_3247_ net1511 net625 _1300_ VPWR VGND sg13g2_nor2_1
Xrebuffer10 net624 net619 VPWR VGND sg13g2_dlygate4sd1_1
X_3178_ _1232_ _1231_ _1233_ VPWR VGND sg13g2_nor2b_1
Xrebuffer76 _1433_ net685 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer87 _0288_ net696 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer98 _0460_ net707 VPWR VGND sg13g2_dlygate4sd1_1
X_5819_ net1912 net1835 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
Xrebuffer111 _0682_ net720 VPWR VGND sg13g2_buf_2
Xrebuffer122 net732 net731 VPWR VGND sg13g2_buf_2
Xrebuffer100 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X
+ net709 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer133 net743 net742 VPWR VGND sg13g2_buf_2
XFILLER_9_4 VPWR VGND sg13g2_fill_2
XFILLER_89_341 VPWR VGND sg13g2_fill_2
XFILLER_17_157 VPWR VGND sg13g2_fill_1
XFILLER_82_20 VPWR VGND sg13g2_fill_2
XFILLER_32_138 VPWR VGND sg13g2_decap_8
X_2480_ _0569_ VPWR _0570_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q
+ _0567_ sg13g2_o21ai_1
X_4150_ _2122_ _2123_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 VPWR VGND sg13g2_mux2_1
X_3101_ _1158_ _1032_ _1034_ VPWR VGND sg13g2_xnor2_1
X_4081_ _2077_ VPWR _2078_ VGND net1693 _0175_ sg13g2_o21ai_1
XFILLER_95_366 VPWR VGND sg13g2_fill_2
X_3032_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q VPWR _1093_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q _1090_ sg13g2_o21ai_1
X_4983_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q _0523_ _0524_
+ VPWR VGND sg13g2_and2_1
X_3934_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q _1937_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X _1944_
+ sg13g2_a21oi_1
X_3865_ _1888_ _1811_ _1810_ VPWR VGND sg13g2_xnor2_1
X_5604_ net1868 net1780 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_2816_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q _0889_ _0890_
+ VPWR VGND sg13g2_nor2_1
X_3796_ _1616_ _1618_ _1825_ VPWR VGND sg13g2_xor2_1
X_5535_ net1858 net1803 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_2747_ _0823_ VPWR _0824_ VGND net33 net1698 sg13g2_o21ai_1
XFILLER_117_254 VPWR VGND sg13g2_fill_1
X_5466_ Tile_X0Y1_UserCLK net598 Tile_X0Y1_DSP_bot.C6 _0013_ _5466_/Q VPWR VGND sg13g2_dfrbp_1
X_2678_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q _0580_
+ _0758_ _0757_ sg13g2_a21oi_1
X_4417_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q net1712 net148
+ net1927 net1565 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q _2338_
+ VPWR VGND sg13g2_mux4_1
X_5397_ net1948 net1830 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_4348_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q net1619 _1699_
+ _1759_ _1091_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q _2279_
+ VPWR VGND sg13g2_mux4_1
X_4279_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q net1570 net643
+ _0966_ net669 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q _2228_
+ VPWR VGND sg13g2_mux4_1
XFILLER_86_344 VPWR VGND sg13g2_fill_1
X_6018_ net1981 net230 VPWR VGND sg13g2_buf_1
XFILLER_100_165 VPWR VGND sg13g2_fill_2
XFILLER_96_108 VPWR VGND sg13g2_fill_2
Xfanout1823 net1825 net1823 VPWR VGND sg13g2_buf_1
Xfanout1812 net1813 net1812 VPWR VGND sg13g2_buf_1
Xfanout1834 net1835 net1834 VPWR VGND sg13g2_buf_1
Xfanout1801 net1803 net1801 VPWR VGND sg13g2_buf_1
Xfanout1845 net1846 net1845 VPWR VGND sg13g2_buf_1
Xfanout1867 Tile_X0Y1_FrameData[4] net1867 VPWR VGND sg13g2_buf_1
Xfanout1856 Tile_X0Y1_FrameData[9] net1856 VPWR VGND sg13g2_buf_1
Xfanout1878 Tile_X0Y1_FrameData[28] net1878 VPWR VGND sg13g2_buf_1
Xfanout1889 Tile_X0Y1_FrameData[23] net1889 VPWR VGND sg13g2_buf_1
XFILLER_92_358 VPWR VGND sg13g2_fill_1
XFILLER_60_200 VPWR VGND sg13g2_fill_1
X_3650_ _1684_ _1686_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q
+ _1687_ VPWR VGND sg13g2_nand3_1
X_3581_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q _0616_ _0723_
+ net1934 net1704 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q _1622_
+ VPWR VGND sg13g2_mux4_1
X_2601_ net147 net1705 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ _0685_ VPWR VGND sg13g2_mux2_1
Xrebuffer1 _0597_ net610 VPWR VGND sg13g2_dlygate4sd1_1
X_5320_ net1983 net1723 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_2532_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q VPWR _0619_ VGND
+ net148 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q sg13g2_o21ai_1
XFILLER_114_213 VPWR VGND sg13g2_fill_2
X_5251_ net1971 net1745 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_4202_ _2168_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q _0232_
+ VPWR VGND sg13g2_nand2_1
X_5182_ net1961 net1766 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_4133_ _2109_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q _0630_
+ VPWR VGND sg13g2_nand2_1
X_4064_ _2061_ net610 net1694 VPWR VGND sg13g2_nand2b_1
XFILLER_95_152 VPWR VGND sg13g2_fill_2
X_3015_ VGND VPWR net1665 _0178_ _1077_ _1076_ sg13g2_a21oi_1
X_4966_ net46 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q
+ _0508_ VPWR VGND sg13g2_mux2_1
X_4897_ net1677 net1594 net1588 net1523 net1540 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q
+ _0443_ VPWR VGND sg13g2_mux4_1
X_3917_ _1927_ _1928_ _1929_ VPWR VGND sg13g2_nor2b_1
X_3848_ _1869_ _1873_ _1875_ VPWR VGND sg13g2_xor2_1
X_3779_ _1808_ _1767_ _1766_ VPWR VGND sg13g2_xnor2_1
X_5518_ net1884 net1804 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput461 net461 Tile_X0Y1_S2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput450 net450 Tile_X0Y1_FrameData_O[6] VPWR VGND sg13g2_buf_1
X_5449_ Tile_X0Y1_UserCLK net581 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X
+ _5449_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[5\] VPWR VGND sg13g2_dfrbp_1
Xoutput483 net483 Tile_X0Y1_S4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput472 net472 Tile_X0Y1_S2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput494 net494 Tile_X0Y1_SS4BEG[13] VPWR VGND sg13g2_buf_8
XFILLER_63_88 VPWR VGND sg13g2_fill_1
XFILLER_111_227 VPWR VGND sg13g2_decap_4
Xfanout1620 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 net1620 VPWR VGND sg13g2_buf_8
Xfanout1642 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q net1642 VPWR
+ VGND sg13g2_buf_1
Xfanout1631 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 net1631 VPWR VGND
+ sg13g2_buf_8
Xfanout1664 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q net1664 VPWR
+ VGND sg13g2_buf_1
Xfanout1653 net1654 net1653 VPWR VGND sg13g2_buf_1
Xfanout1675 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q net1675 VPWR
+ VGND sg13g2_buf_1
Xfanout1686 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q net1686 VPWR
+ VGND sg13g2_buf_1
Xfanout1697 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q net1697 VPWR
+ VGND sg13g2_buf_1
X_4820_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q net1534 net1542
+ net1549 net1557 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q _0369_
+ VPWR VGND sg13g2_mux4_1
X_4751_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q VPWR _0303_ VGND
+ _0299_ _0302_ sg13g2_o21ai_1
X_3702_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q net1706 net106
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 net166 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q
+ _1736_ VPWR VGND sg13g2_mux4_1
X_4682_ net1676 net1597 net1610 net1624 net1632 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q
+ _0236_ VPWR VGND sg13g2_mux4_1
X_3633_ _1449_ _1450_ _1670_ VPWR VGND sg13g2_xor2_1
X_3564_ _1607_ _0138_ _1606_ VPWR VGND sg13g2_nand2_1
XFILLER_52_0 VPWR VGND sg13g2_fill_2
X_6283_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 net495 VPWR VGND sg13g2_buf_1
X_3495_ _1541_ VPWR _1542_ VGND net1669 net1545 sg13g2_o21ai_1
X_2515_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q _0602_
+ _0603_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q sg13g2_a21oi_1
X_5303_ net1956 net1731 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_5234_ net1941 net1751 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_5165_ net1993 net1775 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_4116_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q net690 net694
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 _0647_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 VPWR VGND sg13g2_mux4_1
X_5096_ net1983 net1799 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_4047_ VGND VPWR net1644 _0159_ _2049_ net1649 sg13g2_a21oi_1
XFILLER_71_328 VPWR VGND sg13g2_fill_1
XFILLER_83_177 VPWR VGND sg13g2_fill_1
XFILLER_33_25 VPWR VGND sg13g2_fill_1
XFILLER_24_288 VPWR VGND sg13g2_fill_2
X_4949_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q VPWR _0492_ VGND
+ net1695 net1522 sg13g2_o21ai_1
Xoutput280 net280 Tile_X0Y0_N2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput291 net291 Tile_X0Y0_N2BEGb[6] VPWR VGND sg13g2_buf_1
XFILLER_58_44 VPWR VGND sg13g2_fill_2
XFILLER_58_77 VPWR VGND sg13g2_fill_2
XFILLER_114_61 VPWR VGND sg13g2_fill_2
XFILLER_74_100 VPWR VGND sg13g2_fill_2
XFILLER_62_339 VPWR VGND sg13g2_fill_1
XFILLER_74_54 VPWR VGND sg13g2_decap_4
XFILLER_99_84 VPWR VGND sg13g2_fill_2
X_3280_ net1515 _1331_ _1332_ VPWR VGND sg13g2_nor2b_1
XFILLER_2_192 VPWR VGND sg13g2_fill_2
XFILLER_0_95 VPWR VGND sg13g2_fill_2
XFILLER_80_158 VPWR VGND sg13g2_fill_1
X_5852_ net1915 net1822 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_203 VPWR VGND sg13g2_fill_1
XFILLER_61_350 VPWR VGND sg13g2_fill_1
X_4803_ _0353_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q net1617
+ VPWR VGND sg13g2_nand2b_1
X_5783_ net1904 net1715 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_2995_ _1054_ VPWR _1058_ VGND _1055_ _1057_ sg13g2_o21ai_1
X_4734_ VGND VPWR _0285_ _0286_ _0287_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q
+ sg13g2_a21oi_1
X_4665_ _0220_ VPWR _0221_ VGND _0215_ _0217_ sg13g2_o21ai_1
X_4596_ VPWR _0153_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q VGND
+ sg13g2_inv_1
X_3616_ _1654_ VPWR _1655_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q
+ net1581 sg13g2_o21ai_1
X_3547_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q net1711 net1926
+ net121 net97 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q _1592_
+ VPWR VGND sg13g2_mux4_1
XFILLER_88_214 VPWR VGND sg13g2_fill_2
X_3478_ _1527_ _1526_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q
+ VPWR VGND sg13g2_nand2b_1
X_6266_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 net478 VPWR VGND sg13g2_buf_1
X_6197_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 net409 VPWR VGND sg13g2_buf_1
X_5217_ net1967 net1755 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_5148_ net1958 net1776 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_28_25 VPWR VGND sg13g2_fill_2
X_5079_ net1955 net1810 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_44_35 VPWR VGND sg13g2_fill_1
XFILLER_44_46 VPWR VGND sg13g2_fill_1
XFILLER_12_214 VPWR VGND sg13g2_fill_1
XFILLER_44_79 VPWR VGND sg13g2_fill_1
XFILLER_100_52 VPWR VGND sg13g2_fill_1
XFILLER_60_45 VPWR VGND sg13g2_fill_1
XFILLER_60_56 VPWR VGND sg13g2_decap_8
XFILLER_114_2 VPWR VGND sg13g2_fill_1
XFILLER_109_72 VPWR VGND sg13g2_decap_4
XFILLER_109_94 VPWR VGND sg13g2_fill_2
XFILLER_69_87 VPWR VGND sg13g2_decap_4
XFILLER_62_147 VPWR VGND sg13g2_decap_4
X_2780_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q _0853_
+ _0855_ _0854_ sg13g2_a21oi_1
X_4450_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q net1925 net1704
+ net1528 net1534 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q _2366_
+ VPWR VGND sg13g2_mux4_1
X_4381_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q net1544 net1550
+ net1559 net1565 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q _2307_
+ VPWR VGND sg13g2_mux4_1
X_3401_ _1345_ _1295_ _1452_ _1453_ VPWR VGND sg13g2_nor3_2
X_3332_ _1007_ net1548 _1383_ _1384_ VPWR VGND sg13g2_nor3_1
X_6120_ net76 net341 VPWR VGND sg13g2_buf_1
X_6051_ Tile_X0Y1_FrameStrobe[19] net263 VPWR VGND sg13g2_buf_1
X_3263_ VPWR _1316_ _1315_ VGND sg13g2_inv_1
X_3194_ _1249_ _1247_ _1223_ VPWR VGND sg13g2_nand2b_1
X_5002_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 _0540_ _0542_ _0529_
+ _0535_ VPWR VGND sg13g2_a22oi_1
XFILLER_15_0 VPWR VGND sg13g2_fill_2
X_5835_ net1878 net1825 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_61_180 VPWR VGND sg13g2_fill_1
X_5766_ net1896 net1725 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_2978_ _1039_ _1026_ _1041_ VPWR VGND sg13g2_xor2_1
X_5697_ net1862 net1749 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_4717_ _0269_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q _0270_
+ VPWR VGND sg13g2_nor2b_1
X_4648_ net1657 net117 net133 net1928 net93 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q
+ _0205_ VPWR VGND sg13g2_mux4_1
XFILLER_122_119 VPWR VGND sg13g2_fill_1
X_4579_ VPWR _0136_ _0003_ VGND sg13g2_inv_1
X_6318_ Tile_X0Y1_WW4END[5] net545 VPWR VGND sg13g2_buf_1
X_6249_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 net470 VPWR VGND sg13g2_buf_1
XFILLER_84_250 VPWR VGND sg13g2_fill_1
XFILLER_25_361 VPWR VGND sg13g2_fill_1
X_5453__585 VPWR VGND net585 sg13g2_tiehi
XFILLER_40_375 VPWR VGND sg13g2_fill_2
XFILLER_113_108 VPWR VGND sg13g2_decap_4
XFILLER_35_136 VPWR VGND sg13g2_fill_2
X_3950_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q _1957_
+ _1959_ _1958_ sg13g2_a21oi_1
X_2901_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3
+ net15 net41 net76 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q _0969_
+ VPWR VGND sg13g2_mux4_1
X_3881_ _1829_ _1828_ _1897_ VPWR VGND sg13g2_xor2_1
XFILLER_31_375 VPWR VGND sg13g2_fill_2
X_2832_ _0903_ VPWR _0904_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q
+ _0900_ sg13g2_o21ai_1
X_5620_ net1898 net1773 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_5551_ net1886 net1793 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_2763_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q net73 _0839_
+ VPWR VGND sg13g2_nor2_1
XFILLER_77_2 VPWR VGND sg13g2_fill_1
X_4502_ VPWR _0059_ net20 VGND sg13g2_inv_1
X_5482_ net1876 net1847 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_2694_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q VPWR _0773_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q net642 sg13g2_o21ai_1
X_4433_ _2350_ _2351_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 VPWR VGND sg13g2_mux2_1
XFILLER_116_18 VPWR VGND sg13g2_fill_1
X_4364_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q net1582 _0905_
+ _1130_ _1792_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q _2293_
+ VPWR VGND sg13g2_mux4_1
X_4295_ net1664 net152 _2242_ VPWR VGND sg13g2_nor2b_1
X_3315_ _1363_ _1364_ _1367_ VPWR VGND sg13g2_xor2_1
X_6034_ net1798 net265 VPWR VGND sg13g2_buf_1
X_3246_ net1608 net625 _1299_ VPWR VGND sg13g2_nor2_1
Xrebuffer11 _0597_ net620 VPWR VGND sg13g2_dlygate4sd1_1
X_3177_ _1232_ _1229_ _1230_ VPWR VGND sg13g2_xnor2_1
Xrebuffer33 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 net642 VPWR VGND
+ sg13g2_buf_8
Xrebuffer77 _1804_ net686 VPWR VGND sg13g2_buf_2
Xrebuffer88 _1462_ net697 VPWR VGND sg13g2_buf_1
XFILLER_81_264 VPWR VGND sg13g2_fill_1
Xrebuffer99 _0417_ net708 VPWR VGND sg13g2_dlygate4sd1_1
X_5818_ net1911 net1835 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
Xrebuffer101 _0323_ net710 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer112 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 net721 VPWR VGND sg13g2_buf_2
X_5749_ net1901 net1725 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_41_47 VPWR VGND sg13g2_fill_1
Xrebuffer123 net733 net732 VPWR VGND sg13g2_buf_2
Xrebuffer134 net744 net743 VPWR VGND sg13g2_buf_2
XFILLER_1_257 VPWR VGND sg13g2_fill_2
XFILLER_103_163 VPWR VGND sg13g2_decap_8
XFILLER_57_283 VPWR VGND sg13g2_decap_8
XFILLER_57_294 VPWR VGND sg13g2_fill_1
XFILLER_32_128 VPWR VGND sg13g2_fill_1
X_3100_ _1112_ _1111_ _1156_ _1157_ VPWR VGND sg13g2_a21o_1
X_4080_ _2077_ net1693 net1518 VPWR VGND sg13g2_nand2_1
X_3031_ _1092_ _1058_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_63_231 VPWR VGND sg13g2_decap_8
X_4982_ _0522_ VPWR _0523_ VGND net136 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q
+ sg13g2_o21ai_1
X_3933_ VGND VPWR _0121_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q
+ _1943_ _1939_ _1944_ _1942_ sg13g2_a221oi_1
XFILLER_31_150 VPWR VGND sg13g2_decap_4
X_3864_ _1887_ VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 VGND _1886_ net1652
+ sg13g2_o21ai_1
X_5603_ net1867 net1780 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_2815_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q _0886_
+ _0889_ _0888_ sg13g2_a21oi_1
XFILLER_82_0 VPWR VGND sg13g2_fill_2
X_3795_ VGND VPWR _1671_ _1824_ _1823_ _1822_ sg13g2_a21oi_2
X_5534_ net1856 net1803 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_2746_ _0823_ net1698 net49 VPWR VGND sg13g2_nand2b_1
X_5465_ Tile_X0Y1_UserCLK net597 Tile_X0Y1_DSP_bot.C5 _0015_ _5465_/Q VPWR VGND sg13g2_dfrbp_1
X_2677_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q VPWR _0757_ VGND
+ net167 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q sg13g2_o21ai_1
X_4416_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q net1618 _1699_
+ _1759_ _0805_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q _2337_
+ VPWR VGND sg13g2_mux4_1
X_5396_ net1945 net1830 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_4347_ _2273_ _2278_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A VPWR VGND sg13g2_nor2_1
X_4278_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q net1565 net613
+ _1724_ _1673_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2
+ VPWR VGND sg13g2_mux4_1
X_6017_ net1983 net229 VPWR VGND sg13g2_buf_1
X_3229_ net1640 _1280_ _1281_ _1282_ VPWR VGND sg13g2_a21o_2
XFILLER_54_220 VPWR VGND sg13g2_fill_1
XFILLER_52_68 VPWR VGND sg13g2_fill_1
XFILLER_10_356 VPWR VGND sg13g2_fill_1
XFILLER_108_211 VPWR VGND sg13g2_fill_1
Xfanout1824 net1825 net1824 VPWR VGND sg13g2_buf_1
Xfanout1802 net1803 net1802 VPWR VGND sg13g2_buf_1
Xfanout1813 net1815 net1813 VPWR VGND sg13g2_buf_1
Xfanout1846 net1847 net1846 VPWR VGND sg13g2_buf_1
Xfanout1857 Tile_X0Y1_FrameData[9] net1857 VPWR VGND sg13g2_buf_1
Xfanout1835 Tile_X0Y1_FrameStrobe[10] net1835 VPWR VGND sg13g2_buf_1
Xfanout1868 Tile_X0Y1_FrameData[3] net1868 VPWR VGND sg13g2_buf_1
Xfanout1879 Tile_X0Y1_FrameData[28] net1879 VPWR VGND sg13g2_buf_1
X_5459__591 VPWR VGND net591 sg13g2_tiehi
XFILLER_45_264 VPWR VGND sg13g2_fill_1
Xrebuffer2 net611 net667 VPWR VGND sg13g2_buf_16
XFILLER_42_90 VPWR VGND sg13g2_fill_2
X_3580_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 _0741_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q
+ _1621_ VPWR VGND sg13g2_mux2_1
X_2600_ _0683_ VPWR _0684_ VGND _0682_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ sg13g2_o21ai_1
X_2531_ VGND VPWR _0107_ _0615_ _0618_ _0617_ sg13g2_a21oi_1
X_5250_ net1969 net1745 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_4201_ _2167_ _2166_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 VPWR VGND sg13g2_mux2_1
X_5181_ net1959 net1768 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_4132_ _2107_ VPWR _2108_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q
+ _0868_ sg13g2_o21ai_1
XFILLER_3_95 VPWR VGND sg13g2_fill_1
X_4063_ _2060_ VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 VGND _2059_ net1653
+ sg13g2_o21ai_1
X_3014_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q VPWR _1076_ VGND
+ net1665 net1579 sg13g2_o21ai_1
XFILLER_51_212 VPWR VGND sg13g2_fill_2
XFILLER_51_223 VPWR VGND sg13g2_fill_2
X_4965_ _0507_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 VGND _0489_
+ _0495_ sg13g2_o21ai_1
X_3916_ VGND VPWR _1928_ _1926_ _1903_ sg13g2_or2_1
X_4896_ VPWR _0442_ _0441_ VGND sg13g2_inv_1
XFILLER_22_27 VPWR VGND sg13g2_fill_2
X_3847_ _1873_ _1869_ _1874_ VPWR VGND sg13g2_nor2b_1
X_3778_ VGND VPWR _1788_ _1807_ _1805_ _1806_ sg13g2_a21oi_2
X_2729_ _0785_ VPWR Tile_X0Y1_DSP_bot.A3 VGND _0804_ _0806_ sg13g2_o21ai_1
X_5517_ net1882 net1804 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput451 net451 Tile_X0Y1_FrameData_O[7] VPWR VGND sg13g2_buf_1
Xoutput462 net462 Tile_X0Y1_S2BEG[4] VPWR VGND sg13g2_buf_1
Xoutput440 net440 Tile_X0Y1_FrameData_O[26] VPWR VGND sg13g2_buf_1
X_5448_ Tile_X0Y1_UserCLK net580 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X
+ _5448_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[4\] VPWR VGND sg13g2_dfrbp_1
X_5379_ net1972 net1827 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput484 net484 Tile_X0Y1_S4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput473 net473 Tile_X0Y1_S2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput495 net495 Tile_X0Y1_SS4BEG[14] VPWR VGND sg13g2_buf_1
XFILLER_74_326 VPWR VGND sg13g2_fill_2
XFILLER_103_41 VPWR VGND sg13g2_fill_1
XFILLER_42_234 VPWR VGND sg13g2_decap_8
XFILLER_12_60 VPWR VGND sg13g2_fill_1
XFILLER_12_82 VPWR VGND sg13g2_fill_1
Xfanout1632 net1635 net1632 VPWR VGND sg13g2_buf_1
Xfanout1610 net1611 net1610 VPWR VGND sg13g2_buf_1
Xfanout1621 net1621 net1622 VPWR VGND sg13g2_buf_16
Xfanout1665 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q net1665 VPWR
+ VGND sg13g2_buf_1
Xfanout1643 net1646 net1643 VPWR VGND sg13g2_buf_1
Xfanout1654 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q net1654 VPWR
+ VGND sg13g2_buf_1
Xfanout1676 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q net1676 VPWR
+ VGND sg13g2_buf_1
Xfanout1687 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q net1687 VPWR
+ VGND sg13g2_buf_1
Xfanout1698 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q net1698 VPWR
+ VGND sg13g2_buf_1
XFILLER_18_297 VPWR VGND sg13g2_fill_2
X_4750_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q VPWR _0302_ VGND
+ _0300_ _0301_ sg13g2_o21ai_1
XFILLER_33_289 VPWR VGND sg13g2_fill_1
X_3701_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q net1707 net105
+ net619 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q
+ _1735_ VPWR VGND sg13g2_mux4_1
X_4681_ _0026_ net1650 _0234_ _0235_ VPWR VGND sg13g2_a21o_1
X_3632_ _1620_ VPWR _1669_ VGND _1668_ net1648 sg13g2_o21ai_1
X_3563_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q net1531 net1536
+ net1545 net1552 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q _1606_
+ VPWR VGND sg13g2_mux4_1
X_5302_ net1950 net1731 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_6282_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 net494 VPWR VGND sg13g2_buf_8
XFILLER_45_0 VPWR VGND sg13g2_fill_2
X_3494_ _1541_ net1669 net1552 VPWR VGND sg13g2_nand2b_1
X_2514_ VGND VPWR net1680 net23 _0602_ _0601_ sg13g2_a21oi_1
X_5233_ net1939 net1756 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_5164_ net1991 net1775 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_68_131 VPWR VGND sg13g2_fill_1
X_4115_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q net1630 _0614_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 _0611_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 VPWR VGND sg13g2_mux4_1
X_5095_ net1981 net1798 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_337 VPWR VGND sg13g2_fill_1
X_4046_ _2015_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X
+ VGND _2048_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q sg13g2_o21ai_1
X_5997_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 net209 VPWR VGND sg13g2_buf_1
X_4948_ _0490_ VPWR _0491_ VGND net1695 net1591 sg13g2_o21ai_1
X_4879_ net1574 net1619 net1662 _0426_ VPWR VGND sg13g2_mux2_1
Xoutput270 net270 Tile_X0Y0_FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
Xoutput292 net292 Tile_X0Y0_N2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput281 net281 Tile_X0Y0_N2BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_62_307 VPWR VGND sg13g2_fill_1
XFILLER_74_44 VPWR VGND sg13g2_fill_1
XFILLER_30_237 VPWR VGND sg13g2_decap_8
XFILLER_70_384 VPWR VGND sg13g2_fill_1
XFILLER_97_226 VPWR VGND sg13g2_fill_1
XFILLER_97_248 VPWR VGND sg13g2_decap_8
X_5851_ net1914 net1822 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_2994_ _1057_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q _1056_
+ VPWR VGND sg13g2_nand2_1
X_5782_ net1902 net1715 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_4802_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q net1569
+ _0352_ _0351_ sg13g2_a21oi_1
X_4733_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q _0283_
+ _0286_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q sg13g2_a21oi_1
X_4664_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q _0219_ _0220_
+ VPWR VGND sg13g2_and2_1
X_3615_ _1654_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q _0178_
+ VPWR VGND sg13g2_nand2_1
X_4595_ VPWR _0152_ _0013_ VGND sg13g2_inv_1
X_3546_ _1591_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q _1590_
+ VPWR VGND sg13g2_nand2_1
X_6265_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 net477 VPWR VGND sg13g2_buf_1
X_3477_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q net1516 net2003
+ net1707 net10 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q _1526_
+ VPWR VGND sg13g2_mux4_1
XFILLER_0_119 VPWR VGND sg13g2_fill_2
X_5216_ net1965 net1755 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_6196_ Tile_X0Y1_EE4END[15] net408 VPWR VGND sg13g2_buf_1
X_5147_ net1954 net1779 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_5078_ net1949 net1810 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_96_292 VPWR VGND sg13g2_fill_1
X_4029_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q net1632 net1585
+ net1591 net1520 net1679 _2033_ VPWR VGND sg13g2_mux4_1
XFILLER_52_384 VPWR VGND sg13g2_fill_1
XFILLER_121_301 VPWR VGND sg13g2_fill_1
XFILLER_69_66 VPWR VGND sg13g2_decap_8
XFILLER_79_204 VPWR VGND sg13g2_fill_1
XFILLER_79_226 VPWR VGND sg13g2_decap_8
XFILLER_116_139 VPWR VGND sg13g2_fill_1
X_4380_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q net90 net1704
+ net1529 net1535 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q _2306_
+ VPWR VGND sg13g2_mux4_1
X_3400_ VGND VPWR _1450_ _1370_ _1449_ _1342_ _1452_ _1344_ sg13g2_a221oi_1
X_3331_ _1383_ _1380_ _1382_ VPWR VGND sg13g2_xnor2_1
X_6050_ Tile_X0Y1_FrameStrobe[18] net262 VPWR VGND sg13g2_buf_1
X_3262_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q net142 net97 net44
+ net157 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q _1315_ VPWR VGND
+ sg13g2_mux4_1
X_3193_ net1511 _0808_ _1248_ VPWR VGND sg13g2_nor2_1
XFILLER_85_229 VPWR VGND sg13g2_fill_2
X_5001_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q _0541_
+ _0542_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q sg13g2_a21oi_1
X_5834_ net1876 net1824 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_14_39 VPWR VGND sg13g2_fill_2
X_5765_ net1874 net1724 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_2977_ _1038_ _1027_ _1040_ VPWR VGND sg13g2_nor2_2
X_5696_ net1860 net1749 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_4716_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q _0267_
+ _0269_ _0268_ sg13g2_a21oi_1
X_4647_ _0203_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q _0204_
+ VPWR VGND sg13g2_nor2b_1
X_6317_ Tile_X0Y1_WW4END[4] net538 VPWR VGND sg13g2_buf_1
X_4578_ VPWR _0135_ net1649 VGND sg13g2_inv_1
XFILLER_115_194 VPWR VGND sg13g2_fill_2
X_3529_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q VPWR _1575_ VGND
+ _1571_ _1574_ sg13g2_o21ai_1
XFILLER_103_301 VPWR VGND sg13g2_fill_1
X_6248_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 net469 VPWR VGND sg13g2_buf_1
X_6179_ Tile_X0Y1_E6END[8] net402 VPWR VGND sg13g2_buf_1
XFILLER_25_384 VPWR VGND sg13g2_fill_1
XFILLER_112_0 VPWR VGND sg13g2_fill_1
XFILLER_96_42 VPWR VGND sg13g2_fill_2
XFILLER_96_97 VPWR VGND sg13g2_decap_8
XFILLER_16_384 VPWR VGND sg13g2_fill_1
X_2900_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q _0967_ _0968_
+ VPWR VGND sg13g2_nor2b_1
X_3880_ _1896_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 VGND _1895_
+ net1656 sg13g2_o21ai_1
XFILLER_31_354 VPWR VGND sg13g2_fill_1
X_2831_ _0901_ _0902_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q
+ _0903_ VPWR VGND sg13g2_nand3_1
X_5550_ net1884 net1793 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_2762_ VGND VPWR _0838_ _0646_ _0115_ sg13g2_or2_1
X_5481_ net1872 net1846 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_4501_ VPWR _0058_ net167 VGND sg13g2_inv_1
X_4432_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q net1578 _0905_
+ _1130_ _1751_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q _2351_
+ VPWR VGND sg13g2_mux4_1
X_2693_ _0772_ _0519_ _0769_ VPWR VGND sg13g2_nand2_1
X_4363_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q net1710 net1925
+ _0723_ net1554 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q _2292_
+ VPWR VGND sg13g2_mux4_1
X_4294_ VGND VPWR net116 net1663 _2241_ _2240_ sg13g2_a21oi_1
X_3314_ _1358_ VPWR _1366_ VGND _1355_ _1359_ sg13g2_o21ai_1
X_6033_ net1811 net264 VPWR VGND sg13g2_buf_1
X_3245_ _1298_ _1006_ net1628 VPWR VGND sg13g2_nand2_1
XFILLER_98_376 VPWR VGND sg13g2_fill_1
X_3176_ _1225_ VPWR _1231_ VGND _1151_ _1223_ sg13g2_o21ai_1
Xrebuffer12 _0597_ net621 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer34 _0595_ net643 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer78 _0328_ net687 VPWR VGND sg13g2_buf_8
Xrebuffer89 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 net698 VPWR VGND sg13g2_buf_2
X_5817_ net1909 net1837 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
Xrebuffer113 _0230_ net722 VPWR VGND sg13g2_dlygate4sd1_1
X_5748_ net1899 net1725 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
Xrebuffer102 _2053_ net711 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer135 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 net744 VPWR VGND
+ sg13g2_buf_2
Xrebuffer124 net734 net733 VPWR VGND sg13g2_buf_2
X_5679_ net1886 net1748 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_89_310 VPWR VGND sg13g2_fill_1
X_3030_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q net139 net1935
+ net93 net153 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q _1091_
+ VPWR VGND sg13g2_mux4_1
Xinput170 Tile_X0Y1_WW4END[1] net170 VPWR VGND sg13g2_buf_1
XFILLER_95_368 VPWR VGND sg13g2_fill_1
X_4981_ VGND VPWR _0075_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q
+ _0522_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q sg13g2_a21oi_1
X_3932_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q net16 net77 net42
+ net618 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q _1943_ VPWR
+ VGND sg13g2_mux4_1
X_3863_ _1887_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[4\] net1653 VPWR VGND sg13g2_nand2_1
X_5602_ net1865 net1780 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_2814_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q VPWR _0888_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q _0887_ sg13g2_o21ai_1
X_5533_ net1917 net1803 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_3794_ _1823_ _1669_ _1670_ VPWR VGND sg13g2_xnor2_1
X_2745_ _0822_ _0818_ _0821_ VPWR VGND sg13g2_nand2_1
XFILLER_117_278 VPWR VGND sg13g2_fill_1
X_5464_ Tile_X0Y1_UserCLK net596 Tile_X0Y1_DSP_bot.C4 _0017_ _5464_/Q VPWR VGND sg13g2_dfrbp_1
X_2676_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q _0290_
+ _0756_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q sg13g2_a21oi_1
X_4415_ _2331_ _2336_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 VPWR VGND
+ sg13g2_nor2_1
X_5395_ net1944 net1831 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_4346_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q _2274_
+ _2278_ _2277_ sg13g2_a21oi_1
XFILLER_98_162 VPWR VGND sg13g2_fill_1
X_4277_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q net1559 net689
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 _0362_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 VPWR VGND sg13g2_mux4_1
XFILLER_98_184 VPWR VGND sg13g2_fill_2
X_6016_ net1985 net228 VPWR VGND sg13g2_buf_1
X_3228_ net1640 Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[1\] _1281_ VPWR VGND sg13g2_nor2_1
X_3159_ _1214_ _1213_ VPWR VGND sg13g2_inv_8
XFILLER_54_287 VPWR VGND sg13g2_decap_4
Xfanout1825 net1826 net1825 VPWR VGND sg13g2_buf_1
Xfanout1803 net1811 net1803 VPWR VGND sg13g2_buf_1
Xfanout1814 net1815 net1814 VPWR VGND sg13g2_buf_1
Xfanout1847 net1848 net1847 VPWR VGND sg13g2_buf_1
Xfanout1836 net1838 net1836 VPWR VGND sg13g2_buf_1
Xfanout1858 net1859 net1858 VPWR VGND sg13g2_buf_1
Xfanout1869 Tile_X0Y1_FrameData[3] net1869 VPWR VGND sg13g2_buf_1
Xrebuffer3 net611 net612 VPWR VGND sg13g2_dlygate4sd1_1
X_2530_ net1660 _0099_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q
+ _0617_ VPWR VGND sg13g2_a21o_1
XFILLER_114_215 VPWR VGND sg13g2_fill_1
XFILLER_114_204 VPWR VGND sg13g2_fill_1
X_4200_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2
+ net2003 net1932 net1602 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q
+ _2167_ VPWR VGND sg13g2_mux4_1
X_5180_ net1957 net1768 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_95_121 VPWR VGND sg13g2_fill_2
X_4131_ _2107_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q _1499_
+ VPWR VGND sg13g2_nand2_1
X_4062_ _2060_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[8\] net1653 VPWR VGND sg13g2_nand2_1
X_3013_ VGND VPWR _1074_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q
+ _1073_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q _1075_ _1072_
+ sg13g2_a221oi_1
X_4964_ _0501_ _0506_ _0507_ VPWR VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q
+ sg13g2_nand3b_1
X_3915_ _1903_ _1926_ _1927_ VPWR VGND sg13g2_and2_1
X_4895_ net1677 net1599 net1612 net1605 net1625 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q
+ _0441_ VPWR VGND sg13g2_mux4_1
X_3846_ _1872_ _1871_ _1873_ VPWR VGND sg13g2_xor2_1
X_3777_ _1785_ _1787_ _1806_ VPWR VGND sg13g2_xor2_1
X_2728_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q VPWR _0806_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q _0805_ sg13g2_o21ai_1
X_5516_ net1881 net1804 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_5447_ Tile_X0Y1_UserCLK net579 Tile_X0Y1_DSP_bot.A3 _5447_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[3\]
+ VPWR VGND sg13g2_dfrbp_1
Xoutput452 net452 Tile_X0Y1_FrameData_O[8] VPWR VGND sg13g2_buf_1
Xoutput430 net430 Tile_X0Y1_FrameData_O[17] VPWR VGND sg13g2_buf_1
Xoutput441 net441 Tile_X0Y1_FrameData_O[27] VPWR VGND sg13g2_buf_1
X_2659_ _0740_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q _0734_
+ _0739_ VPWR VGND sg13g2_and3_1
X_5378_ net1969 net1829 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput496 net496 Tile_X0Y1_SS4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput485 net485 Tile_X0Y1_S4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput474 net474 Tile_X0Y1_S4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput463 net463 Tile_X0Y1_S2BEG[5] VPWR VGND sg13g2_buf_1
X_4329_ _1714_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q _2263_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_103_20 VPWR VGND sg13g2_fill_2
XFILLER_63_24 VPWR VGND sg13g2_fill_1
XFILLER_27_298 VPWR VGND sg13g2_fill_2
XFILLER_63_35 VPWR VGND sg13g2_decap_8
Xfanout1622 net1622 net1627 VPWR VGND sg13g2_buf_16
Xfanout1611 net1614 net1611 VPWR VGND sg13g2_buf_1
Xfanout1600 net1601 net1600 VPWR VGND sg13g2_buf_1
Xfanout1633 net1635 net1633 VPWR VGND sg13g2_buf_1
Xfanout1666 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q net1666 VPWR
+ VGND sg13g2_buf_1
Xfanout1655 net1656 net1655 VPWR VGND sg13g2_buf_1
Xfanout1644 net1645 net1644 VPWR VGND sg13g2_buf_1
Xfanout1677 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q net1677 VPWR
+ VGND sg13g2_buf_1
Xfanout1699 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q net1699 VPWR
+ VGND sg13g2_buf_1
XFILLER_19_8 VPWR VGND sg13g2_fill_1
XFILLER_65_338 VPWR VGND sg13g2_fill_2
Xfanout1688 net1689 net1688 VPWR VGND sg13g2_buf_1
XFILLER_33_202 VPWR VGND sg13g2_decap_8
XFILLER_73_382 VPWR VGND sg13g2_fill_2
X_3700_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q net122 net98
+ net1934 net169 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q _1734_
+ VPWR VGND sg13g2_mux4_1
X_4680_ VGND VPWR net1638 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X
+ _0234_ _0233_ sg13g2_a21oi_1
X_3631_ VGND VPWR _1667_ _1668_ _0009_ net1646 sg13g2_a21oi_2
X_3562_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q net1558 net1574
+ net1582 net1616 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q _1605_
+ VPWR VGND sg13g2_mux4_1
XFILLER_52_2 VPWR VGND sg13g2_fill_1
X_2513_ net1680 net136 _0601_ VPWR VGND sg13g2_nor2b_1
X_5301_ net1948 net1731 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_6281_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 net493 VPWR VGND sg13g2_buf_1
X_3493_ VGND VPWR net1670 net1536 _1540_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q
+ sg13g2_a21oi_1
X_5232_ net1937 net1756 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_5163_ net1989 net1775 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_38_0 VPWR VGND sg13g2_decap_8
X_4114_ _2093_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q
+ _2102_ sg13g2_o21ai_1
X_5094_ net1979 net1798 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_4045_ _2030_ VPWR _2048_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q
+ _2047_ sg13g2_o21ai_1
X_5475__607 VPWR VGND net607 sg13g2_tiehi
X_5996_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 net208 VPWR VGND sg13g2_buf_1
X_4947_ _0490_ net1695 net1587 VPWR VGND sg13g2_nand2b_1
X_4878_ _0171_ net1561 net1662 _0425_ VPWR VGND sg13g2_mux2_1
X_3829_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q _1857_
+ _1858_ _0118_ sg13g2_a21oi_1
XFILLER_118_373 VPWR VGND sg13g2_fill_1
Xoutput271 net271 Tile_X0Y0_FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
Xoutput260 net260 Tile_X0Y0_FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
Xoutput293 net293 Tile_X0Y0_N4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput282 net282 Tile_X0Y0_N2BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_59_143 VPWR VGND sg13g2_decap_8
XFILLER_59_154 VPWR VGND sg13g2_fill_2
XFILLER_74_102 VPWR VGND sg13g2_fill_1
XFILLER_55_371 VPWR VGND sg13g2_fill_1
XFILLER_109_384 VPWR VGND sg13g2_fill_1
XFILLER_65_102 VPWR VGND sg13g2_decap_8
XFILLER_65_135 VPWR VGND sg13g2_fill_2
XFILLER_0_97 VPWR VGND sg13g2_fill_1
X_5850_ net1911 net1824 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_5781_ net1900 net1714 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_2993_ _1056_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q net162
+ VPWR VGND sg13g2_nand2_1
X_4801_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q net1563 _0351_
+ VPWR VGND sg13g2_nor2_1
X_4732_ _0285_ _0284_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q
+ VPWR VGND sg13g2_nand2b_1
X_4663_ _0219_ _0218_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q
+ VPWR VGND sg13g2_nand2b_1
X_3614_ _1652_ VPWR _1653_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q
+ net1555 sg13g2_o21ai_1
X_4594_ VPWR _0151_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q VGND
+ sg13g2_inv_1
X_3545_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q _0682_ net44
+ net147 net1705 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q _1590_
+ VPWR VGND sg13g2_mux4_1
X_3476_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q _1523_
+ _1525_ _1524_ sg13g2_a21oi_1
X_6264_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 net476 VPWR VGND sg13g2_buf_1
X_5215_ net1963 net1754 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_6195_ Tile_X0Y1_EE4END[14] net407 VPWR VGND sg13g2_buf_1
X_5146_ net1952 net1779 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_28_27 VPWR VGND sg13g2_fill_1
XFILLER_56_135 VPWR VGND sg13g2_fill_1
XFILLER_56_146 VPWR VGND sg13g2_fill_1
X_5077_ net1948 net1806 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_4028_ VPWR _2032_ _2031_ VGND sg13g2_inv_1
X_5979_ Tile_X0Y0_E6END[9] net202 VPWR VGND sg13g2_buf_1
XFILLER_109_63 VPWR VGND sg13g2_decap_4
XFILLER_43_363 VPWR VGND sg13g2_fill_1
XFILLER_70_182 VPWR VGND sg13g2_decap_8
X_3330_ VPWR _1382_ _1381_ VGND sg13g2_inv_1
XFILLER_112_324 VPWR VGND sg13g2_fill_2
X_3261_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q VPWR _1314_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q _1313_ sg13g2_o21ai_1
X_5000_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q net34 net69 net46
+ net85 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q _0541_ VPWR VGND
+ sg13g2_mux4_1
X_3192_ net1608 _0808_ _1247_ VPWR VGND sg13g2_nor2_2
XFILLER_15_2 VPWR VGND sg13g2_fill_1
XFILLER_38_179 VPWR VGND sg13g2_fill_1
XFILLER_19_382 VPWR VGND sg13g2_fill_2
X_5833_ net1872 net1826 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_5764_ net1868 net1724 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_2976_ _1039_ _0899_ _1023_ VPWR VGND sg13g2_nand2_1
X_5695_ net1859 net1750 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_4715_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q VPWR _0268_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q _0266_ sg13g2_o21ai_1
X_4646_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q _0201_
+ _0203_ _0202_ sg13g2_a21oi_1
X_4577_ VPWR _0134_ net1644 VGND sg13g2_inv_1
X_6316_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 net528 VPWR VGND sg13g2_buf_1
X_3528_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q VPWR _1574_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q _1573_ sg13g2_o21ai_1
X_6247_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 net468 VPWR VGND sg13g2_buf_1
X_3459_ _1295_ VPWR _1508_ VGND _1345_ _1452_ sg13g2_o21ai_1
X_6178_ Tile_X0Y1_E6END[7] net401 VPWR VGND sg13g2_buf_1
X_5129_ net1985 net1787 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_84_230 VPWR VGND sg13g2_fill_1
XFILLER_35_138 VPWR VGND sg13g2_fill_1
XFILLER_16_341 VPWR VGND sg13g2_fill_1
XFILLER_31_300 VPWR VGND sg13g2_fill_1
X_2830_ _0902_ net163 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_43_171 VPWR VGND sg13g2_decap_8
X_2761_ _0836_ _0834_ _0837_ VPWR VGND sg13g2_nor2_2
X_5480_ net1870 net1846 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_2692_ net1515 net1608 _0771_ VPWR VGND sg13g2_nor2_1
X_4500_ net1513 net711 _0057_ VPWR VGND sg13g2_nor2_1
X_4431_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q net1710 net1704
+ _0723_ net1551 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q _2350_
+ VPWR VGND sg13g2_mux4_1
X_4362_ _2285_ _2291_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 VPWR VGND
+ sg13g2_nor2_1
XFILLER_112_110 VPWR VGND sg13g2_fill_2
X_4293_ net1663 net1710 _2240_ VPWR VGND sg13g2_nor2b_1
X_3313_ _1363_ _1364_ _1365_ VPWR VGND sg13g2_nor2_1
X_6101_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 net313 VPWR VGND sg13g2_buf_2
X_3244_ _1243_ _1296_ _1297_ VPWR VGND sg13g2_nor2_1
X_6032_ net1854 net253 VPWR VGND sg13g2_buf_1
XFILLER_100_305 VPWR VGND sg13g2_fill_2
X_3175_ _1230_ _1113_ _1155_ VPWR VGND sg13g2_xnor2_1
Xrebuffer13 _0597_ net622 VPWR VGND sg13g2_buf_8
Xrebuffer24 _0680_ net633 VPWR VGND sg13g2_buf_8
Xrebuffer35 _1804_ net644 VPWR VGND sg13g2_buf_2
Xrebuffer79 net687 net688 VPWR VGND sg13g2_buf_8
XFILLER_81_244 VPWR VGND sg13g2_fill_2
X_5816_ net1907 net1837 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
Xrebuffer103 _0324_ net712 VPWR VGND sg13g2_buf_8
X_5747_ net1894 net1727 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_2959_ _1022_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X
+ VGND _1014_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q sg13g2_o21ai_1
Xrebuffer114 net730 net723 VPWR VGND sg13g2_buf_2
Xrebuffer125 net735 net734 VPWR VGND sg13g2_buf_2
X_5678_ net1885 net1748 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_4629_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q _0185_ _0186_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_1_259 VPWR VGND sg13g2_fill_1
XFILLER_106_20 VPWR VGND sg13g2_fill_1
XFILLER_103_198 VPWR VGND sg13g2_decap_8
XFILLER_32_108 VPWR VGND sg13g2_fill_2
XFILLER_72_288 VPWR VGND sg13g2_fill_2
XFILLER_95_347 VPWR VGND sg13g2_fill_1
Xinput160 Tile_X0Y1_W2MID[1] net160 VPWR VGND sg13g2_buf_1
Xinput171 Tile_X0Y1_WW4END[2] net171 VPWR VGND sg13g2_buf_1
X_4980_ net695 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q _0520_
+ _0521_ VPWR VGND sg13g2_a21o_1
X_3931_ _0121_ _1941_ _1942_ VPWR VGND sg13g2_nor2_1
X_3862_ _1886_ _1813_ _1814_ VPWR VGND sg13g2_xnor2_1
X_5601_ net1863 net1780 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_2813_ net33 net49 net1689 _0887_ VPWR VGND sg13g2_mux2_1
XFILLER_82_2 VPWR VGND sg13g2_fill_1
X_5532_ net1915 net1803 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_3793_ _1694_ VPWR _1822_ VGND _1821_ _1820_ sg13g2_o21ai_1
XFILLER_11_19 VPWR VGND sg13g2_fill_2
X_2744_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q _0820_ _0821_
+ VPWR VGND sg13g2_nor2_1
XFILLER_117_246 VPWR VGND sg13g2_fill_2
X_5463_ Tile_X0Y1_UserCLK net595 Tile_X0Y1_DSP_bot.C3 _0019_ _5463_/Q VPWR VGND sg13g2_dfrbp_1
X_2675_ _0754_ VPWR _0755_ VGND _0742_ _0743_ sg13g2_o21ai_1
X_4414_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q _2334_
+ _2336_ _2335_ sg13g2_a21oi_1
X_5394_ net1941 net1831 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_4345_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q VPWR _2277_
+ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q _2276_ sg13g2_o21ai_1
XFILLER_98_130 VPWR VGND sg13g2_fill_2
X_4276_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q net1551 net693
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 _0308_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 VPWR VGND sg13g2_mux4_1
X_5443__575 VPWR VGND net575 sg13g2_tiehi
XFILLER_100_102 VPWR VGND sg13g2_decap_4
X_6015_ net1988 net227 VPWR VGND sg13g2_buf_1
X_3227_ VPWR Tile_X0Y1_DSP_bot.B1 _1280_ VGND sg13g2_inv_1
XFILLER_86_358 VPWR VGND sg13g2_fill_1
X_3158_ Tile_X0Y1_DSP_bot.A0 Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[0\] net1641 _1213_
+ VPWR VGND sg13g2_mux2_2
XFILLER_94_380 VPWR VGND sg13g2_fill_1
X_3089_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q net119 net95
+ net60 net155 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q _1147_
+ VPWR VGND sg13g2_mux4_1
XFILLER_54_255 VPWR VGND sg13g2_decap_8
XFILLER_54_299 VPWR VGND sg13g2_fill_1
XFILLER_10_325 VPWR VGND sg13g2_fill_2
XFILLER_10_303 VPWR VGND sg13g2_fill_1
XFILLER_123_227 VPWR VGND sg13g2_fill_2
XFILLER_117_85 VPWR VGND sg13g2_fill_1
Xfanout1815 net1816 net1815 VPWR VGND sg13g2_buf_1
Xfanout1804 net1805 net1804 VPWR VGND sg13g2_buf_1
Xfanout1837 net1838 net1837 VPWR VGND sg13g2_buf_1
Xfanout1848 net1850 net1848 VPWR VGND sg13g2_buf_1
Xfanout1826 net1832 net1826 VPWR VGND sg13g2_buf_1
Xfanout1859 Tile_X0Y1_FrameData[8] net1859 VPWR VGND sg13g2_buf_1
XFILLER_92_339 VPWR VGND sg13g2_fill_1
XFILLER_93_44 VPWR VGND sg13g2_fill_1
XFILLER_93_99 VPWR VGND sg13g2_fill_2
XFILLER_45_299 VPWR VGND sg13g2_fill_2
XFILLER_9_134 VPWR VGND sg13g2_fill_2
Xrebuffer4 net611 net613 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_107_290 VPWR VGND sg13g2_decap_4
X_4130_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q _2105_ _2106_
+ VPWR VGND sg13g2_nor2_1
X_4061_ _2059_ _1822_ _1823_ VPWR VGND sg13g2_xnor2_1
X_3012_ VGND VPWR net1665 _0176_ _1074_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q
+ sg13g2_a21oi_1
XFILLER_91_372 VPWR VGND sg13g2_fill_2
XFILLER_36_299 VPWR VGND sg13g2_fill_2
X_4963_ _0503_ _0505_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q
+ _0506_ VPWR VGND sg13g2_nand3_1
XFILLER_51_247 VPWR VGND sg13g2_decap_8
X_3914_ _1904_ VPWR _1926_ VGND net1649 _1925_ sg13g2_o21ai_1
X_4894_ _0437_ _0439_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q
+ _0440_ VPWR VGND sg13g2_nand3_1
X_3845_ _1461_ VPWR _1872_ VGND _1462_ _1171_ sg13g2_o21ai_1
X_3776_ net686 _1434_ _1805_ VPWR VGND sg13g2_nor2_2
X_2727_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q net115 net38 net91
+ net172 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q _0805_ VPWR VGND
+ sg13g2_mux4_1
X_5515_ net1879 net1804 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput420 net420 Tile_X0Y1_EE4BEG[8] VPWR VGND sg13g2_buf_1
X_5446_ Tile_X0Y1_UserCLK net578 Tile_X0Y1_DSP_bot.A2 _5446_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[2\]
+ VPWR VGND sg13g2_dfrbp_1
Xoutput453 net453 Tile_X0Y1_FrameData_O[9] VPWR VGND sg13g2_buf_1
Xoutput442 net442 Tile_X0Y1_FrameData_O[28] VPWR VGND sg13g2_buf_1
Xoutput431 net431 Tile_X0Y1_FrameData_O[18] VPWR VGND sg13g2_buf_1
X_2658_ _0738_ VPWR _0739_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q
+ _0736_ sg13g2_o21ai_1
X_5377_ net1968 net1829 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_2589_ VGND VPWR _0066_ net1658 _0674_ _0673_ sg13g2_a21oi_1
Xoutput486 net486 Tile_X0Y1_S4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput464 net464 Tile_X0Y1_S2BEG[6] VPWR VGND sg13g2_buf_1
Xoutput475 net475 Tile_X0Y1_S4BEG[10] VPWR VGND sg13g2_buf_1
X_4328_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q _1058_
+ _2262_ _2261_ sg13g2_a21oi_1
Xoutput497 net497 Tile_X0Y1_SS4BEG[1] VPWR VGND sg13g2_buf_1
X_4259_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q net2003 net1597
+ net64 net1610 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q _2217_
+ VPWR VGND sg13g2_mux4_1
XFILLER_12_40 VPWR VGND sg13g2_fill_2
Xfanout1601 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 net1601 VPWR VGND
+ sg13g2_buf_8
Xfanout1623 net1627 net1623 VPWR VGND sg13g2_buf_1
Xfanout1612 net1613 net1612 VPWR VGND sg13g2_buf_1
Xfanout1634 net1635 net1634 VPWR VGND sg13g2_buf_1
Xfanout1667 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q net1667 VPWR
+ VGND sg13g2_buf_1
Xfanout1656 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q net1656 VPWR
+ VGND sg13g2_buf_1
Xfanout1645 net1646 net1645 VPWR VGND sg13g2_buf_1
Xfanout1678 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q net1678 VPWR
+ VGND sg13g2_buf_1
XFILLER_65_306 VPWR VGND sg13g2_fill_2
Xfanout1689 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q net1689 VPWR
+ VGND sg13g2_buf_1
XFILLER_18_233 VPWR VGND sg13g2_fill_2
XFILLER_58_380 VPWR VGND sg13g2_fill_1
XFILLER_33_247 VPWR VGND sg13g2_fill_2
XFILLER_53_80 VPWR VGND sg13g2_fill_2
X_3630_ net1643 Tile_X0Y1_DSP_bot.C8 _1667_ VPWR VGND sg13g2_nor2_2
X_3561_ VGND VPWR _0138_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q
+ _1603_ _1599_ _1604_ _1602_ sg13g2_a221oi_1
X_2512_ _0599_ VPWR _0600_ VGND net1680 net610 sg13g2_o21ai_1
X_5300_ net1946 net1731 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_3492_ _1539_ net1531 net1669 VPWR VGND sg13g2_nand2b_1
X_6280_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 net492 VPWR VGND sg13g2_buf_8
XFILLER_45_2 VPWR VGND sg13g2_fill_1
X_5231_ net1998 net1754 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_5162_ net1987 net1775 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_5093_ net1975 net1799 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_4113_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q _2101_ _2099_
+ _2095_ _2097_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q _2102_
+ VPWR VGND sg13g2_mux4_1
X_4044_ net729 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q
+ _2047_ VPWR VGND sg13g2_mux2_1
X_5995_ Tile_X0Y0_EE4END[15] net207 VPWR VGND sg13g2_buf_1
X_4946_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q _0488_ _0489_
+ VPWR VGND sg13g2_nor2_1
X_4877_ VGND VPWR _0423_ _0424_ _0419_ _0421_ sg13g2_a21oi_2
X_3828_ _1856_ VPWR _1857_ VGND net1933 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q
+ sg13g2_o21ai_1
X_3759_ _1789_ net1647 net745 VPWR VGND sg13g2_nand2_1
X_5449__581 VPWR VGND net581 sg13g2_tiehi
Xoutput250 net250 Tile_X0Y0_FrameData_O[7] VPWR VGND sg13g2_buf_1
Xoutput261 net261 Tile_X0Y0_FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
X_5429_ Tile_X0Y1_UserCLK net569 _0043_ _0014_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[5\]
+ VPWR VGND sg13g2_dfrbp_1
Xoutput272 net272 Tile_X0Y0_FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
Xoutput294 net294 Tile_X0Y0_N4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput283 net283 Tile_X0Y0_N2BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_47_317 VPWR VGND sg13g2_fill_1
XFILLER_59_188 VPWR VGND sg13g2_decap_4
XFILLER_23_83 VPWR VGND sg13g2_fill_1
XFILLER_2_162 VPWR VGND sg13g2_fill_2
XFILLER_97_217 VPWR VGND sg13g2_decap_8
XFILLER_38_317 VPWR VGND sg13g2_fill_1
XFILLER_38_328 VPWR VGND sg13g2_fill_2
XFILLER_65_169 VPWR VGND sg13g2_decap_8
X_4800_ _0350_ _0349_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q
+ VPWR VGND sg13g2_nand2b_1
X_2992_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q net638 _1055_
+ VPWR VGND sg13g2_nor2b_1
X_5780_ net1898 net1714 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_4731_ net145 net1 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q _0284_
+ VPWR VGND sg13g2_mux2_1
X_4662_ net1699 net1597 net1610 net1603 net1623 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q
+ _0218_ VPWR VGND sg13g2_mux4_1
X_3613_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q net1564
+ _1652_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q sg13g2_a21oi_1
X_4593_ VPWR _0150_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q VGND
+ sg13g2_inv_1
X_6332_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 net544 VPWR VGND sg13g2_buf_1
X_3544_ VGND VPWR _1585_ _1588_ _1589_ _0141_ sg13g2_a21oi_1
XFILLER_50_0 VPWR VGND sg13g2_decap_8
X_3475_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q VPWR _1524_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q _1521_ sg13g2_o21ai_1
X_6263_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 net475 VPWR VGND sg13g2_buf_1
X_5214_ net1962 net1754 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_6194_ Tile_X0Y1_EE4END[13] net421 VPWR VGND sg13g2_buf_1
X_5145_ net1999 net1789 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_5076_ net1946 net1806 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_4027_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q net1597 net1610
+ net1603 net1624 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q _2031_
+ VPWR VGND sg13g2_mux4_1
XFILLER_37_361 VPWR VGND sg13g2_fill_1
XFILLER_37_383 VPWR VGND sg13g2_fill_2
X_5978_ Tile_X0Y0_E6END[8] net201 VPWR VGND sg13g2_buf_1
X_4929_ _0472_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q _0473_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_18_72 VPWR VGND sg13g2_fill_2
XFILLER_55_191 VPWR VGND sg13g2_fill_2
X_3260_ VGND VPWR net61 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q
+ _1313_ _1312_ sg13g2_a21oi_1
X_3191_ _1246_ _1023_ net1628 VPWR VGND sg13g2_nand2_1
XFILLER_78_261 VPWR VGND sg13g2_fill_1
XFILLER_53_106 VPWR VGND sg13g2_decap_8
X_5832_ net1870 net1826 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_5763_ net1867 net1728 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_61_172 VPWR VGND sg13g2_decap_4
X_2975_ _1038_ _0849_ _1023_ VPWR VGND sg13g2_nand2_1
X_4714_ net1521 net1518 net1683 _0267_ VPWR VGND sg13g2_mux2_1
X_5694_ net1857 net1750 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_4645_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q VPWR _0202_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q _0199_ sg13g2_o21ai_1
X_4576_ VPWR _0133_ _0001_ VGND sg13g2_inv_1
X_6315_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 net527 VPWR VGND sg13g2_buf_1
X_3527_ VGND VPWR net1671 net1561 _1573_ _1572_ sg13g2_a21oi_1
XFILLER_115_163 VPWR VGND sg13g2_fill_2
X_6246_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 net467 VPWR VGND sg13g2_buf_1
X_3458_ _1507_ _1506_ _1504_ VPWR VGND sg13g2_nand2_2
X_6177_ Tile_X0Y1_E6END[6] net400 VPWR VGND sg13g2_buf_1
X_3389_ _1441_ _1439_ _1440_ VPWR VGND sg13g2_nand2b_1
X_5128_ net1984 net1787 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_17_309 VPWR VGND sg13g2_fill_1
X_5059_ net1972 net1808 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_52_194 VPWR VGND sg13g2_decap_4
XFILLER_4_257 VPWR VGND sg13g2_fill_2
XFILLER_106_141 VPWR VGND sg13g2_fill_1
XFILLER_90_267 VPWR VGND sg13g2_decap_4
X_2760_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q VPWR _0836_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q _0835_ sg13g2_o21ai_1
X_2691_ _0462_ _0703_ _0770_ VPWR VGND sg13g2_nor2_1
X_4430_ VGND VPWR _2340_ _2343_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0
+ _2349_ sg13g2_a21oi_1
X_6100_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 net312 VPWR VGND sg13g2_buf_1
X_4361_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q _2289_
+ _2291_ _2290_ sg13g2_a21oi_1
X_4292_ VGND VPWR net108 net1664 _2239_ _2238_ sg13g2_a21oi_1
X_3312_ _1364_ _1335_ _1336_ VPWR VGND sg13g2_xnor2_1
X_6031_ net1952 net245 VPWR VGND sg13g2_buf_1
X_3243_ _1296_ _1213_ _0899_ _1103_ net1575 VPWR VGND sg13g2_a22oi_1
XFILLER_112_188 VPWR VGND sg13g2_fill_1
XFILLER_13_0 VPWR VGND sg13g2_fill_1
X_3174_ _1220_ _1219_ _1228_ _1229_ VPWR VGND sg13g2_a21o_1
Xrebuffer36 _0615_ net645 VPWR VGND sg13g2_buf_2
XFILLER_66_297 VPWR VGND sg13g2_fill_2
Xrebuffer25 net633 net634 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer14 _1943_ net623 VPWR VGND sg13g2_buf_8
Xrebuffer58 net728 net667 VPWR VGND sg13g2_buf_8
X_5815_ net1905 net1837 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
Xrebuffer104 _0323_ net713 VPWR VGND sg13g2_buf_2
X_5746_ net1892 net1727 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_2958_ _1022_ _1019_ _1021_ VPWR VGND sg13g2_nand2b_1
X_5677_ net1882 net1746 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
Xrebuffer115 net723 net724 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer126 net736 net735 VPWR VGND sg13g2_buf_2
X_2889_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q _0957_ _0958_
+ VPWR VGND sg13g2_nor2b_1
X_4628_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q net1516 net8
+ net1708 net20 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q _0185_
+ VPWR VGND sg13g2_mux4_1
X_4559_ VPWR _0116_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q VGND
+ sg13g2_inv_1
X_6229_ net1879 net442 VPWR VGND sg13g2_buf_1
XFILLER_103_144 VPWR VGND sg13g2_fill_2
XFILLER_40_186 VPWR VGND sg13g2_fill_2
XFILLER_31_72 VPWR VGND sg13g2_decap_4
XFILLER_0_260 VPWR VGND sg13g2_fill_1
Xinput150 Tile_X0Y1_W1END[3] net150 VPWR VGND sg13g2_buf_1
Xinput161 Tile_X0Y1_W2MID[2] net161 VPWR VGND sg13g2_buf_1
Xinput172 Tile_X0Y1_WW4END[3] net172 VPWR VGND sg13g2_buf_1
XFILLER_63_245 VPWR VGND sg13g2_fill_2
X_3930_ VGND VPWR net78 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q
+ _1941_ _1940_ sg13g2_a21oi_1
XFILLER_63_289 VPWR VGND sg13g2_fill_1
X_3861_ _1885_ VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 VGND net1652 _1884_
+ sg13g2_o21ai_1
X_5600_ net1861 net1780 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_3792_ _1692_ _1693_ _1821_ VPWR VGND sg13g2_xor2_1
X_2812_ _0885_ VPWR _0886_ VGND net68 net1689 sg13g2_o21ai_1
X_5531_ net1912 net1802 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_2743_ VGND VPWR _0075_ net1697 _0820_ _0819_ sg13g2_a21oi_1
X_5462_ Tile_X0Y1_UserCLK net594 Tile_X0Y1_DSP_bot.C2 _0021_ _5462_/Q VPWR VGND sg13g2_dfrbp_1
X_2674_ VGND VPWR _0125_ _0753_ _0754_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q
+ sg13g2_a21oi_1
X_4413_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q VPWR _2335_
+ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q _2333_ sg13g2_o21ai_1
X_5393_ net1939 net1831 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_4344_ _2275_ VPWR _2276_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q
+ net1615 sg13g2_o21ai_1
X_4275_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q net116 net131
+ net167 net1577 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A
+ VPWR VGND sg13g2_mux4_1
X_6014_ net1990 net226 VPWR VGND sg13g2_buf_1
XFILLER_98_186 VPWR VGND sg13g2_fill_1
X_3226_ _1280_ _1276_ _1279_ _1260_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_39_220 VPWR VGND sg13g2_decap_8
X_3157_ VGND VPWR Tile_X0Y1_DSP_bot.A0 _1209_ _1212_ sg13g2_or2_1
X_3088_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q net140 net108
+ net51 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q
+ _1146_ VPWR VGND sg13g2_mux4_1
X_5729_ net1862 net1735 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_269 VPWR VGND sg13g2_fill_1
Xfanout1805 net1811 net1805 VPWR VGND sg13g2_buf_1
Xfanout1816 net1820 net1816 VPWR VGND sg13g2_buf_1
Xfanout1827 net1830 net1827 VPWR VGND sg13g2_buf_1
Xfanout1838 Tile_X0Y1_FrameStrobe[10] net1838 VPWR VGND sg13g2_buf_1
Xfanout1849 net1850 net1849 VPWR VGND sg13g2_buf_1
Xrebuffer5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 net614 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_54_7 VPWR VGND sg13g2_fill_1
X_5466__598 VPWR VGND net598 sg13g2_tiehi
XFILLER_68_337 VPWR VGND sg13g2_fill_1
X_4060_ _2058_ VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 VGND _2057_ net1652
+ sg13g2_o21ai_1
X_3011_ VGND VPWR _1073_ net1529 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q
+ sg13g2_or2_1
X_4962_ _0505_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q _0504_
+ VPWR VGND sg13g2_nand2_1
X_4893_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q _0082_ _0438_
+ _0439_ VPWR VGND sg13g2_a21o_1
X_3913_ VGND VPWR _1924_ _1925_ _0031_ net1644 sg13g2_a21oi_2
X_3844_ _1871_ _1870_ _1166_ VPWR VGND sg13g2_nand2_2
X_3775_ _1789_ VPWR _1804_ VGND _1803_ _1802_ sg13g2_o21ai_1
X_2726_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q _0800_
+ _0804_ _0803_ sg13g2_a21oi_1
X_5514_ net1877 net1804 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput410 net410 Tile_X0Y1_EE4BEG[13] VPWR VGND sg13g2_buf_1
X_2657_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q _0737_
+ _0738_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q sg13g2_a21oi_1
X_5445_ Tile_X0Y1_UserCLK net577 Tile_X0Y1_DSP_bot.A1 _5445_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[1\]
+ VPWR VGND sg13g2_dfrbp_1
Xoutput421 net421 Tile_X0Y1_EE4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput432 net432 Tile_X0Y1_FrameData_O[19] VPWR VGND sg13g2_buf_1
Xoutput443 net443 Tile_X0Y1_FrameData_O[29] VPWR VGND sg13g2_buf_1
X_5376_ net1966 net1829 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_2588_ net1924 net1659 _0673_ VPWR VGND sg13g2_nor2_1
Xoutput454 net454 Tile_X0Y1_S1BEG[0] VPWR VGND sg13g2_buf_8
Xoutput487 net487 Tile_X0Y1_S4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput465 net465 Tile_X0Y1_S2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput476 net476 Tile_X0Y1_S4BEG[11] VPWR VGND sg13g2_buf_1
X_4327_ _0166_ VPWR _2261_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q
+ net1572 sg13g2_o21ai_1
Xoutput498 net498 Tile_X0Y1_SS4BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_86_101 VPWR VGND sg13g2_fill_1
X_4258_ _2212_ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 VGND _2214_
+ _2216_ sg13g2_o21ai_1
XFILLER_86_134 VPWR VGND sg13g2_fill_2
X_3209_ _1261_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q _1263_
+ _1264_ VPWR VGND sg13g2_a21o_1
XFILLER_103_22 VPWR VGND sg13g2_fill_1
X_4189_ VPWR _2157_ _2156_ VGND sg13g2_inv_1
XFILLER_103_77 VPWR VGND sg13g2_decap_4
XFILLER_42_248 VPWR VGND sg13g2_fill_2
XFILLER_6_149 VPWR VGND sg13g2_fill_2
Xfanout1602 net1607 net1602 VPWR VGND sg13g2_buf_8
Xfanout1613 net1614 net1613 VPWR VGND sg13g2_buf_1
Xfanout1624 net1627 net1624 VPWR VGND sg13g2_buf_1
Xfanout1657 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q net1657 VPWR
+ VGND sg13g2_buf_1
Xfanout1646 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q net1646 VPWR
+ VGND sg13g2_buf_1
XFILLER_77_123 VPWR VGND sg13g2_fill_2
Xfanout1635 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 net1635 VPWR VGND
+ sg13g2_buf_1
Xfanout1679 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q net1679 VPWR
+ VGND sg13g2_buf_1
Xfanout1668 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q net1668 VPWR
+ VGND sg13g2_buf_1
XFILLER_73_340 VPWR VGND sg13g2_fill_1
XFILLER_73_384 VPWR VGND sg13g2_fill_1
XFILLER_53_92 VPWR VGND sg13g2_decap_8
X_3560_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q net1711 net1926
+ net121 net97 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q _1603_
+ VPWR VGND sg13g2_mux4_1
X_2511_ VGND VPWR net124 net1680 _0599_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q
+ sg13g2_a21oi_1
X_3491_ _1509_ _1537_ _1538_ VPWR VGND sg13g2_and2_1
X_5230_ net1996 net1754 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_5161_ net1985 net1778 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_5092_ net1973 net1799 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_4112_ VGND VPWR net136 net1672 _2101_ _2100_ sg13g2_a21oi_1
X_4043_ _2046_ _2035_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 VPWR VGND
+ sg13g2_nor2_2
X_5994_ Tile_X0Y0_EE4END[14] net206 VPWR VGND sg13g2_buf_1
X_4945_ net1695 net1598 net1603 net1623 net1633 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q
+ _0488_ VPWR VGND sg13g2_mux4_1
X_4876_ _0079_ VPWR _0423_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q
+ _0422_ sg13g2_o21ai_1
X_3827_ _1856_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q net1930
+ VPWR VGND sg13g2_nand2b_1
X_3758_ _1785_ _1787_ _1788_ VPWR VGND sg13g2_nor2_1
X_2709_ net1577 net1615 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q
+ _0788_ VPWR VGND sg13g2_mux2_1
X_3689_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q net126 net102
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 net162 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q
+ _1724_ VPWR VGND sg13g2_mux4_1
Xoutput251 net251 Tile_X0Y0_FrameData_O[8] VPWR VGND sg13g2_buf_1
Xoutput262 net262 Tile_X0Y0_FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
Xoutput240 net240 Tile_X0Y0_FrameData_O[27] VPWR VGND sg13g2_buf_1
X_5428_ Tile_X0Y1_UserCLK net570 _0042_ _0016_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[4\]
+ VPWR VGND sg13g2_dfrbp_1
Xoutput273 net273 Tile_X0Y0_N1BEG[0] VPWR VGND sg13g2_buf_1
Xoutput295 net295 Tile_X0Y0_N4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput284 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 Tile_X0Y0_N2BEG[7]
+ VPWR VGND sg13g2_buf_1
X_5359_ net1998 net1839 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_59_156 VPWR VGND sg13g2_fill_1
XFILLER_23_270 VPWR VGND sg13g2_fill_1
XFILLER_24_8 VPWR VGND sg13g2_fill_1
X_2991_ _1053_ VPWR _1054_ VGND _0074_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q
+ sg13g2_o21ai_1
X_4730_ net24 net20 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q _0283_
+ VPWR VGND sg13g2_mux2_1
X_4661_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q VPWR _0217_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q _0216_ sg13g2_o21ai_1
X_3612_ _1651_ _0146_ _1650_ VPWR VGND sg13g2_nand2_1
X_6331_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 net543 VPWR VGND sg13g2_buf_1
X_4592_ VPWR _0149_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q VGND
+ sg13g2_inv_1
X_3543_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q _1587_
+ _1588_ _0140_ sg13g2_a21oi_1
X_3474_ _1522_ VPWR _1523_ VGND net62 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q
+ sg13g2_o21ai_1
XFILLER_43_0 VPWR VGND sg13g2_decap_8
X_6262_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 net489 VPWR VGND sg13g2_buf_1
X_6193_ Tile_X0Y1_EE4END[12] net420 VPWR VGND sg13g2_buf_1
X_5213_ net1959 net1753 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_5144_ net1977 net1789 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_29_307 VPWR VGND sg13g2_fill_2
X_5075_ net1944 net1806 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_4026_ _2030_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q _2029_
+ VPWR VGND sg13g2_nand2_1
X_5977_ Tile_X0Y0_E6END[7] net200 VPWR VGND sg13g2_buf_1
X_4928_ VGND VPWR _0471_ _0472_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q
+ _0470_ sg13g2_a21oi_2
X_4859_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q VPWR _0407_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q _0406_ sg13g2_o21ai_1
XFILLER_109_76 VPWR VGND sg13g2_fill_1
XFILLER_47_159 VPWR VGND sg13g2_fill_1
XFILLER_28_384 VPWR VGND sg13g2_fill_1
XFILLER_43_376 VPWR VGND sg13g2_fill_1
X_3190_ _1245_ _1217_ _1218_ VPWR VGND sg13g2_xnor2_1
XFILLER_78_240 VPWR VGND sg13g2_fill_1
XFILLER_19_384 VPWR VGND sg13g2_fill_1
X_5831_ net1919 net1837 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_5762_ net1865 net1728 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_2974_ _1037_ _0702_ net1575 VPWR VGND sg13g2_nand2_1
X_4713_ _0265_ VPWR _0266_ VGND net1683 net1592 sg13g2_o21ai_1
X_5693_ net1918 net1746 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_4644_ _0200_ VPWR _0201_ VGND net1657 net1577 sg13g2_o21ai_1
X_4575_ VPWR _0132_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q VGND
+ sg13g2_inv_1
XFILLER_115_131 VPWR VGND sg13g2_fill_1
X_6314_ Tile_X0Y1_W6END[11] net537 VPWR VGND sg13g2_buf_1
X_3526_ net1671 net1558 _1572_ VPWR VGND sg13g2_nor2_1
X_6245_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 net466 VPWR VGND sg13g2_buf_1
X_3457_ _1505_ _1454_ _1506_ VPWR VGND sg13g2_xor2_1
X_6176_ Tile_X0Y1_E6END[5] net399 VPWR VGND sg13g2_buf_1
X_3388_ _1440_ _1416_ _1421_ VPWR VGND sg13g2_xnor2_1
X_5127_ net1981 net1787 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_5058_ net1970 net1808 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_84_287 VPWR VGND sg13g2_fill_2
X_4009_ VGND VPWR _2014_ _2012_ _2013_ sg13g2_or2_1
XFILLER_4_214 VPWR VGND sg13g2_fill_2
XFILLER_106_175 VPWR VGND sg13g2_fill_2
XFILLER_45_60 VPWR VGND sg13g2_fill_1
X_2690_ _0703_ _0768_ _0769_ VPWR VGND sg13g2_nor2_2
X_4360_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q VPWR _2290_
+ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q _2287_ sg13g2_o21ai_1
XFILLER_6_76 VPWR VGND sg13g2_fill_2
X_3311_ _1353_ _1362_ _1363_ VPWR VGND sg13g2_nor2_1
X_4291_ net1664 net132 _2238_ VPWR VGND sg13g2_nor2b_1
X_6030_ net1954 net244 VPWR VGND sg13g2_buf_1
X_3242_ _1295_ _1294_ _1293_ VPWR VGND sg13g2_nand2b_1
X_3173_ _1221_ _1227_ _1228_ VPWR VGND sg13g2_nor2b_1
XFILLER_66_210 VPWR VGND sg13g2_fill_2
XFILLER_66_221 VPWR VGND sg13g2_fill_1
Xrebuffer26 net635 net698 VPWR VGND sg13g2_buf_16
Xrebuffer15 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 net624 VPWR VGND
+ sg13g2_buf_8
XFILLER_19_181 VPWR VGND sg13g2_fill_2
Xrebuffer37 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 net646 VPWR VGND
+ sg13g2_dlygate4sd1_1
Xrebuffer59 _0565_ net668 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_81_246 VPWR VGND sg13g2_fill_1
X_5814_ net1902 net1833 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_5745_ net1890 net1727 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_2957_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q VPWR _1021_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q _1020_ sg13g2_o21ai_1
X_2888_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q net118 net134
+ net1927 net94 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q _0957_
+ VPWR VGND sg13g2_mux4_1
X_5676_ net1880 net1746 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
Xrebuffer105 _0929_ net714 VPWR VGND sg13g2_buf_8
Xrebuffer116 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 net725 VPWR VGND
+ sg13g2_dlygate4sd1_1
Xrebuffer127 net737 net736 VPWR VGND sg13g2_buf_2
X_4627_ _0183_ VPWR _0184_ VGND Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q
+ _0181_ sg13g2_o21ai_1
X_4558_ VPWR _0115_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q VGND
+ sg13g2_inv_1
X_4489_ net1512 _2059_ _0046_ VPWR VGND sg13g2_nor2_1
X_3509_ _1555_ VPWR _1556_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q
+ _1552_ sg13g2_o21ai_1
X_6228_ net1881 net441 VPWR VGND sg13g2_buf_1
X_6159_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 net380 VPWR VGND sg13g2_buf_1
XFILLER_57_210 VPWR VGND sg13g2_fill_1
XFILLER_57_298 VPWR VGND sg13g2_fill_1
XFILLER_15_63 VPWR VGND sg13g2_fill_1
XFILLER_31_51 VPWR VGND sg13g2_fill_1
Xinput162 Tile_X0Y1_W2MID[3] net162 VPWR VGND sg13g2_buf_1
Xinput151 Tile_X0Y1_W2END[0] net151 VPWR VGND sg13g2_buf_1
Xinput140 Tile_X0Y1_NN4END[1] net140 VPWR VGND sg13g2_buf_1
XFILLER_48_265 VPWR VGND sg13g2_decap_4
XFILLER_63_224 VPWR VGND sg13g2_decap_8
X_5436__562 VPWR VGND net562 sg13g2_tiehi
X_3860_ _1885_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[0\] net1652 VPWR VGND sg13g2_nand2_1
X_3791_ VGND VPWR _1712_ _1820_ _1818_ _1819_ sg13g2_a21oi_2
X_2811_ _0885_ _0076_ net1689 VPWR VGND sg13g2_nand2_1
X_5530_ net1910 net1802 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_2742_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q VPWR _0819_ VGND
+ net7 net1697 sg13g2_o21ai_1
X_5461_ Tile_X0Y1_UserCLK net593 Tile_X0Y1_DSP_bot.C1 _0023_ _5461_/Q VPWR VGND sg13g2_dfrbp_1
XFILLER_117_259 VPWR VGND sg13g2_fill_2
X_4412_ net1517 _0763_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q
+ _2334_ VPWR VGND sg13g2_mux2_1
X_2673_ _0752_ VPWR _0753_ VGND _0069_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q
+ sg13g2_o21ai_1
X_5392_ net1937 net1831 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_4343_ _2275_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q _1780_
+ VPWR VGND sg13g2_nand2_1
X_4274_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q net115 net134
+ net1703 net1573 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A
+ VPWR VGND sg13g2_mux4_1
XFILLER_98_132 VPWR VGND sg13g2_fill_1
X_3225_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q _1279_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q _1278_ sg13g2_a21oi_2
X_6013_ net1992 net225 VPWR VGND sg13g2_buf_1
X_3156_ VGND VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q net668
+ _1212_ _1211_ sg13g2_a21oi_1
X_3087_ _1145_ VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 VGND _1137_
+ _1135_ sg13g2_o21ai_1
XFILLER_39_298 VPWR VGND sg13g2_fill_2
X_3989_ VGND VPWR net28 net1701 _1994_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q
+ sg13g2_a21oi_1
X_5728_ net1860 net1736 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_5659_ net1912 net1758 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_237 VPWR VGND sg13g2_fill_1
XFILLER_117_76 VPWR VGND sg13g2_fill_1
Xfanout1806 net1808 net1806 VPWR VGND sg13g2_buf_1
Xfanout1828 net1829 net1828 VPWR VGND sg13g2_buf_1
Xfanout1839 net1840 net1839 VPWR VGND sg13g2_buf_1
Xfanout1817 net1818 net1817 VPWR VGND sg13g2_buf_1
XFILLER_45_213 VPWR VGND sg13g2_decap_4
XFILLER_26_95 VPWR VGND sg13g2_fill_2
Xrebuffer6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 net615 VPWR VGND sg13g2_buf_8
X_3010_ net1550 net1559 net1665 _1072_ VPWR VGND sg13g2_mux2_1
X_4961_ net67 net1929 net1695 _0504_ VPWR VGND sg13g2_mux2_1
X_4892_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q VPWR _0438_ VGND
+ net1934 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q sg13g2_o21ai_1
X_3912_ net1645 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X
+ _1924_ VPWR VGND sg13g2_nor2_2
X_3843_ net1515 _0848_ _1870_ VPWR VGND sg13g2_nor2_2
X_3774_ net1636 VPWR _1803_ VGND net1637 _0025_ sg13g2_o21ai_1
X_2725_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q VPWR _0803_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q _0802_ sg13g2_o21ai_1
X_5513_ net1873 net1805 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput400 net400 Tile_X0Y1_E6BEG[4] VPWR VGND sg13g2_buf_1
Xoutput411 net411 Tile_X0Y1_EE4BEG[14] VPWR VGND sg13g2_buf_1
X_5444_ Tile_X0Y1_UserCLK net576 Tile_X0Y1_DSP_bot.A0 _5444_/Q_N Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[0\]
+ VPWR VGND sg13g2_dfrbp_1
X_2656_ net1545 net1552 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ _0737_ VPWR VGND sg13g2_mux2_1
Xoutput444 net444 Tile_X0Y1_FrameData_O[2] VPWR VGND sg13g2_buf_1
Xoutput433 net433 Tile_X0Y1_FrameData_O[1] VPWR VGND sg13g2_buf_1
Xoutput422 net422 Tile_X0Y1_FrameData_O[0] VPWR VGND sg13g2_buf_1
X_2587_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q _0671_ _0665_
+ _0672_ VPWR VGND sg13g2_nand3_1
Xoutput477 net477 Tile_X0Y1_S4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput455 net455 Tile_X0Y1_S1BEG[1] VPWR VGND sg13g2_buf_8
Xoutput466 net466 Tile_X0Y1_S2BEGb[0] VPWR VGND sg13g2_buf_1
X_5375_ net1964 net1828 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_4326_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q _2259_ _2260_
+ VPWR VGND sg13g2_nor2_1
Xoutput499 net499 Tile_X0Y1_SS4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput488 net488 Tile_X0Y1_S4BEG[8] VPWR VGND sg13g2_buf_1
XFILLER_59_305 VPWR VGND sg13g2_fill_1
X_4257_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q VPWR _2216_ VGND
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q _2215_ sg13g2_o21ai_1
XFILLER_86_124 VPWR VGND sg13g2_fill_2
X_3208_ _0128_ VPWR _1263_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q
+ _1262_ sg13g2_o21ai_1
XFILLER_74_319 VPWR VGND sg13g2_fill_1
X_4188_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q net1606 net1634
+ net1626 net1593 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q _2156_
+ VPWR VGND sg13g2_mux4_1
X_3139_ VGND VPWR _1195_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q
+ _1192_ _1190_ _1196_ _1187_ sg13g2_a221oi_1
XFILLER_42_216 VPWR VGND sg13g2_fill_1
XFILLER_12_42 VPWR VGND sg13g2_fill_1
XFILLER_88_46 VPWR VGND sg13g2_fill_2
X_5426__572 VPWR VGND net572 sg13g2_tiehi
Xfanout1614 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 net1614 VPWR VGND
+ sg13g2_buf_8
Xfanout1603 net648 net1603 VPWR VGND sg13g2_buf_1
Xfanout1658 net1659 net1658 VPWR VGND sg13g2_buf_1
Xfanout1647 net1648 net1647 VPWR VGND sg13g2_buf_1
Xfanout1636 _0135_ net1636 VPWR VGND sg13g2_buf_1
Xfanout1625 net1626 net1625 VPWR VGND sg13g2_buf_1
Xfanout1669 net1670 net1669 VPWR VGND sg13g2_buf_1
XFILLER_33_249 VPWR VGND sg13g2_fill_1
X_5433__565 VPWR VGND net565 sg13g2_tiehi
X_3490_ VPWR _1537_ _1536_ VGND sg13g2_inv_1
X_2510_ VPWR _0598_ net621 VGND sg13g2_inv_1
X_5160_ net1983 net1778 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_68_102 VPWR VGND sg13g2_fill_2
X_5091_ net1971 net1799 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_4111_ _0060_ net1672 _2100_ VPWR VGND sg13g2_nor2_1
X_4042_ VGND VPWR _2045_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q
+ _2042_ _2037_ _2046_ _2040_ sg13g2_a221oi_1
X_5440__558 VPWR VGND net558 sg13g2_tiehi
XFILLER_83_116 VPWR VGND sg13g2_fill_1
XFILLER_64_330 VPWR VGND sg13g2_fill_2
X_5993_ Tile_X0Y0_EE4END[13] net220 VPWR VGND sg13g2_buf_1
X_4944_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q _0481_ _0486_
+ _0487_ VPWR VGND sg13g2_nor3_1
X_4875_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q net1713 net1928
+ net115 net107 net1662 _0422_ VPWR VGND sg13g2_mux4_1
X_3826_ _1854_ VPWR _1855_ VGND _0090_ net1678 sg13g2_o21ai_1
X_3757_ _1787_ _1786_ _1435_ VPWR VGND sg13g2_nand2b_1
X_2708_ net1561 net1569 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q
+ _0787_ VPWR VGND sg13g2_mux2_1
X_3688_ VGND VPWR _1721_ _1722_ _1723_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q
+ sg13g2_a21oi_1
Xoutput252 net252 Tile_X0Y0_FrameData_O[9] VPWR VGND sg13g2_buf_1
Xoutput230 net230 Tile_X0Y0_FrameData_O[18] VPWR VGND sg13g2_buf_1
Xoutput241 net241 Tile_X0Y0_FrameData_O[28] VPWR VGND sg13g2_buf_1
X_5427_ Tile_X0Y1_UserCLK net571 _0041_ _0018_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[3\]
+ VPWR VGND sg13g2_dfrbp_1
X_2639_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 _0720_ _0101_ _0711_
+ _0705_ VPWR VGND sg13g2_a22oi_1
Xoutput285 net285 Tile_X0Y0_N2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput274 net274 Tile_X0Y0_N1BEG[1] VPWR VGND sg13g2_buf_1
Xoutput263 net263 Tile_X0Y0_FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
X_5358_ net1995 net1839 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput296 net296 Tile_X0Y0_N4BEG[12] VPWR VGND sg13g2_buf_1
X_4309_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q VPWR _2247_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q net1577 sg13g2_o21ai_1
XFILLER_59_124 VPWR VGND sg13g2_fill_2
X_5289_ net1986 net1729 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_15_216 VPWR VGND sg13g2_fill_1
XFILLER_15_249 VPWR VGND sg13g2_fill_1
XFILLER_15_238 VPWR VGND sg13g2_fill_2
XFILLER_23_260 VPWR VGND sg13g2_fill_2
XFILLER_99_78 VPWR VGND sg13g2_fill_1
XFILLER_3_0 VPWR VGND sg13g2_fill_1
XFILLER_2_164 VPWR VGND sg13g2_fill_1
XFILLER_38_308 VPWR VGND sg13g2_fill_1
XFILLER_46_341 VPWR VGND sg13g2_fill_1
XFILLER_61_333 VPWR VGND sg13g2_fill_1
X_2990_ VGND VPWR net102 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q
+ _1053_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q sg13g2_a21oi_1
X_4660_ net1632 net1585 net1699 _0216_ VPWR VGND sg13g2_mux2_1
X_3611_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q net1532 net1536
+ net1546 net1553 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q _1650_
+ VPWR VGND sg13g2_mux4_1
X_6330_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 net542 VPWR VGND sg13g2_buf_1
X_4591_ VPWR _0148_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q VGND
+ sg13g2_inv_1
XFILLER_115_313 VPWR VGND sg13g2_fill_1
X_3542_ _1586_ VPWR _1587_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q
+ net1581 sg13g2_o21ai_1
X_3473_ _1522_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q net1932
+ VPWR VGND sg13g2_nand2b_1
X_6261_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 net488 VPWR VGND sg13g2_buf_1
X_6192_ Tile_X0Y1_EE4END[11] net419 VPWR VGND sg13g2_buf_1
X_5212_ net1957 net1753 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_36_0 VPWR VGND sg13g2_decap_8
X_5143_ net1955 net1789 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_127 VPWR VGND sg13g2_fill_2
X_5074_ net1942 net1806 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_4025_ VGND VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7
+ _2029_ _2028_ sg13g2_a21oi_1
XFILLER_52_322 VPWR VGND sg13g2_fill_2
X_5976_ Tile_X0Y0_E6END[6] net199 VPWR VGND sg13g2_buf_1
X_4927_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q VPWR _0471_ VGND
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q _0468_ sg13g2_o21ai_1
X_4858_ _0405_ VPWR _0406_ VGND net1685 _0059_ sg13g2_o21ai_1
X_3809_ net138 net22 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q
+ _1838_ VPWR VGND sg13g2_mux2_1
X_4789_ _0338_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q _0339_
+ _0340_ VPWR VGND sg13g2_a21o_1
XFILLER_109_44 VPWR VGND sg13g2_fill_2
XFILLER_47_116 VPWR VGND sg13g2_fill_1
X_5430__568 VPWR VGND net568 sg13g2_tiehi
XFILLER_38_149 VPWR VGND sg13g2_fill_2
XFILLER_46_171 VPWR VGND sg13g2_fill_2
X_5830_ net1896 net1837 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_5761_ net1863 net1726 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_2973_ _1028_ VPWR _1036_ VGND _1025_ _1029_ sg13g2_o21ai_1
X_4712_ _0265_ net1683 net1584 VPWR VGND sg13g2_nand2b_1
X_5692_ net1916 net1746 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_4643_ _0200_ net1657 net1617 VPWR VGND sg13g2_nand2b_1
X_4574_ VPWR _0131_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q VGND
+ sg13g2_inv_1
X_6313_ Tile_X0Y1_W6END[10] net536 VPWR VGND sg13g2_buf_1
X_3525_ VGND VPWR net1671 net1616 _1571_ _1570_ sg13g2_a21oi_1
XFILLER_115_165 VPWR VGND sg13g2_fill_1
X_6244_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 net465 VPWR VGND sg13g2_buf_8
X_3456_ _1505_ _1238_ _1240_ VPWR VGND sg13g2_nand2_1
X_6175_ Tile_X0Y1_E6END[4] net398 VPWR VGND sg13g2_buf_1
X_3387_ _1432_ VPWR _1439_ VGND _1437_ _1436_ sg13g2_o21ai_1
XFILLER_69_230 VPWR VGND sg13g2_fill_2
XFILLER_69_296 VPWR VGND sg13g2_fill_2
X_5126_ net1979 net1787 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_5057_ net1967 net1809 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_4008_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q VPWR _2013_ VGND
+ _1999_ _2011_ sg13g2_o21ai_1
X_5959_ net706 net180 VPWR VGND sg13g2_buf_1
XFILLER_121_135 VPWR VGND sg13g2_fill_1
XFILLER_29_40 VPWR VGND sg13g2_fill_2
XFILLER_29_84 VPWR VGND sg13g2_decap_4
XFILLER_35_108 VPWR VGND sg13g2_fill_2
XFILLER_16_322 VPWR VGND sg13g2_fill_1
XFILLER_16_300 VPWR VGND sg13g2_fill_1
XFILLER_43_141 VPWR VGND sg13g2_fill_1
X_3310_ _1360_ _1361_ _1362_ VPWR VGND sg13g2_nor2b_1
X_4290_ _2232_ _2236_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q
+ _2237_ VPWR VGND sg13g2_nand3_1
X_3241_ _1290_ _1292_ _1241_ _1294_ VPWR VGND sg13g2_nand3_1
X_3172_ _1225_ _1226_ _1227_ VPWR VGND sg13g2_and2_1
Xrebuffer27 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 net636 VPWR VGND sg13g2_buf_2
Xrebuffer16 _0928_ net625 VPWR VGND sg13g2_buf_2
XFILLER_81_203 VPWR VGND sg13g2_decap_4
Xrebuffer38 net716 net647 VPWR VGND sg13g2_buf_8
X_5813_ net1900 net1833 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_5744_ net1888 net1727 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_2956_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q net143 net32 net6
+ net67 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q _1020_ VPWR VGND
+ sg13g2_mux4_1
X_2887_ _0955_ VPWR _0956_ VGND _0954_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q
+ sg13g2_o21ai_1
X_5675_ net1878 net1748 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
Xrebuffer106 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 net715 VPWR VGND
+ sg13g2_buf_8
Xrebuffer128 net738 net737 VPWR VGND sg13g2_buf_2
Xrebuffer117 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 net726 VPWR VGND
+ sg13g2_buf_8
X_4626_ _0183_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q _0182_
+ VPWR VGND sg13g2_nand2b_1
X_4557_ VPWR _0114_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q VGND
+ sg13g2_inv_1
X_4488_ net1514 _1892_ _0045_ VPWR VGND sg13g2_nor2b_1
X_3508_ _0142_ _1554_ _1555_ VPWR VGND sg13g2_nor2_1
X_3439_ VGND VPWR _0116_ _1488_ _1490_ _1489_ sg13g2_a21oi_1
X_6227_ net1883 net440 VPWR VGND sg13g2_buf_1
X_6158_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 net379 VPWR VGND sg13g2_buf_1
XFILLER_66_49 VPWR VGND sg13g2_fill_2
X_5109_ net1947 net1795 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_106_89 VPWR VGND sg13g2_fill_1
X_6089_ Tile_X0Y1_NN4END[9] net316 VPWR VGND sg13g2_buf_1
XFILLER_25_174 VPWR VGND sg13g2_fill_2
XFILLER_40_188 VPWR VGND sg13g2_fill_1
XFILLER_103_0 VPWR VGND sg13g2_fill_2
XFILLER_0_273 VPWR VGND sg13g2_fill_1
Xinput163 Tile_X0Y1_W2MID[4] net163 VPWR VGND sg13g2_buf_1
Xinput152 Tile_X0Y1_W2END[1] net152 VPWR VGND sg13g2_buf_1
Xinput141 Tile_X0Y1_NN4END[2] net141 VPWR VGND sg13g2_buf_1
Xinput130 Tile_X0Y1_N2MID[7] net130 VPWR VGND sg13g2_buf_1
X_3790_ _1819_ _1709_ _1711_ VPWR VGND sg13g2_xnor2_1
X_2810_ _0884_ _0883_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q
+ VPWR VGND sg13g2_nand2b_1
X_2741_ _0817_ VPWR _0818_ VGND net1697 net1527 sg13g2_o21ai_1
X_5460_ Tile_X0Y1_UserCLK net592 Tile_X0Y1_DSP_bot.C0 _0025_ _5460_/Q VPWR VGND sg13g2_dfrbp_1
X_4411_ _2332_ VPWR _2333_ VGND Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q
+ net1615 sg13g2_o21ai_1
X_2672_ _0752_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0
+ VPWR VGND sg13g2_nand2_1
X_5391_ net1998 net1827 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_4342_ _1724_ _1259_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q
+ _2274_ VPWR VGND sg13g2_mux2_1
X_4273_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q net118 net1923
+ net133 net1563 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A
+ VPWR VGND sg13g2_mux4_1
X_3224_ _1277_ _1278_ VPWR VGND sg13g2_inv_4
X_6012_ net1994 net224 VPWR VGND sg13g2_buf_1
.ends

