* NGSPICE file created from RegFile.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_dlhq_1 abstract view
.subckt sg13g2_dlhq_1 D GATE Q VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd1_1 abstract view
.subckt sg13g2_dlygate4sd1_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_16 abstract view
.subckt sg13g2_buf_16 X A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VSS VDD B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_dfrbp_1 abstract view
.subckt sg13g2_dfrbp_1 CLK RESET_B D Q_N Q VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_2 abstract view
.subckt sg13g2_and2_2 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_2 abstract view
.subckt sg13g2_mux2_2 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_16 abstract view
.subckt sg13g2_inv_16 A Y VDD VSS
.ends

.subckt RegFile E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E1END[0] E1END[1] E1END[2] E1END[3]
+ E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3] E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7] E2BEGb[0]
+ E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4] E2BEGb[5] E2BEGb[6] E2BEGb[7] E2END[0] E2END[1]
+ E2END[2] E2END[3] E2END[4] E2END[5] E2END[6] E2END[7] E2MID[0] E2MID[1] E2MID[2]
+ E2MID[3] E2MID[4] E2MID[5] E2MID[6] E2MID[7] E6BEG[0] E6BEG[10] E6BEG[11] E6BEG[1]
+ E6BEG[2] E6BEG[3] E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8] E6BEG[9] E6END[0]
+ E6END[10] E6END[11] E6END[1] E6END[2] E6END[3] E6END[4] E6END[5] E6END[6] E6END[7]
+ E6END[8] E6END[9] EE4BEG[0] EE4BEG[10] EE4BEG[11] EE4BEG[12] EE4BEG[13] EE4BEG[14]
+ EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4] EE4BEG[5] EE4BEG[6] EE4BEG[7]
+ EE4BEG[8] EE4BEG[9] EE4END[0] EE4END[10] EE4END[11] EE4END[12] EE4END[13] EE4END[14]
+ EE4END[15] EE4END[1] EE4END[2] EE4END[3] EE4END[4] EE4END[5] EE4END[6] EE4END[7]
+ EE4END[8] EE4END[9] FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4]
+ N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5]
+ N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6]
+ N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7]
+ N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2]
+ N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12]
+ NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5]
+ NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] NN4END[0] NN4END[10] NN4END[11] NN4END[12]
+ NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3] NN4END[4] NN4END[5]
+ NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S1END[0]
+ S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5]
+ S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6]
+ S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7]
+ S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4BEG[0]
+ S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3]
+ S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] S4END[0] S4END[10] S4END[11]
+ S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5]
+ S4END[6] S4END[7] S4END[8] S4END[9] SS4BEG[0] SS4BEG[10] SS4BEG[11] SS4BEG[12] SS4BEG[13]
+ SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4] SS4BEG[5] SS4BEG[6]
+ SS4BEG[7] SS4BEG[8] SS4BEG[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13]
+ SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6]
+ SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR W1BEG[0] W1BEG[1] W1BEG[2]
+ W1BEG[3] W1END[0] W1END[1] W1END[2] W1END[3] W2BEG[0] W2BEG[1] W2BEG[2] W2BEG[3]
+ W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0] W2BEGb[1] W2BEGb[2] W2BEGb[3] W2BEGb[4]
+ W2BEGb[5] W2BEGb[6] W2BEGb[7] W2END[0] W2END[1] W2END[2] W2END[3] W2END[4] W2END[5]
+ W2END[6] W2END[7] W2MID[0] W2MID[1] W2MID[2] W2MID[3] W2MID[4] W2MID[5] W2MID[6]
+ W2MID[7] W6BEG[0] W6BEG[10] W6BEG[11] W6BEG[1] W6BEG[2] W6BEG[3] W6BEG[4] W6BEG[5]
+ W6BEG[6] W6BEG[7] W6BEG[8] W6BEG[9] W6END[0] W6END[10] W6END[11] W6END[1] W6END[2]
+ W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8] W6END[9] WW4BEG[0] WW4BEG[10]
+ WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15] WW4BEG[1] WW4BEG[2] WW4BEG[3]
+ WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8] WW4BEG[9] WW4END[0] WW4END[10]
+ WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15] WW4END[1] WW4END[2] WW4END[3]
+ WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8] WW4END[9]
X_2106_ _0587_ VPWR _0588_ VGND net1055 net977 sg13g2_o21ai_1
X_3086_ net1210 net1089 Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q VPWR VGND sg13g2_dlhq_1
X_3155_ net1198 net1098 Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q VPWR VGND sg13g2_dlhq_1
X_2037_ net992 Inst_RegFile_32x4.mem\[12\]\[1\] Inst_RegFile_32x4.mem\[13\]\[1\] Inst_RegFile_32x4.mem\[14\]\[1\]
+ Inst_RegFile_32x4.mem\[15\]\[1\] net946 _0525_ VPWR VGND sg13g2_mux4_1
XFILLER_52_18 VPWR VGND sg13g2_fill_2
X_2939_ net1181 net1127 Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q VPWR VGND sg13g2_dlhq_1
Xhold351 Inst_RegFile_32x4.mem\[27\]\[3\] VPWR VGND net849 sg13g2_dlygate4sd3_1
Xhold340 Inst_RegFile_32x4.mem\[21\]\[1\] VPWR VGND net838 sg13g2_dlygate4sd3_1
XFILLER_13_133 VPWR VGND sg13g2_fill_2
XFILLER_5_310 VPWR VGND sg13g2_fill_2
Xrebuffer7 net504 net505 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_47_8 VPWR VGND sg13g2_decap_8
X_2889__433 VPWR VGND net433 sg13g2_tiehi
X_1606_ net60 net68 Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q _1226_ VPWR VGND sg13g2_mux2_1
X_2896__426 VPWR VGND net426 sg13g2_tiehi
X_3773_ WW4END[12] net361 VPWR VGND sg13g2_buf_1
X_2655_ net78 Inst_RegFile_switch_matrix.JW2BEG1 Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q
+ _1070_ VPWR VGND sg13g2_mux2_1
X_2724_ _1033_ _1105_ _1106_ VPWR VGND sg13g2_nor2_2
X_1537_ VPWR _1159_ Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q VGND sg13g2_inv_1
XFILLER_47_29 VPWR VGND sg13g2_fill_2
X_3207_ net1160 net1109 Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q VPWR VGND sg13g2_dlhq_1
X_2586_ Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q net985 _0338_ Inst_RegFile_switch_matrix.E2BEG1
+ net522 Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q Inst_RegFile_switch_matrix.S1BEG2
+ VPWR VGND sg13g2_mux4_1
XFILLER_35_291 VPWR VGND sg13g2_fill_2
X_3138_ net1164 net1093 Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q VPWR VGND sg13g2_dlhq_1
X_3069_ net1176 net1083 Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q VPWR VGND sg13g2_dlhq_1
X_2440_ net1062 net83 _0901_ VPWR VGND sg13g2_nor2b_1
XFILLER_5_173 VPWR VGND sg13g2_fill_2
X_2371_ _0837_ Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q net988 VPWR VGND sg13g2_nand2_1
X_3756_ W6END[5] net340 VPWR VGND sg13g2_buf_1
Xoutput220 net510 N2BEG[6] VPWR VGND sg13g2_buf_1
Xoutput231 net231 N4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput242 net242 N4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput253 net253 NN4BEG[1] VPWR VGND sg13g2_buf_1
X_2569_ Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q VPWR _1012_ VGND _1011_ Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q
+ sg13g2_o21ai_1
Xoutput286 net286 S4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput275 net275 S2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput264 Inst_RegFile_switch_matrix.S1BEG2 S1BEG[2] VPWR VGND sg13g2_buf_1
X_2638_ _1056_ Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q net65 VPWR VGND sg13g2_nand2b_1
X_2707_ net950 net820 _1099_ _0025_ VPWR VGND sg13g2_mux2_1
X_3687_ net511 net269 VPWR VGND sg13g2_buf_1
Xoutput297 net297 S4BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_23_75 VPWR VGND sg13g2_fill_1
XFILLER_11_456 VPWR VGND sg13g2_fill_2
X_2886__436 VPWR VGND net436 sg13g2_tiehi
XFILLER_0_46 VPWR VGND sg13g2_fill_1
X_3610_ net1120 net202 VPWR VGND sg13g2_buf_1
X_1871_ _0365_ VPWR _0366_ VGND _0358_ _0361_ sg13g2_o21ai_1
XFILLER_9_22 VPWR VGND sg13g2_fill_1
X_1940_ VPWR _0432_ _0431_ VGND sg13g2_inv_1
X_2893__429 VPWR VGND net429 sg13g2_tiehi
X_3541_ net14 net123 VPWR VGND sg13g2_buf_1
X_2423_ net999 net1060 _0885_ _0886_ VPWR VGND sg13g2_a21o_1
X_2285_ net718 net970 net1059 _0756_ VPWR VGND sg13g2_mux2_1
X_2354_ VGND VPWR net1046 net999 _0821_ _0820_ sg13g2_a21oi_1
X_3739_ Inst_RegFile_switch_matrix.JW2BEG2 net321 VPWR VGND sg13g2_buf_1
XFILLER_20_231 VPWR VGND sg13g2_decap_4
XFILLER_20_264 VPWR VGND sg13g2_fill_2
XFILLER_47_117 VPWR VGND sg13g2_fill_2
XFILLER_43_301 VPWR VGND sg13g2_decap_4
XFILLER_28_364 VPWR VGND sg13g2_fill_1
XFILLER_7_257 VPWR VGND sg13g2_fill_2
Xfanout1220 net1220 net2 VPWR VGND sg13g2_buf_16
X_2070_ _0556_ _0553_ _0555_ _0551_ _0460_ VPWR VGND sg13g2_a22oi_1
X_2972_ net1179 net1132 Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q VPWR VGND sg13g2_dlhq_1
XFILLER_22_529 VPWR VGND sg13g2_fill_2
X_1854_ VGND VPWR _0349_ _1135_ _0348_ _0343_ _0350_ _0345_ sg13g2_a221oi_1
X_1923_ VGND VPWR net1038 _1166_ _0416_ Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q
+ sg13g2_a21oi_1
X_1785_ VGND VPWR Inst_RegFile_32x4.AD_comb\[1\] _0270_ _0286_ sg13g2_or2_1
X_2406_ net1051 net1070 net1017 net978 net719 Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q
+ _0870_ VPWR VGND sg13g2_mux4_1
X_3386_ UserCLK net494 _0122_ _3386_/Q_N Inst_RegFile_32x4.mem\[11\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_2337_ VGND VPWR _1149_ _0804_ _0805_ _1150_ sg13g2_a21oi_1
XFILLER_57_415 VPWR VGND sg13g2_decap_8
X_2199_ _0674_ _0675_ Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q _0676_ VPWR VGND
+ sg13g2_mux2_1
X_2268_ VGND VPWR _0740_ _0739_ Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q sg13g2_or2_1
XFILLER_56_470 VPWR VGND sg13g2_decap_8
X_1570_ _1191_ net1030 net1048 VPWR VGND sg13g2_nand2b_1
X_3240_ net1158 net1115 Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q VPWR VGND sg13g2_dlhq_1
Xfanout1072 net86 net1072 VPWR VGND sg13g2_buf_1
Xrebuffer17 AD1 net515 VPWR VGND sg13g2_buf_8
X_2122_ Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q net41 net12 net69 net106 Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q
+ _0603_ VPWR VGND sg13g2_mux4_1
Xfanout1061 Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q net1061 VPWR VGND sg13g2_buf_1
XFILLER_39_426 VPWR VGND sg13g2_fill_2
Xfanout1094 net1097 net1094 VPWR VGND sg13g2_buf_1
Xrebuffer39 net538 net537 VPWR VGND sg13g2_dlygate4sd1_1
X_2053_ net990 Inst_RegFile_32x4.mem\[16\]\[3\] Inst_RegFile_32x4.mem\[17\]\[3\] Inst_RegFile_32x4.mem\[18\]\[3\]
+ Inst_RegFile_32x4.mem\[19\]\[3\] net944 _0539_ VPWR VGND sg13g2_mux4_1
Xrebuffer28 net528 net526 VPWR VGND sg13g2_dlygate4sd1_1
X_3171_ net1162 net1098 Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q VPWR VGND sg13g2_dlhq_1
Xfanout1083 net1084 net1083 VPWR VGND sg13g2_buf_1
Xfanout1050 Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q net1050 VPWR VGND sg13g2_buf_1
X_2955_ net26 net1134 Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q VPWR VGND sg13g2_dlhq_1
X_1906_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q _0400_ _0399_ _0398_
+ sg13g2_a21oi_2
X_1768_ VGND VPWR _0269_ _0236_ _0267_ _0263_ _0270_ _0265_ sg13g2_a221oi_1
X_1837_ VGND VPWR net1023 _0331_ _0335_ net955 sg13g2_a21oi_1
X_2886_ UserCLK net436 _0044_ _2886_/Q_N Inst_RegFile_32x4.mem\[23\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_1699_ net1054 net11 net60 net68 net1072 Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q
+ _0205_ VPWR VGND sg13g2_mux4_1
X_3369_ UserCLK net375 _0105_ _3369_/Q_N Inst_RegFile_32x4.mem\[7\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_1_219 VPWR VGND sg13g2_fill_2
XFILLER_53_484 VPWR VGND sg13g2_fill_2
XFILLER_53_440 VPWR VGND sg13g2_fill_2
XFILLER_15_76 VPWR VGND sg13g2_fill_1
XFILLER_0_285 VPWR VGND sg13g2_fill_2
XFILLER_16_131 VPWR VGND sg13g2_fill_1
XFILLER_16_153 VPWR VGND sg13g2_fill_1
X_2671_ Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q _1080_ _1085_ _1086_ VPWR VGND
+ sg13g2_or3_1
X_2740_ net933 net828 _1110_ _0047_ VPWR VGND sg13g2_mux2_1
X_1622_ net9 net24 Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q _0131_ VPWR VGND sg13g2_mux2_1
X_1553_ Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q VPWR _1175_ VGND Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q
+ _1174_ sg13g2_o21ai_1
XFILLER_39_234 VPWR VGND sg13g2_fill_1
X_3223_ net1190 net1111 Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q VPWR VGND sg13g2_dlhq_1
X_2105_ _0587_ net1055 net719 VPWR VGND sg13g2_nand2_1
X_3085_ net1148 net1090 Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q VPWR VGND sg13g2_dlhq_1
XFILLER_35_484 VPWR VGND sg13g2_fill_2
X_2036_ _0524_ _0523_ net1008 VPWR VGND sg13g2_nand2b_1
X_3154_ net1201 net1098 Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q VPWR VGND sg13g2_dlhq_1
X_2938_ net1182 net1130 Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q VPWR VGND sg13g2_dlhq_1
Xhold352 Inst_RegFile_32x4.mem\[25\]\[0\] VPWR VGND net850 sg13g2_dlygate4sd3_1
Xhold341 Inst_RegFile_32x4.mem\[19\]\[2\] VPWR VGND net839 sg13g2_dlygate4sd3_1
Xhold330 Inst_RegFile_32x4.mem\[23\]\[3\] VPWR VGND net828 sg13g2_dlygate4sd3_1
X_2869_ UserCLK net461 _0027_ _2869_/Q_N Inst_RegFile_32x4.mem\[30\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_45_215 VPWR VGND sg13g2_decap_4
XFILLER_45_259 VPWR VGND sg13g2_fill_2
XFILLER_26_451 VPWR VGND sg13g2_fill_1
Xrebuffer8 AD0 net506 VPWR VGND sg13g2_buf_2
XFILLER_3_79 VPWR VGND sg13g2_fill_2
XFILLER_32_487 VPWR VGND sg13g2_fill_1
XFILLER_32_476 VPWR VGND sg13g2_fill_1
X_3772_ WW4END[11] net360 VPWR VGND sg13g2_buf_1
X_2723_ _1025_ _1020_ _1105_ VPWR VGND _1029_ sg13g2_nand3b_1
XFILLER_59_0 VPWR VGND sg13g2_fill_2
X_1605_ net84 net1072 Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q _1225_ VPWR VGND
+ sg13g2_mux2_1
X_2654_ net961 net805 _1062_ _0002_ VPWR VGND sg13g2_mux2_1
X_1536_ VPWR _1158_ Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q VGND sg13g2_inv_1
X_2585_ Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q net1003 _0486_ Inst_RegFile_switch_matrix.E2BEG2
+ _1016_ Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q Inst_RegFile_switch_matrix.S1BEG3
+ VPWR VGND sg13g2_mux4_1
X_3206_ net1166 net1109 Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q VPWR VGND sg13g2_dlhq_1
X_3137_ net1169 net1096 Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q VPWR VGND sg13g2_dlhq_1
XFILLER_42_218 VPWR VGND sg13g2_decap_4
XFILLER_35_270 VPWR VGND sg13g2_decap_8
X_2019_ VGND VPWR _0508_ _0491_ _0506_ _0502_ _0509_ _0504_ sg13g2_a221oi_1
XFILLER_23_465 VPWR VGND sg13g2_fill_2
X_3068_ net1178 net1083 Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q VPWR VGND sg13g2_dlhq_1
XFILLER_58_395 VPWR VGND sg13g2_decap_4
XFILLER_37_96 VPWR VGND sg13g2_fill_2
XFILLER_14_498 VPWR VGND sg13g2_fill_2
XFILLER_52_7 VPWR VGND sg13g2_decap_8
X_2370_ Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q net1072 net1019 AD1 net967 Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q
+ _0836_ VPWR VGND sg13g2_mux4_1
X_3686_ Inst_RegFile_switch_matrix.JS2BEG2 net268 VPWR VGND sg13g2_buf_2
X_3755_ W6END[4] net339 VPWR VGND sg13g2_buf_1
X_2706_ net937 net775 _1099_ _0024_ VPWR VGND sg13g2_mux2_1
Xoutput254 net254 NN4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput210 net210 N1BEG[0] VPWR VGND sg13g2_buf_1
X_1519_ VPWR _1141_ Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q VGND sg13g2_inv_1
Xoutput232 net232 N4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput221 net221 N2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput243 net243 N4BEG[7] VPWR VGND sg13g2_buf_1
X_2568_ VGND VPWR _1010_ _1011_ _0911_ Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q
+ sg13g2_a21oi_2
X_2499_ Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q VPWR _0952_ VGND _0951_ Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q
+ sg13g2_o21ai_1
Xoutput265 Inst_RegFile_switch_matrix.S1BEG3 S1BEG[3] VPWR VGND sg13g2_buf_1
Xoutput276 net276 S2BEGb[2] VPWR VGND sg13g2_buf_1
Xoutput298 net298 SS4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput287 net287 S4BEG[14] VPWR VGND sg13g2_buf_1
X_2637_ VGND VPWR _1054_ _1055_ _1053_ _1163_ sg13g2_a21oi_2
XFILLER_23_251 VPWR VGND sg13g2_fill_2
XFILLER_2_177 VPWR VGND sg13g2_fill_2
XFILLER_46_310 VPWR VGND sg13g2_fill_1
X_1870_ _0364_ Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q _0365_ VPWR VGND sg13g2_nor2b_1
X_3540_ net13 net122 VPWR VGND sg13g2_buf_1
XFILLER_14_284 VPWR VGND sg13g2_fill_1
XFILLER_36_2 VPWR VGND sg13g2_fill_1
X_2353_ Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q VPWR _0820_ VGND net1046 net984
+ sg13g2_o21ai_1
X_2422_ Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q VPWR _0885_ VGND net1060 net984
+ sg13g2_o21ai_1
XFILLER_56_129 VPWR VGND sg13g2_fill_1
X_2284_ _0746_ VPWR Inst_RegFile_switch_matrix.E2BEG1 VGND Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q
+ _0755_ sg13g2_o21ai_1
XFILLER_52_302 VPWR VGND sg13g2_decap_4
X_1999_ VGND VPWR net64 Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q _0489_ _0488_ sg13g2_a21oi_1
X_3669_ NN4END[9] net257 VPWR VGND sg13g2_buf_1
XFILLER_4_409 VPWR VGND sg13g2_fill_1
X_3738_ Inst_RegFile_switch_matrix.JW2BEG1 net320 VPWR VGND sg13g2_buf_1
XFILLER_55_195 VPWR VGND sg13g2_fill_1
XFILLER_43_346 VPWR VGND sg13g2_fill_1
XFILLER_34_20 VPWR VGND sg13g2_fill_2
XFILLER_11_287 VPWR VGND sg13g2_fill_1
X_2892__430 VPWR VGND net430 sg13g2_tiehi
Xfanout1221 net1 net1221 VPWR VGND sg13g2_buf_1
Xfanout1210 net1211 net1210 VPWR VGND sg13g2_buf_1
XFILLER_19_354 VPWR VGND sg13g2_fill_1
X_2971_ net1180 net1132 Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q VPWR VGND sg13g2_dlhq_1
X_1922_ VGND VPWR _0415_ net1038 net109 sg13g2_or2_1
X_1853_ VGND VPWR _1134_ _0349_ _0346_ _1133_ sg13g2_a21oi_2
X_1784_ VGND VPWR net969 _0235_ _0285_ _0275_ _0286_ _0277_ sg13g2_a221oi_1
X_2405_ VGND VPWR _0868_ _0869_ Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q _0865_
+ sg13g2_a21oi_2
X_2336_ net972 net1032 net1042 _0804_ VPWR VGND sg13g2_mux2_1
X_3385_ UserCLK net495 _0121_ _3385_/Q_N Inst_RegFile_32x4.mem\[11\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_41_0 VPWR VGND sg13g2_decap_8
X_2198_ net1044 net1215 net65 net81 net92 Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q
+ _0675_ VPWR VGND sg13g2_mux4_1
XFILLER_37_173 VPWR VGND sg13g2_decap_4
X_2267_ net1050 net1066 net1018 net504 net973 Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q
+ _0739_ VPWR VGND sg13g2_mux4_1
XFILLER_45_63 VPWR VGND sg13g2_fill_2
Xfanout1040 Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q net1040 VPWR VGND sg13g2_buf_1
X_3170_ net1164 net1098 Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q VPWR VGND sg13g2_dlhq_1
Xfanout1051 Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q net1051 VPWR VGND sg13g2_buf_1
X_2121_ VGND VPWR _0601_ _0602_ _0598_ Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q
+ sg13g2_a21oi_2
Xfanout1073 net33 net1073 VPWR VGND sg13g2_buf_1
Xfanout1095 net1096 net1095 VPWR VGND sg13g2_buf_1
Xfanout1062 Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q net1062 VPWR VGND sg13g2_buf_1
Xrebuffer18 net537 net516 VPWR VGND sg13g2_buf_2
X_2052_ VGND VPWR net1004 _0537_ _0538_ _0459_ sg13g2_a21oi_1
Xrebuffer29 net529 net527 VPWR VGND sg13g2_dlygate4sd1_1
Xfanout1084 net1085 net1084 VPWR VGND sg13g2_buf_1
X_1905_ _0399_ net972 net1043 VPWR VGND sg13g2_nand2b_1
X_2954_ net25 net1134 Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q VPWR VGND sg13g2_dlhq_1
X_2885_ UserCLK net437 _0043_ _2885_/Q_N Inst_RegFile_32x4.mem\[22\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_1698_ Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q VPWR _0204_ VGND _0203_ _0200_
+ sg13g2_o21ai_1
X_1836_ _0334_ _0333_ net1023 VPWR VGND sg13g2_nand2b_1
X_1767_ VGND VPWR net983 _0268_ _0269_ _0185_ sg13g2_a21oi_1
XFILLER_57_246 VPWR VGND sg13g2_fill_2
X_3299_ net1162 net1123 Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q VPWR VGND sg13g2_dlhq_1
X_3368_ UserCLK net376 _0104_ _3368_/Q_N Inst_RegFile_32x4.mem\[7\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_2319_ VGND VPWR _0788_ net1041 net1065 sg13g2_or2_1
XFILLER_44_485 VPWR VGND sg13g2_fill_1
XFILLER_31_146 VPWR VGND sg13g2_decap_4
X_1552_ Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q net88 net1019 AD1 net967 Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q
+ _1174_ VPWR VGND sg13g2_mux4_1
X_2670_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q _1083_ _1085_ _1084_ sg13g2_a21oi_1
X_1621_ Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q VPWR _0130_ VGND _1237_ _0129_
+ sg13g2_o21ai_1
X_2104_ _0583_ _0585_ Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q _0586_ VPWR VGND
+ sg13g2_nand3_1
X_3222_ net1192 net1111 Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q VPWR VGND sg13g2_dlhq_1
XFILLER_27_408 VPWR VGND sg13g2_fill_1
X_3153_ net1203 net1099 Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q VPWR VGND sg13g2_dlhq_1
XFILLER_50_422 VPWR VGND sg13g2_fill_2
X_2035_ net995 Inst_RegFile_32x4.mem\[8\]\[1\] Inst_RegFile_32x4.mem\[9\]\[1\] Inst_RegFile_32x4.mem\[10\]\[1\]
+ Inst_RegFile_32x4.mem\[11\]\[1\] net947 _0523_ VPWR VGND sg13g2_mux4_1
X_3084_ net1150 net1090 Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q VPWR VGND sg13g2_dlhq_1
X_2937_ net1184 net1127 Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q VPWR VGND sg13g2_dlhq_1
X_2868_ UserCLK net462 _0026_ _2868_/Q_N Inst_RegFile_32x4.mem\[30\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_2799_ net732 net952 _1123_ _0093_ VPWR VGND sg13g2_mux2_1
X_1819_ net921 Inst_RegFile_32x4.mem\[2\]\[3\] Inst_RegFile_32x4.mem\[3\]\[3\] Inst_RegFile_32x4.mem\[0\]\[3\]
+ Inst_RegFile_32x4.mem\[1\]\[3\] net1022 _0317_ VPWR VGND sg13g2_mux4_1
Xhold320 Inst_RegFile_32x4.mem\[16\]\[3\] VPWR VGND net818 sg13g2_dlygate4sd3_1
Xhold353 Inst_RegFile_32x4.mem\[31\]\[3\] VPWR VGND net851 sg13g2_dlygate4sd3_1
Xhold331 Inst_RegFile_32x4.mem\[31\]\[2\] VPWR VGND net829 sg13g2_dlygate4sd3_1
Xhold342 Inst_RegFile_32x4.mem\[22\]\[2\] VPWR VGND net840 sg13g2_dlygate4sd3_1
XFILLER_53_282 VPWR VGND sg13g2_fill_1
XFILLER_26_43 VPWR VGND sg13g2_fill_1
XFILLER_13_135 VPWR VGND sg13g2_fill_1
XFILLER_13_179 VPWR VGND sg13g2_fill_1
Xrebuffer9 Inst_RegFile_switch_matrix.JW2BEG3 net507 VPWR VGND sg13g2_buf_2
XFILLER_21_190 VPWR VGND sg13g2_fill_2
XFILLER_3_58 VPWR VGND sg13g2_decap_8
XFILLER_3_36 VPWR VGND sg13g2_fill_2
XFILLER_17_463 VPWR VGND sg13g2_fill_1
XFILLER_17_474 VPWR VGND sg13g2_fill_2
X_2722_ net741 net934 _1104_ _0035_ VPWR VGND sg13g2_mux2_1
X_3771_ WW4END[10] net359 VPWR VGND sg13g2_buf_1
X_1604_ net1074 net40 Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q _1224_ VPWR VGND
+ sg13g2_mux2_1
X_1535_ VPWR _1157_ Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q VGND sg13g2_inv_1
X_2653_ Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q _0896_ _0919_ _0486_ _1068_ Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q
+ _1069_ VPWR VGND sg13g2_mux4_1
X_2584_ Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q net1214 net79 net64 net1020 Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q
+ Inst_RegFile_switch_matrix.S4BEG0 VPWR VGND sg13g2_mux4_1
X_3205_ net1188 net1109 Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q VPWR VGND sg13g2_dlhq_1
X_3067_ net1180 net1083 Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q VPWR VGND sg13g2_dlhq_1
X_3136_ net1170 net1096 Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q VPWR VGND sg13g2_dlhq_1
X_2018_ VGND VPWR net1005 _0507_ _0508_ net943 sg13g2_a21oi_1
XFILLER_58_374 VPWR VGND sg13g2_decap_8
Xoutput200 net200 FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
X_3754_ W6END[3] net338 VPWR VGND sg13g2_buf_1
X_3685_ Inst_RegFile_switch_matrix.JS2BEG1 net267 VPWR VGND sg13g2_buf_1
X_2636_ Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q _1031_ _1054_ VPWR VGND sg13g2_and2_1
X_2705_ _1099_ _1090_ _1094_ VPWR VGND sg13g2_nand2_2
Xoutput222 net222 N2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput244 net244 N4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput211 Inst_RegFile_switch_matrix.N1BEG1 N1BEG[1] VPWR VGND sg13g2_buf_1
Xoutput233 net233 N4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput255 net255 NN4BEG[3] VPWR VGND sg13g2_buf_1
X_2567_ Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q net1010 _1010_ VPWR VGND sg13g2_nor2_2
X_2498_ VGND VPWR _0950_ _0951_ _0911_ Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q
+ sg13g2_a21oi_2
X_1518_ VPWR _1140_ Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q VGND sg13g2_inv_1
Xoutput277 net277 S2BEGb[3] VPWR VGND sg13g2_buf_1
Xoutput299 net299 SS4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput266 net266 S2BEG[0] VPWR VGND sg13g2_buf_1
Xoutput288 net288 S4BEG[15] VPWR VGND sg13g2_buf_1
XFILLER_55_388 VPWR VGND sg13g2_decap_8
X_3119_ net1208 net1094 Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q VPWR VGND sg13g2_dlhq_1
XFILLER_15_208 VPWR VGND sg13g2_fill_2
XFILLER_11_458 VPWR VGND sg13g2_fill_1
XFILLER_46_333 VPWR VGND sg13g2_decap_4
XFILLER_34_528 VPWR VGND sg13g2_fill_2
XFILLER_10_491 VPWR VGND sg13g2_fill_1
X_2352_ _0812_ VPWR Inst_RegFile_switch_matrix.JS2BEG7 VGND Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q
+ _0819_ sg13g2_o21ai_1
X_2283_ Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q _0754_ _0752_ _0748_ _0750_ Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q
+ _0755_ VPWR VGND sg13g2_mux4_1
X_2421_ _0883_ VPWR _0884_ VGND net1060 net1029 sg13g2_o21ai_1
XFILLER_37_344 VPWR VGND sg13g2_fill_2
XFILLER_37_311 VPWR VGND sg13g2_fill_2
XFILLER_37_300 VPWR VGND sg13g2_decap_8
XFILLER_20_266 VPWR VGND sg13g2_fill_1
X_3599_ net1181 net173 VPWR VGND sg13g2_buf_1
X_2619_ VGND VPWR net85 Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q _1037_ _1036_ sg13g2_a21oi_1
X_1998_ Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q net36 _0488_ VPWR VGND sg13g2_nor2b_1
X_3668_ NN4END[8] net256 VPWR VGND sg13g2_buf_1
X_3737_ Inst_RegFile_switch_matrix.JW2BEG0 net319 VPWR VGND sg13g2_buf_1
XFILLER_28_377 VPWR VGND sg13g2_fill_1
XFILLER_34_76 VPWR VGND sg13g2_decap_8
XFILLER_11_244 VPWR VGND sg13g2_fill_1
Xfanout1211 FrameData[10] net1211 VPWR VGND sg13g2_buf_1
Xfanout1200 FrameData[15] net1200 VPWR VGND sg13g2_buf_1
X_2970_ net1183 net1133 Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q VPWR VGND sg13g2_dlhq_1
XFILLER_42_380 VPWR VGND sg13g2_fill_1
X_1852_ net999 Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q _0347_ _0348_ VPWR VGND
+ sg13g2_a21o_1
X_1921_ _0413_ VPWR _0414_ VGND net1038 net976 sg13g2_o21ai_1
X_1783_ _0285_ _0283_ _0284_ _0278_ net955 VPWR VGND sg13g2_a22oi_1
X_2404_ Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q VPWR _0868_ VGND Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q
+ _0867_ sg13g2_o21ai_1
X_2335_ VGND VPWR _0802_ _0803_ net987 net1042 sg13g2_a21oi_2
X_3384_ UserCLK net496 _0120_ _3384_/Q_N Inst_RegFile_32x4.mem\[11\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_34_0 VPWR VGND sg13g2_fill_2
X_2266_ _0738_ VPWR Inst_RegFile_switch_matrix.JS2BEG1 VGND _0733_ _0727_ sg13g2_o21ai_1
X_2197_ Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q net37 net8 net1220 net23 Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q
+ _0674_ VPWR VGND sg13g2_mux4_1
XFILLER_25_314 VPWR VGND sg13g2_fill_1
XFILLER_1_80 VPWR VGND sg13g2_fill_2
XFILLER_29_76 VPWR VGND sg13g2_fill_2
XFILLER_29_43 VPWR VGND sg13g2_decap_4
XFILLER_16_347 VPWR VGND sg13g2_fill_2
Xfanout1074 net32 net1074 VPWR VGND sg13g2_buf_1
Xfanout1063 Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q net1063 VPWR VGND sg13g2_buf_1
X_2120_ Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q VPWR _0601_ VGND Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q
+ _0600_ sg13g2_o21ai_1
Xfanout1052 Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q net1052 VPWR VGND sg13g2_buf_1
Xfanout1030 BD0 net1030 VPWR VGND sg13g2_buf_1
Xfanout1041 Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q net1041 VPWR VGND sg13g2_buf_1
Xrebuffer19 Inst_RegFile_switch_matrix.JN2BEG3 net517 VPWR VGND sg13g2_dlygate4sd1_1
Xfanout1096 net1097 net1096 VPWR VGND sg13g2_buf_1
X_2051_ net990 Inst_RegFile_32x4.mem\[28\]\[3\] Inst_RegFile_32x4.mem\[29\]\[3\] Inst_RegFile_32x4.mem\[30\]\[3\]
+ Inst_RegFile_32x4.mem\[31\]\[3\] net944 _0537_ VPWR VGND sg13g2_mux4_1
Xfanout1085 FrameStrobe[8] net1085 VPWR VGND sg13g2_buf_1
X_1904_ _0398_ net1043 net1014 VPWR VGND sg13g2_nand2_2
XFILLER_22_339 VPWR VGND sg13g2_fill_1
X_1835_ VGND VPWR Inst_RegFile_32x4.mem\[23\]\[3\] net923 _0333_ _0332_ sg13g2_a21oi_1
X_2884_ UserCLK net438 _0042_ _2884_/Q_N Inst_RegFile_32x4.mem\[22\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_2953_ net1156 net1131 Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q VPWR VGND sg13g2_dlhq_1
X_1697_ Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q VPWR _0203_ VGND _0201_ _0202_
+ sg13g2_o21ai_1
X_1766_ net931 Inst_RegFile_32x4.mem\[6\]\[1\] Inst_RegFile_32x4.mem\[7\]\[1\] Inst_RegFile_32x4.mem\[4\]\[1\]
+ Inst_RegFile_32x4.mem\[5\]\[1\] net1028 _0268_ VPWR VGND sg13g2_mux4_1
X_3298_ net1165 net1123 Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q VPWR VGND sg13g2_dlhq_1
X_3367_ UserCLK net377 _0103_ _3367_/Q_N Inst_RegFile_32x4.mem\[6\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_2249_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q _0721_ _0723_ _0722_ sg13g2_a21oi_1
X_2318_ net963 net970 net1041 _0787_ VPWR VGND sg13g2_mux2_1
XFILLER_53_475 VPWR VGND sg13g2_fill_1
XFILLER_53_464 VPWR VGND sg13g2_decap_8
XFILLER_31_88 VPWR VGND sg13g2_fill_2
X_3377__367 VPWR VGND net367 sg13g2_tiehi
XFILLER_0_287 VPWR VGND sg13g2_fill_1
Xinput100 W2MID[3] net100 VPWR VGND sg13g2_buf_1
X_1551_ _1172_ _1169_ _1141_ _1173_ VPWR VGND sg13g2_nor3_2
X_1620_ _0128_ Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q _1143_ _0129_ VPWR VGND
+ sg13g2_a21o_1
XFILLER_39_203 VPWR VGND sg13g2_decap_4
X_2103_ _0584_ VPWR _0585_ VGND net1055 net971 sg13g2_o21ai_1
X_3221_ net1194 net1111 Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q VPWR VGND sg13g2_dlhq_1
X_3152_ net1206 net1098 Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q VPWR VGND sg13g2_dlhq_1
X_3083_ net1152 net1088 Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q VPWR VGND sg13g2_dlhq_1
XFILLER_50_434 VPWR VGND sg13g2_fill_2
X_2034_ VGND VPWR net532 _0522_ _0521_ _0519_ sg13g2_a21oi_2
X_2936_ net1186 net1127 Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q VPWR VGND sg13g2_dlhq_1
X_2798_ net726 net940 _1123_ _0092_ VPWR VGND sg13g2_mux2_1
Xhold310 Inst_RegFile_32x4.mem\[29\]\[2\] VPWR VGND net808 sg13g2_dlygate4sd3_1
X_2867_ UserCLK net463 _0025_ _2867_/Q_N Inst_RegFile_32x4.mem\[30\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_1818_ VGND VPWR net956 _0313_ _0316_ net969 sg13g2_a21oi_1
Xhold332 Inst_RegFile_32x4.mem\[25\]\[3\] VPWR VGND net830 sg13g2_dlygate4sd3_1
Xhold321 Inst_RegFile_32x4.mem\[27\]\[2\] VPWR VGND net819 sg13g2_dlygate4sd3_1
Xhold343 Inst_RegFile_32x4.mem\[23\]\[0\] VPWR VGND net841 sg13g2_dlygate4sd3_1
X_1749_ _0253_ Inst_RegFile_32x4.mem\[18\]\[0\] net925 VPWR VGND sg13g2_nand2b_1
XFILLER_21_180 VPWR VGND sg13g2_fill_2
XFILLER_44_294 VPWR VGND sg13g2_decap_4
X_2721_ net753 net960 _1104_ _0034_ VPWR VGND sg13g2_mux2_1
X_3770_ WW4END[9] net358 VPWR VGND sg13g2_buf_1
X_2652_ Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q net51 net1065 net1214 Inst_RegFile_switch_matrix.JS2BEG1
+ Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q _1068_ VPWR VGND sg13g2_mux4_1
XFILLER_59_2 VPWR VGND sg13g2_fill_1
X_1603_ net3 net11 Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q _1223_ VPWR VGND sg13g2_mux2_1
X_1534_ VPWR _1156_ Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q VGND sg13g2_inv_1
X_3204_ net1212 net1109 Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q VPWR VGND sg13g2_dlhq_1
X_2583_ Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q net1216 net65 net80 net979 Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q
+ Inst_RegFile_switch_matrix.S4BEG1 VPWR VGND sg13g2_mux4_1
X_3135_ net1172 net1094 Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q VPWR VGND sg13g2_dlhq_1
X_3367__377 VPWR VGND net377 sg13g2_tiehi
X_2017_ net992 Inst_RegFile_32x4.mem\[20\]\[0\] Inst_RegFile_32x4.mem\[21\]\[0\] Inst_RegFile_32x4.mem\[22\]\[0\]
+ Inst_RegFile_32x4.mem\[23\]\[0\] net945 _0507_ VPWR VGND sg13g2_mux4_1
X_3066_ net1182 net1083 Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q VPWR VGND sg13g2_dlhq_1
XFILLER_50_275 VPWR VGND sg13g2_fill_2
XFILLER_35_250 VPWR VGND sg13g2_fill_1
X_2919_ net1161 net1130 Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q VPWR VGND sg13g2_dlhq_1
XFILLER_23_489 VPWR VGND sg13g2_fill_2
XFILLER_23_467 VPWR VGND sg13g2_fill_1
XFILLER_2_338 VPWR VGND sg13g2_fill_2
XFILLER_46_504 VPWR VGND sg13g2_fill_1
XFILLER_41_242 VPWR VGND sg13g2_fill_1
XFILLER_37_54 VPWR VGND sg13g2_fill_2
XFILLER_37_43 VPWR VGND sg13g2_decap_8
XFILLER_49_320 VPWR VGND sg13g2_decap_4
Xoutput201 net201 FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
Xoutput234 net234 N4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput223 net223 N2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput212 Inst_RegFile_switch_matrix.N1BEG2 N1BEG[2] VPWR VGND sg13g2_buf_1
X_2635_ Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q net44 net99 net15 Inst_RegFile_switch_matrix.E2BEG4
+ Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q _1053_ VPWR VGND sg13g2_mux4_1
X_2704_ net733 net932 _1098_ _0023_ VPWR VGND sg13g2_mux2_1
X_3753_ W6END[2] net335 VPWR VGND sg13g2_buf_1
X_3684_ Inst_RegFile_switch_matrix.JS2BEG0 net266 VPWR VGND sg13g2_buf_1
Xoutput256 net256 NN4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput245 net245 N4BEG[9] VPWR VGND sg13g2_buf_1
X_2566_ _1008_ VPWR _1009_ VGND Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q _0910_
+ sg13g2_o21ai_1
X_2497_ Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q net1010 _0950_ VPWR VGND sg13g2_nor2_2
Xoutput289 net289 S4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput278 net278 S2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput267 net267 S2BEG[1] VPWR VGND sg13g2_buf_1
X_1517_ VPWR _1139_ Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q VGND sg13g2_inv_1
X_3118_ net1211 net1097 Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q VPWR VGND sg13g2_dlhq_1
XFILLER_23_220 VPWR VGND sg13g2_fill_2
X_3049_ net1157 net1085 Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q VPWR VGND sg13g2_dlhq_1
XFILLER_2_179 VPWR VGND sg13g2_fill_1
XFILLER_48_75 VPWR VGND sg13g2_fill_1
XFILLER_46_356 VPWR VGND sg13g2_fill_2
X_3357__387 VPWR VGND net387 sg13g2_tiehi
X_2420_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q _0883_ net1010 net1060
+ sg13g2_a21oi_2
X_2351_ _0818_ VPWR _0819_ VGND Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q _0813_
+ sg13g2_o21ai_1
X_2282_ VGND VPWR net36 net1049 _0754_ _0753_ sg13g2_a21oi_1
X_1997_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q _0486_ _0487_ _1140_ sg13g2_a21oi_1
X_3598_ net1183 net172 VPWR VGND sg13g2_buf_1
X_2549_ Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q net1033 net499 net500 _0994_ Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q
+ _0995_ VPWR VGND sg13g2_mux4_1
X_2618_ Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q net8 _1036_ VPWR VGND sg13g2_nor2b_1
X_3667_ NN4END[7] net255 VPWR VGND sg13g2_buf_1
XFILLER_50_21 VPWR VGND sg13g2_decap_8
XFILLER_3_411 VPWR VGND sg13g2_fill_2
Xfanout1212 FrameData[0] net1212 VPWR VGND sg13g2_buf_1
Xfanout1201 net1202 net1201 VPWR VGND sg13g2_buf_1
X_1851_ Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q VPWR _0347_ VGND Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q
+ net987 sg13g2_o21ai_1
X_1920_ _0413_ net1038 net504 VPWR VGND sg13g2_nand2_1
X_2403_ VGND VPWR net1051 net1031 _0867_ _0866_ sg13g2_a21oi_1
X_3383_ UserCLK net497 _0119_ _3383_/Q_N Inst_RegFile_32x4.mem\[10\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_1782_ VGND VPWR net1023 _0280_ _0284_ net955 sg13g2_a21oi_1
XFILLER_57_429 VPWR VGND sg13g2_decap_8
X_2196_ Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q VPWR _0673_ VGND _0666_ _0667_
+ sg13g2_o21ai_1
X_2334_ net1042 net1014 _0802_ VPWR VGND sg13g2_nor2b_1
XFILLER_27_0 VPWR VGND sg13g2_fill_2
X_2265_ _0737_ VPWR _0738_ VGND Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q _0734_ sg13g2_o21ai_1
XFILLER_52_156 VPWR VGND sg13g2_fill_2
X_3719_ SS4END[7] net307 VPWR VGND sg13g2_buf_1
XFILLER_48_418 VPWR VGND sg13g2_fill_1
XFILLER_45_65 VPWR VGND sg13g2_fill_1
X_3347__397 VPWR VGND net397 sg13g2_tiehi
XFILLER_24_370 VPWR VGND sg13g2_fill_1
Xfanout1042 Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q net1042 VPWR VGND sg13g2_buf_1
Xfanout1064 Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q net1064 VPWR VGND sg13g2_buf_1
Xfanout1075 net1075 net31 VPWR VGND sg13g2_buf_16
Xfanout1053 Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q net1053 VPWR VGND sg13g2_buf_1
X_2050_ _0535_ VPWR _0536_ VGND net1036 _0534_ sg13g2_o21ai_1
Xfanout1097 FrameStrobe[6] net1097 VPWR VGND sg13g2_buf_1
Xfanout1031 BD0 net1031 VPWR VGND sg13g2_buf_1
Xfanout1086 FrameStrobe[8] net1086 VPWR VGND sg13g2_buf_1
Xfanout1020 AD0 net1020 VPWR VGND sg13g2_buf_1
X_2952_ net1158 net1131 Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q VPWR VGND sg13g2_dlhq_1
XFILLER_19_186 VPWR VGND sg13g2_fill_2
X_1903_ Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q VPWR _0397_ VGND net1043 net987
+ sg13g2_o21ai_1
X_1834_ net924 Inst_RegFile_32x4.mem\[22\]\[3\] _0332_ VPWR VGND sg13g2_nor2b_1
X_2883_ UserCLK net447 _0041_ _2883_/Q_N Inst_RegFile_32x4.mem\[22\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_1765_ _0267_ _0143_ _0266_ VPWR VGND sg13g2_nand2_2
X_1696_ Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q VPWR _0202_ VGND net1054 net986
+ sg13g2_o21ai_1
X_3366_ UserCLK net378 _0102_ _3366_/Q_N Inst_RegFile_32x4.mem\[6\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_3297_ net1168 net1123 Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q VPWR VGND sg13g2_dlhq_1
X_2317_ _0786_ VPWR Inst_RegFile_switch_matrix.JW2BEG7 VGND _0775_ _0782_ sg13g2_o21ai_1
X_2179_ Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q net1215 _0657_ VPWR VGND sg13g2_nor2b_1
X_2248_ Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q _0720_ _0722_ VPWR VGND sg13g2_nor2b_1
XFILLER_40_115 VPWR VGND sg13g2_fill_2
XFILLER_25_167 VPWR VGND sg13g2_decap_4
Xinput101 W2MID[4] net101 VPWR VGND sg13g2_buf_1
XFILLER_16_101 VPWR VGND sg13g2_decap_8
X_1550_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q _1172_ _1170_ _1171_
+ sg13g2_a21oi_2
X_3220_ net1196 net1111 Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q VPWR VGND sg13g2_dlhq_1
X_3332__441 VPWR VGND net441 sg13g2_tiehi
X_2102_ VGND VPWR net1055 net1011 _0584_ Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q
+ sg13g2_a21oi_1
X_3151_ net1209 net1100 Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q VPWR VGND sg13g2_dlhq_1
X_2033_ VGND VPWR net1007 _0520_ _0521_ net943 sg13g2_a21oi_1
X_3082_ net1154 net1088 Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q VPWR VGND sg13g2_dlhq_1
X_2935_ net1190 net1129 Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q VPWR VGND sg13g2_dlhq_1
Xhold333 Inst_RegFile_32x4.mem\[9\]\[1\] VPWR VGND net831 sg13g2_dlygate4sd3_1
X_1817_ _0315_ net983 _0314_ VPWR VGND sg13g2_nand2_1
Xhold311 Inst_RegFile_32x4.mem\[29\]\[3\] VPWR VGND net809 sg13g2_dlygate4sd3_1
X_1748_ VGND VPWR Inst_RegFile_32x4.mem\[17\]\[0\] net925 _0252_ _0251_ sg13g2_a21oi_1
Xhold344 Inst_RegFile_32x4.mem\[30\]\[2\] VPWR VGND net842 sg13g2_dlygate4sd3_1
Xhold322 Inst_RegFile_32x4.mem\[30\]\[1\] VPWR VGND net820 sg13g2_dlygate4sd3_1
Xhold300 Inst_RegFile_32x4.mem\[17\]\[0\] VPWR VGND net798 sg13g2_dlygate4sd3_1
X_2866_ UserCLK net464 _0024_ _2866_/Q_N Inst_RegFile_32x4.mem\[30\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_2797_ _1061_ _1122_ _1123_ VPWR VGND sg13g2_and2_2
XFILLER_58_513 VPWR VGND sg13g2_fill_2
X_1679_ _0184_ _0167_ _0185_ VPWR VGND sg13g2_and2_1
X_3349_ UserCLK net395 _0085_ _3349_/Q_N Inst_RegFile_32x4.mem\[31\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_45_229 VPWR VGND sg13g2_fill_2
XFILLER_41_402 VPWR VGND sg13g2_fill_1
XFILLER_42_11 VPWR VGND sg13g2_fill_2
X_1602_ Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q VPWR _1222_ VGND _1219_ _1221_
+ sg13g2_o21ai_1
X_2582_ Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q net62 net1065 net81 net967 Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q
+ Inst_RegFile_switch_matrix.S4BEG2 VPWR VGND sg13g2_mux4_1
X_2651_ net953 net767 _1062_ _0001_ VPWR VGND sg13g2_mux2_1
X_2720_ net751 net951 _1104_ _0033_ VPWR VGND sg13g2_mux2_1
X_3203_ net1163 net1105 Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q VPWR VGND sg13g2_dlhq_1
X_1533_ VPWR _1155_ Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q VGND sg13g2_inv_1
X_3134_ net1175 net1094 Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q VPWR VGND sg13g2_dlhq_1
X_3065_ net1184 net1084 Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q VPWR VGND sg13g2_dlhq_1
X_2016_ _0506_ _0505_ net1005 VPWR VGND sg13g2_nand2b_1
XFILLER_50_287 VPWR VGND sg13g2_fill_2
XFILLER_35_284 VPWR VGND sg13g2_decap_8
XFILLER_31_490 VPWR VGND sg13g2_fill_2
X_2918_ net1167 net1130 Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q VPWR VGND sg13g2_dlhq_1
X_2849_ UserCLK net481 _0007_ _2849_/Q_N Inst_RegFile_32x4.mem\[25\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_53_87 VPWR VGND sg13g2_fill_1
XFILLER_53_21 VPWR VGND sg13g2_fill_2
XFILLER_37_77 VPWR VGND sg13g2_fill_1
XFILLER_5_122 VPWR VGND sg13g2_fill_1
XFILLER_5_133 VPWR VGND sg13g2_fill_2
X_3752_ net104 net334 VPWR VGND sg13g2_buf_1
Xoutput202 net202 FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
Xoutput257 net257 NN4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput246 net246 NN4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput224 net224 N2BEGb[2] VPWR VGND sg13g2_buf_1
Xoutput213 Inst_RegFile_switch_matrix.N1BEG3 N1BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_57_0 VPWR VGND sg13g2_decap_8
Xoutput235 net235 N4BEG[14] VPWR VGND sg13g2_buf_1
X_3373__371 VPWR VGND net371 sg13g2_tiehi
X_2565_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q _0363_ _1008_ _1160_
+ sg13g2_a21oi_1
Xoutput268 net268 S2BEG[2] VPWR VGND sg13g2_buf_1
X_2703_ net745 net959 _1098_ _0022_ VPWR VGND sg13g2_mux2_1
X_1516_ VPWR _1138_ net107 VGND sg13g2_inv_1
X_2634_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q Inst_RegFile_switch_matrix.JN2BEG0
+ _1052_ _1051_ sg13g2_a21oi_1
XFILLER_59_129 VPWR VGND sg13g2_fill_2
X_3117_ net1148 net1095 Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q VPWR VGND sg13g2_dlhq_1
X_2496_ _0948_ VPWR _0949_ VGND Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q _0910_
+ sg13g2_o21ai_1
Xoutput279 net279 S2BEGb[5] VPWR VGND sg13g2_buf_1
X_3380__364 VPWR VGND net364 sg13g2_tiehi
X_3048_ net1159 net1086 Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q VPWR VGND sg13g2_dlhq_1
XFILLER_48_32 VPWR VGND sg13g2_fill_2
XFILLER_48_21 VPWR VGND sg13g2_decap_8
XFILLER_48_54 VPWR VGND sg13g2_fill_1
XFILLER_14_243 VPWR VGND sg13g2_fill_1
XFILLER_50_7 VPWR VGND sg13g2_decap_8
X_2350_ _0817_ VPWR _0818_ VGND Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q _0816_
+ sg13g2_o21ai_1
X_2281_ net1049 net1076 _0753_ VPWR VGND sg13g2_nor2b_1
XFILLER_37_346 VPWR VGND sg13g2_fill_1
XFILLER_33_530 VPWR VGND sg13g2_fill_1
X_1996_ Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q net47 net18 net75 net102 Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q
+ _0486_ VPWR VGND sg13g2_mux4_1
XFILLER_20_224 VPWR VGND sg13g2_fill_2
X_3597_ net1185 net171 VPWR VGND sg13g2_buf_1
X_2617_ net108 Inst_RegFile_switch_matrix.JN2BEG2 Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q
+ _1035_ VPWR VGND sg13g2_mux2_1
X_2548_ Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q net54 net64 net7 net91 Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q
+ _0994_ VPWR VGND sg13g2_mux4_1
X_3666_ NN4END[6] net254 VPWR VGND sg13g2_buf_1
XFILLER_43_305 VPWR VGND sg13g2_fill_1
X_2479_ Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q net34 net62 net5 net109 Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q
+ _0935_ VPWR VGND sg13g2_mux4_1
XFILLER_16_519 VPWR VGND sg13g2_fill_2
XFILLER_51_393 VPWR VGND sg13g2_decap_8
Xfanout1213 FrameData[0] net1213 VPWR VGND sg13g2_buf_1
Xfanout1202 FrameData[14] net1202 VPWR VGND sg13g2_buf_1
X_3363__381 VPWR VGND net381 sg13g2_tiehi
XFILLER_15_530 VPWR VGND sg13g2_fill_1
XFILLER_19_379 VPWR VGND sg13g2_fill_2
XFILLER_42_393 VPWR VGND sg13g2_fill_1
X_1850_ net971 net1013 Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q _0346_ VPWR VGND
+ sg13g2_mux2_1
X_1781_ _0283_ _0282_ net1023 VPWR VGND sg13g2_nand2b_1
X_2402_ net1051 net972 _0866_ VPWR VGND sg13g2_nor2b_1
X_3382_ UserCLK net498 _0118_ _3382_/Q_N Inst_RegFile_32x4.mem\[10\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_34_2 VPWR VGND sg13g2_fill_1
X_2333_ _0801_ VPWR Inst_RegFile_switch_matrix.JW2BEG0 VGND _0796_ _0790_ sg13g2_o21ai_1
X_3370__374 VPWR VGND net374 sg13g2_tiehi
XFILLER_57_408 VPWR VGND sg13g2_decap_8
X_2195_ VGND VPWR _0671_ Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q _0670_ Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q
+ _0672_ _0669_ sg13g2_a221oi_1
XFILLER_1_71 VPWR VGND sg13g2_fill_1
XFILLER_1_82 VPWR VGND sg13g2_fill_1
X_2264_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q _0736_ _0737_ Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q
+ sg13g2_a21oi_1
X_3718_ SS4END[6] net306 VPWR VGND sg13g2_buf_1
X_1979_ VGND VPWR net1052 net1032 _0470_ _0469_ sg13g2_a21oi_1
X_3649_ N4END[5] net237 VPWR VGND sg13g2_buf_1
XFILLER_29_78 VPWR VGND sg13g2_fill_1
XFILLER_56_463 VPWR VGND sg13g2_decap_8
XFILLER_28_154 VPWR VGND sg13g2_fill_2
Xfanout1076 net30 net1076 VPWR VGND sg13g2_buf_1
Xfanout1054 Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q net1054 VPWR VGND sg13g2_buf_1
Xfanout1065 net105 net1065 VPWR VGND sg13g2_buf_1
Xfanout1043 Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q net1043 VPWR VGND sg13g2_buf_1
Xfanout1010 net1010 _1164_ VPWR VGND sg13g2_buf_16
Xfanout1032 BD0 net1032 VPWR VGND sg13g2_buf_8
Xfanout1098 net1102 net1098 VPWR VGND sg13g2_buf_1
Xfanout1087 FrameStrobe[8] net1087 VPWR VGND sg13g2_buf_1
X_1902_ net1003 net1043 _0396_ VPWR VGND sg13g2_nor2b_1
XFILLER_34_157 VPWR VGND sg13g2_decap_4
X_2951_ net1161 net1136 Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q VPWR VGND sg13g2_dlhq_1
XFILLER_15_360 VPWR VGND sg13g2_fill_2
X_1833_ VGND VPWR Inst_RegFile_32x4.mem\[21\]\[3\] net923 _0331_ _0330_ sg13g2_a21oi_1
X_1764_ net921 Inst_RegFile_32x4.mem\[2\]\[1\] Inst_RegFile_32x4.mem\[3\]\[1\] Inst_RegFile_32x4.mem\[0\]\[1\]
+ Inst_RegFile_32x4.mem\[1\]\[1\] net1022 _0266_ VPWR VGND sg13g2_mux4_1
X_2882_ UserCLK net448 _0040_ _2882_/Q_N Inst_RegFile_32x4.mem\[22\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_3296_ net1171 net1123 Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q VPWR VGND sg13g2_dlhq_1
X_1695_ net1002 net1054 _0201_ VPWR VGND sg13g2_nor2b_1
X_2316_ _0786_ _0785_ Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q VPWR VGND sg13g2_nand2b_1
X_3365_ UserCLK net379 _0101_ _3365_/Q_N Inst_RegFile_32x4.mem\[6\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_2178_ net81 net92 Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q _0656_ VPWR VGND sg13g2_mux2_1
XFILLER_25_135 VPWR VGND sg13g2_decap_8
X_2247_ net1040 net64 net80 net83 net91 Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q
+ _0721_ VPWR VGND sg13g2_mux4_1
XFILLER_53_499 VPWR VGND sg13g2_fill_2
X_3353__391 VPWR VGND net391 sg13g2_tiehi
XFILLER_56_65 VPWR VGND sg13g2_fill_1
XFILLER_56_21 VPWR VGND sg13g2_decap_8
Xinput102 W2MID[5] net102 VPWR VGND sg13g2_buf_1
XFILLER_56_293 VPWR VGND sg13g2_fill_1
X_3360__384 VPWR VGND net384 sg13g2_tiehi
X_3150_ net1210 net1100 Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q VPWR VGND sg13g2_dlhq_1
X_2101_ _1165_ net1055 _0582_ _0583_ VPWR VGND sg13g2_a21o_1
X_2032_ net991 Inst_RegFile_32x4.mem\[20\]\[1\] Inst_RegFile_32x4.mem\[21\]\[1\] Inst_RegFile_32x4.mem\[22\]\[1\]
+ Inst_RegFile_32x4.mem\[23\]\[1\] net945 _0520_ VPWR VGND sg13g2_mux4_1
X_3081_ net1156 net1089 Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q VPWR VGND sg13g2_dlhq_1
XFILLER_50_436 VPWR VGND sg13g2_fill_1
X_2865_ UserCLK net465 _0023_ _2865_/Q_N Inst_RegFile_32x4.mem\[2\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_2934_ net1192 net1129 Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q VPWR VGND sg13g2_dlhq_1
Xhold323 Inst_RegFile_32x4.mem\[9\]\[0\] VPWR VGND net821 sg13g2_dlygate4sd3_1
Xhold301 Inst_RegFile_32x4.mem\[24\]\[3\] VPWR VGND net799 sg13g2_dlygate4sd3_1
Xhold312 Inst_RegFile_32x4.mem\[25\]\[1\] VPWR VGND net810 sg13g2_dlygate4sd3_1
X_1816_ net930 Inst_RegFile_32x4.mem\[14\]\[3\] Inst_RegFile_32x4.mem\[15\]\[3\] Inst_RegFile_32x4.mem\[12\]\[3\]
+ Inst_RegFile_32x4.mem\[13\]\[3\] net1026 _0314_ VPWR VGND sg13g2_mux4_1
X_1678_ _0184_ _0182_ _0183_ VPWR VGND sg13g2_nand2_2
Xhold345 Inst_RegFile_32x4.mem\[1\]\[0\] VPWR VGND net843 sg13g2_dlygate4sd3_1
X_1747_ net925 Inst_RegFile_32x4.mem\[16\]\[0\] _0251_ VPWR VGND sg13g2_nor2b_1
Xhold334 Inst_RegFile_32x4.mem\[23\]\[1\] VPWR VGND net832 sg13g2_dlygate4sd3_1
X_2796_ _1033_ _1096_ _1122_ VPWR VGND sg13g2_and2_1
X_3279_ net1208 net1124 Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q VPWR VGND sg13g2_dlhq_1
XFILLER_45_208 VPWR VGND sg13g2_decap_8
X_3348_ UserCLK net396 _0084_ _3348_/Q_N Inst_RegFile_32x4.mem\[31\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_38_260 VPWR VGND sg13g2_fill_1
XFILLER_42_56 VPWR VGND sg13g2_fill_2
XFILLER_42_34 VPWR VGND sg13g2_fill_1
XFILLER_44_241 VPWR VGND sg13g2_fill_2
XFILLER_36_208 VPWR VGND sg13g2_fill_2
XFILLER_29_271 VPWR VGND sg13g2_fill_1
X_1601_ _1220_ Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q _1142_ _1221_ VPWR VGND
+ sg13g2_a21o_1
X_1532_ VPWR _1154_ Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q VGND sg13g2_inv_1
X_2650_ Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q _0484_ _0911_ _0994_ _1066_ Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q
+ _1067_ VPWR VGND sg13g2_mux4_1
X_2581_ Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q net63 net1067 net78 net975 Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q
+ Inst_RegFile_switch_matrix.S4BEG3 VPWR VGND sg13g2_mux4_1
X_3202_ net1164 net1105 Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q VPWR VGND sg13g2_dlhq_1
X_3133_ net1177 net1095 Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q VPWR VGND sg13g2_dlhq_1
X_3064_ net1186 net1084 Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q VPWR VGND sg13g2_dlhq_1
X_2015_ net991 Inst_RegFile_32x4.mem\[16\]\[0\] Inst_RegFile_32x4.mem\[17\]\[0\] Inst_RegFile_32x4.mem\[18\]\[0\]
+ Inst_RegFile_32x4.mem\[19\]\[0\] net945 _0505_ VPWR VGND sg13g2_mux4_1
X_2848_ UserCLK net482 _0006_ _2848_/Q_N Inst_RegFile_32x4.mem\[25\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_2917_ UserCLK net440 _0075_ _2917_/Q_N Inst_RegFile_32x4.mem\[21\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_2779_ net958 net839 _1118_ _0078_ VPWR VGND sg13g2_mux2_1
X_3350__394 VPWR VGND net394 sg13g2_tiehi
XFILLER_58_399 VPWR VGND sg13g2_fill_2
XFILLER_58_388 VPWR VGND sg13g2_decap_8
XFILLER_41_288 VPWR VGND sg13g2_decap_4
XFILLER_41_200 VPWR VGND sg13g2_fill_1
XFILLER_22_491 VPWR VGND sg13g2_fill_2
X_3751_ net103 net333 VPWR VGND sg13g2_buf_1
XFILLER_32_255 VPWR VGND sg13g2_fill_2
X_2702_ net728 net949 _1098_ _0021_ VPWR VGND sg13g2_mux2_1
Xoutput203 net203 FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
Xoutput247 net247 NN4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput258 net258 NN4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput236 net236 N4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput225 net225 N2BEGb[3] VPWR VGND sg13g2_buf_1
Xoutput214 net214 N2BEG[0] VPWR VGND sg13g2_buf_1
X_2564_ _1007_ _1006_ Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q Inst_RegFile_switch_matrix.NN4BEG1
+ VPWR VGND sg13g2_mux2_1
X_2495_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q _0432_ _0948_ _1155_
+ sg13g2_a21oi_1
XFILLER_4_60 VPWR VGND sg13g2_decap_4
X_1515_ VPWR _1137_ Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q VGND sg13g2_inv_1
Xoutput269 net269 S2BEG[3] VPWR VGND sg13g2_buf_1
X_2633_ Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q _0432_ _1051_ VPWR VGND sg13g2_nor2_1
X_3116_ net1150 net1095 Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q VPWR VGND sg13g2_dlhq_1
XFILLER_4_71 VPWR VGND sg13g2_decap_8
XFILLER_4_82 VPWR VGND sg13g2_fill_2
X_3047_ net1161 net1086 Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q VPWR VGND sg13g2_dlhq_1
XFILLER_46_358 VPWR VGND sg13g2_fill_1
X_2280_ VGND VPWR net55 net1049 _0752_ _0751_ sg13g2_a21oi_1
XFILLER_52_306 VPWR VGND sg13g2_fill_1
X_1995_ _0485_ _0484_ Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q VPWR VGND sg13g2_nand2b_1
X_3665_ NN4END[5] net253 VPWR VGND sg13g2_buf_1
X_2616_ _1030_ _1033_ _1034_ VPWR VGND sg13g2_nor2_1
X_3596_ net1187 net170 VPWR VGND sg13g2_buf_1
X_2547_ _0993_ _0992_ Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q Inst_RegFile_switch_matrix.EE4BEG0
+ VPWR VGND sg13g2_mux2_1
X_2478_ _0934_ _0933_ Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q Inst_RegFile_switch_matrix.WW4BEG0
+ VPWR VGND sg13g2_mux2_1
XFILLER_28_325 VPWR VGND sg13g2_fill_2
XFILLER_3_424 VPWR VGND sg13g2_fill_2
XFILLER_3_413 VPWR VGND sg13g2_fill_1
Xfanout1214 E6END[1] net1214 VPWR VGND sg13g2_buf_1
Xfanout1203 net1205 net1203 VPWR VGND sg13g2_buf_1
X_1780_ VGND VPWR Inst_RegFile_32x4.mem\[23\]\[1\] net923 _0282_ _0281_ sg13g2_a21oi_1
X_2401_ _0864_ VPWR _0865_ VGND net1051 net1011 sg13g2_o21ai_1
X_3381_ UserCLK net363 _0117_ _3381_/Q_N Inst_RegFile_32x4.mem\[10\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_27_2 VPWR VGND sg13g2_fill_1
X_2332_ _0800_ VPWR _0801_ VGND Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q _0797_ sg13g2_o21ai_1
X_2194_ VGND VPWR net1044 net1016 _0671_ Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q
+ sg13g2_a21oi_1
XFILLER_37_177 VPWR VGND sg13g2_fill_1
XFILLER_37_111 VPWR VGND sg13g2_fill_2
X_2263_ VPWR _0736_ _0735_ VGND sg13g2_inv_1
XFILLER_52_158 VPWR VGND sg13g2_fill_1
XFILLER_33_383 VPWR VGND sg13g2_fill_1
X_3717_ SS4END[5] net305 VPWR VGND sg13g2_buf_1
X_1978_ net1052 net971 _0469_ VPWR VGND sg13g2_nor2b_1
X_3579_ net1161 net183 VPWR VGND sg13g2_buf_1
X_3648_ N4END[4] net230 VPWR VGND sg13g2_buf_1
XFILLER_20_37 VPWR VGND sg13g2_fill_2
XFILLER_56_442 VPWR VGND sg13g2_decap_8
Xfanout1011 net1011 _1164_ VPWR VGND sg13g2_buf_16
Xfanout1022 net1025 net1022 VPWR VGND sg13g2_buf_1
Xfanout1033 net1034 net1033 VPWR VGND sg13g2_buf_1
Xfanout1044 Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q net1044 VPWR VGND sg13g2_buf_1
Xfanout1055 Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q net1055 VPWR VGND sg13g2_buf_1
Xfanout1077 net1081 net1077 VPWR VGND sg13g2_buf_1
Xfanout1099 net1102 net1099 VPWR VGND sg13g2_buf_1
Xfanout1088 net1092 net1088 VPWR VGND sg13g2_buf_1
Xfanout1066 net1067 net1066 VPWR VGND sg13g2_buf_1
X_1901_ _0393_ _0394_ _0395_ VPWR VGND sg13g2_nor2b_1
X_1832_ net924 Inst_RegFile_32x4.mem\[20\]\[3\] _0330_ VPWR VGND sg13g2_nor2b_1
X_2881_ UserCLK net449 _0039_ _2881_/Q_N Inst_RegFile_32x4.mem\[17\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_2950_ net1167 net1131 Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q VPWR VGND sg13g2_dlhq_1
X_1694_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q _0200_ _0198_ _0199_
+ sg13g2_a21oi_2
X_1763_ VGND VPWR net982 _0264_ _0265_ net969 sg13g2_a21oi_1
X_2315_ _0784_ _0783_ Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q _0785_ VPWR VGND
+ sg13g2_mux2_1
X_3295_ net1173 net1124 Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q VPWR VGND sg13g2_dlhq_1
X_3364_ UserCLK net380 _0100_ _3364_/Q_N Inst_RegFile_32x4.mem\[6\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_2246_ Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q net1076 net7 net36 net1216 net1040
+ _0720_ VPWR VGND sg13g2_mux4_1
XFILLER_53_423 VPWR VGND sg13g2_fill_2
X_2177_ Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q net1075 net37 net56 net8 Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q
+ _0655_ VPWR VGND sg13g2_mux4_1
XFILLER_40_117 VPWR VGND sg13g2_fill_1
XFILLER_33_180 VPWR VGND sg13g2_fill_1
XFILLER_31_14 VPWR VGND sg13g2_fill_2
XFILLER_21_397 VPWR VGND sg13g2_fill_2
XFILLER_56_99 VPWR VGND sg13g2_fill_2
XFILLER_44_423 VPWR VGND sg13g2_fill_1
Xinput103 W2MID[6] net103 VPWR VGND sg13g2_buf_1
XFILLER_31_139 VPWR VGND sg13g2_decap_8
XFILLER_12_397 VPWR VGND sg13g2_fill_2
X_2100_ Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q VPWR _0582_ VGND net1055 net986
+ sg13g2_o21ai_1
X_3080_ net1158 net1089 Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q VPWR VGND sg13g2_dlhq_1
XFILLER_50_415 VPWR VGND sg13g2_decap_8
X_2031_ _0519_ _0518_ net1005 VPWR VGND sg13g2_nand2b_1
X_1815_ net929 Inst_RegFile_32x4.mem\[10\]\[3\] Inst_RegFile_32x4.mem\[11\]\[3\] Inst_RegFile_32x4.mem\[8\]\[3\]
+ Inst_RegFile_32x4.mem\[9\]\[3\] net1027 _0313_ VPWR VGND sg13g2_mux4_1
X_2933_ net1195 net1128 Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q VPWR VGND sg13g2_dlhq_1
X_2795_ net932 net791 _1121_ _0091_ VPWR VGND sg13g2_mux2_1
X_2864_ UserCLK net466 _0022_ _2864_/Q_N Inst_RegFile_32x4.mem\[2\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
Xhold313 Inst_RegFile_32x4.mem\[9\]\[3\] VPWR VGND net811 sg13g2_dlygate4sd3_1
Xhold346 Inst_RegFile_32x4.mem\[24\]\[0\] VPWR VGND net844 sg13g2_dlygate4sd3_1
Xhold335 Inst_RegFile_32x4.mem\[11\]\[2\] VPWR VGND net833 sg13g2_dlygate4sd3_1
XFILLER_7_71 VPWR VGND sg13g2_fill_1
Xhold324 Inst_RegFile_32x4.mem\[17\]\[3\] VPWR VGND net822 sg13g2_dlygate4sd3_1
X_1677_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q _0183_ _0180_ _1144_
+ sg13g2_a21oi_2
Xhold302 Inst_RegFile_32x4.mem\[29\]\[1\] VPWR VGND net800 sg13g2_dlygate4sd3_1
X_1746_ _0248_ _0249_ net982 _0250_ VPWR VGND sg13g2_mux2_1
X_2229_ net1214 net65 net1058 _0704_ VPWR VGND sg13g2_mux2_1
X_3278_ net1211 net1123 Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q VPWR VGND sg13g2_dlhq_1
X_3347_ UserCLK net397 _0083_ _3347_/Q_N Inst_RegFile_32x4.mem\[29\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_41_426 VPWR VGND sg13g2_fill_1
XFILLER_26_69 VPWR VGND sg13g2_decap_4
XFILLER_5_338 VPWR VGND sg13g2_fill_2
XFILLER_12_194 VPWR VGND sg13g2_fill_2
X_1600_ net988 BD3 Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q _1220_ VPWR VGND sg13g2_mux2_1
X_1531_ VPWR _1153_ Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q VGND sg13g2_inv_1
X_2580_ Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q net1012 net512 _1018_ _1017_ Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q
+ Inst_RegFile_switch_matrix.W1BEG0 VPWR VGND sg13g2_mux4_1
X_3201_ net1168 net1105 Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q VPWR VGND sg13g2_dlhq_1
X_3132_ net1179 net1095 Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q VPWR VGND sg13g2_dlhq_1
X_3063_ net1191 net1087 Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q VPWR VGND sg13g2_dlhq_1
X_3339__405 VPWR VGND net405 sg13g2_tiehi
X_2014_ VGND VPWR _0459_ _0504_ _0503_ net1004 sg13g2_a21oi_2
XFILLER_50_289 VPWR VGND sg13g2_fill_1
X_2847_ UserCLK net483 _0005_ _2847_/Q_N Inst_RegFile_32x4.mem\[25\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_2778_ net949 net826 _1118_ _0077_ VPWR VGND sg13g2_mux2_1
XFILLER_12_49 VPWR VGND sg13g2_fill_1
X_2916_ UserCLK net406 _0074_ _2916_/Q_N Inst_RegFile_32x4.mem\[21\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_1729_ VGND VPWR _0231_ _0232_ _0233_ Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q
+ sg13g2_a21oi_1
XFILLER_58_367 VPWR VGND sg13g2_decap_8
XFILLER_37_24 VPWR VGND sg13g2_fill_2
XFILLER_41_223 VPWR VGND sg13g2_fill_2
XFILLER_26_286 VPWR VGND sg13g2_fill_1
XFILLER_49_389 VPWR VGND sg13g2_decap_4
X_2632_ VGND VPWR _1163_ Inst_RegFile_switch_matrix.JS2BEG0 _1050_ _1049_ sg13g2_a21oi_1
X_2701_ net738 net937 _1098_ _0020_ VPWR VGND sg13g2_mux2_1
X_3750_ net102 net332 VPWR VGND sg13g2_buf_1
Xoutput204 net204 FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
Xoutput215 net215 N2BEG[1] VPWR VGND sg13g2_buf_1
Xoutput259 net259 NN4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput237 net237 N4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput248 net248 NN4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput226 net226 N2BEGb[4] VPWR VGND sg13g2_buf_1
X_1514_ VPWR _1136_ Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q VGND sg13g2_inv_1
X_2563_ Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q net1073 net1218 net1068 net718
+ Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q _1007_ VPWR VGND sg13g2_mux4_1
X_2494_ _0947_ _0946_ Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q Inst_RegFile_switch_matrix.SS4BEG1
+ VPWR VGND sg13g2_mux2_2
X_3046_ net1167 net1086 Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q VPWR VGND sg13g2_dlhq_1
XFILLER_28_529 VPWR VGND sg13g2_fill_2
X_3115_ net1152 net1093 Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q VPWR VGND sg13g2_dlhq_1
XFILLER_46_337 VPWR VGND sg13g2_fill_2
XFILLER_46_326 VPWR VGND sg13g2_decap_8
XFILLER_14_212 VPWR VGND sg13g2_fill_2
XFILLER_49_175 VPWR VGND sg13g2_fill_2
XFILLER_49_120 VPWR VGND sg13g2_fill_1
X_1994_ Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q net15 net99 net72 Inst_RegFile_switch_matrix.E2BEG3
+ Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q _0484_ VPWR VGND sg13g2_mux4_1
XFILLER_20_226 VPWR VGND sg13g2_fill_1
X_3595_ net1191 net168 VPWR VGND sg13g2_buf_1
X_3664_ NN4END[4] net246 VPWR VGND sg13g2_buf_1
X_2615_ Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q _0895_ _0922_ _1031_ _1032_ Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q
+ _1033_ VPWR VGND sg13g2_mux4_1
X_2546_ Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q net1074 net1219 net60 net980 Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q
+ _0993_ VPWR VGND sg13g2_mux4_1
X_2477_ Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q net1074 net60 net1070 net978 Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q
+ _0934_ VPWR VGND sg13g2_mux4_1
X_3029_ net1194 net1078 Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q VPWR VGND sg13g2_dlhq_1
XFILLER_28_348 VPWR VGND sg13g2_fill_2
XFILLER_51_384 VPWR VGND sg13g2_decap_4
XFILLER_51_351 VPWR VGND sg13g2_fill_1
Xfanout1204 net1205 net1204 VPWR VGND sg13g2_buf_1
Xfanout1215 E6END[1] net1215 VPWR VGND sg13g2_buf_1
XFILLER_19_337 VPWR VGND sg13g2_fill_1
XFILLER_27_392 VPWR VGND sg13g2_fill_2
X_2400_ _0864_ net1051 net986 VPWR VGND sg13g2_nand2_1
XFILLER_6_274 VPWR VGND sg13g2_fill_1
X_3380_ UserCLK net364 _0116_ _3380_/Q_N Inst_RegFile_32x4.mem\[10\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_2331_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q _0799_ _0800_ Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q
+ sg13g2_a21oi_1
X_2262_ net1045 net64 net80 net91 net107 Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q
+ _0735_ VPWR VGND sg13g2_mux4_1
X_2193_ VGND VPWR _0670_ net1044 net105 sg13g2_or2_1
XFILLER_1_95 VPWR VGND sg13g2_fill_1
X_3716_ SS4END[4] net298 VPWR VGND sg13g2_buf_1
X_1977_ _0467_ VPWR _0468_ VGND Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q _0466_
+ sg13g2_o21ai_1
X_3647_ net49 net229 VPWR VGND sg13g2_buf_1
X_2529_ Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q net1033 net499 net500 _0978_ Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q
+ _0979_ VPWR VGND sg13g2_mux4_1
X_3578_ net1167 net180 VPWR VGND sg13g2_buf_1
XFILLER_56_421 VPWR VGND sg13g2_fill_1
XFILLER_28_156 VPWR VGND sg13g2_fill_1
XFILLER_28_123 VPWR VGND sg13g2_fill_2
XFILLER_29_69 VPWR VGND sg13g2_fill_2
XFILLER_29_58 VPWR VGND sg13g2_fill_2
XFILLER_43_148 VPWR VGND sg13g2_fill_2
XFILLER_43_104 VPWR VGND sg13g2_fill_2
Xfanout1001 net1002 net1001 VPWR VGND sg13g2_buf_1
Xfanout1012 net1012 net1014 VPWR VGND sg13g2_buf_16
Xfanout1034 BD0 net1034 VPWR VGND sg13g2_buf_1
Xfanout1056 net1057 net1056 VPWR VGND sg13g2_buf_1
Xfanout1023 net1024 net1023 VPWR VGND sg13g2_buf_1
Xfanout1045 Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q net1045 VPWR VGND sg13g2_buf_1
XFILLER_10_82 VPWR VGND sg13g2_fill_1
Xfanout1078 net1080 net1078 VPWR VGND sg13g2_buf_1
XFILLER_19_91 VPWR VGND sg13g2_fill_2
XFILLER_19_156 VPWR VGND sg13g2_fill_2
Xfanout1067 W6END[0] net1067 VPWR VGND sg13g2_buf_1
Xfanout1089 net1092 net1089 VPWR VGND sg13g2_buf_1
X_1900_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q _0390_ _0394_ Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q
+ sg13g2_a21oi_1
X_1831_ net921 Inst_RegFile_32x4.mem\[18\]\[3\] Inst_RegFile_32x4.mem\[19\]\[3\] Inst_RegFile_32x4.mem\[16\]\[3\]
+ Inst_RegFile_32x4.mem\[17\]\[3\] net1022 _0329_ VPWR VGND sg13g2_mux4_1
X_2880_ UserCLK net450 _0038_ _2880_/Q_N Inst_RegFile_32x4.mem\[17\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_1693_ _0199_ net973 Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q VPWR VGND sg13g2_nand2b_1
X_3363_ UserCLK net381 _0099_ _3363_/Q_N Inst_RegFile_32x4.mem\[5\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_1762_ net926 Inst_RegFile_32x4.mem\[14\]\[1\] Inst_RegFile_32x4.mem\[15\]\[1\] Inst_RegFile_32x4.mem\[12\]\[1\]
+ Inst_RegFile_32x4.mem\[13\]\[1\] net1024 _0264_ VPWR VGND sg13g2_mux4_1
X_2314_ Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q net1076 net1221 net34 net5 Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q
+ _0784_ VPWR VGND sg13g2_mux4_1
X_2176_ _0648_ _0653_ Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q _0654_ VPWR VGND
+ sg13g2_nand3_1
X_3294_ net1175 net1124 Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q VPWR VGND sg13g2_dlhq_1
X_2245_ _0713_ Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q _0718_ _0719_ VPWR VGND sg13g2_nand3_1
XFILLER_53_457 VPWR VGND sg13g2_decap_8
XFILLER_53_402 VPWR VGND sg13g2_decap_8
XFILLER_15_49 VPWR VGND sg13g2_fill_2
Xinput104 W2MID[7] net104 VPWR VGND sg13g2_buf_1
XFILLER_12_321 VPWR VGND sg13g2_fill_1
XFILLER_39_207 VPWR VGND sg13g2_fill_2
X_2030_ net991 Inst_RegFile_32x4.mem\[16\]\[1\] Inst_RegFile_32x4.mem\[17\]\[1\] Inst_RegFile_32x4.mem\[18\]\[1\]
+ Inst_RegFile_32x4.mem\[19\]\[1\] net945 _0518_ VPWR VGND sg13g2_mux4_1
X_2932_ net1196 net1130 Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q VPWR VGND sg13g2_dlhq_1
XFILLER_35_413 VPWR VGND sg13g2_fill_2
X_2907__415 VPWR VGND net415 sg13g2_tiehi
X_2863_ UserCLK net467 _0021_ _2863_/Q_N Inst_RegFile_32x4.mem\[2\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_2794_ net959 net780 _1121_ _0090_ VPWR VGND sg13g2_mux2_1
XFILLER_15_181 VPWR VGND sg13g2_fill_2
X_1814_ Inst_RegFile_32x4.AD_comb\[2\] Inst_RegFile_32x4.AD_reg\[2\] Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q
+ AD2 VPWR VGND sg13g2_mux2_2
X_1745_ net922 Inst_RegFile_32x4.mem\[30\]\[0\] Inst_RegFile_32x4.mem\[31\]\[0\] Inst_RegFile_32x4.mem\[28\]\[0\]
+ Inst_RegFile_32x4.mem\[29\]\[0\] net1025 _0249_ VPWR VGND sg13g2_mux4_1
Xhold325 Inst_RegFile_32x4.mem\[9\]\[2\] VPWR VGND net823 sg13g2_dlygate4sd3_1
Xhold336 Inst_RegFile_32x4.mem\[17\]\[1\] VPWR VGND net834 sg13g2_dlygate4sd3_1
X_2914__408 VPWR VGND net408 sg13g2_tiehi
Xhold303 Inst_RegFile_32x4.mem\[3\]\[1\] VPWR VGND net801 sg13g2_dlygate4sd3_1
Xhold347 Inst_RegFile_32x4.mem\[16\]\[1\] VPWR VGND net845 sg13g2_dlygate4sd3_1
X_3346_ UserCLK net398 _0082_ _3346_/Q_N Inst_RegFile_32x4.mem\[29\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_1676_ _0182_ Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q _0181_ VPWR VGND sg13g2_nand2_1
Xhold314 Inst_RegFile_32x4.mem\[28\]\[0\] VPWR VGND net812 sg13g2_dlygate4sd3_1
X_2228_ net92 net108 net1058 _0703_ VPWR VGND sg13g2_mux2_1
X_3277_ net1149 net1124 Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q VPWR VGND sg13g2_dlhq_1
X_2159_ VGND VPWR net8 Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q _0638_ _0637_ sg13g2_a21oi_1
XFILLER_44_298 VPWR VGND sg13g2_fill_1
XFILLER_8_188 VPWR VGND sg13g2_fill_2
X_3200_ net1171 net1105 Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q VPWR VGND sg13g2_dlhq_1
X_1530_ VPWR _1152_ Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q VGND sg13g2_inv_1
X_3062_ net1193 net1087 Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q VPWR VGND sg13g2_dlhq_1
XFILLER_35_210 VPWR VGND sg13g2_fill_2
X_3131_ net1180 net1093 Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q VPWR VGND sg13g2_dlhq_1
X_2013_ net992 Inst_RegFile_32x4.mem\[28\]\[0\] Inst_RegFile_32x4.mem\[29\]\[0\] Inst_RegFile_32x4.mem\[30\]\[0\]
+ Inst_RegFile_32x4.mem\[31\]\[0\] net946 _0503_ VPWR VGND sg13g2_mux4_1
XFILLER_23_427 VPWR VGND sg13g2_fill_2
XFILLER_23_405 VPWR VGND sg13g2_fill_2
X_2915_ UserCLK net407 _0073_ _2915_/Q_N Inst_RegFile_32x4.mem\[21\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_2846_ UserCLK net484 _0004_ _2846_/Q_N Inst_RegFile_32x4.mem\[25\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_1728_ VGND VPWR net63 Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q _0232_ Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q
+ sg13g2_a21oi_1
X_2777_ net939 net781 _1118_ _0076_ VPWR VGND sg13g2_mux2_1
XFILLER_58_324 VPWR VGND sg13g2_fill_1
X_3329_ net1169 net1144 Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q VPWR VGND sg13g2_dlhq_1
X_1659_ VGND VPWR _1144_ _0165_ _0166_ _1145_ sg13g2_a21oi_1
XFILLER_5_114 VPWR VGND sg13g2_fill_2
XFILLER_45_530 VPWR VGND sg13g2_fill_1
XFILLER_32_257 VPWR VGND sg13g2_fill_1
XFILLER_17_265 VPWR VGND sg13g2_fill_2
Xoutput205 net205 FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
Xoutput216 net216 N2BEG[2] VPWR VGND sg13g2_buf_1
X_2562_ Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q net986 _0895_ _0896_ _1207_ Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q
+ _1006_ VPWR VGND sg13g2_mux4_1
X_2904__418 VPWR VGND net418 sg13g2_tiehi
X_2631_ Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q Inst_RegFile_switch_matrix.JW2BEG0
+ _1049_ VPWR VGND sg13g2_and2_1
X_2700_ _1090_ _1097_ _1098_ VPWR VGND sg13g2_and2_2
Xoutput249 Inst_RegFile_switch_matrix.NN4BEG0 NN4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput238 net238 N4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput227 net227 N2BEGb[5] VPWR VGND sg13g2_buf_1
X_1513_ VPWR _1135_ Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q VGND sg13g2_inv_1
X_2493_ Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q net1073 net1218 net1069 net505
+ Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q _0947_ VPWR VGND sg13g2_mux4_1
X_3045_ net1188 net1086 Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q VPWR VGND sg13g2_dlhq_1
X_3114_ net1155 net1094 Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q VPWR VGND sg13g2_dlhq_1
XFILLER_23_38 VPWR VGND sg13g2_fill_2
X_2829_ net754 net953 _1129_ _0117_ VPWR VGND sg13g2_mux2_1
XFILLER_58_132 VPWR VGND sg13g2_fill_2
X_3732_ UserCLK net314 VPWR VGND sg13g2_buf_1
X_1993_ Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q _0165_ net516 Inst_RegFile_switch_matrix.JN2BEG6
+ Inst_RegFile_switch_matrix.JW2BEG6 Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q _0483_
+ VPWR VGND sg13g2_mux4_1
XFILLER_55_0 VPWR VGND sg13g2_decap_8
X_3594_ net1193 net167 VPWR VGND sg13g2_buf_1
X_2545_ Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q net1015 _0910_ _0911_ _0603_ Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q
+ _0992_ VPWR VGND sg13g2_mux4_1
X_3663_ Inst_RegFile_switch_matrix.N4BEG3 net236 VPWR VGND sg13g2_buf_1
X_2614_ Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q net55 net22 net79 Inst_RegFile_switch_matrix.JS2BEG2
+ Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q _1032_ VPWR VGND sg13g2_mux4_1
XFILLER_55_102 VPWR VGND sg13g2_fill_1
X_2476_ Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q net1013 _0910_ _0911_ _0408_ Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q
+ _0933_ VPWR VGND sg13g2_mux4_1
X_3028_ net1197 net1078 Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q VPWR VGND sg13g2_dlhq_1
XFILLER_50_58 VPWR VGND sg13g2_fill_1
XFILLER_50_36 VPWR VGND sg13g2_fill_1
XFILLER_50_14 VPWR VGND sg13g2_decap_8
Xfanout1216 E6END[0] net1216 VPWR VGND sg13g2_buf_1
Xfanout1205 FrameData[13] net1205 VPWR VGND sg13g2_buf_1
XFILLER_19_316 VPWR VGND sg13g2_fill_1
X_2192_ _0668_ VPWR _0669_ VGND net1044 net977 sg13g2_o21ai_1
X_2330_ VPWR _0799_ _0798_ VGND sg13g2_inv_1
X_2261_ Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q net36 net7 net1221 net1216 net1045
+ _0734_ VPWR VGND sg13g2_mux4_1
XFILLER_21_503 VPWR VGND sg13g2_fill_2
XFILLER_1_63 VPWR VGND sg13g2_fill_2
X_3342__402 VPWR VGND net402 sg13g2_tiehi
X_1976_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q _0464_ _0467_ Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q
+ sg13g2_a21oi_1
X_3715_ Inst_RegFile_switch_matrix.S4BEG3 net288 VPWR VGND sg13g2_buf_1
X_3646_ net48 net228 VPWR VGND sg13g2_buf_1
X_3577_ net1189 net169 VPWR VGND sg13g2_buf_1
X_2528_ Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q net40 net11 net85 net95 Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q
+ _0978_ VPWR VGND sg13g2_mux4_1
XFILLER_56_477 VPWR VGND sg13g2_fill_1
X_2459_ Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q net38 net66 net21 net93 Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q
+ _0919_ VPWR VGND sg13g2_mux4_1
Xfanout1002 net1003 net1002 VPWR VGND sg13g2_buf_1
Xfanout1013 net1013 net1014 VPWR VGND sg13g2_buf_16
Xfanout1068 net1069 net1068 VPWR VGND sg13g2_buf_1
Xfanout1079 net1080 net1079 VPWR VGND sg13g2_buf_1
Xfanout1057 Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q net1057 VPWR VGND sg13g2_buf_1
Xfanout1046 Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q net1046 VPWR VGND sg13g2_buf_1
Xfanout1024 net1025 net1024 VPWR VGND sg13g2_buf_1
X_1761_ _0263_ net956 _0262_ VPWR VGND sg13g2_nand2_1
X_1830_ VGND VPWR net982 _0327_ _0328_ net969 sg13g2_a21oi_1
X_1692_ _0198_ Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q net1032 VPWR VGND sg13g2_nand2_1
X_2313_ Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q net58 net62 net60 net1072 Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q
+ _0783_ VPWR VGND sg13g2_mux4_1
X_3362_ UserCLK net382 _0098_ _3362_/Q_N Inst_RegFile_32x4.mem\[5\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_2175_ _0652_ VPWR _0653_ VGND Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q _0650_ sg13g2_o21ai_1
X_3293_ net1177 net1124 Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q VPWR VGND sg13g2_dlhq_1
X_2244_ _0717_ _0715_ Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q _0718_ VPWR VGND sg13g2_nand3_1
XFILLER_53_436 VPWR VGND sg13g2_decap_4
XFILLER_21_355 VPWR VGND sg13g2_fill_2
X_1959_ Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q net59 net69 net61 net1068 Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q
+ _0451_ VPWR VGND sg13g2_mux4_1
XFILLER_21_399 VPWR VGND sg13g2_fill_1
XFILLER_29_400 VPWR VGND sg13g2_fill_2
Xinput105 W6END[1] net105 VPWR VGND sg13g2_buf_1
XFILLER_56_35 VPWR VGND sg13g2_fill_1
XFILLER_29_466 VPWR VGND sg13g2_fill_2
XFILLER_16_149 VPWR VGND sg13g2_decap_4
XFILLER_35_469 VPWR VGND sg13g2_fill_1
X_2931_ net1199 net1128 Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q VPWR VGND sg13g2_dlhq_1
X_1744_ net931 Inst_RegFile_32x4.mem\[26\]\[0\] Inst_RegFile_32x4.mem\[27\]\[0\] Inst_RegFile_32x4.mem\[24\]\[0\]
+ Inst_RegFile_32x4.mem\[25\]\[0\] net1028 _0248_ VPWR VGND sg13g2_mux4_1
X_2793_ net949 net801 _1121_ _0089_ VPWR VGND sg13g2_mux2_1
X_2862_ UserCLK net468 _0020_ _2862_/Q_N Inst_RegFile_32x4.mem\[2\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
Xhold304 Inst_RegFile_32x4.mem\[21\]\[2\] VPWR VGND net802 sg13g2_dlygate4sd3_1
X_1813_ VGND VPWR Inst_RegFile_32x4.AD_comb\[2\] _0299_ _0312_ sg13g2_or2_1
Xhold326 Inst_RegFile_32x4.mem\[31\]\[0\] VPWR VGND net824 sg13g2_dlygate4sd3_1
Xhold315 Inst_RegFile_32x4.mem\[12\]\[2\] VPWR VGND net813 sg13g2_dlygate4sd3_1
X_3276_ net1151 net1123 Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q VPWR VGND sg13g2_dlhq_1
Xhold337 Inst_RegFile_32x4.mem\[7\]\[0\] VPWR VGND net835 sg13g2_dlygate4sd3_1
Xhold348 Inst_RegFile_32x4.mem\[18\]\[2\] VPWR VGND net846 sg13g2_dlygate4sd3_1
X_1675_ Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q net43 net14 net71 net98 Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q
+ _0181_ VPWR VGND sg13g2_mux4_1
X_3345_ UserCLK net399 _0081_ _3345_/Q_N Inst_RegFile_32x4.mem\[29\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_2227_ Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q net37 net1220 net53 net8 net1058
+ _0702_ VPWR VGND sg13g2_mux4_1
X_2158_ Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q net53 _0637_ VPWR VGND sg13g2_nor2b_1
X_2089_ VGND VPWR Inst_RegFile_32x4.mem\[9\]\[2\] net994 _0573_ _0572_ sg13g2_a21oi_1
XFILLER_1_524 VPWR VGND sg13g2_fill_2
XFILLER_8_101 VPWR VGND sg13g2_fill_1
XFILLER_8_156 VPWR VGND sg13g2_fill_2
X_3130_ net1182 net1093 Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q VPWR VGND sg13g2_dlhq_1
XFILLER_4_351 VPWR VGND sg13g2_fill_2
X_2012_ _0501_ VPWR _0502_ VGND net1036 _0500_ sg13g2_o21ai_1
X_3061_ net1194 net1085 Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q VPWR VGND sg13g2_dlhq_1
X_2845_ UserCLK net485 _0003_ _2845_/Q_N Inst_RegFile_32x4.mem\[24\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_35_277 VPWR VGND sg13g2_decap_8
X_2914_ UserCLK net408 _0072_ _2914_/Q_N Inst_RegFile_32x4.mem\[21\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_1727_ _0231_ net35 Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q VPWR VGND sg13g2_nand2b_1
X_1658_ Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q net56 net6 net63 net90 Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q
+ _0165_ VPWR VGND sg13g2_mux4_1
X_2776_ _1118_ _1092_ _1106_ VPWR VGND sg13g2_nand2_2
X_3259_ net1181 net1120 Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q VPWR VGND sg13g2_dlhq_1
X_1589_ _1208_ Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q _1209_ VPWR VGND sg13g2_nor2b_1
X_3328_ net1170 net1146 Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q VPWR VGND sg13g2_dlhq_1
XFILLER_53_14 VPWR VGND sg13g2_decap_8
XFILLER_26_222 VPWR VGND sg13g2_fill_2
Xrebuffer220 net965 net718 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_57_380 VPWR VGND sg13g2_decap_8
Xoutput206 net206 FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
Xoutput239 net239 N4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput228 net228 N2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput217 net217 N2BEG[3] VPWR VGND sg13g2_buf_1
X_2561_ _1003_ _1005_ Inst_RegFile_switch_matrix.NN4BEG2 VPWR VGND sg13g2_nor2_1
X_1512_ VPWR _1134_ Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q VGND sg13g2_inv_1
X_2630_ _1048_ _1041_ _1046_ VPWR VGND sg13g2_nand2_1
X_2492_ Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q net985 _0895_ _0896_ _0165_ Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q
+ _0946_ VPWR VGND sg13g2_mux4_1
X_3113_ net1157 net1096 Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q VPWR VGND sg13g2_dlhq_1
X_3044_ net1213 net1087 Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q VPWR VGND sg13g2_dlhq_1
X_2828_ net759 net941 _1129_ _0116_ VPWR VGND sg13g2_mux2_1
XFILLER_48_14 VPWR VGND sg13g2_decap_8
X_2759_ net958 net846 _1114_ _0062_ VPWR VGND sg13g2_mux2_1
XFILLER_45_372 VPWR VGND sg13g2_fill_1
X_2910__412 VPWR VGND net412 sg13g2_tiehi
X_3731_ Inst_RegFile_switch_matrix.SS4BEG3 net304 VPWR VGND sg13g2_buf_1
X_3662_ Inst_RegFile_switch_matrix.N4BEG2 net235 VPWR VGND sg13g2_buf_1
X_1992_ _0475_ VPWR Inst_RegFile_switch_matrix.JN2BEG6 VGND Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q
+ _0482_ sg13g2_o21ai_1
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_3593_ net1195 net166 VPWR VGND sg13g2_buf_1
X_2544_ _0991_ _0990_ Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q Inst_RegFile_switch_matrix.EE4BEG1
+ VPWR VGND sg13g2_mux2_2
X_2613_ Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q net47 net18 net75 net102 Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q
+ _1031_ VPWR VGND sg13g2_mux4_1
X_2475_ _0932_ _0931_ Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q Inst_RegFile_switch_matrix.WW4BEG1
+ VPWR VGND sg13g2_mux2_1
XFILLER_51_320 VPWR VGND sg13g2_fill_2
X_3027_ net1199 net1078 Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q VPWR VGND sg13g2_dlhq_1
XFILLER_59_431 VPWR VGND sg13g2_fill_2
XFILLER_59_420 VPWR VGND sg13g2_decap_8
Xfanout1206 FrameData[12] net1206 VPWR VGND sg13g2_buf_1
Xfanout1217 E6END[0] net1217 VPWR VGND sg13g2_buf_1
XFILLER_46_147 VPWR VGND sg13g2_fill_2
XFILLER_42_353 VPWR VGND sg13g2_fill_1
XFILLER_41_7 VPWR VGND sg13g2_fill_2
X_2191_ _0668_ Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q net971 VPWR VGND sg13g2_nand2_1
XFILLER_37_125 VPWR VGND sg13g2_fill_1
X_2260_ Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q VPWR _0733_ VGND _0732_ _0729_ sg13g2_o21ai_1
XFILLER_52_128 VPWR VGND sg13g2_fill_2
X_3714_ Inst_RegFile_switch_matrix.S4BEG2 net287 VPWR VGND sg13g2_buf_1
X_1975_ VGND VPWR net1052 net506 _0466_ _0465_ sg13g2_a21oi_1
X_3645_ net47 net227 VPWR VGND sg13g2_buf_1
X_2527_ Inst_RegFile_switch_matrix.E6BEG0 _0975_ _0977_ _0970_ _1157_ VPWR VGND sg13g2_a22oi_1
X_2458_ Inst_RegFile_switch_matrix.W6BEG0 _0916_ _0918_ _0909_ _1152_ VPWR VGND sg13g2_a22oi_1
X_3576_ net1213 net158 VPWR VGND sg13g2_buf_1
XFILLER_29_38 VPWR VGND sg13g2_fill_1
XFILLER_56_456 VPWR VGND sg13g2_decap_8
XFILLER_43_106 VPWR VGND sg13g2_fill_1
XFILLER_28_147 VPWR VGND sg13g2_decap_8
XFILLER_28_125 VPWR VGND sg13g2_fill_1
X_2389_ VGND VPWR _0853_ _0854_ _0852_ Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q sg13g2_a21oi_2
XFILLER_16_309 VPWR VGND sg13g2_fill_2
X_2900__422 VPWR VGND net422 sg13g2_tiehi
Xfanout1003 BD3 net1003 VPWR VGND sg13g2_buf_2
Xfanout1058 Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q net1058 VPWR VGND sg13g2_buf_1
Xfanout1047 Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q net1047 VPWR VGND sg13g2_buf_1
Xfanout1014 net1014 BD1 VPWR VGND sg13g2_buf_16
Xfanout1036 _0367_ net1036 VPWR VGND sg13g2_buf_1
Xfanout1025 _1210_ net1025 VPWR VGND sg13g2_buf_1
Xfanout1069 W1END[3] net1069 VPWR VGND sg13g2_buf_1
XFILLER_35_81 VPWR VGND sg13g2_decap_4
XFILLER_30_301 VPWR VGND sg13g2_fill_1
XFILLER_19_93 VPWR VGND sg13g2_fill_1
XFILLER_19_158 VPWR VGND sg13g2_fill_1
X_1691_ VGND VPWR _0196_ Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q _0195_ Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q
+ _0197_ _0194_ sg13g2_a221oi_1
X_1760_ net929 Inst_RegFile_32x4.mem\[10\]\[1\] Inst_RegFile_32x4.mem\[11\]\[1\] Inst_RegFile_32x4.mem\[8\]\[1\]
+ Inst_RegFile_32x4.mem\[9\]\[1\] net1027 _0262_ VPWR VGND sg13g2_mux4_1
XFILLER_7_530 VPWR VGND sg13g2_fill_1
X_2312_ Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q VPWR _0782_ VGND _0778_ _0781_
+ sg13g2_o21ai_1
X_3292_ net1178 net1124 Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q VPWR VGND sg13g2_dlhq_1
X_3361_ UserCLK net383 _0097_ _3361_/Q_N Inst_RegFile_32x4.mem\[5\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_2174_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q _0651_ _0652_ _1147_ sg13g2_a21oi_1
X_2243_ _0716_ VPWR _0717_ VGND net1040 net1029 sg13g2_o21ai_1
X_1889_ _0384_ _0383_ Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q VPWR VGND sg13g2_nand2b_1
X_1958_ _0450_ _0449_ Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q VPWR VGND sg13g2_nand2b_1
X_3628_ Inst_RegFile_switch_matrix.N1BEG0 net210 VPWR VGND sg13g2_buf_8
XFILLER_56_14 VPWR VGND sg13g2_decap_8
Xinput106 WW4END[0] net106 VPWR VGND sg13g2_buf_1
XFILLER_44_448 VPWR VGND sg13g2_fill_2
XFILLER_4_522 VPWR VGND sg13g2_fill_2
XFILLER_47_220 VPWR VGND sg13g2_fill_1
XFILLER_11_8 VPWR VGND sg13g2_fill_2
X_2930_ net1202 net1128 Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q VPWR VGND sg13g2_dlhq_1
X_2861_ UserCLK net469 _0019_ _2861_/Q_N Inst_RegFile_32x4.mem\[28\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
Xhold327 Inst_RegFile_32x4.mem\[12\]\[0\] VPWR VGND net825 sg13g2_dlygate4sd3_1
Xhold305 Inst_RegFile_32x4.mem\[7\]\[2\] VPWR VGND net803 sg13g2_dlygate4sd3_1
X_1743_ _0247_ _0246_ _0241_ VPWR VGND sg13g2_nand2b_1
X_1812_ VGND VPWR net520 _0235_ _0311_ _0303_ _0312_ _0302_ sg13g2_a221oi_1
Xhold338 Inst_RegFile_32x4.mem\[18\]\[1\] VPWR VGND net836 sg13g2_dlygate4sd3_1
X_1674_ Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q net13 net97 net70 Inst_RegFile_switch_matrix.JW2BEG5
+ Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q _0180_ VPWR VGND sg13g2_mux4_1
Xhold316 Inst_RegFile_32x4.mem\[21\]\[3\] VPWR VGND net814 sg13g2_dlygate4sd3_1
X_2792_ net937 net792 _1121_ _0088_ VPWR VGND sg13g2_mux2_1
Xhold349 Inst_RegFile_32x4.mem\[23\]\[2\] VPWR VGND net847 sg13g2_dlygate4sd3_1
X_2226_ _0701_ Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q _0700_ VPWR VGND sg13g2_nand2_1
XFILLER_30_0 VPWR VGND sg13g2_fill_2
X_3275_ net1152 net1121 Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q VPWR VGND sg13g2_dlhq_1
X_3344_ UserCLK net400 _0080_ _3344_/Q_N Inst_RegFile_32x4.mem\[29\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_2088_ net994 Inst_RegFile_32x4.mem\[8\]\[2\] _0572_ VPWR VGND sg13g2_nor2b_1
XFILLER_38_242 VPWR VGND sg13g2_fill_1
X_2157_ net92 Inst_RegFile_switch_matrix.JN2BEG3 Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q
+ _0636_ VPWR VGND sg13g2_mux2_1
XFILLER_21_186 VPWR VGND sg13g2_decap_4
XFILLER_16_72 VPWR VGND sg13g2_fill_2
X_3060_ net1196 net1085 Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q VPWR VGND sg13g2_dlhq_1
X_2011_ VGND VPWR net1036 _0499_ _0501_ net1009 sg13g2_a21oi_1
XFILLER_35_212 VPWR VGND sg13g2_fill_1
X_2844_ UserCLK net486 _0002_ _2844_/Q_N Inst_RegFile_32x4.mem\[24\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_2913_ UserCLK net409 _0071_ _2913_/Q_N Inst_RegFile_32x4.mem\[20\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_16_481 VPWR VGND sg13g2_fill_2
X_1588_ Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q _1207_ _1208_ VPWR VGND sg13g2_nor2_1
X_1726_ _0228_ _0229_ Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q _0230_ VPWR VGND
+ sg13g2_mux2_1
X_2775_ net933 net814 _1117_ _0075_ VPWR VGND sg13g2_mux2_1
X_1657_ Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q VPWR _0164_ VGND Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q
+ _0163_ sg13g2_o21ai_1
X_3258_ net1183 net1120 Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q VPWR VGND sg13g2_dlhq_1
X_2209_ Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q VPWR _0685_ VGND _0679_ _0682_
+ sg13g2_o21ai_1
X_3189_ net1195 net1105 Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q VPWR VGND sg13g2_dlhq_1
X_3327_ net1173 net1144 Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q VPWR VGND sg13g2_dlhq_1
XFILLER_26_267 VPWR VGND sg13g2_fill_2
XFILLER_26_245 VPWR VGND sg13g2_fill_1
Xrebuffer221 net965 net719 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_5_116 VPWR VGND sg13g2_fill_1
XFILLER_17_267 VPWR VGND sg13g2_fill_1
XFILLER_40_292 VPWR VGND sg13g2_decap_4
Xoutput207 net207 FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
Xoutput218 net218 N2BEG[4] VPWR VGND sg13g2_buf_1
Xoutput229 net229 N2BEGb[7] VPWR VGND sg13g2_buf_1
X_2491_ _0943_ _0945_ Inst_RegFile_switch_matrix.SS4BEG2 VPWR VGND sg13g2_nor2_1
X_2560_ Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q _1004_ _1005_ VPWR VGND sg13g2_nor2_2
X_1511_ VPWR _1133_ Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q VGND sg13g2_inv_1
XFILLER_4_31 VPWR VGND sg13g2_fill_2
X_3043_ net1163 net1082 Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q VPWR VGND sg13g2_dlhq_1
XFILLER_4_64 VPWR VGND sg13g2_fill_2
XFILLER_4_53 VPWR VGND sg13g2_decap_8
X_3112_ net1159 net1096 Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q VPWR VGND sg13g2_dlhq_1
X_2827_ _1090_ _1101_ _1129_ VPWR VGND sg13g2_and2_2
XFILLER_31_292 VPWR VGND sg13g2_decap_8
X_2758_ net949 net836 _1114_ _0061_ VPWR VGND sg13g2_mux2_1
X_1709_ VGND VPWR _0214_ net1047 net1068 sg13g2_or2_1
X_2689_ net952 net794 _1093_ _0013_ VPWR VGND sg13g2_mux2_1
XFILLER_54_395 VPWR VGND sg13g2_decap_8
XFILLER_8_0 VPWR VGND sg13g2_fill_1
XFILLER_13_62 VPWR VGND sg13g2_fill_2
Xfanout990 net990 net992 VPWR VGND sg13g2_buf_16
XFILLER_45_362 VPWR VGND sg13g2_fill_2
X_3730_ Inst_RegFile_switch_matrix.SS4BEG2 net303 VPWR VGND sg13g2_buf_8
X_1991_ _0481_ VPWR _0482_ VGND Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q _0476_
+ sg13g2_o21ai_1
X_3592_ net1197 net165 VPWR VGND sg13g2_buf_1
X_3661_ Inst_RegFile_switch_matrix.N4BEG1 net234 VPWR VGND sg13g2_buf_1
X_2612_ _1030_ _1026_ _1029_ VPWR VGND sg13g2_nand2_1
X_2543_ Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q net1073 net1218 net61 net967 Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q
+ _0991_ VPWR VGND sg13g2_mux4_1
X_2878__452 VPWR VGND net452 sg13g2_tiehi
X_2474_ Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q net1073 net61 net1069 net504 Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q
+ _0932_ VPWR VGND sg13g2_mux4_1
X_3026_ net1201 net1078 Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q VPWR VGND sg13g2_dlhq_1
Xfanout1218 net4 net1218 VPWR VGND sg13g2_buf_1
Xfanout1207 FrameData[12] net1207 VPWR VGND sg13g2_buf_1
XFILLER_19_307 VPWR VGND sg13g2_fill_1
X_3335__444 VPWR VGND net444 sg13g2_tiehi
X_2190_ Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q VPWR _0667_ VGND _0662_ _0663_
+ sg13g2_o21ai_1
X_1974_ net1052 net1069 _0465_ VPWR VGND sg13g2_nor2b_1
X_3575_ Inst_RegFile_switch_matrix.EE4BEG3 net148 VPWR VGND sg13g2_buf_1
X_3713_ Inst_RegFile_switch_matrix.S4BEG1 net286 VPWR VGND sg13g2_buf_1
X_3644_ net46 net226 VPWR VGND sg13g2_buf_1
XFILLER_56_413 VPWR VGND sg13g2_fill_2
XFILLER_56_402 VPWR VGND sg13g2_decap_8
X_2526_ VGND VPWR _1157_ _0977_ _1156_ _0976_ sg13g2_a21oi_2
X_2457_ VGND VPWR _1151_ _0917_ _0918_ _1152_ sg13g2_a21oi_1
XFILLER_28_104 VPWR VGND sg13g2_fill_1
X_2388_ Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q VPWR _0853_ VGND Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q
+ _0851_ sg13g2_o21ai_1
XFILLER_56_435 VPWR VGND sg13g2_decap_8
X_3009_ net1168 net1138 Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q VPWR VGND sg13g2_dlhq_1
Xfanout1004 net1006 net1004 VPWR VGND sg13g2_buf_1
Xfanout1037 Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q net1037 VPWR VGND sg13g2_buf_1
Xfanout1026 net1028 net1026 VPWR VGND sg13g2_buf_1
Xfanout1015 net1015 BD1 VPWR VGND sg13g2_buf_16
Xfanout1048 Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q net1048 VPWR VGND sg13g2_buf_1
Xfanout1059 Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q net1059 VPWR VGND sg13g2_buf_1
XFILLER_42_184 VPWR VGND sg13g2_fill_1
X_2868__462 VPWR VGND net462 sg13g2_tiehi
X_1690_ VGND VPWR net1054 net1016 _0196_ Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q
+ sg13g2_a21oi_1
X_3291_ net1181 net1126 Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q VPWR VGND sg13g2_dlhq_1
X_2311_ Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q VPWR _0781_ VGND _0779_ _0780_
+ sg13g2_o21ai_1
XFILLER_32_4 VPWR VGND sg13g2_fill_2
X_3360_ UserCLK net384 _0096_ _3360_/Q_N Inst_RegFile_32x4.mem\[5\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_2875__455 VPWR VGND net455 sg13g2_tiehi
X_2242_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q _0716_ net1010 net1040
+ sg13g2_a21oi_2
XFILLER_53_416 VPWR VGND sg13g2_decap_8
X_2173_ net986 net1002 Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q _0651_ VPWR VGND
+ sg13g2_mux2_1
X_1957_ Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q net33 net41 net4 net12 Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q
+ _0449_ VPWR VGND sg13g2_mux4_1
X_2882__448 VPWR VGND net448 sg13g2_tiehi
XFILLER_21_357 VPWR VGND sg13g2_fill_1
X_3627_ FrameStrobe[19] net200 VPWR VGND sg13g2_buf_1
X_2509_ _0960_ net54 net1063 VPWR VGND sg13g2_nand2b_1
X_1888_ net61 net69 Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q _0383_ VPWR VGND sg13g2_mux2_1
Xinput107 WW4END[1] net107 VPWR VGND sg13g2_buf_1
XFILLER_16_129 VPWR VGND sg13g2_fill_2
XFILLER_8_339 VPWR VGND sg13g2_fill_2
XFILLER_46_92 VPWR VGND sg13g2_decap_4
XFILLER_30_121 VPWR VGND sg13g2_fill_2
X_2860_ UserCLK net470 _0018_ _2860_/Q_N Inst_RegFile_32x4.mem\[28\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_2791_ _1121_ _1092_ _1097_ VPWR VGND sg13g2_nand2_2
X_1811_ _0311_ _0309_ _0310_ _0304_ net955 VPWR VGND sg13g2_a22oi_1
XFILLER_15_151 VPWR VGND sg13g2_decap_8
X_1673_ Inst_RegFile_switch_matrix.JW2BEG5 _0177_ _0179_ _0174_ _0175_ VPWR VGND sg13g2_a22oi_1
Xhold306 Inst_RegFile_32x4.mem\[11\]\[0\] VPWR VGND net804 sg13g2_dlygate4sd3_1
X_1742_ _0245_ VPWR _0246_ VGND net1026 _0242_ sg13g2_o21ai_1
Xhold339 Inst_RegFile_32x4.mem\[18\]\[3\] VPWR VGND net837 sg13g2_dlygate4sd3_1
Xhold328 Inst_RegFile_32x4.mem\[19\]\[1\] VPWR VGND net826 sg13g2_dlygate4sd3_1
Xhold317 Inst_RegFile_32x4.mem\[21\]\[0\] VPWR VGND net815 sg13g2_dlygate4sd3_1
X_2225_ _0699_ VPWR _0700_ VGND Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q _0698_ sg13g2_o21ai_1
X_3343_ UserCLK net401 _0079_ _3343_/Q_N Inst_RegFile_32x4.mem\[19\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_3274_ net1154 net1121 Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q VPWR VGND sg13g2_dlhq_1
XFILLER_53_235 VPWR VGND sg13g2_fill_2
X_2087_ _0571_ net947 _0570_ VPWR VGND sg13g2_nand2_1
X_2156_ _0635_ VPWR Inst_RegFile_switch_matrix.JN2BEG3 VGND _0627_ _0626_ sg13g2_o21ai_1
X_2989_ net1148 net1140 Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q VPWR VGND sg13g2_dlhq_1
XFILLER_1_526 VPWR VGND sg13g2_fill_1
X_2858__472 VPWR VGND net472 sg13g2_tiehi
XFILLER_29_210 VPWR VGND sg13g2_fill_2
XFILLER_52_290 VPWR VGND sg13g2_fill_2
X_2865__465 VPWR VGND net465 sg13g2_tiehi
XFILLER_16_51 VPWR VGND sg13g2_fill_2
XFILLER_32_72 VPWR VGND sg13g2_decap_4
XFILLER_4_353 VPWR VGND sg13g2_fill_1
X_2872__458 VPWR VGND net458 sg13g2_tiehi
X_2010_ Inst_RegFile_32x4.mem\[26\]\[0\] Inst_RegFile_32x4.mem\[27\]\[0\] net998 _0500_
+ VPWR VGND sg13g2_mux2_1
X_2912_ UserCLK net410 _0070_ _2912_/Q_N Inst_RegFile_32x4.mem\[20\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_2843_ UserCLK net487 _0001_ _2843_/Q_N Inst_RegFile_32x4.mem\[24\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_2774_ net958 net802 _1117_ _0074_ VPWR VGND sg13g2_mux2_1
X_1725_ Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q net47 net18 net75 net102 Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q
+ _0229_ VPWR VGND sg13g2_mux4_1
X_1587_ Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q net37 net8 net65 net107 Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q
+ _1207_ VPWR VGND sg13g2_mux4_1
X_3326_ net1174 net1144 Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q VPWR VGND sg13g2_dlhq_1
X_1656_ net24 net78 Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q _0163_ VPWR VGND sg13g2_mux2_1
X_3257_ net1184 net1120 Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q VPWR VGND sg13g2_dlhq_1
X_2208_ Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q _0683_ _0684_ VPWR VGND sg13g2_nor2_1
X_3188_ net1196 net1105 Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q VPWR VGND sg13g2_dlhq_1
X_2139_ VGND VPWR net1056 net1018 _0619_ _0618_ sg13g2_a21oi_1
Xoutput208 net208 FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
X_2490_ Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q _0944_ _0945_ VPWR VGND sg13g2_nor2_1
Xoutput219 Inst_RegFile_switch_matrix.JN2BEG5 N2BEG[5] VPWR VGND sg13g2_buf_1
X_1510_ VPWR _1132_ Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q VGND sg13g2_inv_1
XFILLER_4_10 VPWR VGND sg13g2_fill_1
X_3111_ net1160 net1097 Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q VPWR VGND sg13g2_dlhq_1
X_3042_ net1165 net1082 Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q VPWR VGND sg13g2_dlhq_1
X_2848__482 VPWR VGND net482 sg13g2_tiehi
XFILLER_23_216 VPWR VGND sg13g2_decap_4
X_1708_ _0212_ VPWR _0213_ VGND Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q net976
+ sg13g2_o21ai_1
X_2688_ net942 net807 _1093_ _0012_ VPWR VGND sg13g2_mux2_1
X_2826_ net749 net932 _1128_ _0115_ VPWR VGND sg13g2_mux2_1
X_2757_ net938 net779 _1114_ _0060_ VPWR VGND sg13g2_mux2_1
X_3309_ net1149 net1145 Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q VPWR VGND sg13g2_dlhq_1
X_2855__475 VPWR VGND net475 sg13g2_tiehi
X_1639_ VGND VPWR _0147_ Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q net1067 sg13g2_or2_1
XFILLER_46_319 VPWR VGND sg13g2_decap_8
X_2862__468 VPWR VGND net468 sg13g2_tiehi
XFILLER_1_120 VPWR VGND sg13g2_fill_2
Xfanout980 AD1 net980 VPWR VGND sg13g2_buf_1
Xfanout991 net992 net991 VPWR VGND sg13g2_buf_1
X_1990_ _0480_ VPWR _0481_ VGND Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q _0479_
+ sg13g2_o21ai_1
X_2542_ Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q net988 _0895_ _0896_ _0641_ Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q
+ _0990_ VPWR VGND sg13g2_mux4_1
X_3591_ net1200 net164 VPWR VGND sg13g2_buf_1
X_3660_ Inst_RegFile_switch_matrix.N4BEG0 net233 VPWR VGND sg13g2_buf_1
X_2611_ Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q _1028_ _1018_ _0209_ _1027_ Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q
+ _1029_ VPWR VGND sg13g2_mux4_1
X_2473_ Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q net984 _0895_ _0896_ _0138_ Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q
+ _0931_ VPWR VGND sg13g2_mux4_1
XFILLER_51_322 VPWR VGND sg13g2_fill_1
X_3025_ net1203 net1079 Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q VPWR VGND sg13g2_dlhq_1
XFILLER_51_388 VPWR VGND sg13g2_fill_1
XFILLER_50_28 VPWR VGND sg13g2_decap_4
X_2809_ net746 net952 _1125_ _0101_ VPWR VGND sg13g2_mux2_1
Xfanout1219 net3 net1219 VPWR VGND sg13g2_buf_1
XFILLER_46_149 VPWR VGND sg13g2_fill_1
Xfanout1208 net1209 net1208 VPWR VGND sg13g2_buf_1
X_2845__485 VPWR VGND net485 sg13g2_tiehi
X_1973_ _0463_ VPWR _0464_ VGND net1052 net977 sg13g2_o21ai_1
X_3712_ Inst_RegFile_switch_matrix.S4BEG0 net285 VPWR VGND sg13g2_buf_1
XFILLER_53_0 VPWR VGND sg13g2_decap_8
X_2525_ Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q net1033 net988 net1015 net1003
+ net1064 _0976_ VPWR VGND sg13g2_mux4_1
X_3574_ Inst_RegFile_switch_matrix.EE4BEG2 net147 VPWR VGND sg13g2_buf_2
X_3643_ net45 net225 VPWR VGND sg13g2_buf_1
X_2852__478 VPWR VGND net478 sg13g2_tiehi
X_2456_ Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q net1031 net986 net1013 net1003
+ net1061 _0917_ VPWR VGND sg13g2_mux4_1
X_2387_ net984 net1001 Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q _0852_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_51_152 VPWR VGND sg13g2_fill_2
XFILLER_51_130 VPWR VGND sg13g2_fill_1
X_3008_ net1171 net1138 Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q VPWR VGND sg13g2_dlhq_1
Xfanout1016 _1166_ net1016 VPWR VGND sg13g2_buf_1
Xfanout1027 net1028 net1027 VPWR VGND sg13g2_buf_1
Xfanout1038 Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q net1038 VPWR VGND sg13g2_buf_1
Xfanout1005 net1005 net1006 VPWR VGND sg13g2_buf_16
XFILLER_3_248 VPWR VGND sg13g2_fill_1
XFILLER_19_127 VPWR VGND sg13g2_decap_4
Xfanout1049 Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q net1049 VPWR VGND sg13g2_buf_1
XFILLER_42_196 VPWR VGND sg13g2_fill_1
XFILLER_30_336 VPWR VGND sg13g2_fill_1
X_3290_ net1183 net1126 Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q VPWR VGND sg13g2_dlhq_1
X_2310_ Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q VPWR _0780_ VGND net1037 net1013
+ sg13g2_o21ai_1
X_2172_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q net1013 _0650_ _0649_
+ sg13g2_a21oi_1
X_2241_ net999 net1040 _0714_ _0715_ VPWR VGND sg13g2_a21o_1
XFILLER_38_458 VPWR VGND sg13g2_fill_2
XFILLER_18_160 VPWR VGND sg13g2_fill_1
XFILLER_18_182 VPWR VGND sg13g2_decap_8
X_1887_ net83 net1071 Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q _0382_ VPWR VGND
+ sg13g2_mux2_1
X_1956_ _0447_ Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q _0448_ VPWR VGND sg13g2_and2_1
X_3557_ E6END[11] net141 VPWR VGND sg13g2_buf_1
X_3626_ FrameStrobe[18] net199 VPWR VGND sg13g2_buf_1
X_2508_ Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q _0956_ _0957_ _0959_ _0958_ Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q
+ Inst_RegFile_switch_matrix.E6BEG1 VPWR VGND sg13g2_mux4_1
Xinput108 WW4END[2] net108 VPWR VGND sg13g2_buf_1
X_2439_ VGND VPWR net4 net1062 _0900_ Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q sg13g2_a21oi_1
XFILLER_16_108 VPWR VGND sg13g2_decap_4
XFILLER_24_185 VPWR VGND sg13g2_fill_2
XFILLER_4_524 VPWR VGND sg13g2_fill_1
XFILLER_46_71 VPWR VGND sg13g2_fill_1
X_1741_ VGND VPWR net1026 _0244_ _0245_ net956 sg13g2_a21oi_1
XFILLER_7_32 VPWR VGND sg13g2_fill_2
X_2790_ net932 net851 _1120_ _0087_ VPWR VGND sg13g2_mux2_1
X_1810_ VGND VPWR net1024 _0306_ _0310_ net955 sg13g2_a21oi_1
X_1672_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q _0178_ _0179_ Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q
+ sg13g2_a21oi_1
Xhold307 Inst_RegFile_32x4.mem\[24\]\[2\] VPWR VGND net805 sg13g2_dlygate4sd3_1
Xhold318 Inst_RegFile_32x4.mem\[12\]\[3\] VPWR VGND net816 sg13g2_dlygate4sd3_1
X_3342_ UserCLK net402 _0078_ _3342_/Q_N Inst_RegFile_32x4.mem\[19\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
Xhold329 Inst_RegFile_32x4.mem\[31\]\[1\] VPWR VGND net827 sg13g2_dlygate4sd3_1
X_3387__493 VPWR VGND net493 sg13g2_tiehi
X_2224_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q _0696_ _0699_ Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q
+ sg13g2_a21oi_1
X_2155_ _0634_ VPWR _0635_ VGND Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q _0633_
+ sg13g2_o21ai_1
X_3273_ net1156 net1121 Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q VPWR VGND sg13g2_dlhq_1
XFILLER_38_299 VPWR VGND sg13g2_fill_1
X_2086_ VGND VPWR Inst_RegFile_32x4.mem\[11\]\[2\] net994 _0570_ _0569_ sg13g2_a21oi_1
X_3609_ net1126 net201 VPWR VGND sg13g2_buf_1
X_2988_ net1150 net1140 Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q VPWR VGND sg13g2_dlhq_1
Xinput90 W2END[1] net90 VPWR VGND sg13g2_buf_1
X_1939_ Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q net35 net63 net24 net90 Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q
+ _0431_ VPWR VGND sg13g2_mux4_1
XFILLER_12_166 VPWR VGND sg13g2_fill_1
XFILLER_16_74 VPWR VGND sg13g2_fill_1
X_2911_ UserCLK net411 _0069_ _2911_/Q_N Inst_RegFile_32x4.mem\[20\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_16_483 VPWR VGND sg13g2_fill_1
X_2842_ UserCLK net439 _0000_ _2842_/Q_N Inst_RegFile_32x4.mem\[24\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_1724_ Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q net44 net72 net99 Inst_RegFile_switch_matrix.E2BEG6
+ Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q _0228_ VPWR VGND sg13g2_mux4_1
X_2773_ net951 net838 _1117_ _0073_ VPWR VGND sg13g2_mux2_1
X_3256_ net1187 net1120 Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q VPWR VGND sg13g2_dlhq_1
X_3325_ net1177 net1145 Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q VPWR VGND sg13g2_dlhq_1
X_1586_ _1202_ Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q _1205_ _1206_ VPWR VGND
+ sg13g2_a21o_1
X_1655_ VGND VPWR _0161_ _0162_ Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q Inst_RegFile_switch_matrix.JW2BEG3
+ sg13g2_a21oi_2
X_2207_ Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q net105 net1019 net980 net974 Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q
+ _0683_ VPWR VGND sg13g2_mux4_1
X_3187_ net1199 net1104 Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q VPWR VGND sg13g2_dlhq_1
X_2069_ VGND VPWR net1006 _0554_ _0555_ net943 sg13g2_a21oi_1
X_2138_ net1056 net1066 _0618_ VPWR VGND sg13g2_nor2b_1
Xrebuffer223 Inst_RegFile_switch_matrix.JN2BEG7 net721 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_57_394 VPWR VGND sg13g2_decap_8
Xoutput209 net209 FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
XFILLER_57_7 VPWR VGND sg13g2_decap_8
X_3110_ net1166 net1094 Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q VPWR VGND sg13g2_dlhq_1
X_3384__496 VPWR VGND net496 sg13g2_tiehi
X_3041_ net1169 net1082 Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q VPWR VGND sg13g2_dlhq_1
X_2825_ net742 net959 _1128_ _0114_ VPWR VGND sg13g2_mux2_1
X_1707_ _0212_ net1047 net966 VPWR VGND sg13g2_nand2_1
X_2687_ _1093_ _1092_ _1034_ VPWR VGND sg13g2_nand2_2
X_3391__489 VPWR VGND net489 sg13g2_tiehi
X_2756_ _1114_ _1090_ _1106_ VPWR VGND sg13g2_nand2_2
X_1638_ _0145_ VPWR _0146_ VGND net1039 net976 sg13g2_o21ai_1
XFILLER_48_28 VPWR VGND sg13g2_decap_4
X_3308_ net1150 net1145 Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q VPWR VGND sg13g2_dlhq_1
X_1569_ _1190_ net1048 net1012 VPWR VGND sg13g2_nand2_2
X_3239_ net1160 net1115 Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q VPWR VGND sg13g2_dlhq_1
XFILLER_6_405 VPWR VGND sg13g2_fill_2
XFILLER_6_449 VPWR VGND sg13g2_fill_2
XFILLER_10_489 VPWR VGND sg13g2_fill_2
XFILLER_1_143 VPWR VGND sg13g2_fill_2
Xfanout992 B_ADR0 net992 VPWR VGND sg13g2_buf_8
Xfanout970 net973 net970 VPWR VGND sg13g2_buf_1
XFILLER_45_364 VPWR VGND sg13g2_fill_1
X_2472_ _0928_ _0930_ Inst_RegFile_switch_matrix.WW4BEG2 VPWR VGND sg13g2_nor2_1
X_2541_ _0987_ _0989_ Inst_RegFile_switch_matrix.EE4BEG2 VPWR VGND sg13g2_nor2_1
X_3590_ net1202 net163 VPWR VGND sg13g2_buf_1
X_2610_ Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q net42 net97 net70 net524 Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q
+ _1028_ VPWR VGND sg13g2_mux4_1
X_3024_ net1206 net1078 Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q VPWR VGND sg13g2_dlhq_1
X_2808_ net724 net940 _1125_ _0100_ VPWR VGND sg13g2_mux2_1
Xfanout1209 FrameData[11] net1209 VPWR VGND sg13g2_buf_1
X_2739_ net958 net847 _1110_ _0046_ VPWR VGND sg13g2_mux2_1
XFILLER_27_375 VPWR VGND sg13g2_fill_2
XFILLER_10_242 VPWR VGND sg13g2_fill_1
X_3711_ S4END[15] net284 VPWR VGND sg13g2_buf_1
X_1972_ _0463_ net1053 net966 VPWR VGND sg13g2_nand2_1
X_3642_ net44 net224 VPWR VGND sg13g2_buf_1
X_2524_ _0974_ VPWR _0975_ VGND Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q _0971_
+ sg13g2_o21ai_1
XFILLER_46_0 VPWR VGND sg13g2_decap_8
X_2455_ _0915_ VPWR _0916_ VGND Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q _0912_
+ sg13g2_o21ai_1
XFILLER_56_426 VPWR VGND sg13g2_fill_1
X_2386_ VGND VPWR _0850_ _0851_ net1012 Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q
+ sg13g2_a21oi_2
X_3007_ net1172 net1138 Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q VPWR VGND sg13g2_dlhq_1
XFILLER_3_227 VPWR VGND sg13g2_fill_2
XFILLER_3_205 VPWR VGND sg13g2_fill_1
XFILLER_59_253 VPWR VGND sg13g2_fill_1
Xfanout1017 net1018 net1017 VPWR VGND sg13g2_buf_1
Xfanout1028 _1210_ net1028 VPWR VGND sg13g2_buf_1
Xfanout1006 net1006 net1007 VPWR VGND sg13g2_buf_16
Xfanout1039 Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q net1039 VPWR VGND sg13g2_buf_1
XFILLER_59_275 VPWR VGND sg13g2_fill_2
XFILLER_55_481 VPWR VGND sg13g2_fill_1
XFILLER_27_183 VPWR VGND sg13g2_fill_2
XFILLER_15_323 VPWR VGND sg13g2_fill_1
X_2171_ Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q net1031 _0649_ VPWR VGND sg13g2_nor2b_1
XFILLER_2_271 VPWR VGND sg13g2_fill_2
X_2240_ Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q VPWR _0714_ VGND net1040 net984
+ sg13g2_o21ai_1
XFILLER_53_429 VPWR VGND sg13g2_decap_8
X_3625_ FrameStrobe[17] net198 VPWR VGND sg13g2_buf_1
X_1886_ Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q net1073 net41 net1218 net12 Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q
+ _0381_ VPWR VGND sg13g2_mux4_1
X_1955_ _0447_ _0446_ Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q VPWR VGND sg13g2_nand2b_1
X_3556_ E6END[10] net140 VPWR VGND sg13g2_buf_1
X_2438_ _0899_ net55 net1062 VPWR VGND sg13g2_nand2b_1
X_2507_ Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q net1034 net989 net1015 net1003
+ Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q _0959_ VPWR VGND sg13g2_mux4_1
Xinput109 WW4END[3] net109 VPWR VGND sg13g2_buf_1
XFILLER_56_28 VPWR VGND sg13g2_decap_8
XFILLER_37_492 VPWR VGND sg13g2_fill_2
X_2369_ _0835_ VPWR Inst_RegFile_switch_matrix.JS2BEG0 VGND _0827_ _0826_ sg13g2_o21ai_1
XFILLER_52_462 VPWR VGND sg13g2_decap_8
XFILLER_52_440 VPWR VGND sg13g2_decap_8
X_2898__424 VPWR VGND net424 sg13g2_tiehi
XFILLER_21_20 VPWR VGND sg13g2_fill_1
XFILLER_47_289 VPWR VGND sg13g2_decap_8
XFILLER_46_61 VPWR VGND sg13g2_decap_4
XFILLER_30_112 VPWR VGND sg13g2_fill_1
X_1671_ Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q net58 net68 net60 net1070 Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q
+ _0178_ VPWR VGND sg13g2_mux4_1
X_1740_ VGND VPWR Inst_RegFile_32x4.mem\[5\]\[0\] net930 _0244_ _0243_ sg13g2_a21oi_1
XFILLER_30_123 VPWR VGND sg13g2_fill_1
Xhold308 Inst_RegFile_32x4.mem\[14\]\[1\] VPWR VGND net806 sg13g2_dlygate4sd3_1
Xhold319 Inst_RegFile_32x4.mem\[20\]\[3\] VPWR VGND net817 sg13g2_dlygate4sd3_1
X_3272_ net1158 net1121 Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q VPWR VGND sg13g2_dlhq_1
X_3341_ UserCLK net403 _0077_ _3341_/Q_N Inst_RegFile_32x4.mem\[19\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_2223_ VGND VPWR net1058 net1019 _0698_ _0697_ sg13g2_a21oi_1
X_2085_ net994 Inst_RegFile_32x4.mem\[10\]\[2\] _0569_ VPWR VGND sg13g2_nor2b_1
XFILLER_38_278 VPWR VGND sg13g2_decap_4
X_2154_ Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q _0632_ _0634_ VPWR VGND sg13g2_nor2_1
XFILLER_34_473 VPWR VGND sg13g2_fill_2
X_2987_ net1152 net1137 Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q VPWR VGND sg13g2_dlhq_1
XFILLER_21_145 VPWR VGND sg13g2_fill_1
Xinput80 S4END[2] net80 VPWR VGND sg13g2_buf_1
X_3608_ net1144 net190 VPWR VGND sg13g2_buf_1
X_1869_ Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q _0362_ _0364_ VPWR VGND sg13g2_nor2_1
Xinput91 W2END[2] net91 VPWR VGND sg13g2_buf_1
X_1938_ _0429_ _0430_ VPWR VGND sg13g2_inv_4
X_3539_ Inst_RegFile_switch_matrix.E2BEG7 net121 VPWR VGND sg13g2_buf_2
XFILLER_57_510 VPWR VGND sg13g2_fill_1
XFILLER_12_101 VPWR VGND sg13g2_decap_4
XFILLER_32_41 VPWR VGND sg13g2_decap_8
XFILLER_35_226 VPWR VGND sg13g2_fill_1
XFILLER_43_281 VPWR VGND sg13g2_fill_2
X_2841_ net934 net816 _1131_ _0127_ VPWR VGND sg13g2_mux2_1
X_2910_ UserCLK net412 _0068_ _2910_/Q_N Inst_RegFile_32x4.mem\[20\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_1723_ _0227_ VPWR Inst_RegFile_switch_matrix.E2BEG6 VGND _0223_ _0216_ sg13g2_o21ai_1
X_1654_ Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q VPWR _0161_ VGND _1138_ Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q
+ sg13g2_o21ai_1
X_2772_ net939 net815 _1117_ _0072_ VPWR VGND sg13g2_mux2_1
X_2206_ Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q VPWR _0682_ VGND Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q
+ _0681_ sg13g2_o21ai_1
X_3324_ net1179 net1145 Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q VPWR VGND sg13g2_dlhq_1
X_3255_ net1191 net1117 Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q VPWR VGND sg13g2_dlhq_1
X_1585_ Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q VPWR _1205_ VGND Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q
+ _1204_ sg13g2_o21ai_1
XFILLER_41_218 VPWR VGND sg13g2_fill_1
X_2068_ net991 Inst_RegFile_32x4.mem\[4\]\[3\] Inst_RegFile_32x4.mem\[5\]\[3\] Inst_RegFile_32x4.mem\[6\]\[3\]
+ Inst_RegFile_32x4.mem\[7\]\[3\] net947 _0554_ VPWR VGND sg13g2_mux4_1
X_3186_ net1202 net1104 Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q VPWR VGND sg13g2_dlhq_1
X_2137_ _0616_ VPWR _0617_ VGND net1056 net976 sg13g2_o21ai_1
X_2888__434 VPWR VGND net434 sg13g2_tiehi
XFILLER_34_292 VPWR VGND sg13g2_fill_2
XFILLER_5_108 VPWR VGND sg13g2_fill_1
Xrebuffer224 Inst_RegFile_switch_matrix.JW2BEG6 net722 VPWR VGND sg13g2_dlygate4sd1_1
X_2895__427 VPWR VGND net427 sg13g2_tiehi
XFILLER_57_373 VPWR VGND sg13g2_decap_8
XFILLER_27_96 VPWR VGND sg13g2_fill_2
XFILLER_25_292 VPWR VGND sg13g2_fill_1
XFILLER_13_421 VPWR VGND sg13g2_fill_1
X_3338__488 VPWR VGND net488 sg13g2_tiehi
XFILLER_9_458 VPWR VGND sg13g2_fill_1
XFILLER_4_78 VPWR VGND sg13g2_decap_4
X_3040_ net1170 net1082 Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q VPWR VGND sg13g2_dlhq_1
X_2824_ net735 net949 _1128_ _0113_ VPWR VGND sg13g2_mux2_1
X_2686_ _1047_ _1060_ _1058_ _1092_ VPWR VGND sg13g2_nor3_2
X_1706_ _0211_ Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q _0210_ VPWR VGND sg13g2_nand2_1
X_2755_ net932 net818 _1113_ _0059_ VPWR VGND sg13g2_mux2_1
X_1637_ _0145_ net1039 net963 VPWR VGND sg13g2_nand2_1
X_3169_ net1168 net1101 Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q VPWR VGND sg13g2_dlhq_1
X_1568_ VGND VPWR _1188_ Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q _1187_ Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q
+ _1189_ _1186_ sg13g2_a221oi_1
X_3307_ net1152 net1142 Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q VPWR VGND sg13g2_dlhq_1
X_3238_ net1166 net1115 Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q VPWR VGND sg13g2_dlhq_1
XFILLER_10_446 VPWR VGND sg13g2_fill_2
Xfanout960 net962 net960 VPWR VGND sg13g2_buf_1
Xfanout971 net972 net971 VPWR VGND sg13g2_buf_1
XFILLER_45_332 VPWR VGND sg13g2_decap_4
Xfanout993 net996 net993 VPWR VGND sg13g2_buf_1
Xfanout982 net982 net983 VPWR VGND sg13g2_buf_16
XFILLER_9_244 VPWR VGND sg13g2_fill_1
X_2471_ Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q _0929_ _0930_ VPWR VGND sg13g2_nor2_1
X_2540_ Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q _0988_ _0989_ VPWR VGND sg13g2_nor2_1
X_3390__490 VPWR VGND net490 sg13g2_tiehi
X_3023_ net1208 net1077 Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q VPWR VGND sg13g2_dlhq_1
XFILLER_51_313 VPWR VGND sg13g2_decap_8
XFILLER_51_302 VPWR VGND sg13g2_fill_2
X_2885__437 VPWR VGND net437 sg13g2_tiehi
X_2807_ _1090_ _1122_ _1125_ VPWR VGND sg13g2_and2_1
X_2738_ net951 net832 _1110_ _0045_ VPWR VGND sg13g2_mux2_1
XFILLER_59_413 VPWR VGND sg13g2_decap_8
X_2669_ Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q VPWR _1084_ VGND Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q
+ _1082_ sg13g2_o21ai_1
XFILLER_42_324 VPWR VGND sg13g2_fill_1
XFILLER_10_221 VPWR VGND sg13g2_fill_2
XFILLER_6_0 VPWR VGND sg13g2_fill_2
XFILLER_33_346 VPWR VGND sg13g2_fill_2
X_3710_ S4END[14] net283 VPWR VGND sg13g2_buf_1
X_1971_ _0462_ _0461_ net1008 _0412_ _0371_ VPWR VGND sg13g2_a22oi_1
X_3641_ net43 net223 VPWR VGND sg13g2_buf_1
X_2523_ _1156_ _0973_ _0974_ VPWR VGND sg13g2_nor2_1
X_2454_ _1151_ _0914_ _0915_ VPWR VGND sg13g2_nor2_1
XFILLER_39_0 VPWR VGND sg13g2_decap_4
X_2385_ Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q net1030 _0850_ VPWR VGND sg13g2_nor2b_1
XFILLER_56_449 VPWR VGND sg13g2_decap_8
X_3006_ net1175 net1138 Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q VPWR VGND sg13g2_dlhq_1
Xinput1 E1END[0] net1 VPWR VGND sg13g2_buf_1
XFILLER_10_55 VPWR VGND sg13g2_fill_2
Xfanout1018 net1018 AD0 VPWR VGND sg13g2_buf_16
Xfanout1007 _0409_ net1007 VPWR VGND sg13g2_buf_8
Xoutput360 net360 WW4BEG[7] VPWR VGND sg13g2_buf_1
Xfanout1029 net1030 net1029 VPWR VGND sg13g2_buf_1
XFILLER_19_107 VPWR VGND sg13g2_fill_2
XFILLER_51_62 VPWR VGND sg13g2_fill_1
XFILLER_7_501 VPWR VGND sg13g2_fill_2
X_2170_ _0648_ _1147_ _0647_ VPWR VGND sg13g2_nand2b_1
X_1954_ Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q net107 net1017 net515 net967 Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q
+ _0446_ VPWR VGND sg13g2_mux4_1
X_3555_ E6END[9] net139 VPWR VGND sg13g2_buf_1
X_3624_ FrameStrobe[16] net197 VPWR VGND sg13g2_buf_1
X_1885_ Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q VPWR _0380_ VGND _0379_ _0376_
+ sg13g2_o21ai_1
X_2506_ Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q _0896_ _0895_ net499 net500 Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q
+ _0958_ VPWR VGND sg13g2_mux4_1
X_2437_ Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q _0893_ _0894_ _0898_ _0897_ Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q
+ Inst_RegFile_switch_matrix.W6BEG1 VPWR VGND sg13g2_mux4_1
X_2368_ _0834_ VPWR _0835_ VGND Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q _0828_ sg13g2_o21ai_1
X_2299_ _0769_ VPWR _0770_ VGND Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q _0766_ sg13g2_o21ai_1
XFILLER_21_76 VPWR VGND sg13g2_fill_2
Xoutput190 net190 FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
X_1670_ _0177_ _0176_ Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q VPWR VGND sg13g2_nand2b_1
Xhold309 Inst_RegFile_32x4.mem\[27\]\[0\] VPWR VGND net807 sg13g2_dlygate4sd3_1
X_2222_ net1058 net1065 _0697_ VPWR VGND sg13g2_nor2b_1
X_3271_ net1160 net1121 Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q VPWR VGND sg13g2_dlhq_1
X_3340_ UserCLK net404 _0076_ _3340_/Q_N Inst_RegFile_32x4.mem\[19\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_2084_ VGND VPWR _0567_ net532 _0565_ _0561_ _0568_ _0563_ sg13g2_a221oi_1
X_2153_ net1056 net38 net50 net1219 net9 Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q
+ _0633_ VPWR VGND sg13g2_mux4_1
X_1937_ Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q net54 net1216 net89 Inst_RegFile_switch_matrix.JW2BEG4
+ Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q _0429_ VPWR VGND sg13g2_mux4_1
X_2986_ net1154 net1137 Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q VPWR VGND sg13g2_dlhq_1
X_3607_ net1163 net182 VPWR VGND sg13g2_buf_1
Xinput81 S4END[3] net81 VPWR VGND sg13g2_buf_1
Xinput70 S2MID[0] net70 VPWR VGND sg13g2_buf_1
X_1868_ VPWR _0363_ _0362_ VGND sg13g2_inv_1
X_3538_ Inst_RegFile_switch_matrix.E2BEG6 net120 VPWR VGND sg13g2_buf_1
Xinput92 W2END[3] net92 VPWR VGND sg13g2_buf_1
X_1799_ VGND VPWR net520 _0236_ _0298_ _0288_ _0299_ _0290_ sg13g2_a221oi_1
XFILLER_16_21 VPWR VGND sg13g2_fill_2
X_2840_ net960 net813 _1131_ _0126_ VPWR VGND sg13g2_mux2_1
X_2771_ _1117_ _1108_ _1088_ VPWR VGND sg13g2_nand2_2
X_1722_ _0227_ _0226_ Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q VPWR VGND sg13g2_nand2b_1
X_1584_ VGND VPWR net7 Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q _1204_ _1203_ sg13g2_a21oi_1
X_1653_ _0160_ VPWR Inst_RegFile_switch_matrix.JW2BEG3 VGND _0156_ _0149_ sg13g2_o21ai_1
X_2205_ VGND VPWR _0680_ _0681_ net1015 Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q
+ sg13g2_a21oi_2
X_3254_ net1193 net1117 Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q VPWR VGND sg13g2_dlhq_1
Xfanout1190 net1191 net1190 VPWR VGND sg13g2_buf_1
X_3185_ net1203 net1104 Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q VPWR VGND sg13g2_dlhq_1
X_3323_ net1180 net1142 Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q VPWR VGND sg13g2_dlhq_1
XFILLER_21_0 VPWR VGND sg13g2_fill_2
X_2067_ _0553_ _0552_ net1004 VPWR VGND sg13g2_nand2b_1
X_2136_ _0616_ net1057 net963 VPWR VGND sg13g2_nand2_1
Xrebuffer225 Inst_RegFile_switch_matrix.E2BEG5 net723 VPWR VGND sg13g2_dlygate4sd1_1
X_2969_ net1184 net1133 Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q VPWR VGND sg13g2_dlhq_1
XFILLER_40_296 VPWR VGND sg13g2_fill_2
XFILLER_40_285 VPWR VGND sg13g2_decap_8
XFILLER_40_263 VPWR VGND sg13g2_fill_1
XFILLER_48_374 VPWR VGND sg13g2_fill_2
XFILLER_31_285 VPWR VGND sg13g2_fill_2
X_1705_ Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q Inst_RegFile_switch_matrix.JS2BEG5
+ Inst_RegFile_switch_matrix.JW2BEG5 _0209_ Inst_RegFile_switch_matrix.JN2BEG5 _1146_
+ _0210_ VPWR VGND sg13g2_mux4_1
X_2754_ net958 net848 _1113_ _0058_ VPWR VGND sg13g2_mux2_1
XFILLER_8_481 VPWR VGND sg13g2_fill_2
X_2823_ net739 net937 _1128_ _0112_ VPWR VGND sg13g2_mux2_1
X_1636_ VGND VPWR _1214_ net983 _1213_ net1027 _0144_ _1212_ sg13g2_a221oi_1
X_2685_ net935 net744 _1091_ _0011_ VPWR VGND sg13g2_mux2_1
X_1567_ VGND VPWR net1048 net1016 _1188_ Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q
+ sg13g2_a21oi_1
X_3306_ net1154 net1142 Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q VPWR VGND sg13g2_dlhq_1
X_2119_ VGND VPWR net21 Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q _0600_ _0599_ sg13g2_a21oi_1
X_3168_ net1171 net1101 Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q VPWR VGND sg13g2_dlhq_1
X_3237_ net1188 net1115 Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q VPWR VGND sg13g2_dlhq_1
X_3099_ net1180 net1088 Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q VPWR VGND sg13g2_dlhq_1
XFILLER_6_407 VPWR VGND sg13g2_fill_1
XFILLER_10_469 VPWR VGND sg13g2_fill_1
Xfanout972 net973 net972 VPWR VGND sg13g2_buf_1
Xfanout994 net996 net994 VPWR VGND sg13g2_buf_1
XFILLER_38_41 VPWR VGND sg13g2_decap_8
Xfanout961 net962 net961 VPWR VGND sg13g2_buf_1
Xfanout983 _0142_ net983 VPWR VGND sg13g2_buf_8
Xfanout950 net951 net950 VPWR VGND sg13g2_buf_1
XFILLER_57_193 VPWR VGND sg13g2_fill_2
XFILLER_38_74 VPWR VGND sg13g2_fill_1
XFILLER_13_285 VPWR VGND sg13g2_fill_1
X_2470_ Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q net1076 net58 net1072 net972 Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q
+ _0929_ VPWR VGND sg13g2_mux4_1
XFILLER_55_108 VPWR VGND sg13g2_fill_1
XFILLER_48_160 VPWR VGND sg13g2_fill_1
X_3022_ net1211 net1077 Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q VPWR VGND sg13g2_dlhq_1
XFILLER_36_355 VPWR VGND sg13g2_fill_2
X_2806_ net934 net797 _1124_ _0099_ VPWR VGND sg13g2_mux2_1
X_2668_ net71 net98 Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q _1083_ VPWR VGND sg13g2_mux2_1
X_2737_ net939 net841 _1110_ _0044_ VPWR VGND sg13g2_mux2_1
X_2599_ Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q net970 _0645_ Inst_RegFile_switch_matrix.JW2BEG0
+ net502 Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q Inst_RegFile_switch_matrix.N1BEG1
+ VPWR VGND sg13g2_mux4_1
X_1619_ net985 net1001 Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q _0128_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_27_377 VPWR VGND sg13g2_fill_1
XFILLER_15_528 VPWR VGND sg13g2_fill_2
XFILLER_50_380 VPWR VGND sg13g2_fill_1
XFILLER_24_65 VPWR VGND sg13g2_fill_1
XFILLER_24_10 VPWR VGND sg13g2_fill_1
XFILLER_6_226 VPWR VGND sg13g2_fill_2
XFILLER_10_266 VPWR VGND sg13g2_fill_1
XFILLER_58_491 VPWR VGND sg13g2_fill_1
XFILLER_1_69 VPWR VGND sg13g2_fill_2
X_1970_ net997 Inst_RegFile_32x4.mem\[12\]\[0\] Inst_RegFile_32x4.mem\[13\]\[0\] Inst_RegFile_32x4.mem\[14\]\[0\]
+ Inst_RegFile_32x4.mem\[15\]\[0\] net947 _0461_ VPWR VGND sg13g2_mux4_1
XFILLER_33_336 VPWR VGND sg13g2_fill_1
X_3571_ EE4END[15] net144 VPWR VGND sg13g2_buf_1
X_2522_ VGND VPWR net1063 _0338_ _0973_ _0972_ sg13g2_a21oi_1
X_3640_ net42 net222 VPWR VGND sg13g2_buf_1
X_2453_ VGND VPWR net1062 _0338_ _0914_ _0913_ sg13g2_a21oi_1
X_2891__431 VPWR VGND net431 sg13g2_tiehi
X_2384_ Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q net1065 net504 net979 net970 Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q
+ _0849_ VPWR VGND sg13g2_mux4_1
X_3005_ net1176 net1138 Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q VPWR VGND sg13g2_dlhq_1
Xinput2 net2 E1END[1] VPWR VGND sg13g2_buf_16
Xoutput361 net361 WW4BEG[8] VPWR VGND sg13g2_buf_1
X_3769_ WW4END[8] net357 VPWR VGND sg13g2_buf_1
Xoutput350 net350 WW4BEG[12] VPWR VGND sg13g2_buf_1
Xfanout1019 net1020 net1019 VPWR VGND sg13g2_buf_1
Xfanout1008 net1009 net1008 VPWR VGND sg13g2_buf_1
XFILLER_55_472 VPWR VGND sg13g2_decap_8
XFILLER_15_303 VPWR VGND sg13g2_fill_1
XFILLER_53_409 VPWR VGND sg13g2_decap_8
XFILLER_18_130 VPWR VGND sg13g2_decap_4
X_1884_ _0378_ Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q _1136_ _0379_ VPWR VGND
+ sg13g2_a21o_1
X_1953_ _0444_ _0441_ Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q _0445_ VPWR VGND
+ sg13g2_nand3_1
X_3554_ E6END[8] net138 VPWR VGND sg13g2_buf_1
X_3623_ FrameStrobe[15] net196 VPWR VGND sg13g2_buf_1
XFILLER_51_0 VPWR VGND sg13g2_decap_8
X_2505_ Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q net1020 net967 net980 net974 Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q
+ _0957_ VPWR VGND sg13g2_mux4_1
X_2436_ Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q net1031 net987 net1012 net1001
+ Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q _0898_ VPWR VGND sg13g2_mux4_1
X_2298_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q _0768_ _0769_ Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q
+ sg13g2_a21oi_1
X_2367_ Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q _0833_ _0834_ VPWR VGND sg13g2_nor2_1
XFILLER_37_494 VPWR VGND sg13g2_fill_1
XFILLER_24_166 VPWR VGND sg13g2_decap_8
Xoutput180 net180 FrameData_O[2] VPWR VGND sg13g2_buf_1
Xoutput191 net191 FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
XFILLER_46_96 VPWR VGND sg13g2_fill_2
XFILLER_30_158 VPWR VGND sg13g2_fill_2
XFILLER_15_111 VPWR VGND sg13g2_fill_2
XFILLER_7_57 VPWR VGND sg13g2_fill_2
X_2221_ net980 net974 net1058 _0696_ VPWR VGND sg13g2_mux2_1
X_2152_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q _0630_ _0632_ _0631_
+ sg13g2_a21oi_1
X_3270_ net1166 net1121 Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q VPWR VGND sg13g2_dlhq_1
XFILLER_34_475 VPWR VGND sg13g2_fill_1
XFILLER_34_453 VPWR VGND sg13g2_fill_2
X_2083_ VGND VPWR net1004 _0566_ _0567_ net943 sg13g2_a21oi_1
X_1867_ Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q net37 net8 net82 net92 Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q
+ _0362_ VPWR VGND sg13g2_mux4_1
X_1936_ _0428_ VPWR Inst_RegFile_switch_matrix.JW2BEG4 VGND _0424_ _0417_ sg13g2_o21ai_1
X_2985_ net1157 net1137 Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q VPWR VGND sg13g2_dlhq_1
Xinput82 SS4END[0] net82 VPWR VGND sg13g2_buf_1
Xinput71 S2MID[1] net71 VPWR VGND sg13g2_buf_1
X_3606_ net1165 net181 VPWR VGND sg13g2_buf_1
X_3537_ Inst_RegFile_switch_matrix.E2BEG5 net119 VPWR VGND sg13g2_buf_8
Xinput60 S1END[2] net60 VPWR VGND sg13g2_buf_1
Xinput93 W2END[4] net93 VPWR VGND sg13g2_buf_1
X_1798_ _0298_ _0296_ _0297_ _0291_ net955 VPWR VGND sg13g2_a22oi_1
XFILLER_57_501 VPWR VGND sg13g2_fill_1
X_2419_ _0881_ VPWR _0882_ VGND Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q _0880_ sg13g2_o21ai_1
XFILLER_52_272 VPWR VGND sg13g2_fill_1
XFILLER_25_420 VPWR VGND sg13g2_fill_2
XFILLER_32_76 VPWR VGND sg13g2_fill_2
XFILLER_0_530 VPWR VGND sg13g2_fill_1
X_1721_ _0224_ _0225_ Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q _0226_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_43_283 VPWR VGND sg13g2_fill_1
XFILLER_31_445 VPWR VGND sg13g2_fill_2
X_2770_ net933 net817 _1116_ _0071_ VPWR VGND sg13g2_mux2_1
X_1583_ Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q net56 _1203_ VPWR VGND sg13g2_nor2b_1
X_3322_ net1182 net1142 Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q VPWR VGND sg13g2_dlhq_1
X_1652_ _0160_ _0159_ Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q VPWR VGND sg13g2_nand2b_1
Xfanout1191 FrameData[19] net1191 VPWR VGND sg13g2_buf_1
X_2204_ Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q net1034 _0680_ VPWR VGND sg13g2_nor2b_1
X_2135_ _0615_ VPWR B_ADR0 VGND _0604_ _0602_ sg13g2_o21ai_1
Xfanout1180 net1181 net1180 VPWR VGND sg13g2_buf_1
X_3253_ net1194 net1117 Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q VPWR VGND sg13g2_dlhq_1
X_3184_ net1206 net1103 Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q VPWR VGND sg13g2_dlhq_1
XFILLER_34_294 VPWR VGND sg13g2_fill_1
X_2066_ net990 Inst_RegFile_32x4.mem\[0\]\[3\] Inst_RegFile_32x4.mem\[1\]\[3\] Inst_RegFile_32x4.mem\[2\]\[3\]
+ Inst_RegFile_32x4.mem\[3\]\[3\] net944 _0552_ VPWR VGND sg13g2_mux4_1
X_2968_ net1186 net1133 Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q VPWR VGND sg13g2_dlhq_1
X_1919_ VGND VPWR _0367_ _0411_ _0412_ net1009 sg13g2_a21oi_1
X_2899_ UserCLK net423 _0057_ _2899_/Q_N Inst_RegFile_32x4.mem\[16\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_32_209 VPWR VGND sg13g2_fill_2
XFILLER_27_76 VPWR VGND sg13g2_fill_2
XFILLER_43_97 VPWR VGND sg13g2_decap_8
XFILLER_40_242 VPWR VGND sg13g2_decap_8
XFILLER_48_342 VPWR VGND sg13g2_decap_4
X_2684_ net961 net768 _1091_ _0010_ VPWR VGND sg13g2_mux2_1
XFILLER_31_275 VPWR VGND sg13g2_decap_4
X_1704_ Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q net34 net62 net22 net89 Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q
+ _0209_ VPWR VGND sg13g2_mux4_1
X_2753_ net949 net845 _1113_ _0057_ VPWR VGND sg13g2_mux2_1
X_2822_ _1061_ _1097_ _1128_ VPWR VGND sg13g2_and2_2
X_1566_ VGND VPWR _1187_ net1066 net1048 sg13g2_or2_1
X_3305_ net1156 net1143 Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q VPWR VGND sg13g2_dlhq_1
X_1635_ _1232_ _1230_ _0141_ _0143_ VPWR VGND sg13g2_a21o_2
XFILLER_54_356 VPWR VGND sg13g2_fill_1
X_2118_ Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q net53 _0599_ VPWR VGND sg13g2_nor2b_1
X_3167_ net1172 net1101 Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q VPWR VGND sg13g2_dlhq_1
X_2049_ VGND VPWR net1036 _0533_ _0535_ net1008 sg13g2_a21oi_1
X_3098_ net1182 net1088 Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q VPWR VGND sg13g2_dlhq_1
X_3236_ net1212 net1115 Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q VPWR VGND sg13g2_dlhq_1
XFILLER_10_448 VPWR VGND sg13g2_fill_1
XFILLER_13_23 VPWR VGND sg13g2_fill_1
Xfanout995 net996 net995 VPWR VGND sg13g2_buf_1
Xfanout940 net942 net940 VPWR VGND sg13g2_buf_1
Xfanout973 AD3 net973 VPWR VGND sg13g2_buf_8
Xfanout962 _1069_ net962 VPWR VGND sg13g2_buf_1
Xfanout951 net954 net951 VPWR VGND sg13g2_buf_1
Xfanout984 net985 net984 VPWR VGND sg13g2_buf_1
XFILLER_54_30 VPWR VGND sg13g2_fill_1
XFILLER_55_7 VPWR VGND sg13g2_decap_8
XFILLER_51_304 VPWR VGND sg13g2_fill_1
XFILLER_48_183 VPWR VGND sg13g2_fill_1
X_3021_ net1149 net1077 Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q VPWR VGND sg13g2_dlhq_1
XFILLER_24_529 VPWR VGND sg13g2_fill_2
X_2805_ net962 net764 _1124_ _0098_ VPWR VGND sg13g2_mux2_1
X_2667_ _1081_ VPWR _1082_ VGND net43 Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q sg13g2_o21ai_1
X_2736_ _1110_ _1092_ _1108_ VPWR VGND sg13g2_nand2_2
X_1618_ Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q _1235_ _1236_ _1237_ VPWR VGND
+ sg13g2_nor3_1
X_1549_ _1171_ net974 Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q VPWR VGND sg13g2_nand2b_1
X_3219_ net1199 net1110 Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q VPWR VGND sg13g2_dlhq_1
X_2598_ Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q net1029 _0338_ Inst_RegFile_switch_matrix.JW2BEG1
+ net521 Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q Inst_RegFile_switch_matrix.N1BEG2
+ VPWR VGND sg13g2_mux4_1
Xhold290 Inst_RegFile_32x4.mem\[5\]\[1\] VPWR VGND net788 sg13g2_dlygate4sd3_1
XFILLER_45_175 VPWR VGND sg13g2_fill_2
XFILLER_33_348 VPWR VGND sg13g2_fill_1
X_3379__365 VPWR VGND net365 sg13g2_tiehi
X_3570_ EE4END[14] net143 VPWR VGND sg13g2_buf_1
X_2521_ Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q VPWR _0972_ VGND net1063 _1183_
+ sg13g2_o21ai_1
X_2383_ _0848_ VPWR Inst_RegFile_switch_matrix.E2BEG7 VGND _0842_ _0843_ sg13g2_o21ai_1
X_2452_ Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q VPWR _0913_ VGND net1061 _1183_
+ sg13g2_o21ai_1
XFILLER_36_164 VPWR VGND sg13g2_decap_4
X_3004_ net1178 net1138 Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q VPWR VGND sg13g2_dlhq_1
Xinput3 E1END[2] net3 VPWR VGND sg13g2_buf_1
XFILLER_51_178 VPWR VGND sg13g2_fill_1
X_3768_ WW4END[7] net356 VPWR VGND sg13g2_buf_1
X_3699_ net77 net281 VPWR VGND sg13g2_buf_1
X_2719_ net740 net940 _1104_ _0032_ VPWR VGND sg13g2_mux2_1
Xfanout1009 _0409_ net1009 VPWR VGND sg13g2_buf_1
Xoutput351 Inst_RegFile_switch_matrix.WW4BEG1 WW4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput340 net340 W6BEG[3] VPWR VGND sg13g2_buf_1
Xoutput362 net362 WW4BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_59_289 VPWR VGND sg13g2_fill_1
XFILLER_55_451 VPWR VGND sg13g2_decap_8
XFILLER_19_109 VPWR VGND sg13g2_fill_1
XFILLER_42_189 VPWR VGND sg13g2_decap_8
XFILLER_42_101 VPWR VGND sg13g2_decap_8
XFILLER_35_54 VPWR VGND sg13g2_fill_2
XFILLER_7_503 VPWR VGND sg13g2_fill_1
XFILLER_25_8 VPWR VGND sg13g2_fill_2
X_3622_ FrameStrobe[14] net195 VPWR VGND sg13g2_buf_1
X_1883_ _0377_ VPWR _0378_ VGND Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q net1011
+ sg13g2_o21ai_1
X_1952_ Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q VPWR _0444_ VGND _0443_ _0442_
+ sg13g2_o21ai_1
X_3553_ E6END[7] net137 VPWR VGND sg13g2_buf_1
X_2504_ Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q net57 net85 net1219 net1070 Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q
+ _0956_ VPWR VGND sg13g2_mux4_1
X_2435_ Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q _0896_ _0895_ net499 net500 Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q
+ _0897_ VPWR VGND sg13g2_mux4_1
XFILLER_56_226 VPWR VGND sg13g2_fill_2
X_2297_ VPWR _0768_ _0767_ VGND sg13g2_inv_1
X_2366_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q _0829_ _0833_ _0832_ sg13g2_a21oi_1
XFILLER_52_498 VPWR VGND sg13g2_fill_1
XFILLER_52_487 VPWR VGND sg13g2_fill_2
XFILLER_52_454 VPWR VGND sg13g2_decap_4
XFILLER_21_78 VPWR VGND sg13g2_fill_1
Xoutput192 net192 FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
Xoutput181 net181 FrameData_O[30] VPWR VGND sg13g2_buf_1
Xoutput170 net170 FrameData_O[20] VPWR VGND sg13g2_buf_1
X_3369__375 VPWR VGND net375 sg13g2_tiehi
XFILLER_43_465 VPWR VGND sg13g2_fill_2
X_3376__368 VPWR VGND net368 sg13g2_tiehi
XFILLER_7_69 VPWR VGND sg13g2_fill_2
X_2220_ VGND VPWR _0694_ _0695_ _0691_ Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q sg13g2_a21oi_2
X_2151_ Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q VPWR _0631_ VGND Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q
+ _0629_ sg13g2_o21ai_1
X_2082_ net991 Inst_RegFile_32x4.mem\[20\]\[2\] Inst_RegFile_32x4.mem\[21\]\[2\] Inst_RegFile_32x4.mem\[22\]\[2\]
+ Inst_RegFile_32x4.mem\[23\]\[2\] net945 _0566_ VPWR VGND sg13g2_mux4_1
XFILLER_46_292 VPWR VGND sg13g2_fill_1
X_2984_ net1159 net1139 Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q VPWR VGND sg13g2_dlhq_1
XFILLER_21_115 VPWR VGND sg13g2_decap_8
X_3605_ net1169 net179 VPWR VGND sg13g2_buf_1
Xinput61 S1END[3] net61 VPWR VGND sg13g2_buf_1
Xinput72 S2MID[2] net72 VPWR VGND sg13g2_buf_1
X_1866_ Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q VPWR _0361_ VGND Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q
+ _0360_ sg13g2_o21ai_1
X_1935_ _0428_ _0427_ Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q VPWR VGND sg13g2_nand2b_1
Xinput50 N4END[0] net50 VPWR VGND sg13g2_buf_1
X_1797_ VGND VPWR net1024 _0293_ _0297_ net956 sg13g2_a21oi_1
Xinput83 SS4END[1] net83 VPWR VGND sg13g2_buf_1
X_3536_ Inst_RegFile_switch_matrix.E2BEG4 net118 VPWR VGND sg13g2_buf_1
Xinput94 W2END[5] net94 VPWR VGND sg13g2_buf_1
X_2418_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q _0878_ _0881_ Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q
+ sg13g2_a21oi_1
X_2349_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q _0814_ _0817_ _1150_
+ sg13g2_a21oi_1
XFILLER_40_402 VPWR VGND sg13g2_fill_2
X_1720_ net1047 net22 net59 net61 net69 Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q
+ _0225_ VPWR VGND sg13g2_mux4_1
X_1651_ _0157_ _0158_ Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q _0159_ VPWR VGND
+ sg13g2_mux2_1
X_3252_ net1196 net1117 Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q VPWR VGND sg13g2_dlhq_1
X_1582_ net80 Inst_RegFile_switch_matrix.E2BEG3 Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q
+ _1202_ VPWR VGND sg13g2_mux2_1
X_3321_ net1184 net1143 Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q VPWR VGND sg13g2_dlhq_1
Xfanout1181 FrameData[23] net1181 VPWR VGND sg13g2_buf_1
Xfanout1170 net1171 net1170 VPWR VGND sg13g2_buf_1
X_3183_ net1209 net1108 Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q VPWR VGND sg13g2_dlhq_1
X_2203_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q _1165_ _0679_ _0678_ sg13g2_a21oi_1
X_2134_ Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q _0609_ _0614_ _0615_ VPWR VGND sg13g2_or3_1
Xfanout1192 net1193 net1192 VPWR VGND sg13g2_buf_1
X_2065_ _0551_ _0550_ net1008 _0549_ _0546_ VPWR VGND sg13g2_a22oi_1
XFILLER_21_2 VPWR VGND sg13g2_fill_1
X_2967_ net1191 net1132 Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q VPWR VGND sg13g2_dlhq_1
X_3359__385 VPWR VGND net385 sg13g2_tiehi
X_1918_ VGND VPWR Inst_RegFile_32x4.mem\[9\]\[0\] net995 _0411_ _0410_ sg13g2_a21oi_1
X_1849_ VGND VPWR _1133_ _0344_ _0345_ Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q
+ sg13g2_a21oi_1
X_2898_ UserCLK net424 _0056_ _2898_/Q_N Inst_RegFile_32x4.mem\[16\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_57_343 VPWR VGND sg13g2_fill_1
X_3366__378 VPWR VGND net378 sg13g2_tiehi
XFILLER_57_387 VPWR VGND sg13g2_decap_8
XFILLER_13_402 VPWR VGND sg13g2_fill_2
XFILLER_43_65 VPWR VGND sg13g2_fill_2
XFILLER_4_122 VPWR VGND sg13g2_fill_2
XFILLER_4_155 VPWR VGND sg13g2_fill_2
X_2821_ net748 net935 _1127_ _0111_ VPWR VGND sg13g2_mux2_1
X_1703_ _0208_ VPWR Inst_RegFile_switch_matrix.JN2BEG5 VGND _0204_ _0197_ sg13g2_o21ai_1
X_2683_ net952 net755 _1091_ _0009_ VPWR VGND sg13g2_mux2_1
X_1634_ VGND VPWR _0141_ _0142_ _1232_ _1230_ sg13g2_a21oi_2
XFILLER_8_483 VPWR VGND sg13g2_fill_1
XFILLER_8_494 VPWR VGND sg13g2_fill_2
X_2752_ net938 net774 _1113_ _0056_ VPWR VGND sg13g2_mux2_1
X_3235_ net1163 net1113 Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q VPWR VGND sg13g2_dlhq_1
X_1565_ _1185_ VPWR _1186_ VGND net1048 net976 sg13g2_o21ai_1
X_3304_ net1158 net1143 Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q VPWR VGND sg13g2_dlhq_1
X_2117_ net81 Inst_RegFile_switch_matrix.JN2BEG4 Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q
+ _0598_ VPWR VGND sg13g2_mux2_1
X_3166_ net1174 net1100 Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q VPWR VGND sg13g2_dlhq_1
X_2048_ Inst_RegFile_32x4.mem\[26\]\[3\] Inst_RegFile_32x4.mem\[27\]\[3\] net993 _0534_
+ VPWR VGND sg13g2_mux2_1
X_3097_ net1184 net1091 Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q VPWR VGND sg13g2_dlhq_1
Xfanout974 net974 net975 VPWR VGND sg13g2_buf_16
Xfanout941 net942 net941 VPWR VGND sg13g2_buf_1
Xfanout952 net954 net952 VPWR VGND sg13g2_buf_1
Xfanout996 net997 net996 VPWR VGND sg13g2_buf_1
Xfanout930 net931 net930 VPWR VGND sg13g2_buf_1
Xfanout985 BD2 net985 VPWR VGND sg13g2_buf_8
Xfanout963 net504 net963 VPWR VGND sg13g2_buf_8
XFILLER_41_530 VPWR VGND sg13g2_fill_1
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_5_475 VPWR VGND sg13g2_fill_1
XFILLER_51_327 VPWR VGND sg13g2_fill_2
XFILLER_48_195 VPWR VGND sg13g2_fill_2
X_3020_ net1151 net1078 Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q VPWR VGND sg13g2_dlhq_1
X_3349__395 VPWR VGND net395 sg13g2_tiehi
XFILLER_44_390 VPWR VGND sg13g2_fill_2
XFILLER_32_530 VPWR VGND sg13g2_fill_1
X_2804_ net952 net788 _1124_ _0097_ VPWR VGND sg13g2_mux2_1
X_3356__388 VPWR VGND net388 sg13g2_tiehi
X_2597_ Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q net1013 _0486_ Inst_RegFile_switch_matrix.JW2BEG2
+ _1016_ Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q Inst_RegFile_switch_matrix.N1BEG3
+ VPWR VGND sg13g2_mux4_1
X_2666_ _1081_ Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q net14 VPWR VGND sg13g2_nand2b_1
X_2735_ net933 net795 _1109_ _0043_ VPWR VGND sg13g2_mux2_1
X_1617_ net1012 Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q _1236_ VPWR VGND sg13g2_nor2b_1
XFILLER_59_427 VPWR VGND sg13g2_decap_4
X_1548_ _1170_ Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q net1033 VPWR VGND sg13g2_nand2_1
X_3149_ net1149 net1102 Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q VPWR VGND sg13g2_dlhq_1
XFILLER_27_335 VPWR VGND sg13g2_fill_2
X_3218_ net1202 net1110 Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q VPWR VGND sg13g2_dlhq_1
XFILLER_50_360 VPWR VGND sg13g2_fill_2
Xhold280 Inst_RegFile_32x4.mem\[14\]\[3\] VPWR VGND net778 sg13g2_dlygate4sd3_1
Xhold291 Inst_RegFile_32x4.mem\[28\]\[3\] VPWR VGND net789 sg13g2_dlygate4sd3_1
XFILLER_58_460 VPWR VGND sg13g2_fill_1
XFILLER_1_16 VPWR VGND sg13g2_fill_2
XFILLER_14_530 VPWR VGND sg13g2_fill_1
X_2520_ _0911_ _0910_ net1063 _0971_ VPWR VGND sg13g2_mux2_1
X_2451_ _0911_ _0910_ net1061 _0912_ VPWR VGND sg13g2_mux2_1
X_2382_ _0847_ VPWR _0848_ VGND Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q _0844_
+ sg13g2_o21ai_1
XFILLER_56_419 VPWR VGND sg13g2_fill_2
X_3003_ net1180 net1139 Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q VPWR VGND sg13g2_dlhq_1
Xinput4 E1END[3] net4 VPWR VGND sg13g2_buf_1
XFILLER_51_124 VPWR VGND sg13g2_fill_1
X_3767_ WW4END[6] net355 VPWR VGND sg13g2_buf_1
X_2718_ _1088_ _1103_ _1104_ VPWR VGND sg13g2_and2_2
X_3698_ net76 net280 VPWR VGND sg13g2_buf_1
X_2649_ Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q net23 net96 net80 Inst_RegFile_switch_matrix.E2BEG1
+ Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q _1066_ VPWR VGND sg13g2_mux4_1
Xoutput330 net330 W2BEGb[3] VPWR VGND sg13g2_buf_1
Xoutput352 net352 WW4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput341 net341 W6BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_27_121 VPWR VGND sg13g2_fill_1
XFILLER_51_54 VPWR VGND sg13g2_fill_2
XFILLER_33_135 VPWR VGND sg13g2_fill_2
XFILLER_33_113 VPWR VGND sg13g2_fill_1
X_3346__398 VPWR VGND net398 sg13g2_tiehi
X_3621_ FrameStrobe[13] net194 VPWR VGND sg13g2_buf_1
X_3552_ E6END[6] net136 VPWR VGND sg13g2_buf_1
X_1882_ _0377_ Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q net1002 VPWR VGND sg13g2_nand2_1
X_1951_ Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q BD1 _0443_ VPWR VGND sg13g2_nor2_2
XFILLER_37_0 VPWR VGND sg13g2_fill_2
X_2503_ VGND VPWR _0955_ Inst_RegFile_switch_matrix.SS4BEG0 _0953_ _0949_ sg13g2_a21oi_2
X_2365_ Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q VPWR _0832_ VGND Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q
+ _0831_ sg13g2_o21ai_1
X_2434_ Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q net46 net101 net17 net503 Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q
+ _0896_ VPWR VGND sg13g2_mux4_1
XFILLER_37_463 VPWR VGND sg13g2_fill_2
X_2296_ net1059 net22 net1217 net64 net91 Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q
+ _0767_ VPWR VGND sg13g2_mux4_1
XFILLER_24_102 VPWR VGND sg13g2_decap_8
XFILLER_2_70 VPWR VGND sg13g2_decap_8
XFILLER_52_433 VPWR VGND sg13g2_decap_8
XFILLER_24_113 VPWR VGND sg13g2_fill_2
XFILLER_12_319 VPWR VGND sg13g2_fill_2
XFILLER_4_529 VPWR VGND sg13g2_fill_2
Xoutput193 net193 FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
Xoutput171 net171 FrameData_O[21] VPWR VGND sg13g2_buf_1
Xoutput182 net182 FrameData_O[31] VPWR VGND sg13g2_buf_1
Xoutput160 net160 FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_28_474 VPWR VGND sg13g2_fill_2
XFILLER_11_396 VPWR VGND sg13g2_fill_1
X_2081_ _0565_ _0564_ net1005 VPWR VGND sg13g2_nand2b_1
X_2150_ net93 net109 net1057 _0630_ VPWR VGND sg13g2_mux2_1
XFILLER_34_455 VPWR VGND sg13g2_fill_1
XFILLER_34_444 VPWR VGND sg13g2_fill_1
X_1934_ _0425_ _0426_ Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q _0427_ VPWR VGND
+ sg13g2_mux2_1
X_2983_ net1161 net1139 Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q VPWR VGND sg13g2_dlhq_1
Xinput84 SS4END[2] net84 VPWR VGND sg13g2_buf_1
Xinput62 S2END[0] net62 VPWR VGND sg13g2_buf_1
Xinput73 S2MID[3] net73 VPWR VGND sg13g2_buf_1
X_3604_ net1171 net178 VPWR VGND sg13g2_buf_1
X_1865_ VGND VPWR net84 Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q _0360_ _0359_ sg13g2_a21oi_1
X_3535_ Inst_RegFile_switch_matrix.E2BEG3 net117 VPWR VGND sg13g2_buf_8
Xinput95 W2END[6] net95 VPWR VGND sg13g2_buf_1
Xinput40 N2END[6] net40 VPWR VGND sg13g2_buf_1
Xinput51 N4END[1] net51 VPWR VGND sg13g2_buf_1
X_1796_ _0296_ _0295_ net1024 VPWR VGND sg13g2_nand2b_1
X_2348_ VGND VPWR net62 net1042 _0816_ _0815_ sg13g2_a21oi_1
X_2417_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q net979 _0880_ _0879_ sg13g2_a21oi_1
X_2279_ net1049 net52 _0751_ VPWR VGND sg13g2_nor2b_1
XFILLER_40_425 VPWR VGND sg13g2_fill_2
XFILLER_40_414 VPWR VGND sg13g2_fill_1
XFILLER_57_75 VPWR VGND sg13g2_fill_2
XFILLER_31_447 VPWR VGND sg13g2_fill_1
XFILLER_16_411 VPWR VGND sg13g2_fill_2
XFILLER_16_444 VPWR VGND sg13g2_fill_1
X_1581_ _1201_ VPWR Inst_RegFile_switch_matrix.E2BEG3 VGND _1189_ _1196_ sg13g2_o21ai_1
X_1650_ net1039 net1217 net66 net78 net93 Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q
+ _0158_ VPWR VGND sg13g2_mux4_1
X_2202_ Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q VPWR _0678_ VGND Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q
+ net988 sg13g2_o21ai_1
X_3182_ net1210 net1108 Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q VPWR VGND sg13g2_dlhq_1
X_3251_ net1198 net1116 Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q VPWR VGND sg13g2_dlhq_1
X_3320_ net1186 net1143 Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q VPWR VGND sg13g2_dlhq_1
Xfanout1171 FrameData[28] net1171 VPWR VGND sg13g2_buf_1
Xfanout1182 FrameData[22] net1182 VPWR VGND sg13g2_buf_1
X_2133_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q _0612_ _0614_ _0613_
+ sg13g2_a21oi_1
Xfanout1193 FrameData[18] net1193 VPWR VGND sg13g2_buf_1
X_2064_ net997 Inst_RegFile_32x4.mem\[12\]\[3\] Inst_RegFile_32x4.mem\[13\]\[3\] Inst_RegFile_32x4.mem\[14\]\[3\]
+ Inst_RegFile_32x4.mem\[15\]\[3\] net947 _0550_ VPWR VGND sg13g2_mux4_1
Xfanout1160 FrameData[3] net1160 VPWR VGND sg13g2_buf_1
X_1917_ net995 Inst_RegFile_32x4.mem\[8\]\[0\] _0410_ VPWR VGND sg13g2_nor2b_1
X_2966_ net1193 net1132 Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q VPWR VGND sg13g2_dlhq_1
X_2897_ UserCLK net425 _0055_ _2897_/Q_N Inst_RegFile_32x4.mem\[15\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_22_436 VPWR VGND sg13g2_fill_1
X_1848_ net87 net1017 Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q _0344_ VPWR VGND
+ sg13g2_mux2_1
X_1779_ net923 Inst_RegFile_32x4.mem\[22\]\[1\] _0281_ VPWR VGND sg13g2_nor2b_1
XFILLER_57_366 VPWR VGND sg13g2_decap_8
XFILLER_27_78 VPWR VGND sg13g2_fill_1
XFILLER_25_274 VPWR VGND sg13g2_fill_1
XFILLER_13_447 VPWR VGND sg13g2_fill_2
XFILLER_4_38 VPWR VGND sg13g2_fill_1
XFILLER_4_145 VPWR VGND sg13g2_fill_1
XFILLER_51_509 VPWR VGND sg13g2_fill_2
X_2820_ net730 net960 _1127_ _0110_ VPWR VGND sg13g2_mux2_1
XFILLER_31_299 VPWR VGND sg13g2_fill_2
X_2751_ _1113_ _1061_ _1106_ VPWR VGND sg13g2_nand2_2
X_1702_ _0208_ _0207_ Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q VPWR VGND sg13g2_nand2b_1
X_2682_ net942 net757 _1091_ _0008_ VPWR VGND sg13g2_mux2_1
X_1564_ _1185_ net1048 net504 VPWR VGND sg13g2_nand2_1
X_1633_ VGND VPWR _0140_ _0141_ Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q _0137_
+ sg13g2_a21oi_2
X_3234_ net1165 net1113 Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q VPWR VGND sg13g2_dlhq_1
X_3165_ net1177 net1100 Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q VPWR VGND sg13g2_dlhq_1
X_3303_ net1160 net1144 Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q VPWR VGND sg13g2_dlhq_1
X_2116_ _0593_ VPWR Inst_RegFile_switch_matrix.JN2BEG4 VGND _0597_ Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q
+ sg13g2_o21ai_1
X_2047_ VGND VPWR Inst_RegFile_32x4.mem\[25\]\[3\] net993 _0533_ _0532_ sg13g2_a21oi_1
X_3096_ net1186 net1091 Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q VPWR VGND sg13g2_dlhq_1
X_2949_ net1189 net1136 Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q VPWR VGND sg13g2_dlhq_1
X_3372__372 VPWR VGND net372 sg13g2_tiehi
Xfanout942 _1065_ net942 VPWR VGND sg13g2_buf_1
Xfanout931 A_ADR0 net931 VPWR VGND sg13g2_buf_1
XFILLER_1_126 VPWR VGND sg13g2_fill_1
XFILLER_54_21 VPWR VGND sg13g2_decap_8
Xfanout986 net987 net986 VPWR VGND sg13g2_buf_1
Xfanout953 net954 net953 VPWR VGND sg13g2_buf_1
XFILLER_45_336 VPWR VGND sg13g2_fill_1
Xfanout997 net998 net997 VPWR VGND sg13g2_buf_1
Xfanout975 net975 AD3 VPWR VGND sg13g2_buf_16
XFILLER_36_336 VPWR VGND sg13g2_fill_2
X_2803_ net940 net777 _1124_ _0096_ VPWR VGND sg13g2_mux2_1
X_2734_ net958 net840 _1109_ _0042_ VPWR VGND sg13g2_mux2_1
XFILLER_59_406 VPWR VGND sg13g2_decap_8
X_1547_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q _1165_ _1169_ _1168_
+ sg13g2_a21oi_1
X_2596_ Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q net36 net51 net1214 net1031 Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q
+ Inst_RegFile_switch_matrix.N4BEG0 VPWR VGND sg13g2_mux4_1
X_2665_ VGND VPWR _1079_ Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q _1077_ Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q
+ _1080_ _1076_ sg13g2_a221oi_1
X_1616_ Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q net1029 _1235_ VPWR VGND sg13g2_nor2_1
X_3148_ net1151 net1102 Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q VPWR VGND sg13g2_dlhq_1
XFILLER_39_196 VPWR VGND sg13g2_decap_8
X_3217_ net1203 net1110 Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q VPWR VGND sg13g2_dlhq_1
XFILLER_42_306 VPWR VGND sg13g2_fill_1
XFILLER_35_391 VPWR VGND sg13g2_fill_2
X_3079_ net1160 net1089 Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q VPWR VGND sg13g2_dlhq_1
XFILLER_40_67 VPWR VGND sg13g2_fill_1
XFILLER_49_21 VPWR VGND sg13g2_decap_8
Xhold292 Inst_RegFile_32x4.mem\[11\]\[3\] VPWR VGND net790 sg13g2_dlygate4sd3_1
Xhold270 Inst_RegFile_32x4.mem\[26\]\[2\] VPWR VGND net768 sg13g2_dlygate4sd3_1
Xhold281 Inst_RegFile_32x4.mem\[18\]\[0\] VPWR VGND net779 sg13g2_dlygate4sd3_1
XFILLER_18_303 VPWR VGND sg13g2_fill_2
X_2381_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q _0846_ _0847_ Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q
+ sg13g2_a21oi_1
XFILLER_39_4 VPWR VGND sg13g2_fill_2
X_2450_ Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q net45 net16 net73 net100 Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q
+ _0911_ VPWR VGND sg13g2_mux4_1
XFILLER_56_409 VPWR VGND sg13g2_decap_4
X_3002_ net1182 net1140 Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q VPWR VGND sg13g2_dlhq_1
XFILLER_36_133 VPWR VGND sg13g2_fill_2
Xinput5 E2END[0] net5 VPWR VGND sg13g2_buf_1
X_3362__382 VPWR VGND net382 sg13g2_tiehi
X_3766_ WW4END[5] net354 VPWR VGND sg13g2_buf_1
XFILLER_10_37 VPWR VGND sg13g2_fill_2
X_3697_ net75 net279 VPWR VGND sg13g2_buf_1
X_2717_ _1100_ _1033_ _1103_ VPWR VGND sg13g2_nor2b_1
X_2648_ net942 net844 _1062_ _0000_ VPWR VGND sg13g2_mux2_1
Xoutput320 net320 W2BEG[1] VPWR VGND sg13g2_buf_1
Xoutput331 net331 W2BEGb[4] VPWR VGND sg13g2_buf_1
X_2579_ Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q net43 net14 net71 net98 Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q
+ _1018_ VPWR VGND sg13g2_mux4_1
Xoutput342 net342 W6BEG[5] VPWR VGND sg13g2_buf_1
Xoutput353 net353 WW4BEG[15] VPWR VGND sg13g2_buf_1
XFILLER_35_56 VPWR VGND sg13g2_fill_1
XFILLER_2_265 VPWR VGND sg13g2_fill_1
XFILLER_18_100 VPWR VGND sg13g2_decap_4
X_1950_ BD3 Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q _0442_ VPWR VGND sg13g2_nor2b_1
X_3551_ E6END[5] net135 VPWR VGND sg13g2_buf_1
X_3620_ net1130 net193 VPWR VGND sg13g2_buf_1
X_1881_ Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q _0374_ _0375_ _0376_ VPWR VGND
+ sg13g2_nor3_2
X_2502_ Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q _0954_ _0955_ VPWR VGND sg13g2_nor2_1
X_2433_ Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q net46 net74 net17 Inst_RegFile_switch_matrix.JS2BEG4
+ Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q _0895_ VPWR VGND sg13g2_mux4_1
X_2364_ VGND VPWR net79 net1046 _0831_ _0830_ sg13g2_a21oi_1
X_2295_ Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q net36 net1221 net52 net7 Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q
+ _0766_ VPWR VGND sg13g2_mux4_1
XFILLER_52_489 VPWR VGND sg13g2_fill_1
Xoutput161 net161 FrameData_O[12] VPWR VGND sg13g2_buf_1
Xoutput150 net150 EE4BEG[2] VPWR VGND sg13g2_buf_1
X_3749_ net101 net331 VPWR VGND sg13g2_buf_1
Xoutput194 net194 FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
Xoutput183 net183 FrameData_O[3] VPWR VGND sg13g2_buf_1
Xoutput172 net172 FrameData_O[22] VPWR VGND sg13g2_buf_1
XFILLER_46_33 VPWR VGND sg13g2_fill_2
XFILLER_28_464 VPWR VGND sg13g2_fill_1
XFILLER_15_158 VPWR VGND sg13g2_fill_2
X_2842__439 VPWR VGND net439 sg13g2_tiehi
X_3352__392 VPWR VGND net392 sg13g2_tiehi
XFILLER_34_423 VPWR VGND sg13g2_fill_1
X_2080_ net991 Inst_RegFile_32x4.mem\[16\]\[2\] Inst_RegFile_32x4.mem\[17\]\[2\] Inst_RegFile_32x4.mem\[18\]\[2\]
+ Inst_RegFile_32x4.mem\[19\]\[2\] net945 _0564_ VPWR VGND sg13g2_mux4_1
X_2982_ net1166 net1141 Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q VPWR VGND sg13g2_dlhq_1
X_1933_ Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q net59 net67 net61 net1071 net1038
+ _0426_ VPWR VGND sg13g2_mux4_1
XFILLER_21_139 VPWR VGND sg13g2_fill_2
Xinput85 SS4END[3] net85 VPWR VGND sg13g2_buf_1
Xinput63 S2END[1] net63 VPWR VGND sg13g2_buf_1
Xinput74 S2MID[4] net74 VPWR VGND sg13g2_buf_1
X_3603_ net1173 net177 VPWR VGND sg13g2_buf_1
X_3534_ Inst_RegFile_switch_matrix.E2BEG2 net116 VPWR VGND sg13g2_buf_2
X_1864_ Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q net52 _0359_ VPWR VGND sg13g2_nor2b_1
Xinput30 N1END[0] net30 VPWR VGND sg13g2_buf_1
Xinput41 N2END[7] net41 VPWR VGND sg13g2_buf_1
Xinput52 N4END[2] net52 VPWR VGND sg13g2_buf_1
X_1795_ VGND VPWR Inst_RegFile_32x4.mem\[7\]\[2\] net926 _0295_ _0294_ sg13g2_a21oi_1
Xinput96 W2END[7] net96 VPWR VGND sg13g2_buf_1
X_2347_ net1042 net58 _0815_ VPWR VGND sg13g2_nor2b_1
X_2278_ VGND VPWR net91 net1049 _0750_ _0749_ sg13g2_a21oi_1
X_2416_ net1060 net1065 _0879_ VPWR VGND sg13g2_nor2b_1
XFILLER_52_253 VPWR VGND sg13g2_fill_1
XFILLER_32_35 VPWR VGND sg13g2_fill_2
XFILLER_43_242 VPWR VGND sg13g2_fill_1
X_1580_ _1200_ _1199_ Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q _1201_ VPWR VGND
+ sg13g2_a21o_1
X_2201_ _0677_ VPWR Inst_RegFile_switch_matrix.JS2BEG2 VGND _0673_ _0672_ sg13g2_o21ai_1
X_3181_ net1148 net1108 Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q VPWR VGND sg13g2_dlhq_1
Xfanout1183 FrameData[22] net1183 VPWR VGND sg13g2_buf_1
X_2132_ Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q VPWR _0613_ VGND Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q
+ _0611_ sg13g2_o21ai_1
Xfanout1150 net1151 net1150 VPWR VGND sg13g2_buf_1
Xfanout1172 FrameData[27] net1172 VPWR VGND sg13g2_buf_1
Xfanout1161 FrameData[3] net1161 VPWR VGND sg13g2_buf_1
X_3250_ net1201 net1116 Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q VPWR VGND sg13g2_dlhq_1
Xfanout1194 net1195 net1194 VPWR VGND sg13g2_buf_1
X_2063_ VGND VPWR net1036 _0548_ _0549_ net1008 sg13g2_a21oi_1
XFILLER_19_283 VPWR VGND sg13g2_fill_2
X_2965_ net1194 net1132 Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q VPWR VGND sg13g2_dlhq_1
X_1847_ _0343_ Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q _0342_ VPWR VGND sg13g2_nand2_1
X_1916_ Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q _0388_ _0408_ _0229_ _0407_ Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q
+ _0409_ VPWR VGND sg13g2_mux4_1
X_2896_ UserCLK net426 _0054_ _2896_/Q_N Inst_RegFile_32x4.mem\[15\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_1778_ VGND VPWR Inst_RegFile_32x4.mem\[21\]\[1\] net923 _0280_ _0279_ sg13g2_a21oi_1
X_3379_ UserCLK net365 _0115_ _3379_/Q_N Inst_RegFile_32x4.mem\[0\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_40_256 VPWR VGND sg13g2_decap_8
XFILLER_40_223 VPWR VGND sg13g2_fill_2
XFILLER_40_201 VPWR VGND sg13g2_fill_1
XFILLER_13_404 VPWR VGND sg13g2_fill_1
XFILLER_4_157 VPWR VGND sg13g2_fill_1
X_1701_ _0206_ _0205_ Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q _0207_ VPWR VGND
+ sg13g2_mux2_1
X_2681_ _1091_ _1090_ _1034_ VPWR VGND sg13g2_nand2_2
X_2750_ net736 net934 _1112_ _0055_ VPWR VGND sg13g2_mux2_1
X_1563_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q _1183_ _1184_ Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q
+ sg13g2_a21oi_1
X_3302_ net1167 net1144 Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q VPWR VGND sg13g2_dlhq_1
X_1632_ Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q VPWR _0140_ VGND Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q
+ _0139_ sg13g2_o21ai_1
X_3233_ net1169 net1113 Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q VPWR VGND sg13g2_dlhq_1
X_3164_ net1178 net1100 Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q VPWR VGND sg13g2_dlhq_1
X_2115_ VGND VPWR _0596_ _0597_ _0594_ Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q
+ sg13g2_a21oi_2
X_3095_ net1190 net1091 Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q VPWR VGND sg13g2_dlhq_1
XFILLER_12_0 VPWR VGND sg13g2_fill_1
X_2046_ net993 Inst_RegFile_32x4.mem\[24\]\[3\] _0532_ VPWR VGND sg13g2_nor2b_1
X_2948_ net1213 net1131 Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q VPWR VGND sg13g2_dlhq_1
XFILLER_22_278 VPWR VGND sg13g2_fill_2
X_2879_ UserCLK net451 _0037_ _2879_/Q_N Inst_RegFile_32x4.mem\[17\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
Xfanout965 net965 net513 VPWR VGND sg13g2_buf_16
Xfanout976 _1167_ net976 VPWR VGND sg13g2_buf_8
Xfanout954 _1067_ net954 VPWR VGND sg13g2_buf_1
Xfanout943 _0460_ net943 VPWR VGND sg13g2_buf_8
Xfanout932 net933 net932 VPWR VGND sg13g2_buf_8
Xfanout921 net921 net922 VPWR VGND sg13g2_buf_16
Xfanout998 B_ADR0 net998 VPWR VGND sg13g2_buf_1
Xfanout987 net989 net987 VPWR VGND sg13g2_buf_1
XFILLER_44_392 VPWR VGND sg13g2_fill_1
X_2664_ Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q _1078_ _1079_ VPWR VGND sg13g2_nor2_1
X_2733_ net951 net793 _1109_ _0041_ VPWR VGND sg13g2_mux2_1
X_2802_ _1124_ _1088_ _1122_ VPWR VGND sg13g2_nand2_2
X_1546_ Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q VPWR _1168_ VGND Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q
+ net988 sg13g2_o21ai_1
X_2595_ Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q net37 net52 net1216 net1013 Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q
+ Inst_RegFile_switch_matrix.N4BEG1 VPWR VGND sg13g2_mux4_1
XFILLER_5_71 VPWR VGND sg13g2_fill_1
X_1615_ Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q _1233_ _1234_ VPWR VGND sg13g2_nor2_2
X_3078_ net1166 net1089 Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q VPWR VGND sg13g2_dlhq_1
XFILLER_27_348 VPWR VGND sg13g2_fill_1
XFILLER_27_337 VPWR VGND sg13g2_fill_1
X_3216_ net1206 net1110 Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q VPWR VGND sg13g2_dlhq_1
X_3147_ net1152 net1099 Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q VPWR VGND sg13g2_dlhq_1
X_2029_ _0517_ _0514_ _0516_ VPWR VGND sg13g2_nand2_2
XFILLER_2_425 VPWR VGND sg13g2_fill_1
XFILLER_2_403 VPWR VGND sg13g2_fill_2
Xhold260 Inst_RegFile_32x4.mem\[22\]\[0\] VPWR VGND net758 sg13g2_dlygate4sd3_1
Xhold271 Inst_RegFile_32x4.mem\[28\]\[1\] VPWR VGND net769 sg13g2_dlygate4sd3_1
XFILLER_49_55 VPWR VGND sg13g2_fill_2
Xhold293 Inst_RegFile_32x4.mem\[3\]\[3\] VPWR VGND net791 sg13g2_dlygate4sd3_1
XFILLER_1_18 VPWR VGND sg13g2_fill_1
Xhold282 Inst_RegFile_32x4.mem\[3\]\[2\] VPWR VGND net780 sg13g2_dlygate4sd3_1
XFILLER_41_362 VPWR VGND sg13g2_fill_2
X_2380_ VPWR _0846_ _0845_ VGND sg13g2_inv_1
XFILLER_53_7 VPWR VGND sg13g2_decap_8
X_3001_ net1185 net1140 Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q VPWR VGND sg13g2_dlhq_1
Xinput6 E2END[1] net6 VPWR VGND sg13g2_buf_1
XFILLER_17_370 VPWR VGND sg13g2_fill_2
X_2716_ net935 net811 _1102_ _0031_ VPWR VGND sg13g2_mux2_1
X_2647_ Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q _1063_ _1064_ _0978_ _1016_ Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q
+ _1065_ VPWR VGND sg13g2_mux4_1
Xoutput332 net332 W2BEGb[5] VPWR VGND sg13g2_buf_1
Xoutput321 net321 W2BEG[2] VPWR VGND sg13g2_buf_1
X_3765_ WW4END[4] net347 VPWR VGND sg13g2_buf_1
Xoutput310 net310 SS4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput343 net343 W6BEG[6] VPWR VGND sg13g2_buf_1
X_3696_ net74 net278 VPWR VGND sg13g2_buf_1
X_1529_ VPWR _1151_ Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q VGND sg13g2_inv_1
X_2578_ Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q net52 net96 net7 Inst_RegFile_switch_matrix.E2BEG2
+ Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q _1017_ VPWR VGND sg13g2_mux4_1
Xoutput354 net354 WW4BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_19_47 VPWR VGND sg13g2_fill_1
XFILLER_55_498 VPWR VGND sg13g2_fill_1
XFILLER_55_465 VPWR VGND sg13g2_decap_8
XFILLER_51_56 VPWR VGND sg13g2_fill_1
XFILLER_51_23 VPWR VGND sg13g2_fill_2
X_1880_ net1032 Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q _0375_ VPWR VGND sg13g2_nor2b_1
XFILLER_33_137 VPWR VGND sg13g2_fill_1
XFILLER_14_395 VPWR VGND sg13g2_fill_2
XFILLER_18_189 VPWR VGND sg13g2_fill_1
X_3550_ E6END[4] net134 VPWR VGND sg13g2_buf_1
X_2501_ Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q net1074 net1219 net88 net980 Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q
+ _0954_ VPWR VGND sg13g2_mux4_1
XFILLER_37_2 VPWR VGND sg13g2_fill_1
X_2432_ Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q net1017 net718 net979 net971 Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q
+ _0894_ VPWR VGND sg13g2_mux4_1
X_2294_ Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q VPWR _0765_ VGND _0764_ _0763_ sg13g2_o21ai_1
X_2363_ net1046 net63 _0830_ VPWR VGND sg13g2_nor2b_1
XFILLER_49_281 VPWR VGND sg13g2_fill_1
XFILLER_37_465 VPWR VGND sg13g2_fill_1
X_3748_ net100 net330 VPWR VGND sg13g2_buf_1
XFILLER_32_181 VPWR VGND sg13g2_fill_2
XFILLER_20_310 VPWR VGND sg13g2_fill_1
XFILLER_20_365 VPWR VGND sg13g2_fill_2
Xoutput173 net173 FrameData_O[23] VPWR VGND sg13g2_buf_1
Xoutput195 net195 FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
Xoutput140 net140 E6BEG[8] VPWR VGND sg13g2_buf_1
Xoutput162 net162 FrameData_O[13] VPWR VGND sg13g2_buf_1
Xoutput184 net184 FrameData_O[4] VPWR VGND sg13g2_buf_1
Xoutput151 net151 EE4BEG[3] VPWR VGND sg13g2_buf_1
X_3679_ Inst_RegFile_switch_matrix.NN4BEG3 net252 VPWR VGND sg13g2_buf_1
XFILLER_28_443 VPWR VGND sg13g2_fill_2
XFILLER_55_273 VPWR VGND sg13g2_fill_2
XFILLER_11_321 VPWR VGND sg13g2_fill_1
XFILLER_7_303 VPWR VGND sg13g2_fill_2
XFILLER_7_358 VPWR VGND sg13g2_fill_1
XFILLER_19_421 VPWR VGND sg13g2_fill_1
X_3602_ net1174 net176 VPWR VGND sg13g2_buf_1
X_1863_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q _0356_ _0358_ _0357_
+ sg13g2_a21oi_1
X_1932_ net1038 net1075 net39 net1220 net10 Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q
+ _0425_ VPWR VGND sg13g2_mux4_1
Xinput20 E2MID[7] net20 VPWR VGND sg13g2_buf_1
Xinput31 net31 N1END[1] VPWR VGND sg13g2_buf_16
X_2981_ net1188 net1137 Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q VPWR VGND sg13g2_dlhq_1
Xinput64 S2END[2] net64 VPWR VGND sg13g2_buf_1
Xinput75 S2MID[5] net75 VPWR VGND sg13g2_buf_1
XFILLER_42_0 VPWR VGND sg13g2_decap_8
Xinput97 W2MID[0] net97 VPWR VGND sg13g2_buf_1
Xinput86 W1END[0] net86 VPWR VGND sg13g2_buf_1
Xinput42 N2MID[0] net42 VPWR VGND sg13g2_buf_1
Xinput53 N4END[3] net53 VPWR VGND sg13g2_buf_1
X_2415_ net963 net970 net1060 _0878_ VPWR VGND sg13g2_mux2_1
X_3533_ Inst_RegFile_switch_matrix.E2BEG1 net115 VPWR VGND sg13g2_buf_2
X_1794_ net926 Inst_RegFile_32x4.mem\[6\]\[2\] _0294_ VPWR VGND sg13g2_nor2b_1
X_2346_ net82 net1072 Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q _0814_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_37_240 VPWR VGND sg13g2_fill_2
X_2277_ net1049 net64 _0749_ VPWR VGND sg13g2_nor2b_1
XFILLER_52_232 VPWR VGND sg13g2_fill_2
XFILLER_37_295 VPWR VGND sg13g2_fill_1
XFILLER_57_44 VPWR VGND sg13g2_fill_2
XFILLER_16_413 VPWR VGND sg13g2_fill_1
XFILLER_16_457 VPWR VGND sg13g2_fill_2
Xfanout1184 FrameData[21] net1184 VPWR VGND sg13g2_buf_1
X_3180_ net1150 net1108 Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q VPWR VGND sg13g2_dlhq_1
Xfanout1140 net1141 net1140 VPWR VGND sg13g2_buf_1
X_2200_ _0677_ _0676_ Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q VPWR VGND sg13g2_nand2b_1
Xfanout1162 FrameData[31] net1162 VPWR VGND sg13g2_buf_1
Xfanout1151 FrameData[8] net1151 VPWR VGND sg13g2_buf_1
X_2131_ net77 net104 Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q _0612_ VPWR VGND sg13g2_mux2_1
Xfanout1195 FrameData[17] net1195 VPWR VGND sg13g2_buf_1
X_2062_ VGND VPWR Inst_RegFile_32x4.mem\[9\]\[3\] net995 _0548_ _0547_ sg13g2_a21oi_1
Xfanout1173 FrameData[27] net1173 VPWR VGND sg13g2_buf_1
X_2964_ net1197 net1134 Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q VPWR VGND sg13g2_dlhq_1
XFILLER_34_265 VPWR VGND sg13g2_fill_1
X_1846_ net978 net966 Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q _0342_ VPWR VGND
+ sg13g2_mux2_1
X_1915_ Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q net55 net10 net67 net94 Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q
+ _0408_ VPWR VGND sg13g2_mux4_1
Xrebuffer219 Inst_RegFile_switch_matrix.JN2BEG3 net717 VPWR VGND sg13g2_dlygate4sd1_1
X_2895_ UserCLK net427 _0053_ _2895_/Q_N Inst_RegFile_32x4.mem\[15\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_1777_ net923 Inst_RegFile_32x4.mem\[20\]\[1\] _0279_ VPWR VGND sg13g2_nor2b_1
X_3378_ UserCLK net366 _0114_ _3378_/Q_N Inst_RegFile_32x4.mem\[0\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_2329_ Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q net63 net79 net82 net90 Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q
+ _0798_ VPWR VGND sg13g2_mux4_1
XFILLER_13_449 VPWR VGND sg13g2_fill_1
XFILLER_48_346 VPWR VGND sg13g2_fill_1
XFILLER_0_375 VPWR VGND sg13g2_fill_2
X_1700_ Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q net1074 net56 net40 net1219 net1054
+ _0206_ VPWR VGND sg13g2_mux4_1
X_2680_ _1048_ _1060_ _1058_ _1090_ VPWR VGND sg13g2_nor3_2
XFILLER_31_279 VPWR VGND sg13g2_fill_1
X_1631_ VPWR _0139_ _0138_ VGND sg13g2_inv_1
X_3232_ net1170 net1113 Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q VPWR VGND sg13g2_dlhq_1
X_1562_ VPWR _1183_ _1182_ VGND sg13g2_inv_1
X_3301_ net1188 net1146 Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q VPWR VGND sg13g2_dlhq_1
XFILLER_3_191 VPWR VGND sg13g2_fill_1
X_2114_ Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q _0595_ _0596_ VPWR VGND sg13g2_nor2b_1
X_3094_ net1193 net1091 Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q VPWR VGND sg13g2_dlhq_1
X_2045_ Inst_RegFile_32x4.BD_comb\[1\] Inst_RegFile_32x4.BD_reg\[1\] Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q
+ BD1 VPWR VGND sg13g2_mux2_2
X_3163_ net1180 net1098 Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q VPWR VGND sg13g2_dlhq_1
X_2947_ net1163 net1127 Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q VPWR VGND sg13g2_dlhq_1
XFILLER_10_419 VPWR VGND sg13g2_fill_1
X_1829_ net922 Inst_RegFile_32x4.mem\[30\]\[3\] Inst_RegFile_32x4.mem\[31\]\[3\] Inst_RegFile_32x4.mem\[28\]\[3\]
+ Inst_RegFile_32x4.mem\[29\]\[3\] net1022 _0327_ VPWR VGND sg13g2_mux4_1
X_2878_ UserCLK net452 _0036_ _2878_/Q_N Inst_RegFile_32x4.mem\[17\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_57_110 VPWR VGND sg13g2_fill_1
Xfanout988 net989 net988 VPWR VGND sg13g2_buf_1
Xfanout966 net513 net966 VPWR VGND sg13g2_buf_1
Xfanout977 _1167_ net977 VPWR VGND sg13g2_buf_1
Xfanout999 _1165_ net999 VPWR VGND sg13g2_buf_2
Xfanout922 A_ADR0 net922 VPWR VGND sg13g2_buf_8
Xfanout944 net946 net944 VPWR VGND sg13g2_buf_1
Xfanout933 net936 net933 VPWR VGND sg13g2_buf_8
Xfanout955 _0143_ net955 VPWR VGND sg13g2_buf_1
XFILLER_5_412 VPWR VGND sg13g2_fill_2
XFILLER_17_530 VPWR VGND sg13g2_fill_1
X_2801_ net727 net934 _1123_ _0095_ VPWR VGND sg13g2_mux2_1
X_2594_ Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q net34 net1065 net53 net986 Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q
+ Inst_RegFile_switch_matrix.N4BEG2 VPWR VGND sg13g2_mux4_1
X_2663_ net42 Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q _1078_ VPWR VGND sg13g2_nor2_1
X_2732_ net939 net758 _1109_ _0040_ VPWR VGND sg13g2_mux2_1
X_1614_ Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q net1067 net1018 net979 net504 Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q
+ _1233_ VPWR VGND sg13g2_mux4_1
X_1545_ _1167_ net978 VPWR VGND sg13g2_inv_2
X_3215_ net1209 net1114 Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q VPWR VGND sg13g2_dlhq_1
XFILLER_54_146 VPWR VGND sg13g2_fill_1
X_3077_ net1189 net1090 Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q VPWR VGND sg13g2_dlhq_1
X_2028_ VGND VPWR _0459_ _0516_ _0515_ net1004 sg13g2_a21oi_2
X_3146_ net1154 net1099 Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q VPWR VGND sg13g2_dlhq_1
XFILLER_40_25 VPWR VGND sg13g2_decap_4
Xhold261 Inst_RegFile_32x4.mem\[10\]\[0\] VPWR VGND net759 sg13g2_dlygate4sd3_1
Xhold250 Inst_RegFile_32x4.mem\[8\]\[3\] VPWR VGND net748 sg13g2_dlygate4sd3_1
Xhold272 Inst_RegFile_32x4.mem\[7\]\[1\] VPWR VGND net770 sg13g2_dlygate4sd3_1
Xhold294 Inst_RegFile_32x4.mem\[3\]\[0\] VPWR VGND net792 sg13g2_dlygate4sd3_1
Xhold283 Inst_RegFile_32x4.mem\[19\]\[0\] VPWR VGND net781 sg13g2_dlygate4sd3_1
XFILLER_58_496 VPWR VGND sg13g2_fill_1
XFILLER_18_305 VPWR VGND sg13g2_fill_1
XFILLER_30_80 VPWR VGND sg13g2_fill_2
X_3000_ net1187 net1140 Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q VPWR VGND sg13g2_dlhq_1
XFILLER_36_168 VPWR VGND sg13g2_fill_2
XFILLER_36_113 VPWR VGND sg13g2_fill_2
Xinput7 E2END[2] net7 VPWR VGND sg13g2_buf_1
XFILLER_17_360 VPWR VGND sg13g2_fill_1
XFILLER_32_341 VPWR VGND sg13g2_fill_1
XFILLER_32_330 VPWR VGND sg13g2_fill_2
X_2646_ Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q net49 net20 net77 net104 Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q
+ _1064_ VPWR VGND sg13g2_mux4_1
X_2715_ net961 net823 _1102_ _0030_ VPWR VGND sg13g2_mux2_1
X_3695_ net73 net277 VPWR VGND sg13g2_buf_1
Xoutput322 net507 W2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput355 net355 WW4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput333 net333 W2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput300 net300 SS4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput311 net311 SS4BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_10_39 VPWR VGND sg13g2_fill_1
X_2577_ Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q net984 _0645_ Inst_RegFile_switch_matrix.JS2BEG0
+ net502 Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q Inst_RegFile_switch_matrix.W1BEG1
+ VPWR VGND sg13g2_mux4_1
Xoutput344 net344 W6BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_55_422 VPWR VGND sg13g2_decap_8
X_1528_ VPWR _1150_ Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q VGND sg13g2_inv_1
XFILLER_35_47 VPWR VGND sg13g2_decap_8
X_2909__413 VPWR VGND net413 sg13g2_tiehi
X_3129_ net1185 net1096 Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q VPWR VGND sg13g2_dlhq_1
X_2916__406 VPWR VGND net406 sg13g2_tiehi
X_2431_ Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q net56 net1219 net84 net1070 Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q
+ _0893_ VPWR VGND sg13g2_mux4_1
X_2500_ _0953_ _0952_ VPWR VGND sg13g2_inv_2
X_2293_ _0764_ _0761_ Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q VPWR VGND sg13g2_nand2_2
XFILLER_2_40 VPWR VGND sg13g2_fill_2
X_2362_ net90 net106 net1046 _0829_ VPWR VGND sg13g2_mux2_1
XFILLER_52_469 VPWR VGND sg13g2_fill_1
XFILLER_52_447 VPWR VGND sg13g2_decap_8
XFILLER_17_190 VPWR VGND sg13g2_decap_4
X_3747_ net99 net329 VPWR VGND sg13g2_buf_1
XFILLER_20_399 VPWR VGND sg13g2_fill_2
Xoutput196 net196 FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
Xoutput141 net141 E6BEG[9] VPWR VGND sg13g2_buf_1
Xoutput163 net163 FrameData_O[14] VPWR VGND sg13g2_buf_1
Xoutput174 net174 FrameData_O[24] VPWR VGND sg13g2_buf_1
Xoutput130 net130 E6BEG[0] VPWR VGND sg13g2_buf_1
Xoutput185 net185 FrameData_O[5] VPWR VGND sg13g2_buf_1
X_3678_ Inst_RegFile_switch_matrix.NN4BEG2 net251 VPWR VGND sg13g2_buf_1
Xoutput152 net152 EE4BEG[4] VPWR VGND sg13g2_buf_1
X_2629_ _1041_ _1046_ _1047_ VPWR VGND sg13g2_and2_1
XFILLER_55_263 VPWR VGND sg13g2_fill_1
X_2980_ net1212 net1137 Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q VPWR VGND sg13g2_dlhq_1
X_3601_ net1177 net175 VPWR VGND sg13g2_buf_1
X_1862_ Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q VPWR _0357_ VGND Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q
+ net91 sg13g2_o21ai_1
Xinput21 EE4END[0] net21 VPWR VGND sg13g2_buf_1
X_1931_ Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q VPWR _0424_ VGND _0423_ _0420_
+ sg13g2_o21ai_1
Xinput10 E2END[5] net10 VPWR VGND sg13g2_buf_1
Xinput32 N1END[2] net32 VPWR VGND sg13g2_buf_1
Xinput43 N2MID[1] net43 VPWR VGND sg13g2_buf_1
Xinput54 NN4END[0] net54 VPWR VGND sg13g2_buf_1
X_1793_ VGND VPWR Inst_RegFile_32x4.mem\[5\]\[2\] net926 _0293_ _0292_ sg13g2_a21oi_1
Xinput65 S2END[3] net65 VPWR VGND sg13g2_buf_1
Xinput76 S2MID[6] net76 VPWR VGND sg13g2_buf_1
X_2414_ _0877_ VPWR Inst_RegFile_switch_matrix.JN2BEG7 VGND _0871_ _0869_ sg13g2_o21ai_1
XFILLER_35_0 VPWR VGND sg13g2_fill_1
Xinput87 W1END[1] net87 VPWR VGND sg13g2_buf_8
Xinput98 W2MID[1] net98 VPWR VGND sg13g2_buf_1
XFILLER_6_381 VPWR VGND sg13g2_fill_2
X_3532_ Inst_RegFile_switch_matrix.E2BEG0 net114 VPWR VGND sg13g2_buf_2
X_2345_ Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q net1076 net1221 net34 net5 Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q
+ _0813_ VPWR VGND sg13g2_mux4_1
X_2276_ VGND VPWR net1216 net1049 _0748_ _0747_ sg13g2_a21oi_1
X_2906__416 VPWR VGND net416 sg13g2_tiehi
XFILLER_32_48 VPWR VGND sg13g2_decap_8
XFILLER_57_23 VPWR VGND sg13g2_fill_1
X_2913__409 VPWR VGND net409 sg13g2_tiehi
XFILLER_28_296 VPWR VGND sg13g2_decap_4
XFILLER_22_70 VPWR VGND sg13g2_decap_4
Xfanout1185 FrameData[21] net1185 VPWR VGND sg13g2_buf_1
Xfanout1130 net27 net1130 VPWR VGND sg13g2_buf_1
X_2061_ net995 Inst_RegFile_32x4.mem\[8\]\[3\] _0547_ VPWR VGND sg13g2_nor2b_1
Xfanout1141 FrameStrobe[10] net1141 VPWR VGND sg13g2_buf_1
Xfanout1163 FrameData[31] net1163 VPWR VGND sg13g2_buf_1
X_2130_ _0610_ VPWR _0611_ VGND net49 Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q sg13g2_o21ai_1
Xfanout1174 net1175 net1174 VPWR VGND sg13g2_buf_1
Xfanout1196 net1197 net1196 VPWR VGND sg13g2_buf_1
Xfanout1152 net1153 net1152 VPWR VGND sg13g2_buf_1
X_2963_ net1200 net1134 Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q VPWR VGND sg13g2_dlhq_1
X_1914_ Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q net1215 net79 net109 Inst_RegFile_switch_matrix.JS2BEG4
+ Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q _0407_ VPWR VGND sg13g2_mux4_1
XFILLER_19_285 VPWR VGND sg13g2_fill_1
X_2894_ UserCLK net428 _0052_ _2894_/Q_N Inst_RegFile_32x4.mem\[15\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_1845_ _0340_ VPWR _0341_ VGND Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q _0228_ sg13g2_o21ai_1
XFILLER_8_50 VPWR VGND sg13g2_fill_2
X_1776_ net925 Inst_RegFile_32x4.mem\[18\]\[1\] Inst_RegFile_32x4.mem\[19\]\[1\] Inst_RegFile_32x4.mem\[16\]\[1\]
+ Inst_RegFile_32x4.mem\[17\]\[1\] net1023 _0278_ VPWR VGND sg13g2_mux4_1
XFILLER_57_314 VPWR VGND sg13g2_decap_4
X_3377_ UserCLK net367 _0113_ _3377_/Q_N Inst_RegFile_32x4.mem\[0\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_2328_ net1041 net1073 net35 net6 net1214 Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q
+ _0797_ VPWR VGND sg13g2_mux4_1
X_2259_ _0732_ _0731_ Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q VPWR VGND sg13g2_nand2_2
XFILLER_21_483 VPWR VGND sg13g2_fill_1
X_1630_ Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q net39 net10 net83 net94 Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q
+ _0138_ VPWR VGND sg13g2_mux4_1
XFILLER_12_450 VPWR VGND sg13g2_fill_1
X_3231_ net1172 net1111 Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q VPWR VGND sg13g2_dlhq_1
X_1561_ Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q net45 net16 net73 net100 Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q
+ _1182_ VPWR VGND sg13g2_mux4_1
X_3300_ net1212 net1146 Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q VPWR VGND sg13g2_dlhq_1
X_3162_ net1182 net1098 Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q VPWR VGND sg13g2_dlhq_1
X_3093_ net1195 net1092 Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q VPWR VGND sg13g2_dlhq_1
X_2113_ net1055 net1075 net39 net57 net1220 Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q
+ _0595_ VPWR VGND sg13g2_mux4_1
X_2044_ _0517_ _0522_ _0531_ Inst_RegFile_32x4.BD_comb\[1\] VPWR VGND sg13g2_a21o_1
X_2946_ net1165 net1127 Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q VPWR VGND sg13g2_dlhq_1
X_2877_ UserCLK net453 _0035_ _2877_/Q_N Inst_RegFile_32x4.mem\[13\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_22_247 VPWR VGND sg13g2_fill_2
X_2903__419 VPWR VGND net419 sg13g2_tiehi
X_1828_ _0325_ VPWR _0326_ VGND net1026 _0322_ sg13g2_o21ai_1
X_1759_ Inst_RegFile_32x4.AD_comb\[0\] Inst_RegFile_32x4.AD_reg\[0\] Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q
+ AD0 VPWR VGND sg13g2_mux2_2
Xfanout967 net513 net967 VPWR VGND sg13g2_buf_1
Xfanout978 net979 net978 VPWR VGND sg13g2_buf_8
Xfanout934 net936 net934 VPWR VGND sg13g2_buf_1
Xfanout989 BD2 net989 VPWR VGND sg13g2_buf_1
Xfanout945 net946 net945 VPWR VGND sg13g2_buf_1
Xfanout923 net925 net923 VPWR VGND sg13g2_buf_1
Xfanout956 _0143_ net956 VPWR VGND sg13g2_buf_1
X_3344__400 VPWR VGND net400 sg13g2_tiehi
XFILLER_57_188 VPWR VGND sg13g2_fill_1
X_3780_ Inst_RegFile_switch_matrix.WW4BEG3 net353 VPWR VGND sg13g2_buf_1
X_2731_ _1109_ _1090_ _1108_ VPWR VGND sg13g2_nand2_2
X_2800_ net734 net962 _1123_ _0094_ VPWR VGND sg13g2_mux2_1
X_1544_ VPWR _1166_ net1017 VGND sg13g2_inv_1
X_2593_ Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q net35 net50 net1066 net1001 Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q
+ Inst_RegFile_switch_matrix.N4BEG3 VPWR VGND sg13g2_mux4_1
X_2662_ _1077_ Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q net13 VPWR VGND sg13g2_nand2b_1
X_1613_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q _1231_ _1232_ Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q
+ sg13g2_a21oi_1
X_3214_ net1211 net1112 Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q VPWR VGND sg13g2_dlhq_1
XFILLER_27_317 VPWR VGND sg13g2_fill_1
X_3145_ net1156 net1099 Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q VPWR VGND sg13g2_dlhq_1
XFILLER_54_125 VPWR VGND sg13g2_fill_2
X_3076_ net1213 net1090 Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q VPWR VGND sg13g2_dlhq_1
XFILLER_23_501 VPWR VGND sg13g2_fill_2
X_2027_ net990 Inst_RegFile_32x4.mem\[28\]\[1\] Inst_RegFile_32x4.mem\[29\]\[1\] Inst_RegFile_32x4.mem\[30\]\[1\]
+ Inst_RegFile_32x4.mem\[31\]\[1\] net944 _0515_ VPWR VGND sg13g2_mux4_1
X_2929_ net1203 net1128 Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q VPWR VGND sg13g2_dlhq_1
XFILLER_49_79 VPWR VGND sg13g2_fill_1
XFILLER_49_57 VPWR VGND sg13g2_fill_1
Xhold284 Inst_RegFile_32x4.mem\[25\]\[2\] VPWR VGND net782 sg13g2_dlygate4sd3_1
Xhold262 Inst_RegFile_32x4.mem\[15\]\[0\] VPWR VGND net760 sg13g2_dlygate4sd3_1
Xhold251 Inst_RegFile_32x4.mem\[0\]\[3\] VPWR VGND net749 sg13g2_dlygate4sd3_1
Xhold295 Inst_RegFile_32x4.mem\[22\]\[1\] VPWR VGND net793 sg13g2_dlygate4sd3_1
Xhold240 Inst_RegFile_32x4.mem\[2\]\[0\] VPWR VGND net738 sg13g2_dlygate4sd3_1
Xhold273 Inst_RegFile_32x4.mem\[12\]\[1\] VPWR VGND net771 sg13g2_dlygate4sd3_1
XFILLER_58_453 VPWR VGND sg13g2_decap_8
XFILLER_26_361 VPWR VGND sg13g2_fill_2
Xinput8 E2END[3] net8 VPWR VGND sg13g2_buf_1
XFILLER_17_372 VPWR VGND sg13g2_fill_1
X_3763_ Inst_RegFile_switch_matrix.W6BEG0 net336 VPWR VGND sg13g2_buf_1
X_2714_ net953 net831 _1102_ _0029_ VPWR VGND sg13g2_mux2_1
X_3694_ net72 net276 VPWR VGND sg13g2_buf_1
XFILLER_59_206 VPWR VGND sg13g2_fill_2
X_1527_ VPWR _1149_ Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q VGND sg13g2_inv_1
X_2645_ Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q net48 net76 net103 net517 Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q
+ _1063_ VPWR VGND sg13g2_mux4_1
X_3334__443 VPWR VGND net443 sg13g2_tiehi
Xoutput356 net356 WW4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput323 net323 W2BEG[4] VPWR VGND sg13g2_buf_1
Xoutput334 net334 W2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput301 Inst_RegFile_switch_matrix.SS4BEG0 SS4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput312 net312 SS4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput345 net345 W6BEG[8] VPWR VGND sg13g2_buf_1
X_2576_ Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q net1001 _0338_ Inst_RegFile_switch_matrix.JS2BEG1
+ net522 Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q Inst_RegFile_switch_matrix.W1BEG2
+ VPWR VGND sg13g2_mux4_1
XFILLER_59_239 VPWR VGND sg13g2_fill_2
X_3341__403 VPWR VGND net403 sg13g2_tiehi
X_3128_ net1186 net1096 Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q VPWR VGND sg13g2_dlhq_1
XFILLER_51_25 VPWR VGND sg13g2_fill_1
XFILLER_51_14 VPWR VGND sg13g2_decap_4
X_3059_ net1198 net1085 Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q VPWR VGND sg13g2_dlhq_1
XFILLER_46_445 VPWR VGND sg13g2_fill_2
X_2361_ Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q net35 net6 net1218 net1214 Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q
+ _0828_ VPWR VGND sg13g2_mux4_1
X_2430_ _0888_ VPWR Inst_RegFile_switch_matrix.JN2BEG0 VGND Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q
+ _0892_ sg13g2_o21ai_1
XFILLER_37_423 VPWR VGND sg13g2_fill_2
X_2292_ VGND VPWR net1059 net999 _0763_ _0762_ sg13g2_a21oi_1
XFILLER_2_63 VPWR VGND sg13g2_decap_8
XFILLER_52_426 VPWR VGND sg13g2_decap_8
XFILLER_32_183 VPWR VGND sg13g2_fill_1
X_3746_ net98 net328 VPWR VGND sg13g2_buf_1
XFILLER_20_367 VPWR VGND sg13g2_fill_1
Xoutput197 net197 FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
Xoutput175 net175 FrameData_O[25] VPWR VGND sg13g2_buf_1
Xoutput164 net164 FrameData_O[15] VPWR VGND sg13g2_buf_1
X_2559_ Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q net1076 net1221 net1072 net974
+ Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q _1004_ VPWR VGND sg13g2_mux4_1
Xoutput131 Inst_RegFile_switch_matrix.E6BEG0 E6BEG[10] VPWR VGND sg13g2_buf_1
Xoutput186 net186 FrameData_O[6] VPWR VGND sg13g2_buf_1
Xoutput142 net142 EE4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput153 net153 EE4BEG[5] VPWR VGND sg13g2_buf_1
X_2628_ _1045_ VPWR _1046_ VGND Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q _1042_
+ sg13g2_o21ai_1
Xoutput120 net120 E2BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_46_69 VPWR VGND sg13g2_fill_2
XFILLER_28_445 VPWR VGND sg13g2_fill_1
XFILLER_23_194 VPWR VGND sg13g2_fill_1
X_1930_ Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q VPWR _0423_ VGND _0421_ _0422_
+ sg13g2_o21ai_1
Xinput66 S2END[4] net66 VPWR VGND sg13g2_buf_1
Xinput77 S2MID[7] net77 VPWR VGND sg13g2_buf_1
X_3600_ net1179 net174 VPWR VGND sg13g2_buf_1
X_1861_ _0356_ Inst_RegFile_switch_matrix.E2BEG4 VPWR VGND sg13g2_inv_4
Xinput22 EE4END[1] net22 VPWR VGND sg13g2_buf_1
Xinput11 E2END[6] net11 VPWR VGND sg13g2_buf_1
Xinput88 W1END[2] net88 VPWR VGND sg13g2_buf_1
Xinput33 N1END[3] net33 VPWR VGND sg13g2_buf_1
Xinput44 N2MID[2] net44 VPWR VGND sg13g2_buf_1
Xinput55 NN4END[1] net55 VPWR VGND sg13g2_buf_1
X_1792_ net926 Inst_RegFile_32x4.mem\[4\]\[2\] _0292_ VPWR VGND sg13g2_nor2b_1
X_2344_ Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q _0811_ _0806_ _0812_ VPWR VGND
+ sg13g2_nand3_1
X_2413_ _0877_ _0876_ Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q VPWR VGND sg13g2_nand2b_1
Xinput99 W2MID[2] net99 VPWR VGND sg13g2_buf_1
XFILLER_37_242 VPWR VGND sg13g2_fill_1
X_2275_ net1049 net7 _0747_ VPWR VGND sg13g2_nor2b_1
XFILLER_16_459 VPWR VGND sg13g2_fill_1
Xfanout1120 FrameStrobe[2] net1120 VPWR VGND sg13g2_buf_1
Xfanout1131 net1136 net1131 VPWR VGND sg13g2_buf_1
Xfanout1186 FrameData[20] net1186 VPWR VGND sg13g2_buf_1
Xfanout1164 net1165 net1164 VPWR VGND sg13g2_buf_1
X_2060_ _0546_ net947 _0545_ VPWR VGND sg13g2_nand2_1
Xfanout1175 FrameData[26] net1175 VPWR VGND sg13g2_buf_1
Xfanout1153 net26 net1153 VPWR VGND sg13g2_buf_1
Xfanout1197 FrameData[16] net1197 VPWR VGND sg13g2_buf_1
Xfanout1142 net1143 net1142 VPWR VGND sg13g2_buf_1
X_1913_ _0406_ VPWR Inst_RegFile_switch_matrix.JS2BEG4 VGND _0402_ _0395_ sg13g2_o21ai_1
X_2962_ net1202 net1135 Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q VPWR VGND sg13g2_dlhq_1
X_2893_ UserCLK net429 _0051_ _2893_/Q_N Inst_RegFile_32x4.mem\[14\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_1844_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q _0339_ _0340_ Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q
+ sg13g2_a21oi_1
XFILLER_30_484 VPWR VGND sg13g2_fill_2
X_1775_ VGND VPWR net982 _0276_ _0277_ net969 sg13g2_a21oi_1
X_2912__410 VPWR VGND net410 sg13g2_tiehi
X_2258_ _0730_ VPWR _0731_ VGND net1045 net1029 sg13g2_o21ai_1
X_2327_ Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q VPWR _0796_ VGND _0795_ _0794_ sg13g2_o21ai_1
X_3376_ UserCLK net368 _0112_ _3376_/Q_N Inst_RegFile_32x4.mem\[0\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_2189_ VGND VPWR _0664_ _0665_ _0666_ Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q sg13g2_a21oi_1
XFILLER_56_381 VPWR VGND sg13g2_decap_8
XFILLER_16_256 VPWR VGND sg13g2_fill_2
XFILLER_17_82 VPWR VGND sg13g2_fill_2
XFILLER_33_81 VPWR VGND sg13g2_fill_2
X_1560_ VGND VPWR _1181_ _1180_ Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q sg13g2_or2_1
X_3230_ net1175 net1111 Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q VPWR VGND sg13g2_dlhq_1
XFILLER_39_359 VPWR VGND sg13g2_fill_1
X_2112_ net1055 net10 net59 net67 net1071 Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q
+ _0594_ VPWR VGND sg13g2_mux4_1
X_3161_ net1184 net1099 Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q VPWR VGND sg13g2_dlhq_1
XFILLER_3_160 VPWR VGND sg13g2_fill_1
X_3092_ net1196 net1090 Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q VPWR VGND sg13g2_dlhq_1
X_2043_ VGND VPWR _0530_ _0492_ _0528_ _0524_ _0531_ _0526_ sg13g2_a221oi_1
X_2945_ net1168 net1127 Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q VPWR VGND sg13g2_dlhq_1
X_1827_ VGND VPWR net1027 _0324_ _0325_ net983 sg13g2_a21oi_1
X_2876_ UserCLK net454 _0034_ _2876_/Q_N Inst_RegFile_32x4.mem\[13\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_1689_ VGND VPWR _0195_ net1070 net1054 sg13g2_or2_1
Xfanout924 net925 net924 VPWR VGND sg13g2_buf_1
X_1758_ _0186_ _0192_ _0247_ _0250_ _0261_ _0236_ Inst_RegFile_32x4.AD_comb\[0\] VPWR
+ VGND sg13g2_mux4_1
XFILLER_54_14 VPWR VGND sg13g2_decap_8
Xfanout979 net979 AD1 VPWR VGND sg13g2_buf_16
XFILLER_38_48 VPWR VGND sg13g2_decap_4
Xfanout935 net936 net935 VPWR VGND sg13g2_buf_1
X_3359_ UserCLK net385 _0095_ _3359_/Q_N Inst_RegFile_32x4.mem\[4\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
Xfanout946 _0368_ net946 VPWR VGND sg13g2_buf_1
XFILLER_53_395 VPWR VGND sg13g2_decap_8
XFILLER_53_362 VPWR VGND sg13g2_fill_1
XFILLER_48_189 VPWR VGND sg13g2_fill_1
X_2902__420 VPWR VGND net420 sg13g2_tiehi
X_2661_ net70 net508 Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q _1076_ VPWR VGND sg13g2_mux2_1
X_2730_ _1105_ _1033_ _1108_ VPWR VGND sg13g2_nor2b_2
X_1543_ _1165_ net1003 VPWR VGND sg13g2_inv_2
X_2592_ Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q net975 Inst_RegFile_switch_matrix.JN2BEG3
+ _1018_ _1017_ Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q Inst_RegFile_switch_matrix.E1BEG0
+ VPWR VGND sg13g2_mux4_1
X_1612_ Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q net47 net18 net75 net102 Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q
+ _1231_ VPWR VGND sg13g2_mux4_1
X_3213_ net1148 net1112 Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q VPWR VGND sg13g2_dlhq_1
XFILLER_39_189 VPWR VGND sg13g2_decap_8
X_3075_ net1162 net1084 Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q VPWR VGND sg13g2_dlhq_1
X_3144_ net1158 net1099 Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q VPWR VGND sg13g2_dlhq_1
XFILLER_50_332 VPWR VGND sg13g2_fill_2
X_2026_ _0513_ VPWR _0514_ VGND net948 _0510_ sg13g2_o21ai_1
XFILLER_24_28 VPWR VGND sg13g2_fill_2
X_2928_ net1206 net1128 Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q VPWR VGND sg13g2_dlhq_1
X_2859_ UserCLK net471 _0017_ _2859_/Q_N Inst_RegFile_32x4.mem\[28\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_49_14 VPWR VGND sg13g2_decap_8
Xhold296 Inst_RegFile_32x4.mem\[27\]\[1\] VPWR VGND net794 sg13g2_dlygate4sd3_1
Xhold230 Inst_RegFile_32x4.mem\[2\]\[1\] VPWR VGND net728 sg13g2_dlygate4sd3_1
Xhold285 Inst_RegFile_32x4.mem\[19\]\[3\] VPWR VGND net783 sg13g2_dlygate4sd3_1
Xhold241 Inst_RegFile_32x4.mem\[0\]\[0\] VPWR VGND net739 sg13g2_dlygate4sd3_1
Xhold274 Inst_RegFile_32x4.mem\[29\]\[0\] VPWR VGND net772 sg13g2_dlygate4sd3_1
Xhold263 Inst_RegFile_32x4.mem\[20\]\[2\] VPWR VGND net761 sg13g2_dlygate4sd3_1
Xhold252 Inst_RegFile_32x4.mem\[15\]\[1\] VPWR VGND net750 sg13g2_dlygate4sd3_1
XFILLER_14_61 VPWR VGND sg13g2_fill_2
XFILLER_30_93 VPWR VGND sg13g2_fill_1
XFILLER_30_82 VPWR VGND sg13g2_fill_1
Xinput9 E2END[4] net9 VPWR VGND sg13g2_buf_1
XFILLER_44_192 VPWR VGND sg13g2_fill_1
XFILLER_32_332 VPWR VGND sg13g2_fill_1
X_2713_ net941 net821 _1102_ _0028_ VPWR VGND sg13g2_mux2_1
X_2644_ _1062_ _1061_ _1034_ VPWR VGND sg13g2_nand2_2
X_3693_ net71 net275 VPWR VGND sg13g2_buf_1
X_3762_ W6END[11] net346 VPWR VGND sg13g2_buf_1
XFILLER_58_0 VPWR VGND sg13g2_decap_8
X_1526_ VPWR _1148_ Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q VGND sg13g2_inv_1
X_2575_ Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q net1018 _0486_ Inst_RegFile_switch_matrix.JS2BEG2
+ _1016_ Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q Inst_RegFile_switch_matrix.W1BEG3
+ VPWR VGND sg13g2_mux4_1
Xoutput324 net324 W2BEG[5] VPWR VGND sg13g2_buf_1
Xoutput302 Inst_RegFile_switch_matrix.SS4BEG1 SS4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput313 net313 SS4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput357 net357 WW4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput335 net335 W6BEG[0] VPWR VGND sg13g2_buf_1
Xoutput346 net346 W6BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_55_479 VPWR VGND sg13g2_fill_2
XFILLER_55_402 VPWR VGND sg13g2_fill_2
X_3127_ net1190 net1094 Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q VPWR VGND sg13g2_dlhq_1
X_3058_ net1201 net1085 Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q VPWR VGND sg13g2_dlhq_1
XFILLER_51_48 VPWR VGND sg13g2_fill_1
X_2009_ VGND VPWR Inst_RegFile_32x4.mem\[25\]\[0\] net993 _0499_ _0498_ sg13g2_a21oi_1
XFILLER_46_413 VPWR VGND sg13g2_fill_2
XFILLER_41_81 VPWR VGND sg13g2_fill_1
XFILLER_25_82 VPWR VGND sg13g2_fill_2
XFILLER_51_7 VPWR VGND sg13g2_decap_8
X_2291_ Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q VPWR _0762_ VGND net1059 net987
+ sg13g2_o21ai_1
X_2360_ Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q VPWR _0827_ VGND _0824_ _0821_ sg13g2_o21ai_1
XFILLER_2_42 VPWR VGND sg13g2_fill_1
Xoutput143 net143 EE4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput132 Inst_RegFile_switch_matrix.E6BEG1 E6BEG[11] VPWR VGND sg13g2_buf_1
X_2627_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q _1044_ _1045_ Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q
+ sg13g2_a21oi_1
Xoutput121 net121 E2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput110 Inst_RegFile_switch_matrix.E1BEG0 E1BEG[0] VPWR VGND sg13g2_buf_1
X_3745_ net97 net327 VPWR VGND sg13g2_buf_1
Xoutput187 net187 FrameData_O[7] VPWR VGND sg13g2_buf_1
Xoutput198 net198 FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
Xoutput176 net176 FrameData_O[26] VPWR VGND sg13g2_buf_1
X_2489_ Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q net30 net1 net86 net974 Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q
+ _0944_ VPWR VGND sg13g2_mux4_1
Xoutput165 net165 FrameData_O[16] VPWR VGND sg13g2_buf_1
Xoutput154 net154 EE4BEG[6] VPWR VGND sg13g2_buf_1
X_2558_ _0999_ _1002_ _1003_ VPWR VGND sg13g2_nor2_1
XFILLER_3_512 VPWR VGND sg13g2_fill_2
X_1860_ _0350_ _0355_ _0356_ VPWR VGND sg13g2_nor2_2
Xinput78 S4END[0] net78 VPWR VGND sg13g2_buf_1
Xinput67 S2END[5] net67 VPWR VGND sg13g2_buf_1
Xinput12 E2END[7] net12 VPWR VGND sg13g2_buf_1
Xinput23 EE4END[2] net23 VPWR VGND sg13g2_buf_1
Xinput45 N2MID[3] net45 VPWR VGND sg13g2_buf_1
Xinput34 N2END[0] net34 VPWR VGND sg13g2_buf_1
Xinput56 NN4END[2] net56 VPWR VGND sg13g2_buf_1
X_1791_ net921 Inst_RegFile_32x4.mem\[2\]\[2\] Inst_RegFile_32x4.mem\[3\]\[2\] Inst_RegFile_32x4.mem\[0\]\[2\]
+ Inst_RegFile_32x4.mem\[1\]\[2\] net1022 _0291_ VPWR VGND sg13g2_mux4_1
XFILLER_6_383 VPWR VGND sg13g2_fill_1
Xinput89 W2END[0] net89 VPWR VGND sg13g2_buf_1
X_2343_ _0810_ VPWR _0811_ VGND Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q _0809_
+ sg13g2_o21ai_1
X_2412_ Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q _0875_ _0874_ _0872_ _0873_ Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q
+ _0876_ VPWR VGND sg13g2_mux4_1
X_2274_ _0740_ Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q _0745_ _0746_ VPWR VGND sg13g2_nand3_1
X_1989_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q _0477_ _0480_ _1132_
+ sg13g2_a21oi_1
X_3659_ N4END[15] net232 VPWR VGND sg13g2_buf_1
XFILLER_57_14 VPWR VGND sg13g2_decap_4
Xfanout1165 FrameData[30] net1165 VPWR VGND sg13g2_buf_1
Xfanout1132 net1135 net1132 VPWR VGND sg13g2_buf_1
Xfanout1110 net1114 net1110 VPWR VGND sg13g2_buf_1
Xfanout1143 net1147 net1143 VPWR VGND sg13g2_buf_1
XFILLER_3_342 VPWR VGND sg13g2_fill_2
Xfanout1154 net1155 net1154 VPWR VGND sg13g2_buf_1
Xfanout1121 net1125 net1121 VPWR VGND sg13g2_buf_1
Xfanout1187 FrameData[20] net1187 VPWR VGND sg13g2_buf_1
Xfanout1176 FrameData[25] net1176 VPWR VGND sg13g2_buf_1
XFILLER_34_202 VPWR VGND sg13g2_fill_1
Xfanout1198 net1200 net1198 VPWR VGND sg13g2_buf_1
X_1843_ VPWR _0339_ _0338_ VGND sg13g2_inv_1
X_1912_ _0406_ _0405_ Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q VPWR VGND sg13g2_nand2b_1
X_2961_ net1203 net1132 Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q VPWR VGND sg13g2_dlhq_1
XFILLER_30_496 VPWR VGND sg13g2_fill_1
X_2892_ UserCLK net430 _0050_ _2892_/Q_N Inst_RegFile_32x4.mem\[14\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_8_52 VPWR VGND sg13g2_fill_1
XFILLER_40_0 VPWR VGND sg13g2_decap_8
X_1774_ net922 Inst_RegFile_32x4.mem\[30\]\[1\] Inst_RegFile_32x4.mem\[31\]\[1\] Inst_RegFile_32x4.mem\[28\]\[1\]
+ Inst_RegFile_32x4.mem\[29\]\[1\] net1025 _0276_ VPWR VGND sg13g2_mux4_1
X_3375_ UserCLK net369 _0111_ _3375_/Q_N Inst_RegFile_32x4.mem\[8\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_2326_ _0795_ _0792_ Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q VPWR VGND sg13g2_nand2_2
X_2257_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q _0730_ net1010 net1045
+ sg13g2_a21oi_2
XFILLER_53_511 VPWR VGND sg13g2_fill_1
X_2188_ _0665_ net1031 net1044 VPWR VGND sg13g2_nand2b_1
XFILLER_40_249 VPWR VGND sg13g2_decap_8
XFILLER_29_530 VPWR VGND sg13g2_fill_1
XFILLER_12_441 VPWR VGND sg13g2_fill_1
X_2111_ _0586_ _0592_ Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q _0593_ VPWR VGND
+ sg13g2_nand3_1
XFILLER_39_305 VPWR VGND sg13g2_decap_4
X_3160_ net1186 net1098 Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q VPWR VGND sg13g2_dlhq_1
X_2042_ VGND VPWR net1006 _0529_ _0530_ net943 sg13g2_a21oi_1
X_3091_ net1198 net1088 Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q VPWR VGND sg13g2_dlhq_1
XFILLER_47_360 VPWR VGND sg13g2_fill_2
X_2944_ net1170 net27 Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q VPWR VGND sg13g2_dlhq_1
X_1826_ VGND VPWR Inst_RegFile_32x4.mem\[25\]\[3\] net928 _0324_ _0323_ sg13g2_a21oi_1
X_2875_ UserCLK net455 _0033_ _2875_/Q_N Inst_RegFile_32x4.mem\[13\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_1688_ _0193_ VPWR _0194_ VGND net1054 net976 sg13g2_o21ai_1
Xfanout947 net948 net947 VPWR VGND sg13g2_buf_1
Xfanout958 net962 net958 VPWR VGND sg13g2_buf_1
Xfanout925 net927 net925 VPWR VGND sg13g2_buf_1
Xfanout936 _1087_ net936 VPWR VGND sg13g2_buf_2
X_1757_ _0261_ _0260_ _0255_ VPWR VGND sg13g2_nand2b_1
X_3358_ UserCLK net386 _0094_ _3358_/Q_N Inst_RegFile_32x4.mem\[4\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_3289_ net1185 net1126 Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q VPWR VGND sg13g2_dlhq_1
X_2309_ net986 net1037 _0779_ VPWR VGND sg13g2_nor2b_1
Xfanout969 net520 net969 VPWR VGND sg13g2_buf_8
XFILLER_48_102 VPWR VGND sg13g2_fill_2
XFILLER_32_503 VPWR VGND sg13g2_fill_1
X_1611_ _1230_ _1229_ Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q VPWR VGND sg13g2_nand2b_1
X_2660_ Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q VPWR _1075_ VGND Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q
+ _0935_ sg13g2_o21ai_1
X_3212_ net1150 net1112 Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q VPWR VGND sg13g2_dlhq_1
X_1542_ net1015 _1164_ VPWR VGND sg13g2_inv_16
XFILLER_5_20 VPWR VGND sg13g2_fill_1
X_2591_ Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q net1034 _0645_ Inst_RegFile_switch_matrix.JN2BEG0
+ _0137_ Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q Inst_RegFile_switch_matrix.E1BEG1
+ VPWR VGND sg13g2_mux4_1
XFILLER_54_127 VPWR VGND sg13g2_fill_1
X_2025_ VGND VPWR net948 _0512_ _0513_ net1009 sg13g2_a21oi_1
X_3143_ net1161 net1100 Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q VPWR VGND sg13g2_dlhq_1
X_3074_ net1164 net1083 Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q VPWR VGND sg13g2_dlhq_1
XFILLER_50_311 VPWR VGND sg13g2_decap_8
X_2927_ net1208 net1128 Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q VPWR VGND sg13g2_dlhq_1
XFILLER_40_39 VPWR VGND sg13g2_decap_8
Xhold242 Inst_RegFile_32x4.mem\[13\]\[0\] VPWR VGND net740 sg13g2_dlygate4sd3_1
Xhold231 Inst_RegFile_32x4.mem\[6\]\[2\] VPWR VGND net729 sg13g2_dlygate4sd3_1
X_2877__453 VPWR VGND net453 sg13g2_tiehi
X_2789_ net959 net829 _1120_ _0086_ VPWR VGND sg13g2_mux2_1
X_1809_ _0309_ _0308_ net1024 VPWR VGND sg13g2_nand2b_1
Xhold253 Inst_RegFile_32x4.mem\[13\]\[1\] VPWR VGND net751 sg13g2_dlygate4sd3_1
X_2858_ UserCLK net472 _0016_ _2858_/Q_N Inst_RegFile_32x4.mem\[28\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
Xhold275 Inst_RegFile_32x4.mem\[1\]\[3\] VPWR VGND net773 sg13g2_dlygate4sd3_1
Xhold286 Inst_RegFile_32x4.mem\[1\]\[2\] VPWR VGND net784 sg13g2_dlygate4sd3_1
Xhold297 Inst_RegFile_32x4.mem\[22\]\[3\] VPWR VGND net795 sg13g2_dlygate4sd3_1
Xhold264 Inst_RegFile_32x4.mem\[20\]\[0\] VPWR VGND net762 sg13g2_dlygate4sd3_1
XFILLER_41_322 VPWR VGND sg13g2_fill_2
XFILLER_26_363 VPWR VGND sg13g2_fill_1
XFILLER_55_80 VPWR VGND sg13g2_fill_2
X_3761_ W6END[10] net345 VPWR VGND sg13g2_buf_1
Xoutput314 net314 UserCLKo VPWR VGND sg13g2_buf_1
X_2712_ _1102_ _1088_ _1101_ VPWR VGND sg13g2_nand2_2
X_2643_ _1058_ _1048_ _1059_ _1061_ VPWR VGND sg13g2_nor3_2
X_2574_ Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q net57 net81 net106 Inst_RegFile_switch_matrix.JN2BEG1
+ Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q _1016_ VPWR VGND sg13g2_mux4_1
Xoutput325 net325 W2BEG[6] VPWR VGND sg13g2_buf_1
Xoutput303 net303 SS4BEG[14] VPWR VGND sg13g2_buf_1
X_3692_ net70 net274 VPWR VGND sg13g2_buf_1
XFILLER_59_208 VPWR VGND sg13g2_fill_1
X_1525_ VPWR _1147_ Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q VGND sg13g2_inv_1
Xoutput347 net347 WW4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput358 net358 WW4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput336 net336 W6BEG[10] VPWR VGND sg13g2_buf_1
XFILLER_55_458 VPWR VGND sg13g2_decap_8
XFILLER_42_108 VPWR VGND sg13g2_fill_1
X_2008_ net996 Inst_RegFile_32x4.mem\[24\]\[0\] _0498_ VPWR VGND sg13g2_nor2b_1
X_3126_ net1192 net1094 Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q VPWR VGND sg13g2_dlhq_1
XFILLER_27_127 VPWR VGND sg13g2_fill_1
X_3057_ net1204 net1086 Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q VPWR VGND sg13g2_dlhq_1
XFILLER_41_130 VPWR VGND sg13g2_fill_2
X_2290_ _0760_ VPWR _0761_ VGND net1059 net1031 sg13g2_o21ai_1
XFILLER_37_425 VPWR VGND sg13g2_fill_1
X_3744_ Inst_RegFile_switch_matrix.JW2BEG7 net326 VPWR VGND sg13g2_buf_2
X_2867__463 VPWR VGND net463 sg13g2_tiehi
XFILLER_20_336 VPWR VGND sg13g2_fill_2
Xoutput166 net166 FrameData_O[17] VPWR VGND sg13g2_buf_1
Xoutput177 net177 FrameData_O[27] VPWR VGND sg13g2_buf_1
X_2557_ Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q VPWR _1002_ VGND Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q
+ _1001_ sg13g2_o21ai_1
Xoutput144 net144 EE4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput133 net133 E6BEG[1] VPWR VGND sg13g2_buf_1
X_2874__456 VPWR VGND net456 sg13g2_tiehi
X_2626_ VPWR _1044_ _1043_ VGND sg13g2_inv_1
Xoutput155 net155 EE4BEG[7] VPWR VGND sg13g2_buf_1
X_3675_ NN4END[15] net248 VPWR VGND sg13g2_buf_1
Xoutput111 Inst_RegFile_switch_matrix.E1BEG1 E1BEG[1] VPWR VGND sg13g2_buf_1
Xoutput122 net122 E2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput199 net199 FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
X_2488_ _0939_ _0942_ _0943_ VPWR VGND sg13g2_nor2_1
Xoutput188 net188 FrameData_O[8] VPWR VGND sg13g2_buf_1
X_3109_ net1189 net1095 Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q VPWR VGND sg13g2_dlhq_1
X_2881__449 VPWR VGND net449 sg13g2_tiehi
XFILLER_51_494 VPWR VGND sg13g2_fill_1
XFILLER_36_71 VPWR VGND sg13g2_fill_2
XFILLER_34_428 VPWR VGND sg13g2_fill_1
Xinput13 E2MID[0] net13 VPWR VGND sg13g2_buf_1
X_1790_ VGND VPWR net982 _0289_ _0290_ net969 sg13g2_a21oi_1
Xinput79 S4END[1] net79 VPWR VGND sg13g2_buf_1
Xinput68 S2END[6] net68 VPWR VGND sg13g2_buf_1
X_2411_ net1076 net34 net1051 _0875_ VPWR VGND sg13g2_mux2_1
Xinput24 EE4END[3] net24 VPWR VGND sg13g2_buf_1
X_3391_ UserCLK net489 _0127_ _3391_/Q_N Inst_RegFile_32x4.mem\[12\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
Xinput46 N2MID[4] net46 VPWR VGND sg13g2_buf_1
Xinput35 N2END[1] net35 VPWR VGND sg13g2_buf_1
Xinput57 NN4END[3] net57 VPWR VGND sg13g2_buf_8
X_2342_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q _0807_ _0810_ Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q
+ sg13g2_a21oi_1
XFILLER_37_233 VPWR VGND sg13g2_fill_2
X_2273_ Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q _0744_ _0742_ _0745_ VPWR VGND sg13g2_nand3_1
X_3727_ SS4END[15] net300 VPWR VGND sg13g2_buf_1
X_1988_ VGND VPWR net1053 net61 _0479_ _0478_ sg13g2_a21oi_1
XFILLER_20_111 VPWR VGND sg13g2_fill_2
X_3658_ N4END[14] net231 VPWR VGND sg13g2_buf_1
X_2609_ Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q net50 net1066 net82 Inst_RegFile_switch_matrix.JW2BEG2
+ Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q _1027_ VPWR VGND sg13g2_mux4_1
X_3589_ net1205 net162 VPWR VGND sg13g2_buf_1
XFILLER_3_354 VPWR VGND sg13g2_fill_1
X_2857__473 VPWR VGND net473 sg13g2_tiehi
Xfanout1133 net1135 net1133 VPWR VGND sg13g2_buf_1
Xfanout1177 FrameData[25] net1177 VPWR VGND sg13g2_buf_1
Xfanout1111 net1113 net1111 VPWR VGND sg13g2_buf_1
Xfanout1155 net25 net1155 VPWR VGND sg13g2_buf_1
Xfanout1188 FrameData[1] net1188 VPWR VGND sg13g2_buf_1
Xfanout1100 net1101 net1100 VPWR VGND sg13g2_buf_1
Xfanout1199 net1200 net1199 VPWR VGND sg13g2_buf_1
Xfanout1144 net1146 net1144 VPWR VGND sg13g2_buf_1
XFILLER_0_0 VPWR VGND sg13g2_fill_2
XFILLER_14_8 VPWR VGND sg13g2_fill_1
Xfanout1166 net1167 net1166 VPWR VGND sg13g2_buf_1
Xfanout1122 net1125 net1122 VPWR VGND sg13g2_buf_1
X_2960_ net1207 net1132 Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q VPWR VGND sg13g2_dlhq_1
X_1911_ _0403_ _0404_ Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q _0405_ VPWR VGND
+ sg13g2_mux2_1
X_1842_ Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q net45 net16 net73 net100 Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q
+ _0338_ VPWR VGND sg13g2_mux4_1
X_1773_ _0274_ VPWR _0275_ VGND net1028 _0273_ sg13g2_o21ai_1
X_2864__466 VPWR VGND net466 sg13g2_tiehi
X_2891_ UserCLK net431 _0049_ _2891_/Q_N Inst_RegFile_32x4.mem\[14\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_3374_ UserCLK net370 _0110_ _3374_/Q_N Inst_RegFile_32x4.mem\[8\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_2871__459 VPWR VGND net459 sg13g2_tiehi
X_2187_ _0664_ net1044 net1013 VPWR VGND sg13g2_nand2_1
X_2325_ VGND VPWR net1041 net999 _0794_ _0793_ sg13g2_a21oi_1
X_2256_ VGND VPWR net1045 net999 _0729_ _0728_ sg13g2_a21oi_1
XFILLER_16_258 VPWR VGND sg13g2_fill_1
XFILLER_8_457 VPWR VGND sg13g2_fill_2
X_2110_ _0591_ VPWR _0592_ VGND Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q _0590_
+ sg13g2_o21ai_1
X_2041_ net998 Inst_RegFile_32x4.mem\[4\]\[1\] Inst_RegFile_32x4.mem\[5\]\[1\] Inst_RegFile_32x4.mem\[6\]\[1\]
+ Inst_RegFile_32x4.mem\[7\]\[1\] net948 _0529_ VPWR VGND sg13g2_mux4_1
X_3090_ net1201 net1088 Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q VPWR VGND sg13g2_dlhq_1
X_2943_ net1172 net1130 Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q VPWR VGND sg13g2_dlhq_1
X_1825_ net928 Inst_RegFile_32x4.mem\[24\]\[3\] _0323_ VPWR VGND sg13g2_nor2b_1
X_2874_ UserCLK net456 _0032_ _2874_/Q_N Inst_RegFile_32x4.mem\[13\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_1756_ _0259_ VPWR _0260_ VGND net1024 _0256_ sg13g2_o21ai_1
X_1687_ _0193_ net1054 net966 VPWR VGND sg13g2_nand2_1
X_2308_ VGND VPWR _0776_ _0777_ _0778_ Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q
+ sg13g2_a21oi_1
Xfanout948 _0368_ net948 VPWR VGND sg13g2_buf_1
X_3357_ UserCLK net387 _0093_ _3357_/Q_N Inst_RegFile_32x4.mem\[4\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
Xfanout926 net927 net926 VPWR VGND sg13g2_buf_1
Xfanout937 net938 net937 VPWR VGND sg13g2_buf_1
Xfanout959 net962 net959 VPWR VGND sg13g2_buf_1
X_3288_ net1187 net1126 Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q VPWR VGND sg13g2_dlhq_1
X_2239_ _0712_ VPWR _0713_ VGND Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q _0711_ sg13g2_o21ai_1
X_2847__483 VPWR VGND net483 sg13g2_tiehi
X_2854__476 VPWR VGND net476 sg13g2_tiehi
X_1610_ Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q net46 net101 net74 Inst_RegFile_switch_matrix.JS2BEG5
+ Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q _1229_ VPWR VGND sg13g2_mux4_1
X_2861__469 VPWR VGND net469 sg13g2_tiehi
X_2590_ Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q net1012 _0338_ Inst_RegFile_switch_matrix.JN2BEG1
+ net522 Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q Inst_RegFile_switch_matrix.E1BEG2
+ VPWR VGND sg13g2_mux4_1
X_3142_ net1167 net1100 Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q VPWR VGND sg13g2_dlhq_1
X_3211_ net1153 net1109 Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q VPWR VGND sg13g2_dlhq_1
XFILLER_4_460 VPWR VGND sg13g2_fill_1
X_1541_ VPWR _1163_ Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q VGND sg13g2_inv_1
X_2024_ _0511_ VPWR _0512_ VGND Inst_RegFile_32x4.mem\[26\]\[1\] net998 sg13g2_o21ai_1
X_3073_ net1168 net1084 Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q VPWR VGND sg13g2_dlhq_1
XFILLER_50_334 VPWR VGND sg13g2_fill_1
X_2857_ UserCLK net473 _0015_ _2857_/Q_N Inst_RegFile_32x4.mem\[27\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_2926_ net1211 net1128 Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q VPWR VGND sg13g2_dlhq_1
Xhold232 Inst_RegFile_32x4.mem\[8\]\[2\] VPWR VGND net730 sg13g2_dlygate4sd3_1
X_1739_ net930 Inst_RegFile_32x4.mem\[4\]\[0\] _0243_ VPWR VGND sg13g2_nor2b_1
Xhold243 Inst_RegFile_32x4.mem\[13\]\[3\] VPWR VGND net741 sg13g2_dlygate4sd3_1
X_1808_ VGND VPWR Inst_RegFile_32x4.mem\[23\]\[2\] net923 _0308_ _0307_ sg13g2_a21oi_1
Xhold265 Inst_RegFile_32x4.mem\[20\]\[1\] VPWR VGND net763 sg13g2_dlygate4sd3_1
Xhold287 Inst_RegFile_32x4.mem\[17\]\[2\] VPWR VGND net785 sg13g2_dlygate4sd3_1
Xhold276 Inst_RegFile_32x4.mem\[16\]\[0\] VPWR VGND net774 sg13g2_dlygate4sd3_1
X_2788_ net950 net827 _1120_ _0085_ VPWR VGND sg13g2_mux2_1
Xhold254 Inst_RegFile_32x4.mem\[15\]\[2\] VPWR VGND net752 sg13g2_dlygate4sd3_1
XFILLER_58_489 VPWR VGND sg13g2_fill_2
XFILLER_58_445 VPWR VGND sg13g2_decap_4
XFILLER_58_412 VPWR VGND sg13g2_fill_2
Xhold298 Inst_RegFile_32x4.mem\[11\]\[1\] VPWR VGND net796 sg13g2_dlygate4sd3_1
XFILLER_14_63 VPWR VGND sg13g2_fill_1
XFILLER_49_412 VPWR VGND sg13g2_decap_8
XFILLER_30_73 VPWR VGND sg13g2_decap_8
XFILLER_5_268 VPWR VGND sg13g2_fill_2
XFILLER_39_82 VPWR VGND sg13g2_fill_2
X_3760_ W6END[9] net344 VPWR VGND sg13g2_buf_1
X_2711_ _1033_ _1100_ _1101_ VPWR VGND sg13g2_nor2_1
XFILLER_9_530 VPWR VGND sg13g2_fill_1
X_3691_ Inst_RegFile_switch_matrix.JS2BEG7 net273 VPWR VGND sg13g2_buf_8
X_2573_ VGND VPWR _1015_ Inst_RegFile_switch_matrix.NN4BEG0 _1013_ _1009_ sg13g2_a21oi_2
X_2642_ VPWR _1060_ _1059_ VGND sg13g2_inv_1
X_1524_ VPWR _1146_ Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q VGND sg13g2_inv_1
Xoutput326 net326 W2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput304 net304 SS4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput315 Inst_RegFile_switch_matrix.W1BEG0 W1BEG[0] VPWR VGND sg13g2_buf_1
Xoutput359 net359 WW4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput348 net348 WW4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput337 Inst_RegFile_switch_matrix.W6BEG1 W6BEG[11] VPWR VGND sg13g2_buf_1
XFILLER_55_415 VPWR VGND sg13g2_decap_8
X_3125_ net1195 net1095 Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q VPWR VGND sg13g2_dlhq_1
XFILLER_35_183 VPWR VGND sg13g2_fill_2
X_2007_ _0497_ _0494_ _0496_ _0462_ _0460_ VPWR VGND sg13g2_a22oi_1
X_3056_ net1207 net1086 Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q VPWR VGND sg13g2_dlhq_1
X_2844__486 VPWR VGND net486 sg13g2_tiehi
X_2909_ UserCLK net413 _0067_ _2909_/Q_N Inst_RegFile_32x4.mem\[1\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_3389__491 VPWR VGND net491 sg13g2_tiehi
X_2851__479 VPWR VGND net479 sg13g2_tiehi
XFILLER_33_109 VPWR VGND sg13g2_decap_4
XFILLER_14_301 VPWR VGND sg13g2_fill_1
XFILLER_14_312 VPWR VGND sg13g2_fill_1
XFILLER_2_77 VPWR VGND sg13g2_fill_2
XFILLER_24_109 VPWR VGND sg13g2_fill_1
XFILLER_17_183 VPWR VGND sg13g2_decap_8
XFILLER_17_194 VPWR VGND sg13g2_fill_1
X_3674_ NN4END[14] net247 VPWR VGND sg13g2_buf_1
X_3743_ net722 net325 VPWR VGND sg13g2_buf_8
XFILLER_9_371 VPWR VGND sg13g2_fill_1
Xoutput178 net178 FrameData_O[28] VPWR VGND sg13g2_buf_1
Xoutput189 net189 FrameData_O[9] VPWR VGND sg13g2_buf_1
Xoutput167 net167 FrameData_O[18] VPWR VGND sg13g2_buf_1
X_2556_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q _1182_ _1001_ _1000_
+ sg13g2_a21oi_1
Xoutput145 Inst_RegFile_switch_matrix.EE4BEG0 EE4BEG[12] VPWR VGND sg13g2_buf_1
X_2487_ Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q VPWR _0942_ VGND Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q
+ _0941_ sg13g2_o21ai_1
Xoutput156 net156 EE4BEG[8] VPWR VGND sg13g2_buf_1
X_2625_ Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q net49 net20 net77 net104 Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q
+ _1043_ VPWR VGND sg13g2_mux4_1
Xoutput134 net134 E6BEG[2] VPWR VGND sg13g2_buf_1
Xoutput112 Inst_RegFile_switch_matrix.E1BEG2 E1BEG[2] VPWR VGND sg13g2_buf_1
Xoutput123 net123 E2BEGb[1] VPWR VGND sg13g2_buf_1
X_3108_ net1212 net1095 Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q VPWR VGND sg13g2_dlhq_1
XFILLER_43_407 VPWR VGND sg13g2_fill_1
X_3039_ net1172 net1077 Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q VPWR VGND sg13g2_dlhq_1
XFILLER_34_407 VPWR VGND sg13g2_fill_2
Xinput25 FrameData[6] net25 VPWR VGND sg13g2_buf_1
Xinput14 E2MID[1] net14 VPWR VGND sg13g2_buf_1
Xinput36 N2END[2] net36 VPWR VGND sg13g2_buf_1
Xinput69 S2END[7] net69 VPWR VGND sg13g2_buf_1
X_2341_ VGND VPWR net1042 net506 _0809_ _0808_ sg13g2_a21oi_1
X_2410_ net54 net1221 Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q _0874_ VPWR VGND
+ sg13g2_mux2_1
Xinput58 S1END[0] net58 VPWR VGND sg13g2_buf_1
X_3390_ UserCLK net490 _0126_ _3390_/Q_N Inst_RegFile_32x4.mem\[12\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
Xinput47 N2MID[5] net47 VPWR VGND sg13g2_buf_1
X_2272_ net999 net1050 _0743_ _0744_ VPWR VGND sg13g2_a21o_1
XFILLER_52_248 VPWR VGND sg13g2_fill_1
XFILLER_33_462 VPWR VGND sg13g2_fill_2
XFILLER_18_492 VPWR VGND sg13g2_fill_2
X_3726_ SS4END[14] net299 VPWR VGND sg13g2_buf_1
X_1987_ net1053 net12 _0478_ VPWR VGND sg13g2_nor2b_1
X_2880__450 VPWR VGND net450 sg13g2_tiehi
X_3657_ N4END[13] net245 VPWR VGND sg13g2_buf_1
X_2539_ Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q net1076 net1221 net58 net974 Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q
+ _0988_ VPWR VGND sg13g2_mux4_1
XFILLER_0_528 VPWR VGND sg13g2_fill_2
X_3588_ net1207 net161 VPWR VGND sg13g2_buf_1
X_2608_ _1020_ _1025_ _1026_ VPWR VGND sg13g2_and2_1
X_3386__494 VPWR VGND net494 sg13g2_tiehi
XFILLER_11_123 VPWR VGND sg13g2_fill_2
XFILLER_59_392 VPWR VGND sg13g2_decap_8
Xfanout1112 net1113 net1112 VPWR VGND sg13g2_buf_1
Xfanout1123 net1124 net1123 VPWR VGND sg13g2_buf_1
Xfanout1178 FrameData[24] net1178 VPWR VGND sg13g2_buf_1
Xfanout1189 FrameData[1] net1189 VPWR VGND sg13g2_buf_1
Xfanout1134 net1135 net1134 VPWR VGND sg13g2_buf_1
Xfanout1101 net1102 net1101 VPWR VGND sg13g2_buf_1
Xfanout1145 net1146 net1145 VPWR VGND sg13g2_buf_1
Xfanout1156 net1157 net1156 VPWR VGND sg13g2_buf_1
Xfanout1167 FrameData[2] net1167 VPWR VGND sg13g2_buf_1
XFILLER_47_93 VPWR VGND sg13g2_fill_2
X_1910_ net1043 net59 net67 net85 net1071 Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q
+ _0404_ VPWR VGND sg13g2_mux4_1
X_2890_ UserCLK net432 _0048_ _2890_/Q_N Inst_RegFile_32x4.mem\[14\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_1772_ VGND VPWR net1028 _0272_ _0274_ net983 sg13g2_a21oi_1
X_1841_ Inst_RegFile_32x4.AD_comb\[3\] Inst_RegFile_32x4.AD_reg\[3\] Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q
+ AD3 VPWR VGND sg13g2_mux2_2
X_3373_ UserCLK net371 _0109_ _3373_/Q_N Inst_RegFile_32x4.mem\[8\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_26_0 VPWR VGND sg13g2_fill_1
X_2324_ Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q VPWR _0793_ VGND net1041 net984
+ sg13g2_o21ai_1
X_2186_ Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q VPWR _0663_ VGND net1044 net987
+ sg13g2_o21ai_1
X_2255_ Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q VPWR _0728_ VGND net1045 net984
+ sg13g2_o21ai_1
X_3709_ S4END[13] net297 VPWR VGND sg13g2_buf_1
XFILLER_56_395 VPWR VGND sg13g2_decap_8
X_2870__460 VPWR VGND net460 sg13g2_tiehi
XFILLER_47_384 VPWR VGND sg13g2_fill_2
XFILLER_47_351 VPWR VGND sg13g2_fill_1
X_2040_ _0528_ _0527_ net1006 VPWR VGND sg13g2_nand2b_1
X_2942_ net1174 net27 Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q VPWR VGND sg13g2_dlhq_1
X_2873_ UserCLK net457 _0031_ _2873_/Q_N Inst_RegFile_32x4.mem\[9\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_30_273 VPWR VGND sg13g2_decap_4
X_1824_ Inst_RegFile_32x4.mem\[26\]\[3\] Inst_RegFile_32x4.mem\[27\]\[3\] net928 _0322_
+ VPWR VGND sg13g2_mux2_1
X_1686_ _0192_ _0191_ _0144_ VPWR VGND sg13g2_nand2b_1
X_1755_ VGND VPWR net1024 _0258_ _0259_ net955 sg13g2_a21oi_1
X_2307_ _0777_ net971 net1037 VPWR VGND sg13g2_nand2b_1
Xfanout927 A_ADR0 net927 VPWR VGND sg13g2_buf_1
X_3356_ UserCLK net388 _0092_ _3356_/Q_N Inst_RegFile_32x4.mem\[4\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_3287_ net1191 net1125 Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q VPWR VGND sg13g2_dlhq_1
Xfanout949 net951 net949 VPWR VGND sg13g2_buf_1
X_2238_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q _0709_ _0712_ Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q
+ sg13g2_a21oi_1
Xfanout938 net939 net938 VPWR VGND sg13g2_buf_1
XFILLER_54_28 VPWR VGND sg13g2_fill_2
X_3383__497 VPWR VGND net497 sg13g2_tiehi
X_2169_ Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q net105 net1017 net978 net971 Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q
+ _0647_ VPWR VGND sg13g2_mux4_1
XFILLER_0_111 VPWR VGND sg13g2_fill_2
XFILLER_48_148 VPWR VGND sg13g2_fill_2
XFILLER_44_354 VPWR VGND sg13g2_fill_2
X_1540_ VPWR _1162_ Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q VGND sg13g2_inv_1
X_3141_ net1189 net1102 Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q VPWR VGND sg13g2_dlhq_1
X_3210_ net1155 net1109 Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q VPWR VGND sg13g2_dlhq_1
X_2023_ _0511_ net998 Inst_RegFile_32x4.mem\[27\]\[1\] VPWR VGND sg13g2_nand2b_1
XFILLER_35_310 VPWR VGND sg13g2_fill_2
X_3072_ net1170 net1083 Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q VPWR VGND sg13g2_dlhq_1
X_2856_ UserCLK net474 _0014_ _2856_/Q_N Inst_RegFile_32x4.mem\[27\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_2925_ net1149 net1129 Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q VPWR VGND sg13g2_dlhq_1
X_1807_ net923 Inst_RegFile_32x4.mem\[22\]\[2\] _0307_ VPWR VGND sg13g2_nor2b_1
X_1669_ Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q net32 net40 net3 net11 Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q
+ _0176_ VPWR VGND sg13g2_mux4_1
Xhold233 Inst_RegFile_32x4.mem\[8\]\[0\] VPWR VGND net731 sg13g2_dlygate4sd3_1
XFILLER_49_28 VPWR VGND sg13g2_fill_2
X_1738_ Inst_RegFile_32x4.mem\[6\]\[0\] Inst_RegFile_32x4.mem\[7\]\[0\] net930 _0242_
+ VPWR VGND sg13g2_mux2_1
Xhold299 Inst_RegFile_32x4.mem\[5\]\[3\] VPWR VGND net797 sg13g2_dlygate4sd3_1
Xhold288 Inst_RegFile_32x4.mem\[7\]\[3\] VPWR VGND net786 sg13g2_dlygate4sd3_1
Xhold244 Inst_RegFile_32x4.mem\[0\]\[2\] VPWR VGND net742 sg13g2_dlygate4sd3_1
X_2787_ net937 net824 _1120_ _0084_ VPWR VGND sg13g2_mux2_1
Xhold277 Inst_RegFile_32x4.mem\[30\]\[0\] VPWR VGND net775 sg13g2_dlygate4sd3_1
Xhold266 Inst_RegFile_32x4.mem\[5\]\[2\] VPWR VGND net764 sg13g2_dlygate4sd3_1
Xhold255 Inst_RegFile_32x4.mem\[13\]\[2\] VPWR VGND net753 sg13g2_dlygate4sd3_1
X_3339_ UserCLK net405 Inst_RegFile_32x4.AD_comb\[3\] _3339_/Q_N Inst_RegFile_32x4.AD_reg\[3\]
+ VPWR VGND sg13g2_dfrbp_1
X_2860__470 VPWR VGND net470 sg13g2_tiehi
XFILLER_17_321 VPWR VGND sg13g2_fill_1
XFILLER_17_343 VPWR VGND sg13g2_fill_1
X_3690_ Inst_RegFile_switch_matrix.JS2BEG6 net272 VPWR VGND sg13g2_buf_1
X_2710_ _1100_ _1029_ _1026_ VPWR VGND sg13g2_nand2b_1
X_2572_ Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q _1014_ _1015_ VPWR VGND sg13g2_nor2_1
X_2641_ Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q _1053_ _0997_ _0910_ _1017_ Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q
+ _1059_ VPWR VGND sg13g2_mux4_1
X_1523_ VPWR _1145_ Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q VGND sg13g2_inv_1
Xoutput316 Inst_RegFile_switch_matrix.W1BEG1 W1BEG[1] VPWR VGND sg13g2_buf_1
Xoutput327 net327 W2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput305 net305 SS4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput338 net338 W6BEG[1] VPWR VGND sg13g2_buf_1
Xoutput349 net349 WW4BEG[11] VPWR VGND sg13g2_buf_1
X_3124_ net1197 net1097 Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q VPWR VGND sg13g2_dlhq_1
X_3055_ net1209 net1086 Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q VPWR VGND sg13g2_dlhq_1
XFILLER_51_18 VPWR VGND sg13g2_fill_1
X_2006_ VGND VPWR net1007 _0495_ _0496_ _0460_ sg13g2_a21oi_1
X_2908_ UserCLK net414 _0066_ _2908_/Q_N Inst_RegFile_32x4.mem\[1\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_2839_ net954 net771 _1131_ _0125_ VPWR VGND sg13g2_mux2_1
XFILLER_4_8 VPWR VGND sg13g2_fill_2
XFILLER_2_217 VPWR VGND sg13g2_fill_1
XFILLER_54_460 VPWR VGND sg13g2_decap_8
XFILLER_10_530 VPWR VGND sg13g2_fill_1
XFILLER_41_95 VPWR VGND sg13g2_fill_1
XFILLER_49_221 VPWR VGND sg13g2_fill_1
XFILLER_52_419 VPWR VGND sg13g2_decap_8
XFILLER_32_143 VPWR VGND sg13g2_decap_4
X_2624_ Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q net19 net76 net103 Inst_RegFile_switch_matrix.JN2BEG4
+ Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q _1042_ VPWR VGND sg13g2_mux4_1
X_3673_ NN4END[13] net261 VPWR VGND sg13g2_buf_1
X_3742_ Inst_RegFile_switch_matrix.JW2BEG5 net324 VPWR VGND sg13g2_buf_2
XFILLER_20_338 VPWR VGND sg13g2_fill_1
Xoutput179 net179 FrameData_O[29] VPWR VGND sg13g2_buf_1
X_2555_ Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q _1165_ _1000_ VPWR VGND sg13g2_nor2_1
Xoutput135 net135 E6BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_56_0 VPWR VGND sg13g2_decap_8
Xoutput146 Inst_RegFile_switch_matrix.EE4BEG1 EE4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput168 net168 FrameData_O[19] VPWR VGND sg13g2_buf_1
X_2486_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q _1182_ _0941_ _0940_
+ sg13g2_a21oi_1
Xoutput157 net157 EE4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput113 Inst_RegFile_switch_matrix.E1BEG3 E1BEG[3] VPWR VGND sg13g2_buf_1
Xoutput124 net124 E2BEGb[2] VPWR VGND sg13g2_buf_1
X_2850__480 VPWR VGND net480 sg13g2_tiehi
X_3107_ net1162 net1088 Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q VPWR VGND sg13g2_dlhq_1
X_3038_ net1175 net1077 Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q VPWR VGND sg13g2_dlhq_1
XFILLER_51_430 VPWR VGND sg13g2_decap_4
XFILLER_23_187 VPWR VGND sg13g2_decap_8
XFILLER_11_10 VPWR VGND sg13g2_fill_1
XFILLER_46_213 VPWR VGND sg13g2_fill_1
XFILLER_36_73 VPWR VGND sg13g2_fill_1
Xinput59 S1END[1] net59 VPWR VGND sg13g2_buf_2
X_2897__425 VPWR VGND net425 sg13g2_tiehi
Xinput26 FrameData[7] net26 VPWR VGND sg13g2_buf_1
Xinput15 E2MID[2] net15 VPWR VGND sg13g2_buf_1
Xinput48 N2MID[6] net48 VPWR VGND sg13g2_buf_1
Xinput37 N2END[3] net37 VPWR VGND sg13g2_buf_1
X_2340_ net1042 net1070 _0808_ VPWR VGND sg13g2_nor2b_1
X_2271_ Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q VPWR _0743_ VGND net1050 net985
+ sg13g2_o21ai_1
XFILLER_37_235 VPWR VGND sg13g2_fill_1
XFILLER_18_471 VPWR VGND sg13g2_fill_2
X_1986_ net69 net1071 net1052 _0477_ VPWR VGND sg13g2_mux2_1
X_3725_ SS4END[13] net313 VPWR VGND sg13g2_buf_1
X_3587_ net1209 net160 VPWR VGND sg13g2_buf_1
X_2607_ _1024_ VPWR _1025_ VGND _1021_ _1022_ sg13g2_o21ai_1
X_3656_ N4END[12] net244 VPWR VGND sg13g2_buf_1
X_2469_ _0924_ _0927_ _0928_ VPWR VGND sg13g2_nor2_1
X_2538_ _0983_ _0986_ _0987_ VPWR VGND sg13g2_nor2_1
XFILLER_0_518 VPWR VGND sg13g2_fill_2
Xfanout1113 net1114 net1113 VPWR VGND sg13g2_buf_1
Xfanout1102 net28 net1102 VPWR VGND sg13g2_buf_1
XFILLER_0_2 VPWR VGND sg13g2_fill_1
XFILLER_59_360 VPWR VGND sg13g2_decap_8
Xfanout1168 FrameData[29] net1168 VPWR VGND sg13g2_buf_1
Xfanout1124 net1125 net1124 VPWR VGND sg13g2_buf_1
Xfanout1179 FrameData[24] net1179 VPWR VGND sg13g2_buf_1
Xfanout1135 net1136 net1135 VPWR VGND sg13g2_buf_1
Xfanout1146 net1147 net1146 VPWR VGND sg13g2_buf_1
Xfanout1157 FrameData[5] net1157 VPWR VGND sg13g2_buf_1
XFILLER_19_235 VPWR VGND sg13g2_fill_1
XFILLER_19_257 VPWR VGND sg13g2_fill_1
X_1840_ _0236_ _0337_ _0321_ Inst_RegFile_32x4.AD_comb\[3\] VPWR VGND sg13g2_a21o_1
X_1771_ Inst_RegFile_32x4.mem\[26\]\[1\] Inst_RegFile_32x4.mem\[27\]\[1\] net931 _0273_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_99 VPWR VGND sg13g2_fill_2
X_3372_ UserCLK net372 _0108_ _3372_/Q_N Inst_RegFile_32x4.mem\[8\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_2323_ _0791_ VPWR _0792_ VGND net1041 net1029 sg13g2_o21ai_1
X_2254_ VGND VPWR _0726_ Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q _0725_ Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q
+ _0727_ _0724_ sg13g2_a221oi_1
X_2185_ net1002 net1044 _0662_ VPWR VGND sg13g2_nor2b_1
XFILLER_33_293 VPWR VGND sg13g2_decap_4
X_1969_ _0460_ _0434_ net518 VPWR VGND sg13g2_nand2_2
X_3639_ Inst_RegFile_switch_matrix.JN2BEG7 net221 VPWR VGND sg13g2_buf_1
X_3708_ S4END[12] net296 VPWR VGND sg13g2_buf_1
XFILLER_56_374 VPWR VGND sg13g2_decap_8
X_2887__435 VPWR VGND net435 sg13g2_tiehi
X_2894__428 VPWR VGND net428 sg13g2_tiehi
XFILLER_8_459 VPWR VGND sg13g2_fill_1
XFILLER_12_477 VPWR VGND sg13g2_fill_2
X_2941_ net1176 net1127 Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q VPWR VGND sg13g2_dlhq_1
X_2872_ UserCLK net458 _0030_ _2872_/Q_N Inst_RegFile_32x4.mem\[9\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_1823_ VGND VPWR _0320_ _0236_ _0318_ _0315_ _0321_ _0316_ sg13g2_a221oi_1
XFILLER_15_260 VPWR VGND sg13g2_fill_1
X_1685_ _0190_ VPWR _0191_ VGND net1026 _0187_ sg13g2_o21ai_1
X_1754_ VGND VPWR Inst_RegFile_32x4.mem\[21\]\[0\] net926 _0258_ _0257_ sg13g2_a21oi_1
X_2306_ _0776_ net1037 net1031 VPWR VGND sg13g2_nand2_1
Xfanout928 net931 net928 VPWR VGND sg13g2_buf_1
X_3286_ net1192 net1123 Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q VPWR VGND sg13g2_dlhq_1
X_3355_ UserCLK net389 _0091_ _3355_/Q_N Inst_RegFile_32x4.mem\[3\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_2237_ VGND VPWR net1040 net1018 _0711_ _0710_ sg13g2_a21oi_1
Xfanout939 _1065_ net939 VPWR VGND sg13g2_buf_1
XFILLER_53_388 VPWR VGND sg13g2_decap_8
X_2168_ A_ADR0 _0644_ _0646_ Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q _0642_ VPWR
+ VGND sg13g2_a22oi_1
X_2099_ Inst_RegFile_32x4.BD_comb\[2\] Inst_RegFile_32x4.BD_reg\[2\] Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q
+ BD2 VPWR VGND sg13g2_mux2_1
XFILLER_56_171 VPWR VGND sg13g2_fill_1
XFILLER_29_352 VPWR VGND sg13g2_fill_2
XFILLER_28_96 VPWR VGND sg13g2_fill_2
XFILLER_44_73 VPWR VGND sg13g2_fill_1
XFILLER_8_234 VPWR VGND sg13g2_fill_2
XFILLER_5_89 VPWR VGND sg13g2_fill_2
X_3140_ net1213 net28 Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q VPWR VGND sg13g2_dlhq_1
XFILLER_39_105 VPWR VGND sg13g2_fill_2
X_3071_ net1173 net1083 Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q VPWR VGND sg13g2_dlhq_1
XFILLER_50_325 VPWR VGND sg13g2_decap_8
X_2022_ Inst_RegFile_32x4.mem\[24\]\[1\] Inst_RegFile_32x4.mem\[25\]\[1\] net993 _0510_
+ VPWR VGND sg13g2_mux2_1
X_2855_ UserCLK net475 _0013_ _2855_/Q_N Inst_RegFile_32x4.mem\[27\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_2924_ net1151 net1129 Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q VPWR VGND sg13g2_dlhq_1
X_1806_ VGND VPWR Inst_RegFile_32x4.mem\[21\]\[2\] net924 _0306_ _0305_ sg13g2_a21oi_1
X_2786_ _1120_ _1092_ _1094_ VPWR VGND sg13g2_nand2_2
XFILLER_58_425 VPWR VGND sg13g2_fill_1
X_1668_ Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q _0169_ _0175_ VPWR VGND sg13g2_and2_1
X_1599_ Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q _1217_ _1218_ _1219_ VPWR VGND
+ sg13g2_nor3_1
Xhold256 Inst_RegFile_32x4.mem\[10\]\[1\] VPWR VGND net754 sg13g2_dlygate4sd3_1
Xhold245 Inst_RegFile_32x4.mem\[10\]\[3\] VPWR VGND net743 sg13g2_dlygate4sd3_1
Xhold234 Inst_RegFile_32x4.mem\[4\]\[1\] VPWR VGND net732 sg13g2_dlygate4sd3_1
X_3338_ UserCLK net488 Inst_RegFile_32x4.AD_comb\[2\] _3338_/Q_N Inst_RegFile_32x4.AD_reg\[2\]
+ VPWR VGND sg13g2_dfrbp_1
Xhold267 Inst_RegFile_32x4.mem\[1\]\[1\] VPWR VGND net765 sg13g2_dlygate4sd3_1
Xhold289 Inst_RegFile_32x4.mem\[30\]\[3\] VPWR VGND net787 sg13g2_dlygate4sd3_1
Xhold278 Inst_RegFile_32x4.mem\[28\]\[2\] VPWR VGND net776 sg13g2_dlygate4sd3_1
X_1737_ VGND VPWR _0240_ net982 _0239_ net1022 _0241_ _0238_ sg13g2_a221oi_1
XFILLER_53_130 VPWR VGND sg13g2_fill_2
XFILLER_26_333 VPWR VGND sg13g2_fill_2
X_3269_ net1188 net1121 Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q VPWR VGND sg13g2_dlhq_1
X_2884__438 VPWR VGND net438 sg13g2_tiehi
X_2640_ Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q _1057_ _1055_ _1052_ _1050_ Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q
+ _1058_ VPWR VGND sg13g2_mux4_1
X_2571_ Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q net1074 net1219 net88 net980 Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q
+ _1014_ VPWR VGND sg13g2_mux4_1
Xoutput317 Inst_RegFile_switch_matrix.W1BEG2 W1BEG[2] VPWR VGND sg13g2_buf_1
Xoutput328 net328 W2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput306 net306 SS4BEG[2] VPWR VGND sg13g2_buf_1
X_1522_ VPWR _1144_ Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q VGND sg13g2_inv_1
Xoutput339 net339 W6BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_55_439 VPWR VGND sg13g2_decap_4
X_3054_ net1210 net1086 Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q VPWR VGND sg13g2_dlhq_1
X_2005_ net997 Inst_RegFile_32x4.mem\[4\]\[0\] Inst_RegFile_32x4.mem\[5\]\[0\] Inst_RegFile_32x4.mem\[6\]\[0\]
+ Inst_RegFile_32x4.mem\[7\]\[0\] net947 _0495_ VPWR VGND sg13g2_mux4_1
XFILLER_27_119 VPWR VGND sg13g2_fill_2
X_3123_ net1198 net1093 Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q VPWR VGND sg13g2_dlhq_1
X_2907_ UserCLK net415 _0065_ _2907_/Q_N Inst_RegFile_32x4.mem\[1\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_2838_ net940 net825 _1131_ _0124_ VPWR VGND sg13g2_mux2_1
X_2769_ net958 net761 _1116_ _0070_ VPWR VGND sg13g2_mux2_1
XFILLER_26_152 VPWR VGND sg13g2_decap_8
XFILLER_18_108 VPWR VGND sg13g2_fill_1
XFILLER_45_494 VPWR VGND sg13g2_fill_2
X_3741_ net523 net323 VPWR VGND sg13g2_buf_1
X_2554_ VGND VPWR _1159_ _0339_ _0999_ _0998_ sg13g2_a21oi_1
X_2623_ VGND VPWR _1041_ _1040_ _1039_ sg13g2_or2_1
Xoutput114 net114 E2BEG[0] VPWR VGND sg13g2_buf_1
X_3672_ NN4END[12] net260 VPWR VGND sg13g2_buf_1
Xoutput125 net125 E2BEGb[3] VPWR VGND sg13g2_buf_1
Xoutput169 net169 FrameData_O[1] VPWR VGND sg13g2_buf_1
Xoutput147 net147 EE4BEG[14] VPWR VGND sg13g2_buf_1
X_2485_ Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q _1165_ _0940_ VPWR VGND sg13g2_nor2_1
Xoutput136 net136 E6BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_49_0 VPWR VGND sg13g2_decap_8
Xoutput158 net158 FrameData_O[0] VPWR VGND sg13g2_buf_1
XFILLER_55_236 VPWR VGND sg13g2_fill_2
X_3037_ net1176 net1082 Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q VPWR VGND sg13g2_dlhq_1
X_3106_ net1164 net1088 Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q VPWR VGND sg13g2_dlhq_1
XFILLER_3_505 VPWR VGND sg13g2_fill_2
XFILLER_11_77 VPWR VGND sg13g2_fill_1
XFILLER_36_52 VPWR VGND sg13g2_fill_2
XFILLER_34_409 VPWR VGND sg13g2_fill_1
Xinput16 E2MID[3] net16 VPWR VGND sg13g2_buf_1
Xinput49 N2MID[7] net49 VPWR VGND sg13g2_buf_1
Xinput38 N2END[4] net38 VPWR VGND sg13g2_buf_1
Xinput27 FrameStrobe[12] net27 VPWR VGND sg13g2_buf_1
XFILLER_42_7 VPWR VGND sg13g2_decap_4
X_2270_ _0741_ VPWR _0742_ VGND net1050 net1030 sg13g2_o21ai_1
XFILLER_18_494 VPWR VGND sg13g2_fill_1
X_3724_ SS4END[12] net312 VPWR VGND sg13g2_buf_1
X_1985_ net1052 net33 net41 net55 net4 Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q
+ _0476_ VPWR VGND sg13g2_mux4_1
X_3586_ net1210 net159 VPWR VGND sg13g2_buf_1
X_2537_ Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q VPWR _0986_ VGND Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q
+ _0985_ sg13g2_o21ai_1
X_2606_ VGND VPWR _1162_ _1023_ _1024_ Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q
+ sg13g2_a21oi_1
X_3655_ N4END[11] net243 VPWR VGND sg13g2_buf_1
XFILLER_57_18 VPWR VGND sg13g2_fill_1
X_2468_ Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q VPWR _0927_ VGND Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q
+ _0926_ sg13g2_o21ai_1
X_2399_ _0856_ VPWR Inst_RegFile_switch_matrix.E2BEG0 VGND Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q
+ _0863_ sg13g2_o21ai_1
XFILLER_51_250 VPWR VGND sg13g2_fill_2
XFILLER_43_217 VPWR VGND sg13g2_fill_2
XFILLER_36_280 VPWR VGND sg13g2_fill_1
XFILLER_11_125 VPWR VGND sg13g2_fill_1
Xfanout1125 net1126 net1125 VPWR VGND sg13g2_buf_1
Xfanout1136 FrameStrobe[11] net1136 VPWR VGND sg13g2_buf_1
Xfanout1114 FrameStrobe[3] net1114 VPWR VGND sg13g2_buf_1
Xfanout1103 net1108 net1103 VPWR VGND sg13g2_buf_1
Xfanout1147 FrameStrobe[0] net1147 VPWR VGND sg13g2_buf_1
Xfanout1169 FrameData[29] net1169 VPWR VGND sg13g2_buf_1
Xfanout1158 net1159 net1158 VPWR VGND sg13g2_buf_1
X_1770_ VGND VPWR Inst_RegFile_32x4.mem\[25\]\[1\] net928 _0272_ _0271_ sg13g2_a21oi_1
X_3371_ UserCLK net373 _0107_ _3371_/Q_N Inst_RegFile_32x4.mem\[7\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_2184_ _0654_ VPWR Inst_RegFile_switch_matrix.JW2BEG2 VGND Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q
+ _0661_ sg13g2_o21ai_1
X_2322_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q _0791_ net1010 net1041
+ sg13g2_a21oi_2
X_2253_ VGND VPWR net1045 net1016 _0726_ Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q
+ sg13g2_a21oi_1
X_3707_ S4END[11] net295 VPWR VGND sg13g2_buf_1
X_1899_ Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q _0391_ _0392_ _0393_ VPWR VGND
+ sg13g2_nor3_1
X_1968_ _0458_ _0434_ _0459_ VPWR VGND sg13g2_and2_2
X_3569_ EE4END[13] net157 VPWR VGND sg13g2_buf_1
XFILLER_39_309 VPWR VGND sg13g2_fill_1
XFILLER_47_386 VPWR VGND sg13g2_fill_1
XFILLER_47_342 VPWR VGND sg13g2_fill_1
X_2940_ net1178 net1127 Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q VPWR VGND sg13g2_dlhq_1
X_2871_ UserCLK net459 _0029_ _2871_/Q_N Inst_RegFile_32x4.mem\[9\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_3337__446 VPWR VGND net446 sg13g2_tiehi
XFILLER_7_460 VPWR VGND sg13g2_fill_2
X_1753_ net926 Inst_RegFile_32x4.mem\[20\]\[0\] _0257_ VPWR VGND sg13g2_nor2b_1
X_1822_ VGND VPWR net983 _0319_ _0320_ _0185_ sg13g2_a21oi_1
Xfanout929 net930 net929 VPWR VGND sg13g2_buf_1
X_1684_ VGND VPWR net1026 _0189_ _0190_ net956 sg13g2_a21oi_1
X_3354_ UserCLK net390 _0090_ _3354_/Q_N Inst_RegFile_32x4.mem\[3\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_2305_ VGND VPWR _0774_ Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q _0773_ Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q
+ _0775_ _0772_ sg13g2_a221oi_1
X_2167_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q _0645_ _0646_ Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q
+ sg13g2_a21oi_1
X_2236_ net1040 net1066 _0710_ VPWR VGND sg13g2_nor2b_1
X_3285_ net1194 net1122 Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q VPWR VGND sg13g2_dlhq_1
X_2098_ _0581_ net532 _0568_ Inst_RegFile_32x4.BD_comb\[2\] VPWR VGND sg13g2_a21o_1
XFILLER_0_90 VPWR VGND sg13g2_fill_1
XFILLER_44_356 VPWR VGND sg13g2_fill_1
XFILLER_54_109 VPWR VGND sg13g2_fill_1
XFILLER_35_323 VPWR VGND sg13g2_fill_2
X_3070_ net1174 net1083 Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q VPWR VGND sg13g2_dlhq_1
X_2021_ Inst_RegFile_32x4.BD_comb\[0\] Inst_RegFile_32x4.BD_reg\[0\] Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q
+ BD0 VPWR VGND sg13g2_mux2_2
XFILLER_35_356 VPWR VGND sg13g2_fill_2
XFILLER_23_529 VPWR VGND sg13g2_fill_2
X_2923_ net1152 net1129 Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q VPWR VGND sg13g2_dlhq_1
X_2854_ UserCLK net476 _0012_ _2854_/Q_N Inst_RegFile_32x4.mem\[27\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
Xhold235 Inst_RegFile_32x4.mem\[2\]\[3\] VPWR VGND net733 sg13g2_dlygate4sd3_1
X_2785_ net932 net809 _1119_ _0083_ VPWR VGND sg13g2_mux2_1
X_1736_ VGND VPWR Inst_RegFile_32x4.mem\[3\]\[0\] net921 _0240_ net1022 sg13g2_a21oi_1
X_1805_ net924 Inst_RegFile_32x4.mem\[20\]\[2\] _0305_ VPWR VGND sg13g2_nor2b_1
X_1667_ _0171_ Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q _0173_ _0174_ VPWR VGND
+ sg13g2_a21o_1
X_1598_ net1033 Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q _1218_ VPWR VGND sg13g2_nor2b_1
Xhold257 Inst_RegFile_32x4.mem\[26\]\[1\] VPWR VGND net755 sg13g2_dlygate4sd3_1
Xhold246 Inst_RegFile_32x4.mem\[26\]\[3\] VPWR VGND net744 sg13g2_dlygate4sd3_1
Xhold279 Inst_RegFile_32x4.mem\[5\]\[0\] VPWR VGND net777 sg13g2_dlygate4sd3_1
X_3337_ UserCLK net446 Inst_RegFile_32x4.AD_comb\[1\] _3337_/Q_N Inst_RegFile_32x4.AD_reg\[1\]
+ VPWR VGND sg13g2_dfrbp_1
Xhold268 Inst_RegFile_32x4.mem\[14\]\[2\] VPWR VGND net766 sg13g2_dlygate4sd3_1
X_2219_ Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q VPWR _0694_ VGND Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q
+ _0693_ sg13g2_o21ai_1
X_3199_ net1172 net1106 Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q VPWR VGND sg13g2_dlhq_1
XFILLER_41_315 VPWR VGND sg13g2_decap_8
X_3268_ net1212 net1121 Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q VPWR VGND sg13g2_dlhq_1
XFILLER_44_153 VPWR VGND sg13g2_fill_2
X_2570_ _1013_ _1012_ VPWR VGND sg13g2_inv_2
Xoutput307 net307 SS4BEG[3] VPWR VGND sg13g2_buf_1
X_1521_ VPWR _1143_ Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q VGND sg13g2_inv_1
Xoutput329 net329 W2BEGb[2] VPWR VGND sg13g2_buf_1
Xoutput318 Inst_RegFile_switch_matrix.W1BEG3 W1BEG[3] VPWR VGND sg13g2_buf_1
X_3122_ net1201 net1093 Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q VPWR VGND sg13g2_dlhq_1
XFILLER_55_429 VPWR VGND sg13g2_fill_2
X_3053_ net1148 net1084 Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q VPWR VGND sg13g2_dlhq_1
X_2004_ _0494_ _0493_ net1004 VPWR VGND sg13g2_nand2b_1
X_2906_ UserCLK net416 _0064_ _2906_/Q_N Inst_RegFile_32x4.mem\[1\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_1719_ net1047 net1073 net41 net1218 net12 Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q
+ _0224_ VPWR VGND sg13g2_mux4_1
X_2837_ _1131_ _1061_ _1103_ VPWR VGND sg13g2_nand2_2
X_2768_ net951 net763 _1116_ _0069_ VPWR VGND sg13g2_mux2_1
X_2699_ _1026_ _1029_ _1033_ _1097_ VPWR VGND sg13g2_nor3_1
XFILLER_58_212 VPWR VGND sg13g2_fill_1
X_2890__432 VPWR VGND net432 sg13g2_tiehi
Xrebuffer50 net549 net548 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_25_32 VPWR VGND sg13g2_fill_2
XFILLER_25_10 VPWR VGND sg13g2_fill_1
XFILLER_9_0 VPWR VGND sg13g2_fill_2
Xoutput159 net159 FrameData_O[10] VPWR VGND sg13g2_buf_1
Xoutput137 net137 E6BEG[5] VPWR VGND sg13g2_buf_1
Xoutput148 net148 EE4BEG[15] VPWR VGND sg13g2_buf_1
X_2553_ Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q VPWR _0998_ VGND _1159_ _0997_
+ sg13g2_o21ai_1
X_2622_ Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q VPWR _1040_ VGND Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q
+ _0981_ sg13g2_o21ai_1
Xoutput115 net115 E2BEG[1] VPWR VGND sg13g2_buf_1
X_3671_ NN4END[11] net259 VPWR VGND sg13g2_buf_1
Xoutput126 net126 E2BEGb[4] VPWR VGND sg13g2_buf_1
X_2484_ VGND VPWR _1154_ _0339_ _0939_ _0938_ sg13g2_a21oi_1
X_3105_ net1169 net1089 Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q VPWR VGND sg13g2_dlhq_1
X_3036_ net1179 net1082 Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q VPWR VGND sg13g2_dlhq_1
XFILLER_59_510 VPWR VGND sg13g2_fill_2
XFILLER_46_248 VPWR VGND sg13g2_fill_2
XFILLER_52_63 VPWR VGND sg13g2_fill_2
XFILLER_27_495 VPWR VGND sg13g2_fill_1
Xinput17 E2MID[4] net17 VPWR VGND sg13g2_buf_1
Xinput28 FrameStrobe[5] net28 VPWR VGND sg13g2_buf_1
Xinput39 N2END[5] net39 VPWR VGND sg13g2_buf_2
X_3723_ SS4END[11] net311 VPWR VGND sg13g2_buf_1
X_1984_ _0468_ Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q _0474_ _0475_ VPWR VGND
+ sg13g2_nand3_1
X_3654_ N4END[10] net242 VPWR VGND sg13g2_buf_1
XFILLER_20_159 VPWR VGND sg13g2_fill_2
X_3585_ net1148 net189 VPWR VGND sg13g2_buf_1
X_2467_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q _1182_ _0926_ _0925_ sg13g2_a21oi_1
X_2536_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q _1182_ _0985_ _0984_
+ sg13g2_a21oi_1
X_2605_ net34 net62 Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q _1023_ VPWR VGND sg13g2_mux2_1
X_2398_ _0861_ VPWR _0863_ VGND Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q _0862_ sg13g2_o21ai_1
X_3019_ net1153 net1079 Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q VPWR VGND sg13g2_dlhq_1
XFILLER_24_498 VPWR VGND sg13g2_fill_1
XFILLER_24_454 VPWR VGND sg13g2_fill_2
XFILLER_24_432 VPWR VGND sg13g2_fill_1
XFILLER_11_115 VPWR VGND sg13g2_fill_2
XFILLER_3_314 VPWR VGND sg13g2_fill_2
XFILLER_3_303 VPWR VGND sg13g2_fill_1
Xfanout1126 FrameStrobe[1] net1126 VPWR VGND sg13g2_buf_1
Xfanout1148 net1149 net1148 VPWR VGND sg13g2_buf_1
Xfanout1104 net1108 net1104 VPWR VGND sg13g2_buf_1
Xfanout1159 FrameData[4] net1159 VPWR VGND sg13g2_buf_1
Xfanout1115 net1120 net1115 VPWR VGND sg13g2_buf_1
Xfanout1137 net1141 net1137 VPWR VGND sg13g2_buf_1
XFILLER_15_487 VPWR VGND sg13g2_fill_1
X_3370_ UserCLK net374 _0106_ _3370_/Q_N Inst_RegFile_32x4.mem\[7\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_2321_ VGND VPWR _0789_ Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q _0788_ Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q
+ _0790_ _0787_ sg13g2_a221oi_1
X_2183_ _0660_ VPWR _0661_ VGND Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q _0655_
+ sg13g2_o21ai_1
X_2252_ VGND VPWR _0725_ net1045 net1066 sg13g2_or2_1
XFILLER_53_516 VPWR VGND sg13g2_fill_2
X_3706_ S4END[10] net294 VPWR VGND sg13g2_buf_1
X_1898_ net1018 net1043 _0392_ VPWR VGND sg13g2_nor2b_1
X_1967_ _1139_ VPWR _0458_ VGND _0457_ _0439_ sg13g2_o21ai_1
X_3568_ EE4END[12] net156 VPWR VGND sg13g2_buf_1
X_2519_ VGND VPWR _0968_ _0969_ _0970_ _0964_ sg13g2_a21oi_1
XFILLER_33_87 VPWR VGND sg13g2_fill_1
XFILLER_24_273 VPWR VGND sg13g2_fill_2
X_2870_ UserCLK net460 _0028_ _2870_/Q_N Inst_RegFile_32x4.mem\[9\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_1683_ _0188_ VPWR _0189_ VGND Inst_RegFile_32x4.mem\[12\]\[0\] net930 sg13g2_o21ai_1
X_1821_ net927 Inst_RegFile_32x4.mem\[6\]\[3\] Inst_RegFile_32x4.mem\[7\]\[3\] Inst_RegFile_32x4.mem\[4\]\[3\]
+ Inst_RegFile_32x4.mem\[5\]\[3\] net1026 _0319_ VPWR VGND sg13g2_mux4_1
X_1752_ Inst_RegFile_32x4.mem\[22\]\[0\] Inst_RegFile_32x4.mem\[23\]\[0\] net926 _0256_
+ VPWR VGND sg13g2_mux2_1
X_2304_ VGND VPWR net1037 net1016 _0774_ Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q
+ sg13g2_a21oi_1
X_3284_ net1197 net1123 Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q VPWR VGND sg13g2_dlhq_1
X_3353_ UserCLK net391 _0089_ _3353_/Q_N Inst_RegFile_32x4.mem\[3\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_2166_ Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q net49 net20 net77 net104 Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q
+ _0645_ VPWR VGND sg13g2_mux4_1
X_2097_ _0581_ _0578_ _0580_ _0576_ net943 VPWR VGND sg13g2_a22oi_1
X_2235_ net963 net970 Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q _0709_ VPWR VGND sg13g2_mux2_1
X_2999_ net1191 net1140 Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q VPWR VGND sg13g2_dlhq_1
XFILLER_29_354 VPWR VGND sg13g2_fill_1
XFILLER_28_43 VPWR VGND sg13g2_fill_1
XFILLER_44_324 VPWR VGND sg13g2_fill_2
XFILLER_44_20 VPWR VGND sg13g2_fill_1
XFILLER_28_98 VPWR VGND sg13g2_fill_1
XFILLER_39_107 VPWR VGND sg13g2_fill_1
X_2020_ _0497_ _0491_ _0509_ Inst_RegFile_32x4.BD_comb\[0\] VPWR VGND sg13g2_a21o_1
X_2853_ UserCLK net477 _0011_ _2853_/Q_N Inst_RegFile_32x4.mem\[26\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_31_530 VPWR VGND sg13g2_fill_1
X_2922_ net1154 net1129 Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q VPWR VGND sg13g2_dlhq_1
X_1666_ Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q VPWR _0173_ VGND Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q
+ _0172_ sg13g2_o21ai_1
Xhold269 Inst_RegFile_32x4.mem\[24\]\[1\] VPWR VGND net767 sg13g2_dlygate4sd3_1
Xhold258 Inst_RegFile_32x4.mem\[14\]\[0\] VPWR VGND net756 sg13g2_dlygate4sd3_1
Xhold247 Inst_RegFile_32x4.mem\[2\]\[2\] VPWR VGND net745 sg13g2_dlygate4sd3_1
X_2784_ net959 net808 _1119_ _0082_ VPWR VGND sg13g2_mux2_1
X_1804_ net925 Inst_RegFile_32x4.mem\[18\]\[2\] Inst_RegFile_32x4.mem\[19\]\[2\] Inst_RegFile_32x4.mem\[16\]\[2\]
+ Inst_RegFile_32x4.mem\[17\]\[2\] net1023 _0304_ VPWR VGND sg13g2_mux4_1
X_1735_ _0239_ Inst_RegFile_32x4.mem\[2\]\[0\] net921 VPWR VGND sg13g2_nand2b_1
Xhold236 Inst_RegFile_32x4.mem\[4\]\[2\] VPWR VGND net734 sg13g2_dlygate4sd3_1
XFILLER_58_438 VPWR VGND sg13g2_decap_8
XFILLER_58_405 VPWR VGND sg13g2_decap_8
X_3267_ net1163 net1118 Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q VPWR VGND sg13g2_dlhq_1
X_1597_ Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q net975 _1217_ VPWR VGND sg13g2_nor2_1
X_3336_ UserCLK net445 Inst_RegFile_32x4.AD_comb\[0\] _3336_/Q_N Inst_RegFile_32x4.AD_reg\[0\]
+ VPWR VGND sg13g2_dfrbp_1
XFILLER_53_132 VPWR VGND sg13g2_fill_1
X_2218_ VGND VPWR _0692_ _0693_ net1015 net1058 sg13g2_a21oi_2
X_3198_ net1175 net1106 Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q VPWR VGND sg13g2_dlhq_1
X_2149_ VGND VPWR net66 net1057 _0629_ _0628_ sg13g2_a21oi_1
XFILLER_57_471 VPWR VGND sg13g2_fill_2
XFILLER_39_53 VPWR VGND sg13g2_fill_2
XFILLER_44_176 VPWR VGND sg13g2_fill_2
XFILLER_13_530 VPWR VGND sg13g2_fill_1
X_1520_ VPWR _1142_ Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q VGND sg13g2_inv_1
Xoutput319 net319 W2BEG[0] VPWR VGND sg13g2_buf_1
Xoutput308 net308 SS4BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_4_261 VPWR VGND sg13g2_fill_2
X_3121_ net1204 net1096 Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q VPWR VGND sg13g2_dlhq_1
XFILLER_55_408 VPWR VGND sg13g2_decap_8
X_3052_ net1151 net1084 Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q VPWR VGND sg13g2_dlhq_1
X_2003_ net990 Inst_RegFile_32x4.mem\[0\]\[0\] Inst_RegFile_32x4.mem\[1\]\[0\] Inst_RegFile_32x4.mem\[2\]\[0\]
+ Inst_RegFile_32x4.mem\[3\]\[0\] net944 _0493_ VPWR VGND sg13g2_mux4_1
X_2836_ net935 net790 _1130_ _0123_ VPWR VGND sg13g2_mux2_1
X_2905_ UserCLK net417 _0063_ _2905_/Q_N Inst_RegFile_32x4.mem\[18\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_3378__366 VPWR VGND net366 sg13g2_tiehi
X_1718_ Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q VPWR _0223_ VGND _0219_ _0222_
+ sg13g2_o21ai_1
X_2767_ net939 net762 _1116_ _0068_ VPWR VGND sg13g2_mux2_1
X_1649_ Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q net1074 net38 net57 net9 Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q
+ _0157_ VPWR VGND sg13g2_mux4_1
X_2698_ _1026_ _1029_ _1096_ VPWR VGND sg13g2_nor2_1
X_3319_ net1190 net1146 Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q VPWR VGND sg13g2_dlhq_1
XFILLER_54_496 VPWR VGND sg13g2_fill_2
XFILLER_54_474 VPWR VGND sg13g2_decap_4
Xrebuffer51 net550 net549 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer40 net539 net538 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_41_87 VPWR VGND sg13g2_fill_2
XFILLER_49_202 VPWR VGND sg13g2_fill_2
XFILLER_49_279 VPWR VGND sg13g2_fill_2
XFILLER_45_496 VPWR VGND sg13g2_fill_1
XFILLER_45_430 VPWR VGND sg13g2_fill_2
XFILLER_32_113 VPWR VGND sg13g2_decap_4
XFILLER_17_176 VPWR VGND sg13g2_decap_8
X_3670_ NN4END[10] net258 VPWR VGND sg13g2_buf_1
XFILLER_9_320 VPWR VGND sg13g2_fill_1
XFILLER_20_308 VPWR VGND sg13g2_fill_2
Xoutput138 net138 E6BEG[6] VPWR VGND sg13g2_buf_1
X_2483_ Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q VPWR _0938_ VGND _1154_ _0209_
+ sg13g2_o21ai_1
X_2621_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q _1035_ _1039_ _1038_ sg13g2_a21oi_1
Xoutput127 net127 E2BEGb[5] VPWR VGND sg13g2_buf_1
X_2552_ Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q net36 net64 net7 net108 Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q
+ _0997_ VPWR VGND sg13g2_mux4_1
Xoutput116 net116 E2BEG[2] VPWR VGND sg13g2_buf_1
Xoutput149 net149 EE4BEG[1] VPWR VGND sg13g2_buf_1
X_3035_ net1180 net1080 Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q VPWR VGND sg13g2_dlhq_1
X_3104_ net1170 net1089 Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q VPWR VGND sg13g2_dlhq_1
XFILLER_51_400 VPWR VGND sg13g2_decap_4
X_2819_ net747 net952 _1127_ _0109_ VPWR VGND sg13g2_mux2_1
XFILLER_3_518 VPWR VGND sg13g2_fill_1
XFILLER_3_507 VPWR VGND sg13g2_fill_1
XFILLER_19_419 VPWR VGND sg13g2_fill_2
Xinput18 E2MID[5] net18 VPWR VGND sg13g2_buf_1
Xinput29 FrameStrobe[9] net29 VPWR VGND sg13g2_buf_1
XFILLER_6_356 VPWR VGND sg13g2_fill_2
XFILLER_10_363 VPWR VGND sg13g2_fill_1
XFILLER_10_374 VPWR VGND sg13g2_fill_1
XFILLER_37_216 VPWR VGND sg13g2_fill_2
X_3368__376 VPWR VGND net376 sg13g2_tiehi
XFILLER_33_433 VPWR VGND sg13g2_fill_2
XFILLER_18_441 VPWR VGND sg13g2_fill_1
X_3722_ SS4END[10] net310 VPWR VGND sg13g2_buf_1
X_3375__369 VPWR VGND net369 sg13g2_tiehi
X_1983_ _0473_ VPWR _0474_ VGND Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q _0470_
+ sg13g2_o21ai_1
X_2604_ Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q VPWR _1022_ VGND _1161_ _1231_
+ sg13g2_o21ai_1
X_3653_ N4END[9] net241 VPWR VGND sg13g2_buf_1
XFILLER_54_0 VPWR VGND sg13g2_decap_8
X_3584_ net1150 net188 VPWR VGND sg13g2_buf_1
X_2466_ Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q _1165_ _0925_ VPWR VGND sg13g2_nor2_1
X_2535_ Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q _1165_ _0984_ VPWR VGND sg13g2_nor2_1
X_3018_ net1155 net1079 Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q VPWR VGND sg13g2_dlhq_1
X_2397_ Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q net1073 net35 net51 net54 Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q
+ _0862_ VPWR VGND sg13g2_mux4_1
XFILLER_59_385 VPWR VGND sg13g2_decap_8
Xfanout1105 net1107 net1105 VPWR VGND sg13g2_buf_1
XFILLER_47_42 VPWR VGND sg13g2_decap_8
XFILLER_47_31 VPWR VGND sg13g2_fill_1
Xfanout1127 net1128 net1127 VPWR VGND sg13g2_buf_1
Xfanout1149 FrameData[9] net1149 VPWR VGND sg13g2_buf_1
Xfanout1116 net1120 net1116 VPWR VGND sg13g2_buf_1
XFILLER_19_205 VPWR VGND sg13g2_decap_8
XFILLER_19_216 VPWR VGND sg13g2_fill_2
Xfanout1138 net1141 net1138 VPWR VGND sg13g2_buf_1
XFILLER_42_296 VPWR VGND sg13g2_decap_4
XFILLER_42_274 VPWR VGND sg13g2_fill_1
X_2251_ net963 net970 Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q _0724_ VPWR VGND sg13g2_mux2_1
X_2320_ VGND VPWR net1041 net976 _0789_ Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q
+ sg13g2_a21oi_1
X_2182_ _0659_ VPWR _0660_ VGND Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q _0658_ sg13g2_o21ai_1
XFILLER_38_514 VPWR VGND sg13g2_fill_1
XFILLER_33_274 VPWR VGND sg13g2_fill_2
XFILLER_21_436 VPWR VGND sg13g2_fill_2
X_1966_ VGND VPWR _0456_ Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q _0455_ _0454_ _0457_
+ Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q sg13g2_a221oi_1
X_3705_ S4END[9] net293 VPWR VGND sg13g2_buf_1
X_3567_ EE4END[11] net155 VPWR VGND sg13g2_buf_1
X_3636_ Inst_RegFile_switch_matrix.JN2BEG4 net218 VPWR VGND sg13g2_buf_1
X_1897_ net1068 net1043 _0391_ VPWR VGND sg13g2_nor2_1
X_2518_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q _0966_ _0969_ _1156_
+ sg13g2_a21oi_1
X_2449_ Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q net45 net16 net73 net100 Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q
+ _0910_ VPWR VGND sg13g2_mux4_1
XFILLER_56_388 VPWR VGND sg13g2_decap_8
XFILLER_33_77 VPWR VGND sg13g2_decap_4
XFILLER_33_55 VPWR VGND sg13g2_fill_1
X_3358__386 VPWR VGND net386 sg13g2_tiehi
XFILLER_3_123 VPWR VGND sg13g2_fill_2
XFILLER_47_333 VPWR VGND sg13g2_fill_1
XFILLER_47_300 VPWR VGND sg13g2_decap_4
X_3365__379 VPWR VGND net379 sg13g2_tiehi
X_1820_ _0318_ _0143_ _0317_ VPWR VGND sg13g2_nand2_1
X_1682_ _0188_ net930 Inst_RegFile_32x4.mem\[13\]\[0\] VPWR VGND sg13g2_nand2b_1
XFILLER_30_299 VPWR VGND sg13g2_fill_2
XFILLER_30_277 VPWR VGND sg13g2_fill_1
X_1751_ VGND VPWR _0254_ net982 _0253_ net1023 _0255_ _0252_ sg13g2_a221oi_1
XFILLER_57_108 VPWR VGND sg13g2_fill_2
X_2303_ VGND VPWR _0773_ net1037 net106 sg13g2_or2_1
X_2234_ _0708_ VPWR Inst_RegFile_switch_matrix.JN2BEG2 VGND _0701_ _0695_ sg13g2_o21ai_1
X_3352_ UserCLK net392 _0088_ _3352_/Q_N Inst_RegFile_32x4.mem\[3\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_3283_ net1198 net1122 Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q VPWR VGND sg13g2_dlhq_1
X_2165_ _0644_ _0643_ Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q VPWR VGND sg13g2_nand2b_1
X_2096_ VGND VPWR net1007 _0579_ _0580_ net943 sg13g2_a21oi_1
X_2998_ net1193 net1141 Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q VPWR VGND sg13g2_dlhq_1
X_1949_ VGND VPWR _0441_ _0440_ Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q sg13g2_or2_1
X_3619_ net1134 net192 VPWR VGND sg13g2_buf_1
XFILLER_28_77 VPWR VGND sg13g2_fill_2
XFILLER_5_26 VPWR VGND sg13g2_fill_1
XFILLER_35_325 VPWR VGND sg13g2_fill_1
XFILLER_43_380 VPWR VGND sg13g2_fill_2
X_2852_ UserCLK net478 _0010_ _2852_/Q_N Inst_RegFile_32x4.mem\[26\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_2921_ net1157 net1129 Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q VPWR VGND sg13g2_dlhq_1
X_2783_ net950 net800 _1119_ _0081_ VPWR VGND sg13g2_mux2_1
X_1803_ VGND VPWR net956 _0300_ _0303_ net969 sg13g2_a21oi_1
X_1665_ net975 net1034 Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q _0172_ VPWR VGND
+ sg13g2_mux2_1
X_1596_ Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q _1215_ _1216_ VPWR VGND sg13g2_nor2_1
Xhold259 Inst_RegFile_32x4.mem\[26\]\[0\] VPWR VGND net757 sg13g2_dlygate4sd3_1
Xhold248 Inst_RegFile_32x4.mem\[6\]\[1\] VPWR VGND net746 sg13g2_dlygate4sd3_1
Xhold226 Inst_RegFile_32x4.mem\[6\]\[0\] VPWR VGND net724 sg13g2_dlygate4sd3_1
Xhold237 Inst_RegFile_32x4.mem\[0\]\[1\] VPWR VGND net735 sg13g2_dlygate4sd3_1
X_1734_ VGND VPWR Inst_RegFile_32x4.mem\[1\]\[0\] net921 _0238_ _0237_ sg13g2_a21oi_1
X_3266_ net1165 net1118 Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q VPWR VGND sg13g2_dlhq_1
X_2217_ net1058 net1033 _0692_ VPWR VGND sg13g2_nor2b_1
X_3197_ net1176 net1106 Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q VPWR VGND sg13g2_dlhq_1
X_3335_ UserCLK net444 Inst_RegFile_32x4.BD_comb\[3\] _3335_/Q_N Inst_RegFile_32x4.BD_reg\[3\]
+ VPWR VGND sg13g2_dfrbp_1
X_3348__396 VPWR VGND net396 sg13g2_tiehi
XFILLER_53_199 VPWR VGND sg13g2_fill_1
XFILLER_38_174 VPWR VGND sg13g2_fill_1
X_2079_ VGND VPWR _0459_ _0563_ _0562_ net1004 sg13g2_a21oi_2
X_2148_ net1056 net1216 _0628_ VPWR VGND sg13g2_nor2b_1
XFILLER_14_509 VPWR VGND sg13g2_fill_1
X_3355__389 VPWR VGND net389 sg13g2_tiehi
XFILLER_1_402 VPWR VGND sg13g2_fill_2
XFILLER_57_450 VPWR VGND sg13g2_decap_8
XFILLER_17_314 VPWR VGND sg13g2_fill_2
XFILLER_58_7 VPWR VGND sg13g2_decap_4
Xoutput309 net309 SS4BEG[5] VPWR VGND sg13g2_buf_1
X_3051_ net1153 net1084 Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q VPWR VGND sg13g2_dlhq_1
X_3120_ net1207 net1093 Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q VPWR VGND sg13g2_dlhq_1
X_2002_ _0483_ Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q _0490_ _0492_ VPWR VGND sg13g2_a21o_1
X_2835_ net961 net833 _1130_ _0122_ VPWR VGND sg13g2_mux2_1
X_2904_ UserCLK net418 _0062_ _2904_/Q_N Inst_RegFile_32x4.mem\[18\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_2766_ _1116_ _1061_ _1108_ VPWR VGND sg13g2_nand2_2
X_1717_ Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q VPWR _0222_ VGND _0220_ _0221_
+ sg13g2_o21ai_1
X_3318_ net1192 net1146 Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q VPWR VGND sg13g2_dlhq_1
X_1579_ _1200_ Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q _1198_ VPWR VGND sg13g2_nand2_1
XFILLER_6_91 VPWR VGND sg13g2_fill_1
X_2697_ net933 net789 _1095_ _0019_ VPWR VGND sg13g2_mux2_1
X_1648_ Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q VPWR _0156_ VGND _0155_ _0152_
+ sg13g2_o21ai_1
XFILLER_54_453 VPWR VGND sg13g2_decap_8
XFILLER_54_420 VPWR VGND sg13g2_decap_8
Xrebuffer52 net551 net550 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer41 net540 net539 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer30 net530 net528 VPWR VGND sg13g2_dlygate4sd1_1
X_3249_ net1203 net1116 Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q VPWR VGND sg13g2_dlhq_1
XFILLER_25_78 VPWR VGND sg13g2_decap_4
XFILLER_25_34 VPWR VGND sg13g2_fill_1
XFILLER_9_2 VPWR VGND sg13g2_fill_1
X_2620_ Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q VPWR _1038_ VGND Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q
+ _1037_ sg13g2_o21ai_1
XFILLER_9_398 VPWR VGND sg13g2_fill_2
Xoutput139 net139 E6BEG[7] VPWR VGND sg13g2_buf_1
X_2482_ _0937_ _0936_ Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q Inst_RegFile_switch_matrix.SS4BEG3
+ VPWR VGND sg13g2_mux2_1
X_2551_ _0996_ _0995_ Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q Inst_RegFile_switch_matrix.NN4BEG3
+ VPWR VGND sg13g2_mux2_1
Xoutput128 net128 E2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput117 net117 E2BEG[3] VPWR VGND sg13g2_buf_1
X_3034_ net1182 net1080 Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q VPWR VGND sg13g2_dlhq_1
X_3103_ net1173 net1091 Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q VPWR VGND sg13g2_dlhq_1
XFILLER_51_423 VPWR VGND sg13g2_decap_8
X_3345__399 VPWR VGND net399 sg13g2_tiehi
X_2818_ net731 net941 _1127_ _0108_ VPWR VGND sg13g2_mux2_1
X_2749_ net752 net960 _1112_ _0054_ VPWR VGND sg13g2_mux2_1
XFILLER_59_512 VPWR VGND sg13g2_fill_1
XFILLER_46_206 VPWR VGND sg13g2_decap_8
XFILLER_14_125 VPWR VGND sg13g2_fill_1
XFILLER_52_65 VPWR VGND sg13g2_fill_1
XFILLER_42_489 VPWR VGND sg13g2_fill_2
Xinput19 E2MID[6] net19 VPWR VGND sg13g2_buf_1
XFILLER_14_147 VPWR VGND sg13g2_fill_2
X_1982_ VGND VPWR _1132_ _0473_ Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q _0472_
+ sg13g2_a21oi_2
XFILLER_45_261 VPWR VGND sg13g2_fill_1
X_3721_ SS4END[9] net309 VPWR VGND sg13g2_buf_1
X_3583_ net26 net187 VPWR VGND sg13g2_buf_1
X_2534_ VGND VPWR _1158_ _0339_ _0983_ _0982_ sg13g2_a21oi_1
X_2603_ Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q _1180_ _1021_ VPWR VGND sg13g2_nor2_1
X_3652_ N4END[8] net240 VPWR VGND sg13g2_buf_1
X_2465_ VGND VPWR _1153_ _0339_ _0924_ _0923_ sg13g2_a21oi_1
XFILLER_3_81 VPWR VGND sg13g2_fill_1
X_2396_ _0859_ Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q _0860_ _0861_ VPWR VGND sg13g2_a21o_1
X_3017_ net1156 net1077 Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q VPWR VGND sg13g2_dlhq_1
XFILLER_11_117 VPWR VGND sg13g2_fill_1
XFILLER_3_316 VPWR VGND sg13g2_fill_1
XFILLER_59_353 VPWR VGND sg13g2_fill_2
Xfanout1106 net1107 net1106 VPWR VGND sg13g2_buf_1
Xfanout1117 net1119 net1117 VPWR VGND sg13g2_buf_1
Xfanout1139 net1140 net1139 VPWR VGND sg13g2_buf_1
Xfanout1128 net1130 net1128 VPWR VGND sg13g2_buf_1
XFILLER_27_294 VPWR VGND sg13g2_fill_2
X_3374__370 VPWR VGND net370 sg13g2_tiehi
XFILLER_40_7 VPWR VGND sg13g2_fill_1
X_2250_ _0719_ VPWR Inst_RegFile_switch_matrix.JW2BEG1 VGND Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q
+ _0723_ sg13g2_o21ai_1
XFILLER_53_518 VPWR VGND sg13g2_fill_1
X_3381__363 VPWR VGND net363 sg13g2_tiehi
X_2181_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q _0656_ _0659_ _1147_ sg13g2_a21oi_1
X_3704_ S4END[8] net292 VPWR VGND sg13g2_buf_1
XFILLER_21_448 VPWR VGND sg13g2_fill_1
X_1965_ VGND VPWR net42 _1137_ _0456_ Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q sg13g2_a21oi_1
X_3566_ EE4END[10] net154 VPWR VGND sg13g2_buf_1
X_2517_ _0967_ VPWR _0968_ VGND net1063 _1166_ sg13g2_o21ai_1
X_1896_ _0389_ VPWR _0390_ VGND Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q net976
+ sg13g2_o21ai_1
X_3635_ net717 net217 VPWR VGND sg13g2_buf_1
X_2379_ Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q net21 net60 net58 net62 Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q
+ _0845_ VPWR VGND sg13g2_mux4_1
X_2448_ VGND VPWR _0907_ _0908_ _0909_ _0903_ sg13g2_a21oi_1
XFILLER_24_275 VPWR VGND sg13g2_fill_1
XFILLER_12_448 VPWR VGND sg13g2_fill_2
XFILLER_30_234 VPWR VGND sg13g2_fill_1
X_1750_ VGND VPWR Inst_RegFile_32x4.mem\[19\]\[0\] net925 _0254_ net1023 sg13g2_a21oi_1
X_1681_ Inst_RegFile_32x4.mem\[14\]\[0\] Inst_RegFile_32x4.mem\[15\]\[0\] net930 _0187_
+ VPWR VGND sg13g2_mux2_1
X_3351_ UserCLK net393 _0087_ _3351_/Q_N Inst_RegFile_32x4.mem\[31\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_2302_ _0771_ VPWR _0772_ VGND net1037 net977 sg13g2_o21ai_1
X_2233_ _0707_ VPWR _0708_ VGND Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q _0702_
+ sg13g2_o21ai_1
X_2164_ Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q net48 net19 net103 Inst_RegFile_switch_matrix.JN2BEG5
+ Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q _0643_ VPWR VGND sg13g2_mux4_1
X_3282_ net1201 net1122 Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q VPWR VGND sg13g2_dlhq_1
X_2095_ net991 Inst_RegFile_32x4.mem\[4\]\[2\] Inst_RegFile_32x4.mem\[5\]\[2\] Inst_RegFile_32x4.mem\[6\]\[2\]
+ Inst_RegFile_32x4.mem\[7\]\[2\] net945 _0579_ VPWR VGND sg13g2_mux4_1
X_1879_ Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q net972 _0374_ VPWR VGND sg13g2_nor2_1
X_1948_ net973 net1033 Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q _0440_ VPWR VGND
+ sg13g2_mux2_1
X_2997_ net1194 net1137 Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q VPWR VGND sg13g2_dlhq_1
X_3618_ net1140 net191 VPWR VGND sg13g2_buf_1
X_3549_ E6END[3] net133 VPWR VGND sg13g2_buf_1
XFILLER_44_326 VPWR VGND sg13g2_fill_1
XFILLER_29_334 VPWR VGND sg13g2_fill_2
X_3364__380 VPWR VGND net380 sg13g2_tiehi
X_3371__373 VPWR VGND net373 sg13g2_tiehi
XFILLER_50_318 VPWR VGND sg13g2_decap_8
X_2920_ net1159 net1129 Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q VPWR VGND sg13g2_dlhq_1
X_2851_ UserCLK net479 _0009_ _2851_/Q_N Inst_RegFile_32x4.mem\[26\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_1733_ net922 Inst_RegFile_32x4.mem\[0\]\[0\] _0237_ VPWR VGND sg13g2_nor2b_1
X_2782_ net937 net772 _1119_ _0080_ VPWR VGND sg13g2_mux2_1
X_1802_ _0302_ net982 _0301_ VPWR VGND sg13g2_nand2_2
X_1664_ _0170_ VPWR _0171_ VGND Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q net989
+ sg13g2_o21ai_1
X_1595_ Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q net1070 net1019 net980 net967 Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q
+ _1215_ VPWR VGND sg13g2_mux4_1
Xhold249 Inst_RegFile_32x4.mem\[8\]\[1\] VPWR VGND net747 sg13g2_dlygate4sd3_1
Xhold227 Inst_RegFile_32x4.mem\[10\]\[2\] VPWR VGND net725 sg13g2_dlygate4sd3_1
Xhold238 Inst_RegFile_32x4.mem\[15\]\[3\] VPWR VGND net736 sg13g2_dlygate4sd3_1
X_3334_ UserCLK net443 Inst_RegFile_32x4.BD_comb\[2\] _3334_/Q_N Inst_RegFile_32x4.BD_reg\[2\]
+ VPWR VGND sg13g2_dfrbp_1
XFILLER_58_418 VPWR VGND sg13g2_decap_8
X_3265_ net1168 net1118 Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q VPWR VGND sg13g2_dlhq_1
X_2216_ net988 BD3 Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q _0691_ VPWR VGND sg13g2_mux2_1
X_3196_ net1178 net1106 Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q VPWR VGND sg13g2_dlhq_1
X_2147_ _0627_ Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q _0621_ VPWR VGND sg13g2_nand2_1
X_2078_ net990 Inst_RegFile_32x4.mem\[28\]\[2\] Inst_RegFile_32x4.mem\[29\]\[2\] Inst_RegFile_32x4.mem\[30\]\[2\]
+ Inst_RegFile_32x4.mem\[31\]\[2\] net944 _0562_ VPWR VGND sg13g2_mux4_1
XFILLER_55_32 VPWR VGND sg13g2_fill_2
XFILLER_55_21 VPWR VGND sg13g2_decap_8
XFILLER_29_175 VPWR VGND sg13g2_fill_2
X_2001_ VGND VPWR _0490_ _0491_ Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q _0483_ sg13g2_a21oi_2
X_3050_ net1154 net1085 Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q VPWR VGND sg13g2_dlhq_1
X_2903_ UserCLK net419 _0061_ _2903_/Q_N Inst_RegFile_32x4.mem\[18\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_2834_ net953 net796 _1130_ _0121_ VPWR VGND sg13g2_mux2_1
X_1716_ Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q VPWR _0221_ VGND net1047 net1015
+ sg13g2_o21ai_1
X_2765_ net932 net773 _1115_ _0067_ VPWR VGND sg13g2_mux2_1
X_3354__390 VPWR VGND net390 sg13g2_tiehi
X_2696_ net959 net776 _1095_ _0018_ VPWR VGND sg13g2_mux2_1
X_3317_ net1195 net1144 Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q VPWR VGND sg13g2_dlhq_1
X_1578_ _1199_ _1197_ Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q VPWR VGND sg13g2_nand2b_1
X_1647_ Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q VPWR _0155_ VGND _0153_ _0154_
+ sg13g2_o21ai_1
XFILLER_54_498 VPWR VGND sg13g2_fill_1
Xrebuffer53 Inst_RegFile_switch_matrix.JS2BEG6 net551 VPWR VGND sg13g2_buf_2
X_3361__383 VPWR VGND net383 sg13g2_tiehi
X_3179_ net1153 net1103 Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q VPWR VGND sg13g2_dlhq_1
XFILLER_26_145 VPWR VGND sg13g2_decap_8
Xrebuffer42 net541 net540 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer20 _0458_ net518 VPWR VGND sg13g2_buf_2
Xrebuffer31 net531 net529 VPWR VGND sg13g2_buf_2
X_3248_ net1206 net1116 Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q VPWR VGND sg13g2_dlhq_1
XFILLER_22_351 VPWR VGND sg13g2_fill_1
XFILLER_10_502 VPWR VGND sg13g2_fill_2
XFILLER_41_89 VPWR VGND sg13g2_fill_1
X_2550_ Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q net1075 net1220 net1071 net1019
+ Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q _0996_ VPWR VGND sg13g2_mux4_1
Xoutput129 net129 E2BEGb[7] VPWR VGND sg13g2_buf_1
X_2481_ Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q net31 net2 net1071 net1020 Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q
+ _0937_ VPWR VGND sg13g2_mux4_1
Xoutput118 net118 E2BEG[4] VPWR VGND sg13g2_buf_1
X_3033_ net1185 net29 Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q VPWR VGND sg13g2_dlhq_1
X_3102_ net1174 net1091 Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q VPWR VGND sg13g2_dlhq_1
XFILLER_51_446 VPWR VGND sg13g2_fill_2
X_2679_ net935 net830 _1089_ _0007_ VPWR VGND sg13g2_mux2_1
X_2817_ _1061_ _1101_ _1127_ VPWR VGND sg13g2_and2_2
XFILLER_11_59 VPWR VGND sg13g2_fill_1
X_2748_ net750 net951 _1112_ _0053_ VPWR VGND sg13g2_mux2_1
XFILLER_54_284 VPWR VGND sg13g2_fill_2
XFILLER_54_240 VPWR VGND sg13g2_fill_2
XFILLER_36_45 VPWR VGND sg13g2_decap_8
XFILLER_6_358 VPWR VGND sg13g2_fill_1
X_3720_ SS4END[8] net308 VPWR VGND sg13g2_buf_1
X_1981_ _0471_ VPWR _0472_ VGND net1052 net1011 sg13g2_o21ai_1
X_2533_ Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q VPWR _0982_ VGND _1158_ _0981_
+ sg13g2_o21ai_1
X_3582_ net25 net186 VPWR VGND sg13g2_buf_1
X_2602_ _1020_ Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q _1019_ VPWR VGND sg13g2_nand2b_1
X_3651_ N4END[7] net239 VPWR VGND sg13g2_buf_1
X_2464_ Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q VPWR _0923_ VGND _1153_ _0922_ sg13g2_o21ai_1
X_3351__393 VPWR VGND net393 sg13g2_tiehi
X_2395_ Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q VPWR _0860_ VGND Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q
+ _0858_ sg13g2_o21ai_1
X_3016_ net1158 net1077 Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q VPWR VGND sg13g2_dlhq_1
XFILLER_11_129 VPWR VGND sg13g2_fill_2
Xfanout1118 net1119 net1118 VPWR VGND sg13g2_buf_1
Xfanout1107 net1108 net1107 VPWR VGND sg13g2_buf_1
Xfanout1129 net1130 net1129 VPWR VGND sg13g2_buf_1
XFILLER_47_22 VPWR VGND sg13g2_decap_8
X_2180_ VGND VPWR net65 Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q _0658_ _0657_ sg13g2_a21oi_1
X_3703_ S4END[7] net291 VPWR VGND sg13g2_buf_1
X_1895_ _0389_ net1043 net966 VPWR VGND sg13g2_nand2_1
X_3634_ Inst_RegFile_switch_matrix.JN2BEG2 net216 VPWR VGND sg13g2_buf_8
X_1964_ _0455_ net13 Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q VPWR VGND sg13g2_nand2_1
X_3565_ EE4END[9] net153 VPWR VGND sg13g2_buf_1
X_2516_ VGND VPWR net1063 net978 _0967_ Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q
+ sg13g2_a21oi_1
X_2447_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q _0905_ _0908_ _1151_
+ sg13g2_a21oi_1
XFILLER_56_346 VPWR VGND sg13g2_fill_1
X_2378_ Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q net30 net1221 net34 net5 Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q
+ _0844_ VPWR VGND sg13g2_mux4_1
XFILLER_3_125 VPWR VGND sg13g2_fill_1
Xoutput290 net290 S4BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_15_210 VPWR VGND sg13g2_fill_1
X_2301_ _0771_ net1037 net719 VPWR VGND sg13g2_nand2_1
X_3350_ UserCLK net394 _0086_ _3350_/Q_N Inst_RegFile_32x4.mem\[31\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_1680_ _0186_ _0184_ _0167_ VPWR VGND sg13g2_nand2_2
X_2232_ VGND VPWR _0705_ _0706_ _0707_ Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q
+ sg13g2_a21oi_1
X_2163_ _0640_ VPWR _0642_ VGND Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q _0641_
+ sg13g2_o21ai_1
X_3281_ net1203 net1122 Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q VPWR VGND sg13g2_dlhq_1
XFILLER_34_530 VPWR VGND sg13g2_fill_1
X_2094_ _0578_ _0577_ net1004 VPWR VGND sg13g2_nand2b_1
X_1878_ Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q _0372_ _0373_ VPWR VGND sg13g2_nor2_2
X_3617_ net1082 net209 VPWR VGND sg13g2_buf_1
X_1947_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q _0436_ _0439_ _0438_
+ sg13g2_a21oi_1
X_2996_ net1196 net1137 Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q VPWR VGND sg13g2_dlhq_1
X_3548_ E6END[2] net130 VPWR VGND sg13g2_buf_1
XFILLER_56_198 VPWR VGND sg13g2_fill_2
XFILLER_47_176 VPWR VGND sg13g2_fill_2
X_2850_ UserCLK net480 _0008_ _2850_/Q_N Inst_RegFile_32x4.mem\[26\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_35_316 VPWR VGND sg13g2_decap_8
XFILLER_31_511 VPWR VGND sg13g2_fill_2
XFILLER_16_530 VPWR VGND sg13g2_fill_1
X_1663_ _0170_ Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q net1003 VPWR VGND sg13g2_nand2b_1
X_1732_ _0236_ _0234_ _0211_ VPWR VGND sg13g2_nand2_2
X_1801_ net921 Inst_RegFile_32x4.mem\[30\]\[2\] Inst_RegFile_32x4.mem\[31\]\[2\] Inst_RegFile_32x4.mem\[28\]\[2\]
+ Inst_RegFile_32x4.mem\[29\]\[2\] net1022 _0301_ VPWR VGND sg13g2_mux4_1
X_2781_ _1119_ _1088_ _1094_ VPWR VGND sg13g2_nand2_2
X_3264_ net1171 net1118 Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q VPWR VGND sg13g2_dlhq_1
X_1594_ VGND VPWR Inst_RegFile_32x4.mem\[11\]\[0\] net928 _1214_ net1027 sg13g2_a21oi_1
Xhold228 Inst_RegFile_32x4.mem\[4\]\[0\] VPWR VGND net726 sg13g2_dlygate4sd3_1
X_3333_ UserCLK net442 Inst_RegFile_32x4.BD_comb\[1\] _3333_/Q_N Inst_RegFile_32x4.BD_reg\[1\]
+ VPWR VGND sg13g2_dfrbp_1
Xhold239 Inst_RegFile_32x4.mem\[6\]\[3\] VPWR VGND net737 sg13g2_dlygate4sd3_1
X_3195_ net1181 net1107 Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q VPWR VGND sg13g2_dlhq_1
X_2215_ _0686_ VPWR Inst_RegFile_switch_matrix.E2BEG2 VGND Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q
+ _0690_ sg13g2_o21ai_1
XFILLER_38_110 VPWR VGND sg13g2_fill_1
X_2077_ _0560_ VPWR _0561_ VGND net1036 _0559_ sg13g2_o21ai_1
X_2146_ VGND VPWR _0625_ _0626_ _0624_ Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q
+ sg13g2_a21oi_2
X_2979_ net1162 net1131 Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q VPWR VGND sg13g2_dlhq_1
XFILLER_1_404 VPWR VGND sg13g2_fill_1
XFILLER_49_419 VPWR VGND sg13g2_fill_1
XFILLER_39_23 VPWR VGND sg13g2_fill_2
XFILLER_55_55 VPWR VGND sg13g2_fill_2
XFILLER_17_316 VPWR VGND sg13g2_fill_1
XFILLER_40_341 VPWR VGND sg13g2_fill_1
XFILLER_35_135 VPWR VGND sg13g2_fill_2
X_2000_ VGND VPWR _1140_ Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q _0489_ _0485_ _0490_
+ _0487_ sg13g2_a221oi_1
X_2833_ net941 net804 _1130_ _0120_ VPWR VGND sg13g2_mux2_1
X_2902_ UserCLK net420 _0060_ _2902_/Q_N Inst_RegFile_32x4.mem\[18\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
X_1715_ net1002 net1047 _0220_ VPWR VGND sg13g2_nor2b_1
X_2764_ net959 net784 _1115_ _0066_ VPWR VGND sg13g2_mux2_1
X_1646_ Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q VPWR _0154_ VGND net1039 net985
+ sg13g2_o21ai_1
X_2695_ net950 net769 _1095_ _0017_ VPWR VGND sg13g2_mux2_1
X_3247_ net1208 net1119 Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q VPWR VGND sg13g2_dlhq_1
X_3316_ net1197 net1144 Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q VPWR VGND sg13g2_dlhq_1
X_1577_ Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q net1217 net66 net85 net93 Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q
+ _1198_ VPWR VGND sg13g2_mux4_1
X_2129_ _0610_ Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q net20 VPWR VGND sg13g2_nand2b_1
Xrebuffer65 Inst_RegFile_switch_matrix.JS2BEG6 net563 VPWR VGND sg13g2_buf_2
X_3178_ net1155 net1103 Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q VPWR VGND sg13g2_dlhq_1
Xrebuffer43 net542 net541 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer21 _0491_ net519 VPWR VGND sg13g2_buf_2
Xrebuffer10 net526 net508 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer32 Inst_RegFile_switch_matrix.JW2BEG3 net530 VPWR VGND sg13g2_buf_2
XFILLER_41_79 VPWR VGND sg13g2_fill_2
X_3333__442 VPWR VGND net442 sg13g2_tiehi
XFILLER_45_411 VPWR VGND sg13g2_fill_1
XFILLER_17_135 VPWR VGND sg13g2_fill_2
X_2480_ Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q net1034 net499 net500 _0935_ Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q
+ _0936_ VPWR VGND sg13g2_mux4_1
XFILLER_31_90 VPWR VGND sg13g2_fill_1
Xoutput119 net119 E2BEG[5] VPWR VGND sg13g2_buf_8
X_3101_ net1177 net1090 Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q VPWR VGND sg13g2_dlhq_1
X_3032_ net1187 net1082 Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q VPWR VGND sg13g2_dlhq_1
XFILLER_36_477 VPWR VGND sg13g2_fill_2
XFILLER_31_193 VPWR VGND sg13g2_fill_2
X_2816_ net934 net786 _1126_ _0107_ VPWR VGND sg13g2_mux2_1
X_2678_ net961 net782 _1089_ _0006_ VPWR VGND sg13g2_mux2_1
X_2747_ net760 net940 _1112_ _0052_ VPWR VGND sg13g2_mux2_1
X_1629_ Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q net51 net93 net83 Inst_RegFile_switch_matrix.JS2BEG3
+ Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q _0137_ VPWR VGND sg13g2_mux4_1
X_1980_ _0471_ net1053 net1002 VPWR VGND sg13g2_nand2_1
X_3650_ N4END[6] net238 VPWR VGND sg13g2_buf_1
XFILLER_9_164 VPWR VGND sg13g2_fill_2
X_2532_ Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q net57 net11 net68 net95 Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q
+ _0981_ VPWR VGND sg13g2_mux4_1
X_2601_ _1161_ Inst_RegFile_switch_matrix.JW2BEG7 Inst_RegFile_switch_matrix.JS2BEG7
+ net721 _0935_ _1162_ _1019_ VPWR VGND sg13g2_mux4_1
X_2463_ Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q net38 net9 net84 net93 Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q
+ _0922_ VPWR VGND sg13g2_mux4_1
Xrebuffer1 _1229_ net499 VPWR VGND sg13g2_dlygate4sd1_1
X_3581_ net1157 net185 VPWR VGND sg13g2_buf_1
XFILLER_56_506 VPWR VGND sg13g2_fill_1
XFILLER_3_72 VPWR VGND sg13g2_decap_8
X_2394_ net63 net90 Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q _0859_ VPWR VGND sg13g2_mux2_1
X_3015_ net1160 net1077 Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q VPWR VGND sg13g2_dlhq_1
XFILLER_11_108 VPWR VGND sg13g2_decap_8
X_3779_ Inst_RegFile_switch_matrix.WW4BEG2 net352 VPWR VGND sg13g2_buf_1
XFILLER_59_355 VPWR VGND sg13g2_fill_1
Xfanout1119 net1120 net1119 VPWR VGND sg13g2_buf_1
Xfanout1108 FrameStrobe[4] net1108 VPWR VGND sg13g2_buf_1
XFILLER_59_399 VPWR VGND sg13g2_decap_8
XFILLER_47_89 VPWR VGND sg13g2_decap_4
XFILLER_10_130 VPWR VGND sg13g2_fill_1
XFILLER_10_152 VPWR VGND sg13g2_fill_1
XFILLER_6_112 VPWR VGND sg13g2_fill_1
XFILLER_53_509 VPWR VGND sg13g2_fill_2
X_3702_ S4END[6] net290 VPWR VGND sg13g2_buf_1
X_1894_ Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q net17 net74 net101 net563 Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q
+ _0388_ VPWR VGND sg13g2_mux4_1
X_1963_ _0453_ VPWR _0454_ VGND Inst_RegFile_switch_matrix.JW2BEG6 _1137_ sg13g2_o21ai_1
XFILLER_14_480 VPWR VGND sg13g2_fill_2
X_3633_ Inst_RegFile_switch_matrix.JN2BEG1 net215 VPWR VGND sg13g2_buf_2
X_3564_ EE4END[8] net152 VPWR VGND sg13g2_buf_1
XFILLER_52_0 VPWR VGND sg13g2_decap_8
X_2515_ VGND VPWR net1064 net972 _0966_ _0965_ sg13g2_a21oi_1
X_2446_ _0906_ VPWR _0907_ VGND net1061 net1016 sg13g2_o21ai_1
X_2377_ Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q VPWR _0843_ VGND Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q
+ _0836_ sg13g2_o21ai_1
XFILLER_52_520 VPWR VGND sg13g2_fill_2
XFILLER_12_439 VPWR VGND sg13g2_fill_2
XFILLER_3_104 VPWR VGND sg13g2_fill_2
Xoutput291 net291 S4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput280 net280 S2BEGb[6] VPWR VGND sg13g2_buf_1
XFILLER_11_450 VPWR VGND sg13g2_fill_1
X_2231_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q _0703_ _0706_ _1148_ sg13g2_a21oi_1
X_2300_ _0770_ VPWR Inst_RegFile_switch_matrix.JN2BEG1 VGND _0765_ _0759_ sg13g2_o21ai_1
X_3280_ net1206 net1122 Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q VPWR VGND sg13g2_dlhq_1
X_2162_ Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q net41 net69 net23 net96 Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q
+ _0641_ VPWR VGND sg13g2_mux4_1
X_2093_ net990 Inst_RegFile_32x4.mem\[0\]\[2\] Inst_RegFile_32x4.mem\[1\]\[2\] Inst_RegFile_32x4.mem\[2\]\[2\]
+ Inst_RegFile_32x4.mem\[3\]\[2\] net944 _0577_ VPWR VGND sg13g2_mux4_1
XFILLER_46_391 VPWR VGND sg13g2_fill_1
X_2995_ net1198 net1137 Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q VPWR VGND sg13g2_dlhq_1
X_1877_ Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q net1068 net1017 net978 net965 Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q
+ _0372_ VPWR VGND sg13g2_mux4_1
X_3547_ net20 net129 VPWR VGND sg13g2_buf_1
X_3616_ net1087 net208 VPWR VGND sg13g2_buf_1
X_1946_ Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q VPWR _0438_ VGND Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q
+ _0437_ sg13g2_o21ai_1
XFILLER_29_336 VPWR VGND sg13g2_fill_1
XFILLER_28_36 VPWR VGND sg13g2_decap_8
X_2429_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q _0890_ _0892_ _0891_ sg13g2_a21oi_1
XFILLER_8_207 VPWR VGND sg13g2_fill_2
X_1800_ net928 Inst_RegFile_32x4.mem\[26\]\[2\] Inst_RegFile_32x4.mem\[27\]\[2\] Inst_RegFile_32x4.mem\[24\]\[2\]
+ Inst_RegFile_32x4.mem\[25\]\[2\] net1027 _0300_ VPWR VGND sg13g2_mux4_1
X_1662_ _0169_ _0168_ Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q VPWR VGND sg13g2_nand2b_1
Xhold229 Inst_RegFile_32x4.mem\[4\]\[3\] VPWR VGND net727 sg13g2_dlygate4sd3_1
X_1731_ _0211_ _0234_ _0235_ VPWR VGND sg13g2_and2_1
X_2780_ net933 net783 _1118_ _0079_ VPWR VGND sg13g2_mux2_1
X_3194_ net1183 net1107 Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q VPWR VGND sg13g2_dlhq_1
X_3263_ net1172 net1117 Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q VPWR VGND sg13g2_dlhq_1
X_2214_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q _0688_ _0690_ _0689_
+ sg13g2_a21oi_1
X_1593_ _1213_ Inst_RegFile_32x4.mem\[10\]\[0\] net928 VPWR VGND sg13g2_nand2b_1
X_3332_ UserCLK net441 Inst_RegFile_32x4.BD_comb\[0\] _3332_/Q_N Inst_RegFile_32x4.BD_reg\[0\]
+ VPWR VGND sg13g2_dfrbp_1
X_2076_ VGND VPWR net1036 _0558_ _0560_ net1008 sg13g2_a21oi_1
XFILLER_34_361 VPWR VGND sg13g2_fill_1
X_2145_ Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q VPWR _0625_ VGND Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q
+ _0623_ sg13g2_o21ai_1
X_1929_ Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q VPWR _0422_ VGND net1038 net987
+ sg13g2_o21ai_1
X_2978_ net1164 net1131 Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q VPWR VGND sg13g2_dlhq_1
XFILLER_57_464 VPWR VGND sg13g2_decap_8
XFILLER_39_46 VPWR VGND sg13g2_decap_8
XFILLER_29_177 VPWR VGND sg13g2_fill_1
XFILLER_25_350 VPWR VGND sg13g2_fill_1
XFILLER_35_125 VPWR VGND sg13g2_fill_2
XFILLER_43_191 VPWR VGND sg13g2_decap_4
X_2832_ _1130_ _1092_ _1101_ VPWR VGND sg13g2_nand2_2
XFILLER_31_375 VPWR VGND sg13g2_fill_2
X_2763_ net949 net765 _1115_ _0065_ VPWR VGND sg13g2_mux2_1
X_2901_ UserCLK net421 _0059_ _2901_/Q_N Inst_RegFile_32x4.mem\[16\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_1714_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q _0219_ _0218_ _0217_
+ sg13g2_a21oi_2
X_1576_ Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q net1074 net38 net50 net9 Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q
+ _1197_ VPWR VGND sg13g2_mux4_1
X_1645_ net1001 net1039 _0153_ VPWR VGND sg13g2_nor2b_1
X_2694_ net937 net812 _1095_ _0016_ VPWR VGND sg13g2_mux2_1
XFILLER_58_217 VPWR VGND sg13g2_fill_1
X_3246_ net1211 net1119 Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q VPWR VGND sg13g2_dlhq_1
XFILLER_39_475 VPWR VGND sg13g2_fill_2
X_3315_ net1198 net1142 Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q VPWR VGND sg13g2_dlhq_1
Xrebuffer11 net527 net509 VPWR VGND sg13g2_buf_2
X_3177_ net1157 net1103 Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q VPWR VGND sg13g2_dlhq_1
XFILLER_54_478 VPWR VGND sg13g2_fill_2
XFILLER_54_467 VPWR VGND sg13g2_decap_8
XFILLER_54_434 VPWR VGND sg13g2_decap_4
X_2059_ VGND VPWR Inst_RegFile_32x4.mem\[11\]\[3\] net994 _0545_ _0544_ sg13g2_a21oi_1
X_2128_ VGND VPWR _0608_ Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q _0606_ Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q
+ _0609_ _0605_ sg13g2_a221oi_1
Xrebuffer44 net543 net542 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer33 Inst_RegFile_switch_matrix.JW2BEG3 net531 VPWR VGND sg13g2_buf_2
Xrebuffer22 _0186_ net520 VPWR VGND sg13g2_buf_8
XFILLER_41_36 VPWR VGND sg13g2_fill_1
XFILLER_40_194 VPWR VGND sg13g2_decap_8
XFILLER_40_183 VPWR VGND sg13g2_fill_1
XFILLER_32_117 VPWR VGND sg13g2_fill_1
X_2908__414 VPWR VGND net414 sg13g2_tiehi
XFILLER_56_7 VPWR VGND sg13g2_decap_8
X_3100_ net1179 net1090 Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q VPWR VGND sg13g2_dlhq_1
X_3031_ net1190 net1081 Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q VPWR VGND sg13g2_dlhq_1
X_2915__407 VPWR VGND net407 sg13g2_tiehi
XFILLER_51_448 VPWR VGND sg13g2_fill_1
XFILLER_51_404 VPWR VGND sg13g2_fill_1
XFILLER_36_456 VPWR VGND sg13g2_fill_1
XFILLER_36_412 VPWR VGND sg13g2_fill_2
XFILLER_31_150 VPWR VGND sg13g2_fill_1
X_2746_ _1092_ _1103_ _1112_ VPWR VGND sg13g2_and2_2
X_2815_ net960 net803 _1126_ _0106_ VPWR VGND sg13g2_mux2_1
X_2677_ net952 net810 _1089_ _0005_ VPWR VGND sg13g2_mux2_1
X_1559_ Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q net44 net72 net15 net723 Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q
+ _1180_ VPWR VGND sg13g2_mux4_1
X_1628_ _0136_ VPWR Inst_RegFile_switch_matrix.JS2BEG3 VGND _0130_ _1234_ sg13g2_o21ai_1
X_3229_ net1176 net1111 Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q VPWR VGND sg13g2_dlhq_1
XFILLER_42_437 VPWR VGND sg13g2_fill_1
XFILLER_22_172 VPWR VGND sg13g2_decap_8
XFILLER_18_401 VPWR VGND sg13g2_fill_2
XFILLER_45_297 VPWR VGND sg13g2_fill_1
XFILLER_45_231 VPWR VGND sg13g2_fill_1
Xrebuffer2 _0388_ net500 VPWR VGND sg13g2_dlygate4sd1_1
X_2600_ Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q net963 net509 _1018_ _1017_ Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q
+ Inst_RegFile_switch_matrix.N1BEG0 VPWR VGND sg13g2_mux4_1
X_3580_ net1159 net184 VPWR VGND sg13g2_buf_1
XFILLER_9_132 VPWR VGND sg13g2_fill_2
X_2531_ _0980_ _0979_ Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q Inst_RegFile_switch_matrix.EE4BEG3
+ VPWR VGND sg13g2_mux2_1
X_2462_ _0921_ _0920_ Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q Inst_RegFile_switch_matrix.WW4BEG3
+ VPWR VGND sg13g2_mux2_1
X_2393_ VGND VPWR net1214 Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q _0858_ _0857_
+ sg13g2_a21oi_1
X_3014_ net1166 net1078 Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q VPWR VGND sg13g2_dlhq_1
XFILLER_36_231 VPWR VGND sg13g2_fill_2
XFILLER_36_220 VPWR VGND sg13g2_fill_2
XFILLER_28_209 VPWR VGND sg13g2_fill_2
XFILLER_32_470 VPWR VGND sg13g2_fill_1
X_2729_ net936 net822 _1107_ _0039_ VPWR VGND sg13g2_mux2_1
XFILLER_59_367 VPWR VGND sg13g2_fill_2
XFILLER_47_529 VPWR VGND sg13g2_fill_2
Xfanout1109 net1114 net1109 VPWR VGND sg13g2_buf_1
X_2905__417 VPWR VGND net417 sg13g2_tiehi
XFILLER_38_529 VPWR VGND sg13g2_fill_2
X_1962_ VGND VPWR _0453_ net97 Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q sg13g2_or2_1
X_3701_ S4END[5] net289 VPWR VGND sg13g2_buf_1
X_3563_ EE4END[7] net151 VPWR VGND sg13g2_buf_1
X_1893_ _0387_ VPWR Inst_RegFile_switch_matrix.JS2BEG6 VGND _0380_ _0373_ sg13g2_o21ai_1
X_3632_ Inst_RegFile_switch_matrix.JN2BEG0 net214 VPWR VGND sg13g2_buf_8
X_2376_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q _0838_ _0842_ _0841_
+ sg13g2_a21oi_1
X_2514_ net1064 net967 _0965_ VPWR VGND sg13g2_nor2b_1
X_2445_ VGND VPWR net1061 net978 _0906_ Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q
+ sg13g2_a21oi_1
XFILLER_45_0 VPWR VGND sg13g2_decap_4
XFILLER_17_38 VPWR VGND sg13g2_fill_2
Xoutput270 net270 S2BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_59_175 VPWR VGND sg13g2_fill_1
XFILLER_47_326 VPWR VGND sg13g2_decap_8
XFILLER_47_304 VPWR VGND sg13g2_fill_1
Xoutput292 net292 S4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput281 net281 S2BEGb[7] VPWR VGND sg13g2_buf_1
XFILLER_55_381 VPWR VGND sg13g2_decap_8
X_2230_ _0705_ _0704_ Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q VPWR VGND sg13g2_nand2b_1
X_2161_ _0636_ Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q _0639_ _0640_ VPWR VGND
+ sg13g2_a21o_1
X_2092_ _0576_ _0575_ net1008 _0574_ _0571_ VPWR VGND sg13g2_a22oi_1
X_2994_ net1202 net1139 Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q VPWR VGND sg13g2_dlhq_1
X_1945_ net43 net14 Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q _0437_ VPWR VGND sg13g2_mux2_1
X_3546_ net19 net128 VPWR VGND sg13g2_buf_1
X_3615_ net1090 net207 VPWR VGND sg13g2_buf_1
X_1876_ _0371_ net948 _0370_ VPWR VGND sg13g2_nand2_1
XFILLER_56_101 VPWR VGND sg13g2_fill_1
X_2428_ Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q _0889_ _0891_ VPWR VGND sg13g2_nor2b_1
X_2359_ Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q _0825_ _0826_ VPWR VGND sg13g2_nor2_1
XFILLER_47_156 VPWR VGND sg13g2_fill_2
X_3343__401 VPWR VGND net401 sg13g2_tiehi
X_1661_ Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q net108 net1019 net980 net514 Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q
+ _0168_ VPWR VGND sg13g2_mux4_1
X_1592_ VGND VPWR Inst_RegFile_32x4.mem\[9\]\[0\] net929 _1212_ _1211_ sg13g2_a21oi_1
X_1730_ _0233_ VPWR _0234_ VGND _1146_ _0230_ sg13g2_o21ai_1
X_3331_ net1162 net1142 Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q VPWR VGND sg13g2_dlhq_1
X_3193_ net1184 net1107 Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q VPWR VGND sg13g2_dlhq_1
X_3262_ net1174 net1117 Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q VPWR VGND sg13g2_dlhq_1
X_2213_ Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q _0687_ _0689_ VPWR VGND sg13g2_nor2b_1
X_2144_ net985 net1001 net1056 _0624_ VPWR VGND sg13g2_mux2_1
X_2075_ Inst_RegFile_32x4.mem\[26\]\[2\] Inst_RegFile_32x4.mem\[27\]\[2\] net993 _0559_
+ VPWR VGND sg13g2_mux2_1
XFILLER_19_381 VPWR VGND sg13g2_fill_1
X_1859_ _0352_ _0354_ _0355_ VPWR VGND sg13g2_nor2_1
X_1928_ net1002 net1038 _0421_ VPWR VGND sg13g2_nor2b_1
X_2977_ net1168 net1131 Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q VPWR VGND sg13g2_dlhq_1
XFILLER_14_39 VPWR VGND sg13g2_fill_2
XFILLER_57_443 VPWR VGND sg13g2_decap_8
XFILLER_55_57 VPWR VGND sg13g2_fill_1
XFILLER_25_362 VPWR VGND sg13g2_fill_2
XFILLER_25_340 VPWR VGND sg13g2_fill_2
XFILLER_4_222 VPWR VGND sg13g2_fill_1
X_2900_ UserCLK net422 _0058_ _2900_/Q_N Inst_RegFile_32x4.mem\[16\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
X_2831_ net743 net935 _1129_ _0119_ VPWR VGND sg13g2_mux2_1
X_1713_ _0218_ net972 net1047 VPWR VGND sg13g2_nand2b_1
XFILLER_31_332 VPWR VGND sg13g2_fill_1
X_2762_ net937 net843 _1115_ _0064_ VPWR VGND sg13g2_mux2_1
X_1575_ Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q VPWR _1196_ VGND _1195_ _1192_
+ sg13g2_o21ai_1
X_3314_ net1201 net1142 Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q VPWR VGND sg13g2_dlhq_1
X_1644_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q _0152_ _0150_ _0151_
+ sg13g2_a21oi_2
X_2693_ _1095_ _1061_ _1094_ VPWR VGND sg13g2_nand2_2
XFILLER_54_446 VPWR VGND sg13g2_decap_8
XFILLER_54_413 VPWR VGND sg13g2_decap_8
XFILLER_54_402 VPWR VGND sg13g2_decap_8
X_3245_ net1149 net1119 Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q VPWR VGND sg13g2_dlhq_1
X_2127_ Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q _0607_ _0608_ VPWR VGND sg13g2_nor2_1
Xrebuffer12 Inst_RegFile_switch_matrix.JN2BEG6 net510 VPWR VGND sg13g2_buf_8
Xrebuffer45 net544 net543 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_26_115 VPWR VGND sg13g2_fill_2
Xrebuffer34 _0491_ net532 VPWR VGND sg13g2_buf_8
X_3176_ net1159 net1104 Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q VPWR VGND sg13g2_dlhq_1
Xrebuffer23 _0429_ net521 VPWR VGND sg13g2_dlygate4sd1_1
X_2058_ net994 Inst_RegFile_32x4.mem\[10\]\[3\] _0544_ VPWR VGND sg13g2_nor2b_1
X_3340__404 VPWR VGND net404 sg13g2_tiehi
XFILLER_17_137 VPWR VGND sg13g2_fill_1
XFILLER_53_490 VPWR VGND sg13g2_fill_1
XFILLER_13_332 VPWR VGND sg13g2_fill_1
XFILLER_49_7 VPWR VGND sg13g2_decap_8
X_3030_ net1192 net1081 Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q VPWR VGND sg13g2_dlhq_1
XFILLER_51_416 VPWR VGND sg13g2_decap_8
X_2676_ net942 net850 _1089_ _0004_ VPWR VGND sg13g2_mux2_1
X_2814_ net952 net770 _1126_ _0105_ VPWR VGND sg13g2_mux2_1
X_2745_ net934 net778 _1111_ _0051_ VPWR VGND sg13g2_mux2_1
XFILLER_59_505 VPWR VGND sg13g2_fill_1
X_1558_ _1179_ VPWR Inst_RegFile_switch_matrix.E2BEG5 VGND _1175_ _1173_ sg13g2_o21ai_1
X_1627_ _0136_ _0135_ Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q VPWR VGND sg13g2_nand2b_1
X_3228_ net1178 net1111 Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q VPWR VGND sg13g2_dlhq_1
X_3159_ net1190 net1101 Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q VPWR VGND sg13g2_dlhq_1
XFILLER_27_435 VPWR VGND sg13g2_fill_2
XFILLER_14_118 VPWR VGND sg13g2_fill_2
XFILLER_52_14 VPWR VGND sg13g2_decap_4
XFILLER_9_100 VPWR VGND sg13g2_fill_2
Xrebuffer3 Inst_RegFile_switch_matrix.JS2BEG5 net501 VPWR VGND sg13g2_dlygate4sd1_1
X_2530_ Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q net1075 net1220 net59 net1019
+ Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q _0980_ VPWR VGND sg13g2_mux4_1
XFILLER_9_166 VPWR VGND sg13g2_fill_1
X_2461_ Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q net1075 net59 net1071 net1018 Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q
+ _0921_ VPWR VGND sg13g2_mux4_1
X_2392_ Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q net6 _0857_ VPWR VGND sg13g2_nor2b_1
X_3013_ net1188 net1078 Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q VPWR VGND sg13g2_dlhq_1
X_3777_ Inst_RegFile_switch_matrix.WW4BEG0 net350 VPWR VGND sg13g2_buf_1
X_2659_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q _1070_ _1074_ _1073_ sg13g2_a21oi_1
X_2728_ net958 net785 _1107_ _0038_ VPWR VGND sg13g2_mux2_1
XFILLER_15_438 VPWR VGND sg13g2_fill_2
XFILLER_15_449 VPWR VGND sg13g2_fill_2
XFILLER_5_0 VPWR VGND sg13g2_fill_2
XFILLER_19_8 VPWR VGND sg13g2_fill_2
XFILLER_18_265 VPWR VGND sg13g2_fill_1
X_3700_ S4END[4] net282 VPWR VGND sg13g2_buf_1
X_1892_ _0386_ VPWR _0387_ VGND Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q _0381_
+ sg13g2_o21ai_1
X_1961_ Inst_RegFile_switch_matrix.JW2BEG6 _0450_ _0452_ _0448_ _0445_ VPWR VGND sg13g2_a22oi_1
XFILLER_14_482 VPWR VGND sg13g2_fill_1
X_3562_ EE4END[6] net150 VPWR VGND sg13g2_buf_1
X_2513_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q
+ _0963_ _0960_ _0964_ _0961_ sg13g2_a221oi_1
X_2375_ Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q VPWR _0841_ VGND Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q
+ _0840_ sg13g2_o21ai_1
X_2444_ VGND VPWR net1061 net971 _0905_ _0904_ sg13g2_a21oi_1
XFILLER_38_0 VPWR VGND sg13g2_fill_2
XFILLER_52_522 VPWR VGND sg13g2_fill_1
Xoutput260 net260 NN4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput293 net293 S4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput282 net282 S4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput271 net271 S2BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_47_338 VPWR VGND sg13g2_decap_4
X_2911__411 VPWR VGND net411 sg13g2_tiehi
XFILLER_11_485 VPWR VGND sg13g2_fill_1
X_2160_ Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q VPWR _0639_ VGND Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q
+ _0638_ sg13g2_o21ai_1
X_2091_ net997 Inst_RegFile_32x4.mem\[12\]\[2\] Inst_RegFile_32x4.mem\[13\]\[2\] Inst_RegFile_32x4.mem\[14\]\[2\]
+ Inst_RegFile_32x4.mem\[15\]\[2\] net947 _0575_ VPWR VGND sg13g2_mux4_1
X_3614_ net1095 net206 VPWR VGND sg13g2_buf_1
X_1875_ VGND VPWR Inst_RegFile_32x4.mem\[11\]\[0\] net994 _0370_ _0369_ sg13g2_a21oi_1
X_1944_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q net98 _0436_ _0435_ sg13g2_a21oi_1
XFILLER_21_238 VPWR VGND sg13g2_fill_1
X_2993_ net1205 net1139 Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q VPWR VGND sg13g2_dlhq_1
X_2427_ net1060 net21 net1214 net63 net90 Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q
+ _0890_ VPWR VGND sg13g2_mux4_1
X_3545_ net18 net127 VPWR VGND sg13g2_buf_1
X_2289_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q _0760_ net1011 net1059
+ sg13g2_a21oi_2
X_2358_ Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q net1065 net963 net979 net970 net1046
+ _0825_ VPWR VGND sg13g2_mux4_1
XFILLER_47_124 VPWR VGND sg13g2_fill_2
X_1591_ net929 Inst_RegFile_32x4.mem\[8\]\[0\] _1211_ VPWR VGND sg13g2_nor2b_1
X_3330_ net1164 net1142 Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q VPWR VGND sg13g2_dlhq_1
X_1660_ _0166_ VPWR _0167_ VGND _0164_ _0162_ sg13g2_o21ai_1
X_3192_ net1186 net1107 Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q VPWR VGND sg13g2_dlhq_1
X_2212_ Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q net1215 net65 net84 net92 Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q
+ _0688_ VPWR VGND sg13g2_mux4_1
X_3261_ net1176 net1117 Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q VPWR VGND sg13g2_dlhq_1
X_2143_ VGND VPWR net1056 net1012 _0623_ _0622_ sg13g2_a21oi_1
X_2074_ VGND VPWR Inst_RegFile_32x4.mem\[25\]\[2\] net993 _0558_ _0557_ sg13g2_a21oi_1
XFILLER_34_396 VPWR VGND sg13g2_fill_1
X_1858_ _1135_ VPWR _0354_ VGND _1134_ _0353_ sg13g2_o21ai_1
X_1927_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q _0420_ _0419_ _0418_
+ sg13g2_a21oi_2
X_2976_ net1170 net1131 Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q VPWR VGND sg13g2_dlhq_1
X_2901__421 VPWR VGND net421 sg13g2_tiehi
X_1789_ net927 Inst_RegFile_32x4.mem\[14\]\[2\] Inst_RegFile_32x4.mem\[15\]\[2\] Inst_RegFile_32x4.mem\[12\]\[2\]
+ Inst_RegFile_32x4.mem\[13\]\[2\] net1026 _0289_ VPWR VGND sg13g2_mux4_1
XFILLER_57_422 VPWR VGND sg13g2_decap_8
XFILLER_55_14 VPWR VGND sg13g2_decap_8
X_2830_ net725 net961 _1129_ _0118_ VPWR VGND sg13g2_mux2_1
X_1712_ _0217_ net1047 net1032 VPWR VGND sg13g2_nand2_2
XFILLER_31_377 VPWR VGND sg13g2_fill_1
X_2761_ _1115_ _1088_ _1097_ VPWR VGND sg13g2_nand2_2
X_1643_ _0151_ net1030 net1039 VPWR VGND sg13g2_nand2b_1
X_2692_ _1030_ _1033_ _1094_ VPWR VGND sg13g2_nor2b_1
X_3244_ net1151 net1119 Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q VPWR VGND sg13g2_dlhq_1
X_1574_ Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q VPWR _1195_ VGND _1193_ _1194_
+ sg13g2_o21ai_1
XFILLER_6_63 VPWR VGND sg13g2_fill_1
X_3313_ net1204 net1143 Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q VPWR VGND sg13g2_dlhq_1
X_2126_ net48 Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q _0607_ VPWR VGND sg13g2_nor2_1
Xfanout1090 net1092 net1090 VPWR VGND sg13g2_buf_1
XFILLER_39_477 VPWR VGND sg13g2_fill_1
Xrebuffer46 net545 net544 VPWR VGND sg13g2_dlygate4sd1_1
X_2057_ VGND VPWR _0540_ net519 _0542_ _0536_ _0543_ _0538_ sg13g2_a221oi_1
XFILLER_26_127 VPWR VGND sg13g2_fill_1
Xrebuffer35 AD2 net533 VPWR VGND sg13g2_buf_8
Xrebuffer24 _0429_ net522 VPWR VGND sg13g2_dlygate4sd1_1
X_3175_ net1160 net1103 Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q VPWR VGND sg13g2_dlhq_1
XFILLER_20_0 VPWR VGND sg13g2_fill_2
Xrebuffer13 Inst_RegFile_switch_matrix.JS2BEG3 net511 VPWR VGND sg13g2_dlygate4sd1_1
X_2959_ net1208 net1132 Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q VPWR VGND sg13g2_dlhq_1
XFILLER_34_182 VPWR VGND sg13g2_fill_2
XFILLER_1_259 VPWR VGND sg13g2_fill_2
XFILLER_45_458 VPWR VGND sg13g2_fill_1
XFILLER_25_171 VPWR VGND sg13g2_fill_2
XFILLER_56_90 VPWR VGND sg13g2_fill_1
XFILLER_36_414 VPWR VGND sg13g2_fill_1
X_2813_ net940 net835 _1126_ _0104_ VPWR VGND sg13g2_mux2_1
XFILLER_16_171 VPWR VGND sg13g2_fill_1
X_2675_ _1089_ _1088_ _1034_ VPWR VGND sg13g2_nand2_2
X_2744_ net960 net766 _1111_ _0050_ VPWR VGND sg13g2_mux2_1
X_1626_ Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q _0132_ _0134_ _0131_ _0133_ Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q
+ _0135_ VPWR VGND sg13g2_mux4_1
XFILLER_59_517 VPWR VGND sg13g2_fill_2
X_3227_ net1181 net1112 Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q VPWR VGND sg13g2_dlhq_1
X_1557_ _1179_ _1178_ Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q VPWR VGND sg13g2_nand2b_1
X_2109_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q _0588_ _0591_ Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q
+ sg13g2_a21oi_1
X_3158_ net1192 net1101 Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q VPWR VGND sg13g2_dlhq_1
X_3089_ net1204 net1091 Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q VPWR VGND sg13g2_dlhq_1
XFILLER_22_141 VPWR VGND sg13g2_fill_2
XFILLER_2_513 VPWR VGND sg13g2_fill_1
XFILLER_7_4 VPWR VGND sg13g2_fill_2
X_2460_ Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q net1030 net499 net500 _0919_ Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q
+ _0920_ VPWR VGND sg13g2_mux4_1
XFILLER_5_340 VPWR VGND sg13g2_fill_1
Xrebuffer4 _0137_ net502 VPWR VGND sg13g2_dlygate4sd1_1
X_2391_ _0855_ VPWR _0856_ VGND Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q _0849_ sg13g2_o21ai_1
X_3012_ net1212 net1079 Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q VPWR VGND sg13g2_dlhq_1
XFILLER_36_233 VPWR VGND sg13g2_fill_1
XFILLER_36_222 VPWR VGND sg13g2_fill_1
X_3776_ WW4END[15] net349 VPWR VGND sg13g2_buf_1
X_1609_ _1228_ VPWR Inst_RegFile_switch_matrix.JS2BEG5 VGND _1222_ _1216_ sg13g2_o21ai_1
X_2589_ Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q net988 _0486_ Inst_RegFile_switch_matrix.JN2BEG2
+ _1016_ Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q Inst_RegFile_switch_matrix.E1BEG3
+ VPWR VGND sg13g2_mux4_1
X_2658_ Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q VPWR _1073_ VGND Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q
+ _1072_ sg13g2_o21ai_1
X_2727_ net949 net834 _1107_ _0037_ VPWR VGND sg13g2_mux2_1
XFILLER_47_15 VPWR VGND sg13g2_decap_8
XFILLER_15_428 VPWR VGND sg13g2_fill_2
XFILLER_2_376 VPWR VGND sg13g2_fill_1
X_1891_ VGND VPWR _0384_ _0385_ _0386_ Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q
+ sg13g2_a21oi_1
X_1960_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q _0451_ _0452_ Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q
+ sg13g2_a21oi_1
X_3561_ EE4END[5] net149 VPWR VGND sg13g2_buf_1
X_2512_ VGND VPWR net1068 net1063 _0963_ _0962_ sg13g2_a21oi_1
X_2443_ net1061 net719 _0904_ VPWR VGND sg13g2_nor2b_1
X_2374_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q net1033 _0840_ _0839_
+ sg13g2_a21oi_1
X_3759_ W6END[8] net343 VPWR VGND sg13g2_buf_1
XFILLER_59_100 VPWR VGND sg13g2_fill_2
Xoutput261 net261 NN4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput250 Inst_RegFile_switch_matrix.NN4BEG1 NN4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput272 net272 S2BEG[6] VPWR VGND sg13g2_buf_1
Xoutput283 net283 S4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput294 net294 S4BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_23_61 VPWR VGND sg13g2_fill_2
XFILLER_15_258 VPWR VGND sg13g2_fill_2
XFILLER_2_140 VPWR VGND sg13g2_fill_1
X_2879__451 VPWR VGND net451 sg13g2_tiehi
XFILLER_38_339 VPWR VGND sg13g2_decap_4
X_2090_ VGND VPWR net1036 _0573_ _0574_ net1008 sg13g2_a21oi_1
XFILLER_31_8 VPWR VGND sg13g2_fill_2
X_2992_ net1207 net1139 Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q VPWR VGND sg13g2_dlhq_1
X_1874_ net994 Inst_RegFile_32x4.mem\[10\]\[0\] _0369_ VPWR VGND sg13g2_nor2b_1
X_3613_ net1102 net205 VPWR VGND sg13g2_buf_1
X_1943_ Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q net71 _0435_ VPWR VGND sg13g2_nor2b_1
XFILLER_50_0 VPWR VGND sg13g2_decap_8
X_2426_ net1060 net35 net51 net1218 net6 Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q
+ _0889_ VPWR VGND sg13g2_mux4_1
X_3544_ net17 net126 VPWR VGND sg13g2_buf_1
XFILLER_29_306 VPWR VGND sg13g2_fill_2
X_2288_ VGND VPWR _0758_ Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q _0757_ Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q
+ _0759_ _0756_ sg13g2_a221oi_1
X_2357_ _0824_ _0823_ Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q VPWR VGND sg13g2_nand2_2
XFILLER_47_158 VPWR VGND sg13g2_fill_1
XFILLER_28_350 VPWR VGND sg13g2_fill_1
XFILLER_7_210 VPWR VGND sg13g2_fill_1
X_3260_ net1178 net1117 Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q VPWR VGND sg13g2_dlhq_1
X_1590_ _1210_ _1206_ _1209_ _1184_ _1181_ VPWR VGND sg13g2_a22oi_1
X_2211_ Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q net31 net37 net53 net8 Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q
+ _0687_ VPWR VGND sg13g2_mux4_1
X_3191_ net1190 net1105 Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q VPWR VGND sg13g2_dlhq_1
X_2073_ net993 Inst_RegFile_32x4.mem\[24\]\[2\] _0557_ VPWR VGND sg13g2_nor2b_1
X_2142_ net1056 net1029 _0622_ VPWR VGND sg13g2_nor2b_1
X_2975_ net1173 net1134 Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q VPWR VGND sg13g2_dlhq_1
X_1857_ Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q net24 net59 net61 net67 Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q
+ _0353_ VPWR VGND sg13g2_mux4_1
X_1926_ _0419_ net973 Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q VPWR VGND sg13g2_nand2b_1
X_1788_ _0288_ net956 _0287_ VPWR VGND sg13g2_nand2_1
XFILLER_57_401 VPWR VGND sg13g2_decap_8
X_2409_ net62 net1072 net1051 _0873_ VPWR VGND sg13g2_mux2_1
X_3389_ UserCLK net491 _0125_ _3389_/Q_N Inst_RegFile_32x4.mem\[12\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_2869__461 VPWR VGND net461 sg13g2_tiehi
X_2917__440 VPWR VGND net440 sg13g2_tiehi
X_2876__454 VPWR VGND net454 sg13g2_tiehi
XFILLER_35_106 VPWR VGND sg13g2_fill_2
XFILLER_29_71 VPWR VGND sg13g2_fill_1
XFILLER_29_60 VPWR VGND sg13g2_fill_1
XFILLER_43_150 VPWR VGND sg13g2_fill_1
X_2883__447 VPWR VGND net447 sg13g2_tiehi
X_1711_ VGND VPWR _0215_ Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q _0214_ Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q
+ _0216_ _0213_ sg13g2_a221oi_1
X_2691_ net935 net849 _1093_ _0015_ VPWR VGND sg13g2_mux2_1
X_2760_ net932 net837 _1114_ _0063_ VPWR VGND sg13g2_mux2_1
X_1642_ _0150_ net1039 net1012 VPWR VGND sg13g2_nand2_2
X_1573_ Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q VPWR _1194_ VGND net1048 net985
+ sg13g2_o21ai_1
X_3243_ net1152 net1115 Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q VPWR VGND sg13g2_dlhq_1
X_3312_ net1206 net1143 Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q VPWR VGND sg13g2_dlhq_1
X_2125_ _0606_ Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q net19 VPWR VGND sg13g2_nand2b_1
XFILLER_39_456 VPWR VGND sg13g2_fill_2
Xfanout1080 net1081 net1080 VPWR VGND sg13g2_buf_1
XFILLER_34_150 VPWR VGND sg13g2_decap_8
Xrebuffer47 net546 net545 VPWR VGND sg13g2_dlygate4sd1_1
X_2056_ VGND VPWR net943 _0542_ _0541_ net1005 sg13g2_a21oi_2
Xrebuffer25 Inst_RegFile_switch_matrix.JW2BEG4 net523 VPWR VGND sg13g2_dlygate4sd1_1
X_3174_ net1166 net1103 Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q VPWR VGND sg13g2_dlhq_1
XFILLER_13_0 VPWR VGND sg13g2_fill_1
Xrebuffer14 Inst_RegFile_switch_matrix.JS2BEG3 net512 VPWR VGND sg13g2_dlygate4sd1_1
Xfanout1091 net1092 net1091 VPWR VGND sg13g2_buf_1
X_2958_ net1210 net1135 Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q VPWR VGND sg13g2_dlhq_1
X_1909_ Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q net1075 net39 net1220 net10 Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q
+ _0403_ VPWR VGND sg13g2_mux4_1
X_2889_ UserCLK net433 _0047_ _2889_/Q_N Inst_RegFile_32x4.mem\[23\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_48_264 VPWR VGND sg13g2_fill_2
X_2812_ _1126_ _1092_ _1122_ VPWR VGND sg13g2_nand2_2
X_2743_ net954 net806 _1111_ _0049_ VPWR VGND sg13g2_mux2_1
X_1556_ _1176_ _1177_ _1141_ _1178_ VPWR VGND sg13g2_mux2_1
X_2674_ _1058_ _1047_ _1059_ _1088_ VPWR VGND sg13g2_nor3_2
X_2859__471 VPWR VGND net471 sg13g2_tiehi
X_1625_ net1217 net66 Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q _0134_ VPWR VGND
+ sg13g2_mux2_1
X_3226_ net1183 net1112 Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q VPWR VGND sg13g2_dlhq_1
X_3157_ net1194 net1100 Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q VPWR VGND sg13g2_dlhq_1
X_2108_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q net1017 _0590_ _0589_
+ sg13g2_a21oi_1
XFILLER_27_437 VPWR VGND sg13g2_fill_1
X_3088_ net1207 net1091 Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q VPWR VGND sg13g2_dlhq_1
XFILLER_22_120 VPWR VGND sg13g2_decap_4
X_2039_ net990 Inst_RegFile_32x4.mem\[0\]\[1\] Inst_RegFile_32x4.mem\[1\]\[1\] Inst_RegFile_32x4.mem\[2\]\[1\]
+ Inst_RegFile_32x4.mem\[3\]\[1\] net944 _0527_ VPWR VGND sg13g2_mux4_1
X_2866__464 VPWR VGND net464 sg13g2_tiehi
XFILLER_52_49 VPWR VGND sg13g2_fill_1
XFILLER_6_319 VPWR VGND sg13g2_fill_2
X_2873__457 VPWR VGND net457 sg13g2_tiehi
XFILLER_33_407 VPWR VGND sg13g2_fill_1
XFILLER_9_102 VPWR VGND sg13g2_fill_1
XFILLER_13_153 VPWR VGND sg13g2_decap_4
XFILLER_54_7 VPWR VGND sg13g2_decap_8
Xrebuffer5 Inst_RegFile_switch_matrix.JS2BEG3 net503 VPWR VGND sg13g2_dlygate4sd1_1
X_3011_ net1162 net1138 Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q VPWR VGND sg13g2_dlhq_1
XFILLER_3_65 VPWR VGND sg13g2_decap_8
X_2390_ _0854_ Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q _0855_ VPWR VGND sg13g2_nor2b_1
X_3775_ WW4END[14] net348 VPWR VGND sg13g2_buf_1
X_2726_ net938 net798 _1107_ _0036_ VPWR VGND sg13g2_mux2_1
X_1608_ _1228_ _1227_ Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q VPWR VGND sg13g2_nand2b_1
X_1539_ VPWR _1161_ Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q VGND sg13g2_inv_1
X_2588_ Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q net1030 Inst_RegFile_switch_matrix.E2BEG3
+ _1018_ _1017_ Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q Inst_RegFile_switch_matrix.S1BEG0
+ VPWR VGND sg13g2_mux4_1
X_2657_ VGND VPWR net1216 Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q _1072_ _1071_
+ sg13g2_a21oi_1
XFILLER_47_49 VPWR VGND sg13g2_fill_1
X_3209_ net1156 net1109 Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q VPWR VGND sg13g2_dlhq_1
XFILLER_42_237 VPWR VGND sg13g2_fill_2
XFILLER_5_2 VPWR VGND sg13g2_fill_1
XFILLER_58_381 VPWR VGND sg13g2_decap_8
X_2849__481 VPWR VGND net481 sg13g2_tiehi
X_3560_ EE4END[4] net142 VPWR VGND sg13g2_buf_1
X_1890_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q _0382_ _0385_ _1136_
+ sg13g2_a21oi_1
XFILLER_41_292 VPWR VGND sg13g2_fill_2
XFILLER_41_281 VPWR VGND sg13g2_decap_8
X_2373_ Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q net974 _0839_ VPWR VGND sg13g2_nor2b_1
X_2511_ net1063 net82 _0962_ VPWR VGND sg13g2_nor2b_1
X_2442_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q
+ _0902_ _0899_ _0903_ _0900_ sg13g2_a221oi_1
XFILLER_38_2 VPWR VGND sg13g2_fill_1
X_2856__474 VPWR VGND net474 sg13g2_tiehi
XFILLER_32_292 VPWR VGND sg13g2_fill_1
XFILLER_24_204 VPWR VGND sg13g2_fill_1
X_2863__467 VPWR VGND net467 sg13g2_tiehi
X_3689_ net501 net271 VPWR VGND sg13g2_buf_1
X_3758_ W6END[7] net342 VPWR VGND sg13g2_buf_1
X_2709_ net933 net787 _1099_ _0027_ VPWR VGND sg13g2_mux2_1
XFILLER_59_156 VPWR VGND sg13g2_fill_2
Xoutput240 net240 N4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput251 net251 NN4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput284 net284 S4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput295 net295 S4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput273 net273 S2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput262 Inst_RegFile_switch_matrix.S1BEG0 S1BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_55_395 VPWR VGND sg13g2_decap_8
XFILLER_23_73 VPWR VGND sg13g2_fill_2
XFILLER_23_40 VPWR VGND sg13g2_fill_1
XFILLER_24_8 VPWR VGND sg13g2_fill_2
XFILLER_0_44 VPWR VGND sg13g2_fill_2
XFILLER_0_88 VPWR VGND sg13g2_fill_2
XFILLER_9_20 VPWR VGND sg13g2_fill_2
X_1942_ _0430_ Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q _0433_ _0434_ VPWR VGND sg13g2_a21o_1
X_2991_ net1209 net1139 Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q VPWR VGND sg13g2_dlhq_1
X_3612_ net1108 net204 VPWR VGND sg13g2_buf_1
X_3543_ net16 net125 VPWR VGND sg13g2_buf_1
X_1873_ _0368_ _0341_ _0366_ VPWR VGND sg13g2_nand2_1
XFILLER_43_0 VPWR VGND sg13g2_decap_4
X_2356_ _0822_ VPWR _0823_ VGND net1046 net1029 sg13g2_o21ai_1
X_2425_ _0882_ Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q _0887_ _0888_ VPWR VGND sg13g2_nand3_1
X_2287_ VGND VPWR net1059 _1166_ _0758_ Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q
+ sg13g2_a21oi_1
XFILLER_18_62 VPWR VGND sg13g2_fill_1
XFILLER_28_362 VPWR VGND sg13g2_fill_2
XFILLER_18_73 VPWR VGND sg13g2_fill_1
X_2846__484 VPWR VGND net484 sg13g2_tiehi
XFILLER_34_83 VPWR VGND sg13g2_decap_8
X_2210_ VGND VPWR _0686_ _0685_ _0684_ sg13g2_or2_1
X_3190_ net1192 net1105 Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q VPWR VGND sg13g2_dlhq_1
XFILLER_53_118 VPWR VGND sg13g2_fill_2
X_2853__477 VPWR VGND net477 sg13g2_tiehi
X_2072_ Inst_RegFile_32x4.BD_comb\[3\] Inst_RegFile_32x4.BD_reg\[3\] Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q
+ BD3 VPWR VGND sg13g2_mux2_2
X_2141_ _0620_ VPWR _0621_ VGND Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q _0619_
+ sg13g2_o21ai_1
XFILLER_15_4 VPWR VGND sg13g2_fill_2
X_2974_ net1174 net1134 Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q VPWR VGND sg13g2_dlhq_1
X_1925_ _0418_ Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q net1014 VPWR VGND sg13g2_nand2_1
X_1787_ net929 Inst_RegFile_32x4.mem\[10\]\[2\] Inst_RegFile_32x4.mem\[11\]\[2\] Inst_RegFile_32x4.mem\[8\]\[2\]
+ Inst_RegFile_32x4.mem\[9\]\[2\] net1027 _0287_ VPWR VGND sg13g2_mux4_1
X_1856_ Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q _0351_ _0352_ VPWR VGND sg13g2_nor2_1
X_2408_ net5 net58 net1051 _0872_ VPWR VGND sg13g2_mux2_1
XFILLER_57_457 VPWR VGND sg13g2_decap_8
X_2339_ net979 net966 net1042 _0807_ VPWR VGND sg13g2_mux2_1
X_3388_ UserCLK net492 _0124_ _3388_/Q_N Inst_RegFile_32x4.mem\[12\]\[0\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_43_195 VPWR VGND sg13g2_fill_1
X_1710_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q net1016 _0215_ Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q
+ sg13g2_a21oi_1
X_2690_ net960 net819 _1093_ _0014_ VPWR VGND sg13g2_mux2_1
X_1572_ net1001 net1048 _1193_ VPWR VGND sg13g2_nor2b_1
X_3311_ net1208 net1147 Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q VPWR VGND sg13g2_dlhq_1
X_1641_ VGND VPWR _0148_ Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q _0147_ _0146_
+ _0149_ Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q sg13g2_a221oi_1
Xfanout1070 net88 net1070 VPWR VGND sg13g2_buf_1
X_2124_ net76 net510 Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q _0605_ VPWR VGND sg13g2_mux2_1
Xfanout1081 net29 net1081 VPWR VGND sg13g2_buf_1
X_3242_ net1154 net1115 Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q VPWR VGND sg13g2_dlhq_1
Xfanout1092 FrameStrobe[7] net1092 VPWR VGND sg13g2_buf_1
X_3173_ net1188 net1103 Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q VPWR VGND sg13g2_dlhq_1
XFILLER_20_2 VPWR VGND sg13g2_fill_1
XFILLER_54_427 VPWR VGND sg13g2_decap_8
XFILLER_34_184 VPWR VGND sg13g2_fill_1
Xrebuffer48 net547 net546 VPWR VGND sg13g2_dlygate4sd1_1
Xrebuffer26 Inst_RegFile_switch_matrix.JW2BEG4 net524 VPWR VGND sg13g2_dlygate4sd1_1
X_2055_ net991 Inst_RegFile_32x4.mem\[20\]\[3\] Inst_RegFile_32x4.mem\[21\]\[3\] Inst_RegFile_32x4.mem\[22\]\[3\]
+ Inst_RegFile_32x4.mem\[23\]\[3\] net945 _0541_ VPWR VGND sg13g2_mux4_1
Xrebuffer15 net513 net533 VPWR VGND sg13g2_buf_16
X_2957_ net1148 net1133 Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q VPWR VGND sg13g2_dlhq_1
X_1908_ Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q VPWR _0402_ VGND _0401_ _0400_
+ sg13g2_o21ai_1
XFILLER_41_29 VPWR VGND sg13g2_decap_8
X_1839_ _0337_ _0336_ net969 _0328_ _0326_ VPWR VGND sg13g2_a22oi_1
X_2888_ UserCLK net434 _0046_ _2888_/Q_N Inst_RegFile_32x4.mem\[23\]\[2\] VPWR VGND
+ sg13g2_dfrbp_1
XFILLER_53_471 VPWR VGND sg13g2_decap_4
XFILLER_15_74 VPWR VGND sg13g2_fill_2
X_2843__487 VPWR VGND net487 sg13g2_tiehi
X_3388__492 VPWR VGND net492 sg13g2_tiehi
X_2742_ net940 net756 _1111_ _0048_ VPWR VGND sg13g2_mux2_1
X_2811_ net737 net934 _1125_ _0103_ VPWR VGND sg13g2_mux2_1
X_1555_ Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q net32 net40 net3 net11 Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q
+ _1177_ VPWR VGND sg13g2_mux4_1
X_2673_ net935 net799 _1062_ _0003_ VPWR VGND sg13g2_mux2_1
X_1624_ net78 net93 Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q _0133_ VPWR VGND sg13g2_mux2_1
X_3225_ net1185 net1112 Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q VPWR VGND sg13g2_dlhq_1
X_2107_ Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q net1068 _0589_ VPWR VGND sg13g2_nor2b_1
X_3156_ net1196 net1102 Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q VPWR VGND sg13g2_dlhq_1
XFILLER_39_298 VPWR VGND sg13g2_decap_8
X_3087_ net1208 net1089 Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q VPWR VGND sg13g2_dlhq_1
X_2038_ VGND VPWR net1006 _0525_ _0526_ _0459_ sg13g2_a21oi_1
XFILLER_22_165 VPWR VGND sg13g2_decap_8
XFILLER_22_143 VPWR VGND sg13g2_fill_1
Xhold350 Inst_RegFile_32x4.mem\[16\]\[2\] VPWR VGND net848 sg13g2_dlygate4sd3_1
XFILLER_42_94 VPWR VGND sg13g2_decap_8
Xrebuffer6 net525 net504 VPWR VGND sg13g2_buf_8
X_3010_ net1164 net1138 Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q VPWR VGND sg13g2_dlhq_1
X_3774_ WW4END[13] net362 VPWR VGND sg13g2_buf_1
X_2656_ Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q net50 _1071_ VPWR VGND sg13g2_nor2b_1
X_2725_ _1107_ _1088_ _1106_ VPWR VGND sg13g2_nand2_2
XFILLER_59_338 VPWR VGND sg13g2_fill_2
X_1607_ Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q _1224_ _1226_ _1223_ _1225_ Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q
+ _1227_ VPWR VGND sg13g2_mux4_1
X_1538_ VPWR _1160_ Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q VGND sg13g2_inv_1
X_2587_ Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q net1015 _0645_ Inst_RegFile_switch_matrix.E2BEG0
+ _0137_ Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q Inst_RegFile_switch_matrix.S1BEG1
+ VPWR VGND sg13g2_mux4_1
X_3139_ net1162 net1093 Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q VPWR VGND sg13g2_dlhq_1
X_3208_ net1158 net1109 Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q VPWR VGND sg13g2_dlhq_1
XFILLER_10_179 VPWR VGND sg13g2_fill_1
X_3385__495 VPWR VGND net495 sg13g2_tiehi
XFILLER_37_50 VPWR VGND sg13g2_decap_4
XFILLER_33_227 VPWR VGND sg13g2_fill_1
X_2510_ VGND VPWR net1218 net1064 _0961_ Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q
+ sg13g2_a21oi_1
X_2372_ _0837_ VPWR _0838_ VGND Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q net1011
+ sg13g2_o21ai_1
X_2441_ VGND VPWR net1068 net1061 _0902_ _0901_ sg13g2_a21oi_1
XFILLER_45_4 VPWR VGND sg13g2_fill_1
XFILLER_5_150 VPWR VGND sg13g2_fill_1
XFILLER_52_503 VPWR VGND sg13g2_fill_1
XFILLER_49_393 VPWR VGND sg13g2_fill_2
Xoutput252 net252 NN4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput241 net241 N4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput230 net230 N4BEG[0] VPWR VGND sg13g2_buf_1
X_3688_ Inst_RegFile_switch_matrix.JS2BEG4 net270 VPWR VGND sg13g2_buf_1
X_3757_ W6END[6] net341 VPWR VGND sg13g2_buf_1
X_2708_ net959 net842 _1099_ _0026_ VPWR VGND sg13g2_mux2_1
X_2639_ _1056_ VPWR _1057_ VGND net37 Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q sg13g2_o21ai_1
XFILLER_59_102 VPWR VGND sg13g2_fill_1
Xoutput263 Inst_RegFile_switch_matrix.S1BEG1 S1BEG[1] VPWR VGND sg13g2_buf_1
Xoutput296 net296 S4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput274 net274 S2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput285 net285 S4BEG[12] VPWR VGND sg13g2_buf_1
X_1872_ _0341_ _0366_ _0367_ VPWR VGND sg13g2_and2_1
X_1941_ Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q VPWR _0433_ VGND Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q
+ _0431_ sg13g2_o21ai_1
XFILLER_14_282 VPWR VGND sg13g2_fill_2
X_2990_ net1210 net1139 Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q VPWR VGND sg13g2_dlhq_1
X_3611_ net1112 net203 VPWR VGND sg13g2_buf_1
X_3542_ net15 net124 VPWR VGND sg13g2_buf_1
XFILLER_56_127 VPWR VGND sg13g2_fill_2
XFILLER_36_0 VPWR VGND sg13g2_fill_2
XFILLER_29_308 VPWR VGND sg13g2_fill_1
X_2286_ VGND VPWR _0757_ net1059 net1066 sg13g2_or2_1
X_2355_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q _0822_ net1010 net1046
+ sg13g2_a21oi_2
X_2424_ Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q _0886_ _0884_ _0887_ VPWR VGND sg13g2_nand3_1
XFILLER_37_330 VPWR VGND sg13g2_decap_4
XFILLER_25_503 VPWR VGND sg13g2_fill_2
XFILLER_52_399 VPWR VGND sg13g2_decap_4
X_3336__445 VPWR VGND net445 sg13g2_tiehi
X_3382__498 VPWR VGND net498 sg13g2_tiehi
XFILLER_43_322 VPWR VGND sg13g2_decap_8
XFILLER_7_201 VPWR VGND sg13g2_fill_2
X_2140_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q _0617_ _0620_ Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q
+ sg13g2_a21oi_1
XFILLER_46_160 VPWR VGND sg13g2_fill_2
XFILLER_34_333 VPWR VGND sg13g2_fill_2
X_2071_ _0556_ net519 _0543_ Inst_RegFile_32x4.BD_comb\[3\] VPWR VGND sg13g2_a21o_1
XFILLER_19_352 VPWR VGND sg13g2_fill_2
X_2973_ net1176 net1134 Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q VPWR VGND sg13g2_dlhq_1
X_1855_ Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q net1075 net39 net1220 net10 Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q
+ _0351_ VPWR VGND sg13g2_mux4_1
X_1924_ VGND VPWR _0416_ Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q _0415_ Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q
+ _0417_ _0414_ sg13g2_a221oi_1
X_1786_ Inst_RegFile_32x4.AD_comb\[1\] Inst_RegFile_32x4.AD_reg\[1\] Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q
+ AD1 VPWR VGND sg13g2_mux2_2
X_2338_ _0805_ VPWR _0806_ VGND _0803_ _1149_ sg13g2_o21ai_1
XFILLER_57_436 VPWR VGND sg13g2_decap_8
X_2407_ Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q VPWR _0871_ VGND Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q
+ _0870_ sg13g2_o21ai_1
XFILLER_55_28 VPWR VGND sg13g2_decap_4
X_3387_ UserCLK net493 _0123_ _3387_/Q_N Inst_RegFile_32x4.mem\[11\]\[3\] VPWR VGND
+ sg13g2_dfrbp_1
X_2269_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q _0741_ net1010 net1050
+ sg13g2_a21oi_2
XFILLER_16_311 VPWR VGND sg13g2_fill_1
X_1571_ VGND VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q _1192_ _1190_ _1191_
+ sg13g2_a21oi_2
X_3310_ net1210 net1147 Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q VPWR VGND sg13g2_dlhq_1
XFILLER_6_44 VPWR VGND sg13g2_fill_2
X_1640_ VGND VPWR net1039 net1016 _0148_ Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q
+ sg13g2_a21oi_1
Xrebuffer16 net513 net514 VPWR VGND sg13g2_dlygate4sd1_1
X_2123_ Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q VPWR _0604_ VGND Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q
+ _0603_ sg13g2_o21ai_1
Xfanout1071 net87 net1071 VPWR VGND sg13g2_buf_8
Xfanout1082 net29 net1082 VPWR VGND sg13g2_buf_1
Xrebuffer27 AD2 net525 VPWR VGND sg13g2_buf_2
Xfanout1093 net1094 net1093 VPWR VGND sg13g2_buf_1
X_3241_ net1156 net1115 Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q VPWR VGND sg13g2_dlhq_1
X_3172_ net1212 net1103 Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q VPWR VGND sg13g2_dlhq_1
Xfanout1060 Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q net1060 VPWR VGND sg13g2_buf_1
Xrebuffer49 net548 net547 VPWR VGND sg13g2_dlygate4sd1_1
X_2054_ _0540_ _0539_ net1005 VPWR VGND sg13g2_nand2b_1
X_2956_ net1150 net1133 Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q VPWR VGND sg13g2_dlhq_1
X_1907_ Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q VPWR _0401_ VGND _0396_ _0397_
+ sg13g2_o21ai_1
X_2899__423 VPWR VGND net423 sg13g2_tiehi
X_1838_ _0336_ _0334_ _0335_ _0329_ net955 VPWR VGND sg13g2_a22oi_1
X_2887_ UserCLK net435 _0045_ _2887_/Q_N Inst_RegFile_32x4.mem\[23\]\[1\] VPWR VGND
+ sg13g2_dfrbp_1
X_1769_ net928 Inst_RegFile_32x4.mem\[24\]\[1\] _0271_ VPWR VGND sg13g2_nor2b_1
XFILLER_53_450 VPWR VGND sg13g2_decap_8
XFILLER_9_318 VPWR VGND sg13g2_fill_2
XFILLER_48_266 VPWR VGND sg13g2_fill_1
XFILLER_51_409 VPWR VGND sg13g2_decap_8
XFILLER_44_483 VPWR VGND sg13g2_fill_2
XFILLER_44_450 VPWR VGND sg13g2_fill_1
X_2810_ net729 net960 _1125_ _0102_ VPWR VGND sg13g2_mux2_1
X_2672_ _1086_ VPWR _1087_ VGND _1074_ _1075_ sg13g2_o21ai_1
X_2741_ _1111_ _1090_ _1103_ VPWR VGND sg13g2_nand2_2
X_3224_ net1187 net1112 Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q VPWR VGND sg13g2_dlhq_1
X_1554_ Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q net23 net58 net60 net68 Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q
+ _1176_ VPWR VGND sg13g2_mux4_1
X_1623_ net38 net1219 Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q _0132_ VPWR VGND
+ sg13g2_mux2_1
.ends

