magic
tech sky130A
magscale 1 2
timestamp 1740383427
<< viali >>
rect 1501 8585 1535 8619
rect 3893 8585 3927 8619
rect 6469 8585 6503 8619
rect 8585 8585 8619 8619
rect 10885 8585 10919 8619
rect 13185 8585 13219 8619
rect 15485 8585 15519 8619
rect 17693 8585 17727 8619
rect 19993 8585 20027 8619
rect 22293 8585 22327 8619
rect 24593 8585 24627 8619
rect 27077 8585 27111 8619
rect 29193 8585 29227 8619
rect 31493 8585 31527 8619
rect 33793 8585 33827 8619
rect 36093 8585 36127 8619
rect 38393 8585 38427 8619
rect 40693 8585 40727 8619
rect 42993 8585 43027 8619
rect 45293 8585 45327 8619
rect 45845 8585 45879 8619
rect 46213 8585 46247 8619
rect 46949 8585 46983 8619
rect 1685 8449 1719 8483
rect 4077 8449 4111 8483
rect 6653 8449 6687 8483
rect 8401 8449 8435 8483
rect 10701 8449 10735 8483
rect 13001 8449 13035 8483
rect 15301 8449 15335 8483
rect 17877 8449 17911 8483
rect 20177 8449 20211 8483
rect 22477 8449 22511 8483
rect 24777 8449 24811 8483
rect 27261 8449 27295 8483
rect 29377 8449 29411 8483
rect 31677 8449 31711 8483
rect 33977 8449 34011 8483
rect 36289 8449 36323 8483
rect 38577 8449 38611 8483
rect 40877 8449 40911 8483
rect 43177 8449 43211 8483
rect 45477 8449 45511 8483
rect 45661 8449 45695 8483
rect 46029 8449 46063 8483
rect 46397 8449 46431 8483
rect 46765 8449 46799 8483
rect 47133 8449 47167 8483
rect 46581 8313 46615 8347
rect 47317 8313 47351 8347
rect 8309 8041 8343 8075
rect 10241 8041 10275 8075
rect 19533 8041 19567 8075
rect 20545 8041 20579 8075
rect 20637 8041 20671 8075
rect 21741 8041 21775 8075
rect 22109 8041 22143 8075
rect 23489 8041 23523 8075
rect 23949 8041 23983 8075
rect 26065 8041 26099 8075
rect 26525 8041 26559 8075
rect 29837 8041 29871 8075
rect 37841 8041 37875 8075
rect 46673 8041 46707 8075
rect 2237 7905 2271 7939
rect 2053 7837 2087 7871
rect 8033 7837 8067 7871
rect 8125 7837 8159 7871
rect 10057 7837 10091 7871
rect 11989 7837 12023 7871
rect 15945 7837 15979 7871
rect 19349 7837 19383 7871
rect 19625 7837 19659 7871
rect 20361 7837 20395 7871
rect 20821 7837 20855 7871
rect 20913 7837 20947 7871
rect 21833 7837 21867 7871
rect 21925 7837 21959 7871
rect 23305 7837 23339 7871
rect 23673 7837 23707 7871
rect 23765 7837 23799 7871
rect 24041 7837 24075 7871
rect 25605 7837 25639 7871
rect 25973 7837 26007 7871
rect 26249 7837 26283 7871
rect 26341 7837 26375 7871
rect 29561 7837 29595 7871
rect 30021 7837 30055 7871
rect 35265 7837 35299 7871
rect 35357 7837 35391 7871
rect 38025 7837 38059 7871
rect 39589 7837 39623 7871
rect 40325 7837 40359 7871
rect 40601 7837 40635 7871
rect 45385 7837 45419 7871
rect 45661 7837 45695 7871
rect 46029 7837 46063 7871
rect 46121 7837 46155 7871
rect 46489 7837 46523 7871
rect 46857 7837 46891 7871
rect 47225 7837 47259 7871
rect 8033 7701 8067 7735
rect 12173 7701 12207 7735
rect 16129 7701 16163 7735
rect 21097 7701 21131 7735
rect 29745 7701 29779 7735
rect 35173 7701 35207 7735
rect 35541 7701 35575 7735
rect 39405 7701 39439 7735
rect 40233 7701 40267 7735
rect 40417 7701 40451 7735
rect 45293 7701 45327 7735
rect 45477 7701 45511 7735
rect 45845 7701 45879 7735
rect 46305 7701 46339 7735
rect 47041 7701 47075 7735
rect 47409 7701 47443 7735
rect 12265 7497 12299 7531
rect 15025 7497 15059 7531
rect 17877 7497 17911 7531
rect 38117 7497 38151 7531
rect 38761 7497 38795 7531
rect 39589 7497 39623 7531
rect 40785 7497 40819 7531
rect 46673 7497 46707 7531
rect 46949 7497 46983 7531
rect 11621 7429 11655 7463
rect 11805 7361 11839 7395
rect 11989 7361 12023 7395
rect 12081 7361 12115 7395
rect 14841 7361 14875 7395
rect 18061 7361 18095 7395
rect 23029 7361 23063 7395
rect 23121 7361 23155 7395
rect 33149 7361 33183 7395
rect 33241 7361 33275 7395
rect 38209 7361 38243 7395
rect 38853 7361 38887 7395
rect 39773 7361 39807 7395
rect 40969 7361 41003 7395
rect 46489 7361 46523 7395
rect 46765 7361 46799 7395
rect 47133 7361 47167 7395
rect 11989 7157 12023 7191
rect 22937 7157 22971 7191
rect 23305 7157 23339 7191
rect 33149 7157 33183 7191
rect 33425 7157 33459 7191
rect 47317 7157 47351 7191
rect 46213 6953 46247 6987
rect 27077 6885 27111 6919
rect 18429 6817 18463 6851
rect 26709 6817 26743 6851
rect 26065 6749 26099 6783
rect 26157 6749 26191 6783
rect 26801 6749 26835 6783
rect 26893 6749 26927 6783
rect 40233 6749 40267 6783
rect 41521 6749 41555 6783
rect 44741 6749 44775 6783
rect 46029 6749 46063 6783
rect 46397 6749 46431 6783
rect 46673 6749 46707 6783
rect 46857 6749 46891 6783
rect 47225 6749 47259 6783
rect 15577 6681 15611 6715
rect 15853 6681 15887 6715
rect 18521 6681 18555 6715
rect 18705 6681 18739 6715
rect 18889 6681 18923 6715
rect 15945 6613 15979 6647
rect 25973 6613 26007 6647
rect 26341 6613 26375 6647
rect 40049 6613 40083 6647
rect 41337 6613 41371 6647
rect 44557 6613 44591 6647
rect 46489 6613 46523 6647
rect 47041 6613 47075 6647
rect 47409 6613 47443 6647
rect 42441 6409 42475 6443
rect 47317 6409 47351 6443
rect 22017 6273 22051 6307
rect 33609 6273 33643 6307
rect 33793 6273 33827 6307
rect 42625 6273 42659 6307
rect 43545 6273 43579 6307
rect 46581 6273 46615 6307
rect 47041 6273 47075 6307
rect 47133 6273 47167 6307
rect 43361 6137 43395 6171
rect 22201 6069 22235 6103
rect 33977 6069 34011 6103
rect 46765 6069 46799 6103
rect 46949 6069 46983 6103
rect 8677 5865 8711 5899
rect 17969 5865 18003 5899
rect 19533 5865 19567 5899
rect 18429 5797 18463 5831
rect 47409 5797 47443 5831
rect 8493 5661 8527 5695
rect 14565 5661 14599 5695
rect 18061 5661 18095 5695
rect 18245 5661 18279 5695
rect 19625 5661 19659 5695
rect 19717 5661 19751 5695
rect 32781 5661 32815 5695
rect 32965 5661 32999 5695
rect 46857 5661 46891 5695
rect 47225 5661 47259 5695
rect 14749 5525 14783 5559
rect 19901 5525 19935 5559
rect 33149 5525 33183 5559
rect 47041 5525 47075 5559
rect 8585 5321 8619 5355
rect 17693 5321 17727 5355
rect 22017 5321 22051 5355
rect 23857 5321 23891 5355
rect 25145 5321 25179 5355
rect 47317 5321 47351 5355
rect 8125 5185 8159 5219
rect 8401 5185 8435 5219
rect 9229 5185 9263 5219
rect 10425 5185 10459 5219
rect 11161 5185 11195 5219
rect 12357 5185 12391 5219
rect 12725 5185 12759 5219
rect 13763 5185 13797 5219
rect 15301 5185 15335 5219
rect 16313 5185 16347 5219
rect 17049 5185 17083 5219
rect 17509 5185 17543 5219
rect 21833 5209 21867 5243
rect 23581 5185 23615 5219
rect 23673 5185 23707 5219
rect 23949 5185 23983 5219
rect 24961 5185 24995 5219
rect 26985 5185 27019 5219
rect 27261 5185 27295 5219
rect 27445 5185 27479 5219
rect 46765 5185 46799 5219
rect 47133 5185 47167 5219
rect 22109 5117 22143 5151
rect 23305 5117 23339 5151
rect 12541 5049 12575 5083
rect 16497 5049 16531 5083
rect 8309 4981 8343 5015
rect 9413 4981 9447 5015
rect 10609 4981 10643 5015
rect 11345 4981 11379 5015
rect 12909 4981 12943 5015
rect 13921 4981 13955 5015
rect 15485 4981 15519 5015
rect 17233 4981 17267 5015
rect 23213 4981 23247 5015
rect 23489 4981 23523 5015
rect 24133 4981 24167 5015
rect 27169 4981 27203 5015
rect 27629 4981 27663 5015
rect 46949 4981 46983 5015
rect 4169 4777 4203 4811
rect 2881 4709 2915 4743
rect 47409 4709 47443 4743
rect 2421 4573 2455 4607
rect 2697 4573 2731 4607
rect 3985 4573 4019 4607
rect 4261 4573 4295 4607
rect 4813 4573 4847 4607
rect 5549 4573 5583 4607
rect 6285 4573 6319 4607
rect 19257 4573 19291 4607
rect 21189 4573 21223 4607
rect 26801 4573 26835 4607
rect 26893 4573 26927 4607
rect 46857 4573 46891 4607
rect 47225 4573 47259 4607
rect 2605 4437 2639 4471
rect 4445 4437 4479 4471
rect 4997 4437 5031 4471
rect 5733 4437 5767 4471
rect 6469 4437 6503 4471
rect 19441 4437 19475 4471
rect 21373 4437 21407 4471
rect 26709 4437 26743 4471
rect 27077 4437 27111 4471
rect 47041 4437 47075 4471
rect 2237 4165 2271 4199
rect 18429 4165 18463 4199
rect 18705 4165 18739 4199
rect 7389 4097 7423 4131
rect 8493 4097 8527 4131
rect 8769 4097 8803 4131
rect 18889 4097 18923 4131
rect 40049 4097 40083 4131
rect 40233 4097 40267 4131
rect 42441 4097 42475 4131
rect 42717 4097 42751 4131
rect 46397 4097 46431 4131
rect 46489 4097 46523 4131
rect 46765 4097 46799 4131
rect 47133 4097 47167 4131
rect 2421 4029 2455 4063
rect 40417 3961 40451 3995
rect 47317 3961 47351 3995
rect 7573 3893 7607 3927
rect 8677 3893 8711 3927
rect 8953 3893 8987 3927
rect 42625 3893 42659 3927
rect 46305 3893 46339 3927
rect 46673 3893 46707 3927
rect 46949 3893 46983 3927
rect 46029 3689 46063 3723
rect 23949 3621 23983 3655
rect 29837 3621 29871 3655
rect 32965 3621 32999 3655
rect 46397 3621 46431 3655
rect 23765 3485 23799 3519
rect 24409 3485 24443 3519
rect 28549 3485 28583 3519
rect 28641 3485 28675 3519
rect 29193 3485 29227 3519
rect 29653 3485 29687 3519
rect 30113 3485 30147 3519
rect 30573 3485 30607 3519
rect 30665 3485 30699 3519
rect 31309 3485 31343 3519
rect 31861 3485 31895 3519
rect 32505 3485 32539 3519
rect 33057 3485 33091 3519
rect 33149 3485 33183 3519
rect 46121 3485 46155 3519
rect 46213 3485 46247 3519
rect 46489 3485 46523 3519
rect 46765 3485 46799 3519
rect 46949 3485 46983 3519
rect 24593 3349 24627 3383
rect 28457 3349 28491 3383
rect 28825 3349 28859 3383
rect 29377 3349 29411 3383
rect 30297 3349 30331 3383
rect 30481 3349 30515 3383
rect 30849 3349 30883 3383
rect 31493 3349 31527 3383
rect 32045 3349 32079 3383
rect 32689 3349 32723 3383
rect 33333 3349 33367 3383
rect 46673 3349 46707 3383
rect 47133 3349 47167 3383
rect 14105 3145 14139 3179
rect 17785 3145 17819 3179
rect 18153 3145 18187 3179
rect 47317 3145 47351 3179
rect 14197 3077 14231 3111
rect 14381 3077 14415 3111
rect 14565 3077 14599 3111
rect 17877 3009 17911 3043
rect 18061 3009 18095 3043
rect 19441 3009 19475 3043
rect 19625 3009 19659 3043
rect 21925 3009 21959 3043
rect 24777 3009 24811 3043
rect 25973 3009 26007 3043
rect 26065 3009 26099 3043
rect 28089 3009 28123 3043
rect 28181 3009 28215 3043
rect 29929 3009 29963 3043
rect 30665 3009 30699 3043
rect 31125 3009 31159 3043
rect 33701 3009 33735 3043
rect 36553 3009 36587 3043
rect 38853 3009 38887 3043
rect 46397 3009 46431 3043
rect 46765 3009 46799 3043
rect 47133 3009 47167 3043
rect 19349 2941 19383 2975
rect 25881 2941 25915 2975
rect 19809 2873 19843 2907
rect 26249 2873 26283 2907
rect 28365 2873 28399 2907
rect 46581 2873 46615 2907
rect 22109 2805 22143 2839
rect 24961 2805 24995 2839
rect 27997 2805 28031 2839
rect 30113 2805 30147 2839
rect 30849 2805 30883 2839
rect 31309 2805 31343 2839
rect 33885 2805 33919 2839
rect 36369 2805 36403 2839
rect 39037 2805 39071 2839
rect 46949 2805 46983 2839
rect 28641 2601 28675 2635
rect 29929 2601 29963 2635
rect 31217 2601 31251 2635
rect 33793 2601 33827 2635
rect 36369 2601 36403 2635
rect 38577 2601 38611 2635
rect 47317 2601 47351 2635
rect 27905 2533 27939 2567
rect 29653 2533 29687 2567
rect 31493 2533 31527 2567
rect 33425 2533 33459 2567
rect 35265 2533 35299 2567
rect 36645 2533 36679 2567
rect 37841 2533 37875 2567
rect 39313 2533 39347 2567
rect 40417 2533 40451 2567
rect 20637 2397 20671 2431
rect 21005 2397 21039 2431
rect 21373 2397 21407 2431
rect 22109 2397 22143 2431
rect 22477 2397 22511 2431
rect 22845 2397 22879 2431
rect 23213 2397 23247 2431
rect 23581 2397 23615 2431
rect 23949 2397 23983 2431
rect 24501 2397 24535 2431
rect 24869 2397 24903 2431
rect 25237 2397 25271 2431
rect 25605 2397 25639 2431
rect 25973 2397 26007 2431
rect 26341 2397 26375 2431
rect 26985 2397 27019 2431
rect 27353 2397 27387 2431
rect 27721 2397 27755 2431
rect 28089 2397 28123 2431
rect 28457 2397 28491 2431
rect 28825 2397 28859 2431
rect 29837 2397 29871 2431
rect 29929 2397 29963 2431
rect 30205 2397 30239 2431
rect 30297 2397 30331 2431
rect 30849 2397 30883 2431
rect 31033 2397 31067 2431
rect 31677 2397 31711 2431
rect 31769 2397 31803 2431
rect 32137 2397 32171 2431
rect 32505 2397 32539 2431
rect 32873 2397 32907 2431
rect 33241 2397 33275 2431
rect 33609 2397 33643 2431
rect 33977 2397 34011 2431
rect 34713 2397 34747 2431
rect 35081 2397 35115 2431
rect 35449 2397 35483 2431
rect 35817 2397 35851 2431
rect 36185 2397 36219 2431
rect 36829 2397 36863 2431
rect 37565 2397 37599 2431
rect 37682 2397 37716 2431
rect 38025 2397 38059 2431
rect 38393 2397 38427 2431
rect 38761 2397 38795 2431
rect 39129 2397 39163 2431
rect 39865 2397 39899 2431
rect 40233 2397 40267 2431
rect 45661 2397 45695 2431
rect 46029 2397 46063 2431
rect 46397 2397 46431 2431
rect 46765 2397 46799 2431
rect 47133 2397 47167 2431
rect 20821 2261 20855 2295
rect 21189 2261 21223 2295
rect 21557 2261 21591 2295
rect 22293 2261 22327 2295
rect 22661 2261 22695 2295
rect 23029 2261 23063 2295
rect 23397 2261 23431 2295
rect 23765 2261 23799 2295
rect 24133 2261 24167 2295
rect 24685 2261 24719 2295
rect 25053 2261 25087 2295
rect 25421 2261 25455 2295
rect 25789 2261 25823 2295
rect 26157 2261 26191 2295
rect 26525 2261 26559 2295
rect 27169 2261 27203 2295
rect 27537 2261 27571 2295
rect 28273 2261 28307 2295
rect 29009 2261 29043 2295
rect 30113 2261 30147 2295
rect 30481 2261 30515 2295
rect 31769 2261 31803 2295
rect 32321 2261 32355 2295
rect 32689 2261 32723 2295
rect 33057 2261 33091 2295
rect 34161 2261 34195 2295
rect 34897 2261 34931 2295
rect 35633 2261 35667 2295
rect 36001 2261 36035 2295
rect 37381 2261 37415 2295
rect 38209 2261 38243 2295
rect 38945 2261 38979 2295
rect 40049 2261 40083 2295
rect 45845 2261 45879 2295
rect 46213 2261 46247 2295
rect 46581 2261 46615 2295
rect 46949 2261 46983 2295
<< metal1 >>
rect 33870 9188 33876 9240
rect 33928 9228 33934 9240
rect 38562 9228 38568 9240
rect 33928 9200 38568 9228
rect 33928 9188 33934 9200
rect 38562 9188 38568 9200
rect 38620 9188 38626 9240
rect 19518 9120 19524 9172
rect 19576 9160 19582 9172
rect 46014 9160 46020 9172
rect 19576 9132 46020 9160
rect 19576 9120 19582 9132
rect 46014 9120 46020 9132
rect 46072 9120 46078 9172
rect 33962 9052 33968 9104
rect 34020 9092 34026 9104
rect 40402 9092 40408 9104
rect 34020 9064 40408 9092
rect 34020 9052 34026 9064
rect 40402 9052 40408 9064
rect 40460 9052 40466 9104
rect 37274 9024 37280 9036
rect 4080 8996 37280 9024
rect 4080 8832 4108 8996
rect 37274 8984 37280 8996
rect 37332 8984 37338 9036
rect 6638 8916 6644 8968
rect 6696 8956 6702 8968
rect 38746 8956 38752 8968
rect 6696 8928 38752 8956
rect 6696 8916 6702 8928
rect 38746 8916 38752 8928
rect 38804 8916 38810 8968
rect 23934 8848 23940 8900
rect 23992 8888 23998 8900
rect 46382 8888 46388 8900
rect 23992 8860 46388 8888
rect 23992 8848 23998 8860
rect 46382 8848 46388 8860
rect 46440 8848 46446 8900
rect 4062 8780 4068 8832
rect 4120 8780 4126 8832
rect 26510 8780 26516 8832
rect 26568 8820 26574 8832
rect 41230 8820 41236 8832
rect 26568 8792 41236 8820
rect 26568 8780 26574 8792
rect 41230 8780 41236 8792
rect 41288 8780 41294 8832
rect 1104 8730 47840 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 39010 8730
rect 39062 8678 39074 8730
rect 39126 8678 39138 8730
rect 39190 8678 39202 8730
rect 39254 8678 39266 8730
rect 39318 8678 45010 8730
rect 45062 8678 45074 8730
rect 45126 8678 45138 8730
rect 45190 8678 45202 8730
rect 45254 8678 45266 8730
rect 45318 8678 47840 8730
rect 1104 8656 47840 8678
rect 1394 8576 1400 8628
rect 1452 8616 1458 8628
rect 1489 8619 1547 8625
rect 1489 8616 1501 8619
rect 1452 8588 1501 8616
rect 1452 8576 1458 8588
rect 1489 8585 1501 8588
rect 1535 8585 1547 8619
rect 1489 8579 1547 8585
rect 3694 8576 3700 8628
rect 3752 8616 3758 8628
rect 3881 8619 3939 8625
rect 3881 8616 3893 8619
rect 3752 8588 3893 8616
rect 3752 8576 3758 8588
rect 3881 8585 3893 8588
rect 3927 8585 3939 8619
rect 3881 8579 3939 8585
rect 4062 8576 4068 8628
rect 4120 8576 4126 8628
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 6457 8619 6515 8625
rect 6457 8616 6469 8619
rect 6052 8588 6469 8616
rect 6052 8576 6058 8588
rect 6457 8585 6469 8588
rect 6503 8585 6515 8619
rect 6457 8579 6515 8585
rect 8294 8576 8300 8628
rect 8352 8616 8358 8628
rect 8573 8619 8631 8625
rect 8573 8616 8585 8619
rect 8352 8588 8585 8616
rect 8352 8576 8358 8588
rect 8573 8585 8585 8588
rect 8619 8585 8631 8619
rect 8573 8579 8631 8585
rect 10594 8576 10600 8628
rect 10652 8616 10658 8628
rect 10873 8619 10931 8625
rect 10873 8616 10885 8619
rect 10652 8588 10885 8616
rect 10652 8576 10658 8588
rect 10873 8585 10885 8588
rect 10919 8585 10931 8619
rect 10873 8579 10931 8585
rect 12894 8576 12900 8628
rect 12952 8616 12958 8628
rect 13173 8619 13231 8625
rect 13173 8616 13185 8619
rect 12952 8588 13185 8616
rect 12952 8576 12958 8588
rect 13173 8585 13185 8588
rect 13219 8585 13231 8619
rect 13173 8579 13231 8585
rect 15378 8576 15384 8628
rect 15436 8616 15442 8628
rect 15473 8619 15531 8625
rect 15473 8616 15485 8619
rect 15436 8588 15485 8616
rect 15436 8576 15442 8588
rect 15473 8585 15485 8588
rect 15519 8585 15531 8619
rect 15473 8579 15531 8585
rect 17494 8576 17500 8628
rect 17552 8616 17558 8628
rect 17681 8619 17739 8625
rect 17681 8616 17693 8619
rect 17552 8588 17693 8616
rect 17552 8576 17558 8588
rect 17681 8585 17693 8588
rect 17727 8585 17739 8619
rect 17681 8579 17739 8585
rect 19794 8576 19800 8628
rect 19852 8616 19858 8628
rect 19981 8619 20039 8625
rect 19981 8616 19993 8619
rect 19852 8588 19993 8616
rect 19852 8576 19858 8588
rect 19981 8585 19993 8588
rect 20027 8585 20039 8619
rect 19981 8579 20039 8585
rect 22094 8576 22100 8628
rect 22152 8616 22158 8628
rect 22281 8619 22339 8625
rect 22281 8616 22293 8619
rect 22152 8588 22293 8616
rect 22152 8576 22158 8588
rect 22281 8585 22293 8588
rect 22327 8585 22339 8619
rect 22281 8579 22339 8585
rect 24394 8576 24400 8628
rect 24452 8616 24458 8628
rect 24581 8619 24639 8625
rect 24581 8616 24593 8619
rect 24452 8588 24593 8616
rect 24452 8576 24458 8588
rect 24581 8585 24593 8588
rect 24627 8585 24639 8619
rect 24581 8579 24639 8585
rect 26694 8576 26700 8628
rect 26752 8616 26758 8628
rect 27065 8619 27123 8625
rect 27065 8616 27077 8619
rect 26752 8588 27077 8616
rect 26752 8576 26758 8588
rect 27065 8585 27077 8588
rect 27111 8585 27123 8619
rect 27065 8579 27123 8585
rect 28994 8576 29000 8628
rect 29052 8616 29058 8628
rect 29181 8619 29239 8625
rect 29181 8616 29193 8619
rect 29052 8588 29193 8616
rect 29052 8576 29058 8588
rect 29181 8585 29193 8588
rect 29227 8585 29239 8619
rect 29181 8579 29239 8585
rect 31294 8576 31300 8628
rect 31352 8616 31358 8628
rect 31481 8619 31539 8625
rect 31481 8616 31493 8619
rect 31352 8588 31493 8616
rect 31352 8576 31358 8588
rect 31481 8585 31493 8588
rect 31527 8585 31539 8619
rect 31481 8579 31539 8585
rect 33594 8576 33600 8628
rect 33652 8616 33658 8628
rect 33781 8619 33839 8625
rect 33781 8616 33793 8619
rect 33652 8588 33793 8616
rect 33652 8576 33658 8588
rect 33781 8585 33793 8588
rect 33827 8585 33839 8619
rect 33781 8579 33839 8585
rect 34054 8576 34060 8628
rect 34112 8576 34118 8628
rect 35894 8576 35900 8628
rect 35952 8616 35958 8628
rect 36081 8619 36139 8625
rect 36081 8616 36093 8619
rect 35952 8588 36093 8616
rect 35952 8576 35958 8588
rect 36081 8585 36093 8588
rect 36127 8585 36139 8619
rect 36081 8579 36139 8585
rect 38194 8576 38200 8628
rect 38252 8616 38258 8628
rect 38381 8619 38439 8625
rect 38381 8616 38393 8619
rect 38252 8588 38393 8616
rect 38252 8576 38258 8588
rect 38381 8585 38393 8588
rect 38427 8585 38439 8619
rect 38381 8579 38439 8585
rect 40494 8576 40500 8628
rect 40552 8616 40558 8628
rect 40681 8619 40739 8625
rect 40681 8616 40693 8619
rect 40552 8588 40693 8616
rect 40552 8576 40558 8588
rect 40681 8585 40693 8588
rect 40727 8585 40739 8619
rect 40681 8579 40739 8585
rect 42794 8576 42800 8628
rect 42852 8616 42858 8628
rect 42981 8619 43039 8625
rect 42981 8616 42993 8619
rect 42852 8588 42993 8616
rect 42852 8576 42858 8588
rect 42981 8585 42993 8588
rect 43027 8585 43039 8619
rect 42981 8579 43039 8585
rect 45281 8619 45339 8625
rect 45281 8585 45293 8619
rect 45327 8616 45339 8619
rect 45370 8616 45376 8628
rect 45327 8588 45376 8616
rect 45327 8585 45339 8588
rect 45281 8579 45339 8585
rect 45370 8576 45376 8588
rect 45428 8576 45434 8628
rect 45830 8576 45836 8628
rect 45888 8576 45894 8628
rect 46198 8576 46204 8628
rect 46256 8576 46262 8628
rect 46937 8619 46995 8625
rect 46937 8585 46949 8619
rect 46983 8616 46995 8619
rect 47394 8616 47400 8628
rect 46983 8588 47400 8616
rect 46983 8585 46995 8588
rect 46937 8579 46995 8585
rect 47394 8576 47400 8588
rect 47452 8576 47458 8628
rect 4080 8489 4108 8576
rect 22186 8508 22192 8560
rect 22244 8548 22250 8560
rect 34072 8548 34100 8576
rect 22244 8520 34100 8548
rect 22244 8508 22250 8520
rect 34238 8508 34244 8560
rect 34296 8548 34302 8560
rect 34296 8520 45692 8548
rect 34296 8508 34302 8520
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8449 1731 8483
rect 1673 8443 1731 8449
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 1688 8412 1716 8443
rect 6638 8440 6644 8492
rect 6696 8440 6702 8492
rect 8386 8440 8392 8492
rect 8444 8440 8450 8492
rect 10686 8440 10692 8492
rect 10744 8440 10750 8492
rect 12986 8440 12992 8492
rect 13044 8440 13050 8492
rect 15289 8483 15347 8489
rect 15289 8449 15301 8483
rect 15335 8480 15347 8483
rect 15378 8480 15384 8492
rect 15335 8452 15384 8480
rect 15335 8449 15347 8452
rect 15289 8443 15347 8449
rect 15378 8440 15384 8452
rect 15436 8440 15442 8492
rect 17862 8440 17868 8492
rect 17920 8440 17926 8492
rect 20165 8483 20223 8489
rect 20165 8449 20177 8483
rect 20211 8480 20223 8483
rect 20622 8480 20628 8492
rect 20211 8452 20628 8480
rect 20211 8449 20223 8452
rect 20165 8443 20223 8449
rect 20622 8440 20628 8452
rect 20680 8440 20686 8492
rect 22465 8483 22523 8489
rect 22465 8449 22477 8483
rect 22511 8480 22523 8483
rect 23474 8480 23480 8492
rect 22511 8452 23480 8480
rect 22511 8449 22523 8452
rect 22465 8443 22523 8449
rect 23474 8440 23480 8452
rect 23532 8440 23538 8492
rect 24765 8483 24823 8489
rect 24765 8449 24777 8483
rect 24811 8480 24823 8483
rect 25866 8480 25872 8492
rect 24811 8452 25872 8480
rect 24811 8449 24823 8452
rect 24765 8443 24823 8449
rect 25866 8440 25872 8452
rect 25924 8440 25930 8492
rect 27249 8483 27307 8489
rect 27249 8449 27261 8483
rect 27295 8480 27307 8483
rect 29270 8480 29276 8492
rect 27295 8452 29276 8480
rect 27295 8449 27307 8452
rect 27249 8443 27307 8449
rect 29270 8440 29276 8452
rect 29328 8440 29334 8492
rect 29362 8440 29368 8492
rect 29420 8440 29426 8492
rect 31665 8483 31723 8489
rect 31665 8449 31677 8483
rect 31711 8480 31723 8483
rect 33870 8480 33876 8492
rect 31711 8452 33876 8480
rect 31711 8449 31723 8452
rect 31665 8443 31723 8449
rect 33870 8440 33876 8452
rect 33928 8440 33934 8492
rect 33962 8440 33968 8492
rect 34020 8440 34026 8492
rect 36277 8483 36335 8489
rect 36277 8449 36289 8483
rect 36323 8480 36335 8483
rect 37182 8480 37188 8492
rect 36323 8452 37188 8480
rect 36323 8449 36335 8452
rect 36277 8443 36335 8449
rect 37182 8440 37188 8452
rect 37240 8440 37246 8492
rect 38565 8483 38623 8489
rect 38565 8449 38577 8483
rect 38611 8480 38623 8483
rect 39574 8480 39580 8492
rect 38611 8452 39580 8480
rect 38611 8449 38623 8452
rect 38565 8443 38623 8449
rect 39574 8440 39580 8452
rect 39632 8440 39638 8492
rect 40862 8440 40868 8492
rect 40920 8440 40926 8492
rect 43162 8440 43168 8492
rect 43220 8440 43226 8492
rect 45462 8440 45468 8492
rect 45520 8440 45526 8492
rect 45664 8489 45692 8520
rect 45649 8483 45707 8489
rect 45649 8449 45661 8483
rect 45695 8449 45707 8483
rect 45649 8443 45707 8449
rect 46014 8440 46020 8492
rect 46072 8440 46078 8492
rect 46382 8440 46388 8492
rect 46440 8440 46446 8492
rect 46750 8440 46756 8492
rect 46808 8440 46814 8492
rect 47121 8483 47179 8489
rect 47121 8449 47133 8483
rect 47167 8449 47179 8483
rect 47121 8443 47179 8449
rect 37826 8412 37832 8424
rect 1688 8384 22094 8412
rect 22066 8344 22094 8384
rect 29380 8384 37832 8412
rect 29380 8344 29408 8384
rect 37826 8372 37832 8384
rect 37884 8372 37890 8424
rect 41230 8372 41236 8424
rect 41288 8412 41294 8424
rect 47136 8412 47164 8443
rect 41288 8384 47164 8412
rect 41288 8372 41294 8384
rect 39942 8344 39948 8356
rect 22066 8316 29408 8344
rect 38626 8316 39948 8344
rect 29270 8236 29276 8288
rect 29328 8276 29334 8288
rect 38626 8276 38654 8316
rect 39942 8304 39948 8316
rect 40000 8304 40006 8356
rect 46569 8347 46627 8353
rect 46569 8313 46581 8347
rect 46615 8344 46627 8347
rect 47210 8344 47216 8356
rect 46615 8316 47216 8344
rect 46615 8313 46627 8316
rect 46569 8307 46627 8313
rect 47210 8304 47216 8316
rect 47268 8304 47274 8356
rect 47302 8304 47308 8356
rect 47360 8304 47366 8356
rect 29328 8248 38654 8276
rect 29328 8236 29334 8248
rect 1104 8186 47840 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 37950 8186
rect 38002 8134 38014 8186
rect 38066 8134 38078 8186
rect 38130 8134 38142 8186
rect 38194 8134 38206 8186
rect 38258 8134 43950 8186
rect 44002 8134 44014 8186
rect 44066 8134 44078 8186
rect 44130 8134 44142 8186
rect 44194 8134 44206 8186
rect 44258 8134 47840 8186
rect 1104 8112 47840 8134
rect 8297 8075 8355 8081
rect 8297 8041 8309 8075
rect 8343 8072 8355 8075
rect 8386 8072 8392 8084
rect 8343 8044 8392 8072
rect 8343 8041 8355 8044
rect 8297 8035 8355 8041
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 10229 8075 10287 8081
rect 10229 8041 10241 8075
rect 10275 8072 10287 8075
rect 10686 8072 10692 8084
rect 10275 8044 10692 8072
rect 10275 8041 10287 8044
rect 10229 8035 10287 8041
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 19518 8032 19524 8084
rect 19576 8032 19582 8084
rect 20530 8032 20536 8084
rect 20588 8032 20594 8084
rect 20622 8032 20628 8084
rect 20680 8032 20686 8084
rect 21726 8032 21732 8084
rect 21784 8032 21790 8084
rect 22097 8075 22155 8081
rect 22097 8041 22109 8075
rect 22143 8072 22155 8075
rect 22186 8072 22192 8084
rect 22143 8044 22192 8072
rect 22143 8041 22155 8044
rect 22097 8035 22155 8041
rect 22186 8032 22192 8044
rect 22244 8032 22250 8084
rect 23474 8032 23480 8084
rect 23532 8032 23538 8084
rect 23934 8032 23940 8084
rect 23992 8032 23998 8084
rect 25866 8032 25872 8084
rect 25924 8072 25930 8084
rect 26053 8075 26111 8081
rect 26053 8072 26065 8075
rect 25924 8044 26065 8072
rect 25924 8032 25930 8044
rect 26053 8041 26065 8044
rect 26099 8041 26111 8075
rect 26053 8035 26111 8041
rect 26510 8032 26516 8084
rect 26568 8032 26574 8084
rect 29362 8032 29368 8084
rect 29420 8072 29426 8084
rect 29825 8075 29883 8081
rect 29825 8072 29837 8075
rect 29420 8044 29837 8072
rect 29420 8032 29426 8044
rect 29825 8041 29837 8044
rect 29871 8041 29883 8075
rect 29825 8035 29883 8041
rect 37826 8032 37832 8084
rect 37884 8032 37890 8084
rect 43806 8032 43812 8084
rect 43864 8072 43870 8084
rect 43864 8044 46612 8072
rect 43864 8032 43870 8044
rect 7558 7964 7564 8016
rect 7616 8004 7622 8016
rect 11606 8004 11612 8016
rect 7616 7976 11612 8004
rect 7616 7964 7622 7976
rect 11606 7964 11612 7976
rect 11664 7964 11670 8016
rect 11790 7964 11796 8016
rect 11848 8004 11854 8016
rect 46584 8004 46612 8044
rect 46658 8032 46664 8084
rect 46716 8032 46722 8084
rect 11848 7976 46520 8004
rect 46584 7976 46888 8004
rect 11848 7964 11854 7976
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7936 2283 7939
rect 2271 7908 41414 7936
rect 2271 7905 2283 7908
rect 2225 7899 2283 7905
rect 1026 7828 1032 7880
rect 1084 7868 1090 7880
rect 2041 7871 2099 7877
rect 2041 7868 2053 7871
rect 1084 7840 2053 7868
rect 1084 7828 1090 7840
rect 2041 7837 2053 7840
rect 2087 7837 2099 7871
rect 2041 7831 2099 7837
rect 8021 7871 8079 7877
rect 8021 7837 8033 7871
rect 8067 7868 8079 7871
rect 8113 7871 8171 7877
rect 8113 7868 8125 7871
rect 8067 7840 8125 7868
rect 8067 7837 8079 7840
rect 8021 7831 8079 7837
rect 8113 7837 8125 7840
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 10042 7828 10048 7880
rect 10100 7828 10106 7880
rect 10134 7828 10140 7880
rect 10192 7868 10198 7880
rect 11977 7871 12035 7877
rect 11977 7868 11989 7871
rect 10192 7840 11989 7868
rect 10192 7828 10198 7840
rect 11977 7837 11989 7840
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 14182 7828 14188 7880
rect 14240 7868 14246 7880
rect 15933 7871 15991 7877
rect 15933 7868 15945 7871
rect 14240 7840 15945 7868
rect 14240 7828 14246 7840
rect 15933 7837 15945 7840
rect 15979 7837 15991 7871
rect 15933 7831 15991 7837
rect 19334 7828 19340 7880
rect 19392 7868 19398 7880
rect 19613 7871 19671 7877
rect 19613 7868 19625 7871
rect 19392 7840 19625 7868
rect 19392 7828 19398 7840
rect 19613 7837 19625 7840
rect 19659 7837 19671 7871
rect 19613 7831 19671 7837
rect 20346 7828 20352 7880
rect 20404 7828 20410 7880
rect 20806 7828 20812 7880
rect 20864 7828 20870 7880
rect 20901 7871 20959 7877
rect 20901 7837 20913 7871
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 21821 7871 21879 7877
rect 21821 7837 21833 7871
rect 21867 7868 21879 7871
rect 21913 7871 21971 7877
rect 21913 7868 21925 7871
rect 21867 7840 21925 7868
rect 21867 7837 21879 7840
rect 21821 7831 21879 7837
rect 21913 7837 21925 7840
rect 21959 7837 21971 7871
rect 21913 7831 21971 7837
rect 23293 7871 23351 7877
rect 23293 7837 23305 7871
rect 23339 7868 23351 7871
rect 23661 7871 23719 7877
rect 23661 7868 23673 7871
rect 23339 7840 23673 7868
rect 23339 7837 23351 7840
rect 23293 7831 23351 7837
rect 23661 7837 23673 7840
rect 23707 7837 23719 7871
rect 23661 7831 23719 7837
rect 3786 7760 3792 7812
rect 3844 7800 3850 7812
rect 20916 7800 20944 7831
rect 23382 7800 23388 7812
rect 3844 7772 20944 7800
rect 21100 7772 23388 7800
rect 3844 7760 3850 7772
rect 8021 7735 8079 7741
rect 8021 7701 8033 7735
rect 8067 7732 8079 7735
rect 11882 7732 11888 7744
rect 8067 7704 11888 7732
rect 8067 7701 8079 7704
rect 8021 7695 8079 7701
rect 11882 7692 11888 7704
rect 11940 7692 11946 7744
rect 12161 7735 12219 7741
rect 12161 7701 12173 7735
rect 12207 7732 12219 7735
rect 16022 7732 16028 7744
rect 12207 7704 16028 7732
rect 12207 7701 12219 7704
rect 12161 7695 12219 7701
rect 16022 7692 16028 7704
rect 16080 7692 16086 7744
rect 16117 7735 16175 7741
rect 16117 7701 16129 7735
rect 16163 7732 16175 7735
rect 20714 7732 20720 7744
rect 16163 7704 20720 7732
rect 16163 7701 16175 7704
rect 16117 7695 16175 7701
rect 20714 7692 20720 7704
rect 20772 7692 20778 7744
rect 21100 7741 21128 7772
rect 23382 7760 23388 7772
rect 23440 7760 23446 7812
rect 23676 7800 23704 7831
rect 23750 7828 23756 7880
rect 23808 7868 23814 7880
rect 24029 7871 24087 7877
rect 24029 7868 24041 7871
rect 23808 7840 24041 7868
rect 23808 7828 23814 7840
rect 24029 7837 24041 7840
rect 24075 7837 24087 7871
rect 24029 7831 24087 7837
rect 25590 7828 25596 7880
rect 25648 7828 25654 7880
rect 25961 7871 26019 7877
rect 25961 7837 25973 7871
rect 26007 7868 26019 7871
rect 26007 7864 26188 7868
rect 26234 7864 26240 7880
rect 26007 7840 26240 7864
rect 26007 7837 26019 7840
rect 25961 7831 26019 7837
rect 26160 7836 26240 7840
rect 26234 7828 26240 7836
rect 26292 7828 26298 7880
rect 26326 7828 26332 7880
rect 26384 7828 26390 7880
rect 26510 7828 26516 7880
rect 26568 7868 26574 7880
rect 29549 7871 29607 7877
rect 29549 7868 29561 7871
rect 26568 7840 29561 7868
rect 26568 7828 26574 7840
rect 29549 7837 29561 7840
rect 29595 7837 29607 7871
rect 29549 7831 29607 7837
rect 29914 7828 29920 7880
rect 29972 7868 29978 7880
rect 30009 7871 30067 7877
rect 30009 7868 30021 7871
rect 29972 7840 30021 7868
rect 29972 7828 29978 7840
rect 30009 7837 30021 7840
rect 30055 7837 30067 7871
rect 30009 7831 30067 7837
rect 35253 7871 35311 7877
rect 35253 7837 35265 7871
rect 35299 7868 35311 7871
rect 35345 7871 35403 7877
rect 35345 7868 35357 7871
rect 35299 7840 35357 7868
rect 35299 7837 35311 7840
rect 35253 7831 35311 7837
rect 35345 7837 35357 7840
rect 35391 7837 35403 7871
rect 35345 7831 35403 7837
rect 38013 7871 38071 7877
rect 38013 7837 38025 7871
rect 38059 7837 38071 7871
rect 38013 7831 38071 7837
rect 39577 7871 39635 7877
rect 39577 7837 39589 7871
rect 39623 7868 39635 7871
rect 39666 7868 39672 7880
rect 39623 7840 39672 7868
rect 39623 7837 39635 7840
rect 39577 7831 39635 7837
rect 24946 7800 24952 7812
rect 23676 7772 24952 7800
rect 24946 7760 24952 7772
rect 25004 7760 25010 7812
rect 36538 7800 36544 7812
rect 26528 7772 36544 7800
rect 21085 7735 21143 7741
rect 21085 7701 21097 7735
rect 21131 7701 21143 7735
rect 21085 7695 21143 7701
rect 24670 7692 24676 7744
rect 24728 7732 24734 7744
rect 26528 7732 26556 7772
rect 36538 7760 36544 7772
rect 36596 7760 36602 7812
rect 38028 7800 38056 7831
rect 39666 7828 39672 7840
rect 39724 7828 39730 7880
rect 40313 7871 40371 7877
rect 40313 7837 40325 7871
rect 40359 7868 40371 7871
rect 40589 7871 40647 7877
rect 40589 7868 40601 7871
rect 40359 7840 40601 7868
rect 40359 7837 40371 7840
rect 40313 7831 40371 7837
rect 40589 7837 40601 7840
rect 40635 7837 40647 7871
rect 40589 7831 40647 7837
rect 39850 7800 39856 7812
rect 38028 7772 39856 7800
rect 39850 7760 39856 7772
rect 39908 7760 39914 7812
rect 41386 7800 41414 7908
rect 45373 7871 45431 7877
rect 45373 7837 45385 7871
rect 45419 7868 45431 7871
rect 45649 7871 45707 7877
rect 45649 7868 45661 7871
rect 45419 7840 45661 7868
rect 45419 7837 45431 7840
rect 45373 7831 45431 7837
rect 45649 7837 45661 7840
rect 45695 7837 45707 7871
rect 45649 7831 45707 7837
rect 46014 7828 46020 7880
rect 46072 7828 46078 7880
rect 46106 7828 46112 7880
rect 46164 7828 46170 7880
rect 46492 7877 46520 7976
rect 46860 7877 46888 7976
rect 46477 7871 46535 7877
rect 46477 7837 46489 7871
rect 46523 7837 46535 7871
rect 46477 7831 46535 7837
rect 46845 7871 46903 7877
rect 46845 7837 46857 7871
rect 46891 7837 46903 7871
rect 46845 7831 46903 7837
rect 47210 7828 47216 7880
rect 47268 7828 47274 7880
rect 46566 7800 46572 7812
rect 41386 7772 46572 7800
rect 46566 7760 46572 7772
rect 46624 7760 46630 7812
rect 24728 7704 26556 7732
rect 24728 7692 24734 7704
rect 29730 7692 29736 7744
rect 29788 7692 29794 7744
rect 30466 7692 30472 7744
rect 30524 7732 30530 7744
rect 35161 7735 35219 7741
rect 35161 7732 35173 7735
rect 30524 7704 35173 7732
rect 30524 7692 30530 7704
rect 35161 7701 35173 7704
rect 35207 7701 35219 7735
rect 35161 7695 35219 7701
rect 35529 7735 35587 7741
rect 35529 7701 35541 7735
rect 35575 7732 35587 7735
rect 36170 7732 36176 7744
rect 35575 7704 36176 7732
rect 35575 7701 35587 7704
rect 35529 7695 35587 7701
rect 36170 7692 36176 7704
rect 36228 7692 36234 7744
rect 36814 7692 36820 7744
rect 36872 7732 36878 7744
rect 39393 7735 39451 7741
rect 39393 7732 39405 7735
rect 36872 7704 39405 7732
rect 36872 7692 36878 7704
rect 39393 7701 39405 7704
rect 39439 7701 39451 7735
rect 39393 7695 39451 7701
rect 40126 7692 40132 7744
rect 40184 7732 40190 7744
rect 40221 7735 40279 7741
rect 40221 7732 40233 7735
rect 40184 7704 40233 7732
rect 40184 7692 40190 7704
rect 40221 7701 40233 7704
rect 40267 7701 40279 7735
rect 40221 7695 40279 7701
rect 40310 7692 40316 7744
rect 40368 7732 40374 7744
rect 40405 7735 40463 7741
rect 40405 7732 40417 7735
rect 40368 7704 40417 7732
rect 40368 7692 40374 7704
rect 40405 7701 40417 7704
rect 40451 7701 40463 7735
rect 40405 7695 40463 7701
rect 44818 7692 44824 7744
rect 44876 7732 44882 7744
rect 45281 7735 45339 7741
rect 45281 7732 45293 7735
rect 44876 7704 45293 7732
rect 44876 7692 44882 7704
rect 45281 7701 45293 7704
rect 45327 7701 45339 7735
rect 45281 7695 45339 7701
rect 45370 7692 45376 7744
rect 45428 7732 45434 7744
rect 45465 7735 45523 7741
rect 45465 7732 45477 7735
rect 45428 7704 45477 7732
rect 45428 7692 45434 7704
rect 45465 7701 45477 7704
rect 45511 7701 45523 7735
rect 45465 7695 45523 7701
rect 45833 7735 45891 7741
rect 45833 7701 45845 7735
rect 45879 7732 45891 7735
rect 45922 7732 45928 7744
rect 45879 7704 45928 7732
rect 45879 7701 45891 7704
rect 45833 7695 45891 7701
rect 45922 7692 45928 7704
rect 45980 7692 45986 7744
rect 46290 7692 46296 7744
rect 46348 7692 46354 7744
rect 47026 7692 47032 7744
rect 47084 7692 47090 7744
rect 47394 7692 47400 7744
rect 47452 7692 47458 7744
rect 1104 7642 47840 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 39010 7642
rect 39062 7590 39074 7642
rect 39126 7590 39138 7642
rect 39190 7590 39202 7642
rect 39254 7590 39266 7642
rect 39318 7590 45010 7642
rect 45062 7590 45074 7642
rect 45126 7590 45138 7642
rect 45190 7590 45202 7642
rect 45254 7590 45266 7642
rect 45318 7590 47840 7642
rect 1104 7568 47840 7590
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 12253 7531 12311 7537
rect 4212 7500 11744 7528
rect 4212 7488 4218 7500
rect 1578 7420 1584 7472
rect 1636 7460 1642 7472
rect 1636 7432 10824 7460
rect 1636 7420 1642 7432
rect 10042 7352 10048 7404
rect 10100 7392 10106 7404
rect 10100 7364 10732 7392
rect 10100 7352 10106 7364
rect 1854 7284 1860 7336
rect 1912 7324 1918 7336
rect 10134 7324 10140 7336
rect 1912 7296 10140 7324
rect 1912 7284 1918 7296
rect 10134 7284 10140 7296
rect 10192 7284 10198 7336
rect 10704 7256 10732 7364
rect 10796 7324 10824 7432
rect 11606 7420 11612 7472
rect 11664 7420 11670 7472
rect 11716 7460 11744 7500
rect 12253 7497 12265 7531
rect 12299 7528 12311 7531
rect 12986 7528 12992 7540
rect 12299 7500 12992 7528
rect 12299 7497 12311 7500
rect 12253 7491 12311 7497
rect 12986 7488 12992 7500
rect 13044 7488 13050 7540
rect 15013 7531 15071 7537
rect 15013 7497 15025 7531
rect 15059 7528 15071 7531
rect 15378 7528 15384 7540
rect 15059 7500 15384 7528
rect 15059 7497 15071 7500
rect 15013 7491 15071 7497
rect 15378 7488 15384 7500
rect 15436 7488 15442 7540
rect 17862 7488 17868 7540
rect 17920 7488 17926 7540
rect 20530 7488 20536 7540
rect 20588 7528 20594 7540
rect 23566 7528 23572 7540
rect 20588 7500 23572 7528
rect 20588 7488 20594 7500
rect 23566 7488 23572 7500
rect 23624 7488 23630 7540
rect 29730 7488 29736 7540
rect 29788 7528 29794 7540
rect 36446 7528 36452 7540
rect 29788 7500 36452 7528
rect 29788 7488 29794 7500
rect 36446 7488 36452 7500
rect 36504 7488 36510 7540
rect 37274 7488 37280 7540
rect 37332 7528 37338 7540
rect 38105 7531 38163 7537
rect 38105 7528 38117 7531
rect 37332 7500 38117 7528
rect 37332 7488 37338 7500
rect 38105 7497 38117 7500
rect 38151 7497 38163 7531
rect 38105 7491 38163 7497
rect 38746 7488 38752 7540
rect 38804 7488 38810 7540
rect 39574 7488 39580 7540
rect 39632 7488 39638 7540
rect 40773 7531 40831 7537
rect 40773 7497 40785 7531
rect 40819 7528 40831 7531
rect 40862 7528 40868 7540
rect 40819 7500 40868 7528
rect 40819 7497 40831 7500
rect 40773 7491 40831 7497
rect 40862 7488 40868 7500
rect 40920 7488 40926 7540
rect 43438 7488 43444 7540
rect 43496 7528 43502 7540
rect 45370 7528 45376 7540
rect 43496 7500 45376 7528
rect 43496 7488 43502 7500
rect 45370 7488 45376 7500
rect 45428 7488 45434 7540
rect 46661 7531 46719 7537
rect 46661 7497 46673 7531
rect 46707 7528 46719 7531
rect 46750 7528 46756 7540
rect 46707 7500 46756 7528
rect 46707 7497 46719 7500
rect 46661 7491 46719 7497
rect 46750 7488 46756 7500
rect 46808 7488 46814 7540
rect 46934 7488 46940 7540
rect 46992 7488 46998 7540
rect 20346 7460 20352 7472
rect 11716 7432 20352 7460
rect 20346 7420 20352 7432
rect 20404 7420 20410 7472
rect 20806 7420 20812 7472
rect 20864 7460 20870 7472
rect 31202 7460 31208 7472
rect 20864 7432 31208 7460
rect 20864 7420 20870 7432
rect 31202 7420 31208 7432
rect 31260 7420 31266 7472
rect 36538 7420 36544 7472
rect 36596 7460 36602 7472
rect 36596 7432 47164 7460
rect 36596 7420 36602 7432
rect 11790 7352 11796 7404
rect 11848 7352 11854 7404
rect 11977 7395 12035 7401
rect 11977 7361 11989 7395
rect 12023 7392 12035 7395
rect 12069 7395 12127 7401
rect 12069 7392 12081 7395
rect 12023 7364 12081 7392
rect 12023 7361 12035 7364
rect 11977 7355 12035 7361
rect 12069 7361 12081 7364
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 14829 7395 14887 7401
rect 14829 7361 14841 7395
rect 14875 7361 14887 7395
rect 14829 7355 14887 7361
rect 14182 7324 14188 7336
rect 10796 7296 14188 7324
rect 14182 7284 14188 7296
rect 14240 7284 14246 7336
rect 14844 7324 14872 7355
rect 18046 7352 18052 7404
rect 18104 7352 18110 7404
rect 23017 7395 23075 7401
rect 23017 7361 23029 7395
rect 23063 7392 23075 7395
rect 23109 7395 23167 7401
rect 23109 7392 23121 7395
rect 23063 7364 23121 7392
rect 23063 7361 23075 7364
rect 23017 7355 23075 7361
rect 23109 7361 23121 7364
rect 23155 7361 23167 7395
rect 23109 7355 23167 7361
rect 33137 7395 33195 7401
rect 33137 7361 33149 7395
rect 33183 7392 33195 7395
rect 33229 7395 33287 7401
rect 33229 7392 33241 7395
rect 33183 7364 33241 7392
rect 33183 7361 33195 7364
rect 33137 7355 33195 7361
rect 33229 7361 33241 7364
rect 33275 7361 33287 7395
rect 33229 7355 33287 7361
rect 38197 7395 38255 7401
rect 38197 7361 38209 7395
rect 38243 7361 38255 7395
rect 38197 7355 38255 7361
rect 38841 7395 38899 7401
rect 38841 7361 38853 7395
rect 38887 7361 38899 7395
rect 38841 7355 38899 7361
rect 39761 7395 39819 7401
rect 39761 7361 39773 7395
rect 39807 7361 39819 7395
rect 39761 7355 39819 7361
rect 40957 7395 41015 7401
rect 40957 7361 40969 7395
rect 41003 7392 41015 7395
rect 45922 7392 45928 7404
rect 41003 7364 45928 7392
rect 41003 7361 41015 7364
rect 40957 7355 41015 7361
rect 33778 7324 33784 7336
rect 14844 7296 33784 7324
rect 33778 7284 33784 7296
rect 33836 7284 33842 7336
rect 38212 7256 38240 7355
rect 38856 7256 38884 7355
rect 38930 7284 38936 7336
rect 38988 7324 38994 7336
rect 39574 7324 39580 7336
rect 38988 7296 39580 7324
rect 38988 7284 38994 7296
rect 39574 7284 39580 7296
rect 39632 7284 39638 7336
rect 39776 7324 39804 7355
rect 45922 7352 45928 7364
rect 45980 7352 45986 7404
rect 46477 7395 46535 7401
rect 46477 7361 46489 7395
rect 46523 7361 46535 7395
rect 46477 7355 46535 7361
rect 45738 7324 45744 7336
rect 39776 7296 45744 7324
rect 45738 7284 45744 7296
rect 45796 7284 45802 7336
rect 46492 7324 46520 7355
rect 46566 7352 46572 7404
rect 46624 7392 46630 7404
rect 47136 7401 47164 7432
rect 46753 7395 46811 7401
rect 46753 7392 46765 7395
rect 46624 7364 46765 7392
rect 46624 7352 46630 7364
rect 46753 7361 46765 7364
rect 46799 7361 46811 7395
rect 46753 7355 46811 7361
rect 47121 7395 47179 7401
rect 47121 7361 47133 7395
rect 47167 7361 47179 7395
rect 47121 7355 47179 7361
rect 47486 7324 47492 7336
rect 46492 7296 47492 7324
rect 47486 7284 47492 7296
rect 47544 7284 47550 7336
rect 40586 7256 40592 7268
rect 10704 7228 37504 7256
rect 38212 7228 38792 7256
rect 38856 7228 40592 7256
rect 11974 7148 11980 7200
rect 12032 7148 12038 7200
rect 22922 7148 22928 7200
rect 22980 7148 22986 7200
rect 23290 7148 23296 7200
rect 23348 7148 23354 7200
rect 27614 7148 27620 7200
rect 27672 7188 27678 7200
rect 33137 7191 33195 7197
rect 33137 7188 33149 7191
rect 27672 7160 33149 7188
rect 27672 7148 27678 7160
rect 33137 7157 33149 7160
rect 33183 7157 33195 7191
rect 33137 7151 33195 7157
rect 33413 7191 33471 7197
rect 33413 7157 33425 7191
rect 33459 7188 33471 7191
rect 37366 7188 37372 7200
rect 33459 7160 37372 7188
rect 33459 7157 33471 7160
rect 33413 7151 33471 7157
rect 37366 7148 37372 7160
rect 37424 7148 37430 7200
rect 37476 7188 37504 7228
rect 38654 7188 38660 7200
rect 37476 7160 38660 7188
rect 38654 7148 38660 7160
rect 38712 7148 38718 7200
rect 38764 7188 38792 7228
rect 40586 7216 40592 7228
rect 40644 7216 40650 7268
rect 40218 7188 40224 7200
rect 38764 7160 40224 7188
rect 40218 7148 40224 7160
rect 40276 7148 40282 7200
rect 47302 7148 47308 7200
rect 47360 7148 47366 7200
rect 1104 7098 47840 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 37950 7098
rect 38002 7046 38014 7098
rect 38066 7046 38078 7098
rect 38130 7046 38142 7098
rect 38194 7046 38206 7098
rect 38258 7046 43950 7098
rect 44002 7046 44014 7098
rect 44066 7046 44078 7098
rect 44130 7046 44142 7098
rect 44194 7046 44206 7098
rect 44258 7046 47840 7098
rect 1104 7024 47840 7046
rect 23290 6944 23296 6996
rect 23348 6984 23354 6996
rect 43714 6984 43720 6996
rect 23348 6956 43720 6984
rect 23348 6944 23354 6956
rect 43714 6944 43720 6956
rect 43772 6944 43778 6996
rect 46014 6944 46020 6996
rect 46072 6984 46078 6996
rect 46201 6987 46259 6993
rect 46201 6984 46213 6987
rect 46072 6956 46213 6984
rect 46072 6944 46078 6956
rect 46201 6953 46213 6956
rect 46247 6953 46259 6987
rect 46201 6947 46259 6953
rect 27065 6919 27123 6925
rect 27065 6885 27077 6919
rect 27111 6885 27123 6919
rect 27065 6879 27123 6885
rect 12342 6808 12348 6860
rect 12400 6848 12406 6860
rect 18417 6851 18475 6857
rect 18417 6848 18429 6851
rect 12400 6820 18429 6848
rect 12400 6808 12406 6820
rect 18417 6817 18429 6820
rect 18463 6817 18475 6851
rect 26697 6851 26755 6857
rect 26697 6848 26709 6851
rect 18417 6811 18475 6817
rect 22066 6820 26709 6848
rect 1302 6740 1308 6792
rect 1360 6780 1366 6792
rect 22066 6780 22094 6820
rect 26697 6817 26709 6820
rect 26743 6817 26755 6851
rect 27080 6848 27108 6879
rect 36446 6876 36452 6928
rect 36504 6916 36510 6928
rect 44358 6916 44364 6928
rect 36504 6888 44364 6916
rect 36504 6876 36510 6888
rect 44358 6876 44364 6888
rect 44416 6876 44422 6928
rect 43806 6848 43812 6860
rect 27080 6820 43812 6848
rect 26697 6811 26755 6817
rect 43806 6808 43812 6820
rect 43864 6808 43870 6860
rect 46290 6848 46296 6860
rect 44744 6820 46296 6848
rect 1360 6752 22094 6780
rect 26053 6783 26111 6789
rect 1360 6740 1366 6752
rect 26053 6749 26065 6783
rect 26099 6780 26111 6783
rect 26145 6783 26203 6789
rect 26145 6780 26157 6783
rect 26099 6752 26157 6780
rect 26099 6749 26111 6752
rect 26053 6743 26111 6749
rect 26145 6749 26157 6752
rect 26191 6749 26203 6783
rect 26145 6743 26203 6749
rect 26789 6783 26847 6789
rect 26789 6749 26801 6783
rect 26835 6780 26847 6783
rect 26881 6783 26939 6789
rect 26881 6780 26893 6783
rect 26835 6752 26893 6780
rect 26835 6749 26847 6752
rect 26789 6743 26847 6749
rect 26881 6749 26893 6752
rect 26927 6749 26939 6783
rect 26881 6743 26939 6749
rect 40221 6783 40279 6789
rect 40221 6749 40233 6783
rect 40267 6780 40279 6783
rect 41509 6783 41567 6789
rect 40267 6752 41460 6780
rect 40267 6749 40279 6752
rect 40221 6743 40279 6749
rect 12250 6672 12256 6724
rect 12308 6712 12314 6724
rect 15565 6715 15623 6721
rect 15565 6712 15577 6715
rect 12308 6684 15577 6712
rect 12308 6672 12314 6684
rect 15565 6681 15577 6684
rect 15611 6712 15623 6715
rect 15841 6715 15899 6721
rect 15841 6712 15853 6715
rect 15611 6684 15853 6712
rect 15611 6681 15623 6684
rect 15565 6675 15623 6681
rect 15841 6681 15853 6684
rect 15887 6681 15899 6715
rect 15841 6675 15899 6681
rect 18509 6715 18567 6721
rect 18509 6681 18521 6715
rect 18555 6712 18567 6715
rect 18693 6715 18751 6721
rect 18693 6712 18705 6715
rect 18555 6684 18705 6712
rect 18555 6681 18567 6684
rect 18509 6675 18567 6681
rect 18693 6681 18705 6684
rect 18739 6681 18751 6715
rect 18693 6675 18751 6681
rect 18877 6715 18935 6721
rect 18877 6681 18889 6715
rect 18923 6712 18935 6715
rect 36538 6712 36544 6724
rect 18923 6684 36544 6712
rect 18923 6681 18935 6684
rect 18877 6675 18935 6681
rect 36538 6672 36544 6684
rect 36596 6672 36602 6724
rect 38562 6672 38568 6724
rect 38620 6712 38626 6724
rect 38620 6684 41368 6712
rect 38620 6672 38626 6684
rect 15933 6647 15991 6653
rect 15933 6613 15945 6647
rect 15979 6644 15991 6647
rect 18966 6644 18972 6656
rect 15979 6616 18972 6644
rect 15979 6613 15991 6616
rect 15933 6607 15991 6613
rect 18966 6604 18972 6616
rect 19024 6604 19030 6656
rect 25866 6604 25872 6656
rect 25924 6644 25930 6656
rect 25961 6647 26019 6653
rect 25961 6644 25973 6647
rect 25924 6616 25973 6644
rect 25924 6604 25930 6616
rect 25961 6613 25973 6616
rect 26007 6613 26019 6647
rect 25961 6607 26019 6613
rect 26326 6604 26332 6656
rect 26384 6604 26390 6656
rect 39942 6604 39948 6656
rect 40000 6644 40006 6656
rect 41340 6653 41368 6684
rect 40037 6647 40095 6653
rect 40037 6644 40049 6647
rect 40000 6616 40049 6644
rect 40000 6604 40006 6616
rect 40037 6613 40049 6616
rect 40083 6613 40095 6647
rect 40037 6607 40095 6613
rect 41325 6647 41383 6653
rect 41325 6613 41337 6647
rect 41371 6613 41383 6647
rect 41432 6644 41460 6752
rect 41509 6749 41521 6783
rect 41555 6780 41567 6783
rect 44634 6780 44640 6792
rect 41555 6752 44640 6780
rect 41555 6749 41567 6752
rect 41509 6743 41567 6749
rect 44634 6740 44640 6752
rect 44692 6740 44698 6792
rect 44744 6789 44772 6820
rect 46290 6808 46296 6820
rect 46348 6808 46354 6860
rect 44729 6783 44787 6789
rect 44729 6749 44741 6783
rect 44775 6749 44787 6783
rect 44729 6743 44787 6749
rect 46014 6740 46020 6792
rect 46072 6780 46078 6792
rect 46385 6783 46443 6789
rect 46385 6780 46397 6783
rect 46072 6752 46397 6780
rect 46072 6740 46078 6752
rect 46385 6749 46397 6752
rect 46431 6749 46443 6783
rect 46385 6743 46443 6749
rect 46658 6740 46664 6792
rect 46716 6740 46722 6792
rect 46845 6783 46903 6789
rect 46845 6749 46857 6783
rect 46891 6749 46903 6783
rect 46845 6743 46903 6749
rect 42702 6672 42708 6724
rect 42760 6712 42766 6724
rect 46860 6712 46888 6743
rect 47118 6740 47124 6792
rect 47176 6780 47182 6792
rect 47213 6783 47271 6789
rect 47213 6780 47225 6783
rect 47176 6752 47225 6780
rect 47176 6740 47182 6752
rect 47213 6749 47225 6752
rect 47259 6749 47271 6783
rect 47213 6743 47271 6749
rect 42760 6684 46888 6712
rect 42760 6672 42766 6684
rect 42794 6644 42800 6656
rect 41432 6616 42800 6644
rect 41325 6607 41383 6613
rect 42794 6604 42800 6616
rect 42852 6604 42858 6656
rect 43162 6604 43168 6656
rect 43220 6644 43226 6656
rect 44545 6647 44603 6653
rect 44545 6644 44557 6647
rect 43220 6616 44557 6644
rect 43220 6604 43226 6616
rect 44545 6613 44557 6616
rect 44591 6613 44603 6647
rect 44545 6607 44603 6613
rect 45462 6604 45468 6656
rect 45520 6644 45526 6656
rect 46477 6647 46535 6653
rect 46477 6644 46489 6647
rect 45520 6616 46489 6644
rect 45520 6604 45526 6616
rect 46477 6613 46489 6616
rect 46523 6613 46535 6647
rect 46477 6607 46535 6613
rect 47026 6604 47032 6656
rect 47084 6604 47090 6656
rect 47394 6604 47400 6656
rect 47452 6604 47458 6656
rect 1104 6554 47840 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 39010 6554
rect 39062 6502 39074 6554
rect 39126 6502 39138 6554
rect 39190 6502 39202 6554
rect 39254 6502 39266 6554
rect 39318 6502 45010 6554
rect 45062 6502 45074 6554
rect 45126 6502 45138 6554
rect 45190 6502 45202 6554
rect 45254 6502 45266 6554
rect 45318 6502 47840 6554
rect 1104 6480 47840 6502
rect 8662 6400 8668 6452
rect 8720 6440 8726 6452
rect 23290 6440 23296 6452
rect 8720 6412 23296 6440
rect 8720 6400 8726 6412
rect 23290 6400 23296 6412
rect 23348 6400 23354 6452
rect 26326 6400 26332 6452
rect 26384 6440 26390 6452
rect 40034 6440 40040 6452
rect 26384 6412 40040 6440
rect 26384 6400 26390 6412
rect 40034 6400 40040 6412
rect 40092 6400 40098 6452
rect 40402 6400 40408 6452
rect 40460 6440 40466 6452
rect 42429 6443 42487 6449
rect 42429 6440 42441 6443
rect 40460 6412 42441 6440
rect 40460 6400 40466 6412
rect 42429 6409 42441 6412
rect 42475 6409 42487 6443
rect 42429 6403 42487 6409
rect 47302 6400 47308 6452
rect 47360 6400 47366 6452
rect 18046 6332 18052 6384
rect 18104 6372 18110 6384
rect 30926 6372 30932 6384
rect 18104 6344 30932 6372
rect 18104 6332 18110 6344
rect 30926 6332 30932 6344
rect 30984 6332 30990 6384
rect 36538 6332 36544 6384
rect 36596 6372 36602 6384
rect 47210 6372 47216 6384
rect 36596 6344 47216 6372
rect 36596 6332 36602 6344
rect 47210 6332 47216 6344
rect 47268 6332 47274 6384
rect 3418 6264 3424 6316
rect 3476 6304 3482 6316
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 3476 6276 22017 6304
rect 3476 6264 3482 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 30374 6264 30380 6316
rect 30432 6304 30438 6316
rect 33597 6307 33655 6313
rect 33597 6304 33609 6307
rect 30432 6276 33609 6304
rect 30432 6264 30438 6276
rect 33597 6273 33609 6276
rect 33643 6304 33655 6307
rect 33781 6307 33839 6313
rect 33781 6304 33793 6307
rect 33643 6276 33793 6304
rect 33643 6273 33655 6276
rect 33597 6267 33655 6273
rect 33781 6273 33793 6276
rect 33827 6273 33839 6307
rect 33781 6267 33839 6273
rect 42613 6307 42671 6313
rect 42613 6273 42625 6307
rect 42659 6273 42671 6307
rect 42613 6267 42671 6273
rect 43533 6307 43591 6313
rect 43533 6273 43545 6307
rect 43579 6304 43591 6307
rect 45370 6304 45376 6316
rect 43579 6276 45376 6304
rect 43579 6273 43591 6276
rect 43533 6267 43591 6273
rect 1302 6196 1308 6248
rect 1360 6236 1366 6248
rect 26510 6236 26516 6248
rect 1360 6208 26516 6236
rect 1360 6196 1366 6208
rect 26510 6196 26516 6208
rect 26568 6196 26574 6248
rect 42628 6236 42656 6267
rect 45370 6264 45376 6276
rect 45428 6264 45434 6316
rect 46566 6264 46572 6316
rect 46624 6264 46630 6316
rect 47029 6307 47087 6313
rect 47029 6273 47041 6307
rect 47075 6304 47087 6307
rect 47121 6307 47179 6313
rect 47121 6304 47133 6307
rect 47075 6276 47133 6304
rect 47075 6273 47087 6276
rect 47029 6267 47087 6273
rect 47121 6273 47133 6276
rect 47167 6273 47179 6307
rect 47121 6267 47179 6273
rect 44910 6236 44916 6248
rect 42628 6208 44916 6236
rect 44910 6196 44916 6208
rect 44968 6196 44974 6248
rect 474 6128 480 6180
rect 532 6168 538 6180
rect 27614 6168 27620 6180
rect 532 6140 27620 6168
rect 532 6128 538 6140
rect 27614 6128 27620 6140
rect 27672 6128 27678 6180
rect 37182 6128 37188 6180
rect 37240 6168 37246 6180
rect 43349 6171 43407 6177
rect 43349 6168 43361 6171
rect 37240 6140 43361 6168
rect 37240 6128 37246 6140
rect 43349 6137 43361 6140
rect 43395 6137 43407 6171
rect 43349 6131 43407 6137
rect 22189 6103 22247 6109
rect 22189 6069 22201 6103
rect 22235 6100 22247 6103
rect 24762 6100 24768 6112
rect 22235 6072 24768 6100
rect 22235 6069 22247 6072
rect 22189 6063 22247 6069
rect 24762 6060 24768 6072
rect 24820 6060 24826 6112
rect 33965 6103 34023 6109
rect 33965 6069 33977 6103
rect 34011 6100 34023 6103
rect 35434 6100 35440 6112
rect 34011 6072 35440 6100
rect 34011 6069 34023 6072
rect 33965 6063 34023 6069
rect 35434 6060 35440 6072
rect 35492 6060 35498 6112
rect 46750 6060 46756 6112
rect 46808 6060 46814 6112
rect 46934 6060 46940 6112
rect 46992 6060 46998 6112
rect 1104 6010 47840 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 37950 6010
rect 38002 5958 38014 6010
rect 38066 5958 38078 6010
rect 38130 5958 38142 6010
rect 38194 5958 38206 6010
rect 38258 5958 43950 6010
rect 44002 5958 44014 6010
rect 44066 5958 44078 6010
rect 44130 5958 44142 6010
rect 44194 5958 44206 6010
rect 44258 5958 47840 6010
rect 1104 5936 47840 5958
rect 8662 5856 8668 5908
rect 8720 5856 8726 5908
rect 12158 5856 12164 5908
rect 12216 5896 12222 5908
rect 17957 5899 18015 5905
rect 17957 5896 17969 5899
rect 12216 5868 17969 5896
rect 12216 5856 12222 5868
rect 17957 5865 17969 5868
rect 18003 5865 18015 5899
rect 17957 5859 18015 5865
rect 19242 5856 19248 5908
rect 19300 5896 19306 5908
rect 19521 5899 19579 5905
rect 19521 5896 19533 5899
rect 19300 5868 19533 5896
rect 19300 5856 19306 5868
rect 19521 5865 19533 5868
rect 19567 5865 19579 5899
rect 19521 5859 19579 5865
rect 20714 5856 20720 5908
rect 20772 5896 20778 5908
rect 20772 5868 31754 5896
rect 20772 5856 20778 5868
rect 18417 5831 18475 5837
rect 18417 5797 18429 5831
rect 18463 5828 18475 5831
rect 24670 5828 24676 5840
rect 18463 5800 24676 5828
rect 18463 5797 18475 5800
rect 18417 5791 18475 5797
rect 24670 5788 24676 5800
rect 24728 5788 24734 5840
rect 31726 5828 31754 5868
rect 42794 5856 42800 5908
rect 42852 5896 42858 5908
rect 43806 5896 43812 5908
rect 42852 5868 43812 5896
rect 42852 5856 42858 5868
rect 43806 5856 43812 5868
rect 43864 5856 43870 5908
rect 46934 5828 46940 5840
rect 31726 5800 46940 5828
rect 46934 5788 46940 5800
rect 46992 5788 46998 5840
rect 47394 5788 47400 5840
rect 47452 5788 47458 5840
rect 18966 5720 18972 5772
rect 19024 5760 19030 5772
rect 46106 5760 46112 5772
rect 19024 5732 46112 5760
rect 19024 5720 19030 5732
rect 46106 5720 46112 5732
rect 46164 5720 46170 5772
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 12618 5692 12624 5704
rect 8527 5664 12624 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 12618 5652 12624 5664
rect 12676 5652 12682 5704
rect 14553 5695 14611 5701
rect 14553 5661 14565 5695
rect 14599 5692 14611 5695
rect 15930 5692 15936 5704
rect 14599 5664 15936 5692
rect 14599 5661 14611 5664
rect 14553 5655 14611 5661
rect 15930 5652 15936 5664
rect 15988 5652 15994 5704
rect 18049 5695 18107 5701
rect 18049 5661 18061 5695
rect 18095 5692 18107 5695
rect 18233 5695 18291 5701
rect 18233 5692 18245 5695
rect 18095 5664 18245 5692
rect 18095 5661 18107 5664
rect 18049 5655 18107 5661
rect 18233 5661 18245 5664
rect 18279 5661 18291 5695
rect 18233 5655 18291 5661
rect 19613 5695 19671 5701
rect 19613 5661 19625 5695
rect 19659 5692 19671 5695
rect 19705 5695 19763 5701
rect 19705 5692 19717 5695
rect 19659 5664 19717 5692
rect 19659 5661 19671 5664
rect 19613 5655 19671 5661
rect 19705 5661 19717 5664
rect 19751 5661 19763 5695
rect 19705 5655 19763 5661
rect 22002 5652 22008 5704
rect 22060 5692 22066 5704
rect 27522 5692 27528 5704
rect 22060 5664 27528 5692
rect 22060 5652 22066 5664
rect 27522 5652 27528 5664
rect 27580 5652 27586 5704
rect 32766 5652 32772 5704
rect 32824 5692 32830 5704
rect 32953 5695 33011 5701
rect 32953 5692 32965 5695
rect 32824 5664 32965 5692
rect 32824 5652 32830 5664
rect 32953 5661 32965 5664
rect 32999 5661 33011 5695
rect 32953 5655 33011 5661
rect 45554 5652 45560 5704
rect 45612 5692 45618 5704
rect 46845 5695 46903 5701
rect 46845 5692 46857 5695
rect 45612 5664 46857 5692
rect 45612 5652 45618 5664
rect 46845 5661 46857 5664
rect 46891 5661 46903 5695
rect 46845 5655 46903 5661
rect 47210 5652 47216 5704
rect 47268 5652 47274 5704
rect 18966 5584 18972 5636
rect 19024 5624 19030 5636
rect 30466 5624 30472 5636
rect 19024 5596 30472 5624
rect 19024 5584 19030 5596
rect 30466 5584 30472 5596
rect 30524 5584 30530 5636
rect 47118 5624 47124 5636
rect 31726 5596 47124 5624
rect 14737 5559 14795 5565
rect 14737 5525 14749 5559
rect 14783 5556 14795 5559
rect 14918 5556 14924 5568
rect 14783 5528 14924 5556
rect 14783 5525 14795 5528
rect 14737 5519 14795 5525
rect 14918 5516 14924 5528
rect 14976 5516 14982 5568
rect 19889 5559 19947 5565
rect 19889 5525 19901 5559
rect 19935 5556 19947 5559
rect 31726 5556 31754 5596
rect 47118 5584 47124 5596
rect 47176 5584 47182 5636
rect 19935 5528 31754 5556
rect 33137 5559 33195 5565
rect 19935 5525 19947 5528
rect 19889 5519 19947 5525
rect 33137 5525 33149 5559
rect 33183 5556 33195 5559
rect 46198 5556 46204 5568
rect 33183 5528 46204 5556
rect 33183 5525 33195 5528
rect 33137 5519 33195 5525
rect 46198 5516 46204 5528
rect 46256 5516 46262 5568
rect 47026 5516 47032 5568
rect 47084 5516 47090 5568
rect 1104 5466 47840 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 39010 5466
rect 39062 5414 39074 5466
rect 39126 5414 39138 5466
rect 39190 5414 39202 5466
rect 39254 5414 39266 5466
rect 39318 5414 45010 5466
rect 45062 5414 45074 5466
rect 45126 5414 45138 5466
rect 45190 5414 45202 5466
rect 45254 5414 45266 5466
rect 45318 5414 47840 5466
rect 1104 5392 47840 5414
rect 8573 5355 8631 5361
rect 8573 5321 8585 5355
rect 8619 5352 8631 5355
rect 11422 5352 11428 5364
rect 8619 5324 11428 5352
rect 8619 5321 8631 5324
rect 8573 5315 8631 5321
rect 11422 5312 11428 5324
rect 11480 5312 11486 5364
rect 11514 5312 11520 5364
rect 11572 5352 11578 5364
rect 17681 5355 17739 5361
rect 11572 5324 17632 5352
rect 11572 5312 11578 5324
rect 11054 5284 11060 5296
rect 8128 5256 11060 5284
rect 8128 5225 8156 5256
rect 11054 5244 11060 5256
rect 11112 5244 11118 5296
rect 15470 5284 15476 5296
rect 11164 5256 12664 5284
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5185 8171 5219
rect 8113 5179 8171 5185
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5185 8447 5219
rect 8389 5179 8447 5185
rect 9217 5219 9275 5225
rect 9217 5185 9229 5219
rect 9263 5185 9275 5219
rect 9217 5179 9275 5185
rect 8404 5080 8432 5179
rect 9232 5148 9260 5179
rect 10410 5176 10416 5228
rect 10468 5176 10474 5228
rect 11164 5225 11192 5256
rect 11149 5219 11207 5225
rect 11149 5185 11161 5219
rect 11195 5185 11207 5219
rect 11149 5179 11207 5185
rect 12342 5176 12348 5228
rect 12400 5176 12406 5228
rect 12636 5148 12664 5256
rect 12728 5256 15476 5284
rect 12728 5225 12756 5256
rect 15470 5244 15476 5256
rect 15528 5244 15534 5296
rect 12713 5219 12771 5225
rect 12713 5185 12725 5219
rect 12759 5185 12771 5219
rect 12713 5179 12771 5185
rect 13751 5219 13809 5225
rect 13751 5185 13763 5219
rect 13797 5216 13809 5219
rect 15289 5219 15347 5225
rect 13797 5188 15240 5216
rect 13797 5185 13809 5188
rect 13751 5179 13809 5185
rect 14274 5148 14280 5160
rect 9232 5120 12296 5148
rect 12636 5120 14280 5148
rect 11882 5080 11888 5092
rect 8404 5052 11888 5080
rect 11882 5040 11888 5052
rect 11940 5040 11946 5092
rect 8297 5015 8355 5021
rect 8297 4981 8309 5015
rect 8343 5012 8355 5015
rect 8478 5012 8484 5024
rect 8343 4984 8484 5012
rect 8343 4981 8355 4984
rect 8297 4975 8355 4981
rect 8478 4972 8484 4984
rect 8536 4972 8542 5024
rect 9401 5015 9459 5021
rect 9401 4981 9413 5015
rect 9447 5012 9459 5015
rect 10502 5012 10508 5024
rect 9447 4984 10508 5012
rect 9447 4981 9459 4984
rect 9401 4975 9459 4981
rect 10502 4972 10508 4984
rect 10560 4972 10566 5024
rect 10594 4972 10600 5024
rect 10652 4972 10658 5024
rect 11330 4972 11336 5024
rect 11388 4972 11394 5024
rect 12268 5012 12296 5120
rect 14274 5108 14280 5120
rect 14332 5108 14338 5160
rect 15212 5148 15240 5188
rect 15289 5185 15301 5219
rect 15335 5216 15347 5219
rect 16206 5216 16212 5228
rect 15335 5188 16212 5216
rect 15335 5185 15347 5188
rect 15289 5179 15347 5185
rect 16206 5176 16212 5188
rect 16264 5176 16270 5228
rect 16301 5219 16359 5225
rect 16301 5185 16313 5219
rect 16347 5216 16359 5219
rect 16666 5216 16672 5228
rect 16347 5188 16672 5216
rect 16347 5185 16359 5188
rect 16301 5179 16359 5185
rect 16666 5176 16672 5188
rect 16724 5176 16730 5228
rect 17034 5176 17040 5228
rect 17092 5176 17098 5228
rect 17402 5176 17408 5228
rect 17460 5216 17466 5228
rect 17497 5219 17555 5225
rect 17497 5216 17509 5219
rect 17460 5188 17509 5216
rect 17460 5176 17466 5188
rect 17497 5185 17509 5188
rect 17543 5185 17555 5219
rect 17604 5216 17632 5324
rect 17681 5321 17693 5355
rect 17727 5321 17739 5355
rect 17681 5315 17739 5321
rect 17696 5284 17724 5315
rect 22002 5312 22008 5364
rect 22060 5312 22066 5364
rect 23845 5355 23903 5361
rect 23845 5321 23857 5355
rect 23891 5352 23903 5355
rect 25133 5355 25191 5361
rect 23891 5324 25084 5352
rect 23891 5321 23903 5324
rect 23845 5315 23903 5321
rect 21634 5284 21640 5296
rect 17696 5256 21640 5284
rect 21634 5244 21640 5256
rect 21692 5244 21698 5296
rect 25056 5284 25084 5324
rect 25133 5321 25145 5355
rect 25179 5352 25191 5355
rect 46566 5352 46572 5364
rect 25179 5324 46572 5352
rect 25179 5321 25191 5324
rect 25133 5315 25191 5321
rect 46566 5312 46572 5324
rect 46624 5312 46630 5364
rect 47302 5312 47308 5364
rect 47360 5312 47366 5364
rect 26602 5284 26608 5296
rect 25056 5256 26608 5284
rect 21821 5243 21879 5249
rect 26602 5244 26608 5256
rect 26660 5244 26666 5296
rect 45646 5244 45652 5296
rect 45704 5284 45710 5296
rect 47210 5284 47216 5296
rect 45704 5256 47216 5284
rect 45704 5244 45710 5256
rect 47210 5244 47216 5256
rect 47268 5244 47274 5296
rect 21726 5216 21732 5228
rect 17604 5188 21732 5216
rect 17497 5179 17555 5185
rect 21726 5176 21732 5188
rect 21784 5176 21790 5228
rect 21821 5209 21833 5243
rect 21867 5240 21879 5243
rect 21867 5212 22048 5240
rect 21867 5209 21879 5212
rect 21821 5203 21879 5209
rect 15562 5148 15568 5160
rect 15212 5120 15568 5148
rect 15562 5108 15568 5120
rect 15620 5108 15626 5160
rect 22020 5148 22048 5212
rect 23569 5219 23627 5225
rect 23569 5185 23581 5219
rect 23615 5216 23627 5219
rect 23661 5219 23719 5225
rect 23661 5216 23673 5219
rect 23615 5188 23673 5216
rect 23615 5185 23627 5188
rect 23569 5179 23627 5185
rect 23661 5185 23673 5188
rect 23707 5185 23719 5219
rect 23661 5179 23719 5185
rect 23937 5219 23995 5225
rect 23937 5185 23949 5219
rect 23983 5185 23995 5219
rect 23937 5179 23995 5185
rect 22097 5151 22155 5157
rect 22097 5148 22109 5151
rect 16408 5120 22109 5148
rect 12526 5040 12532 5092
rect 12584 5040 12590 5092
rect 13722 5040 13728 5092
rect 13780 5080 13786 5092
rect 16408 5080 16436 5120
rect 22097 5117 22109 5120
rect 22143 5117 22155 5151
rect 22097 5111 22155 5117
rect 23293 5151 23351 5157
rect 23293 5117 23305 5151
rect 23339 5148 23351 5151
rect 23952 5148 23980 5179
rect 24026 5176 24032 5228
rect 24084 5216 24090 5228
rect 24949 5219 25007 5225
rect 24949 5216 24961 5219
rect 24084 5188 24961 5216
rect 24084 5176 24090 5188
rect 24949 5185 24961 5188
rect 24995 5185 25007 5219
rect 24949 5179 25007 5185
rect 26970 5176 26976 5228
rect 27028 5216 27034 5228
rect 27249 5219 27307 5225
rect 27249 5216 27261 5219
rect 27028 5188 27261 5216
rect 27028 5176 27034 5188
rect 27249 5185 27261 5188
rect 27295 5185 27307 5219
rect 27249 5179 27307 5185
rect 27433 5219 27491 5225
rect 27433 5185 27445 5219
rect 27479 5185 27491 5219
rect 27433 5179 27491 5185
rect 23339 5120 23980 5148
rect 23339 5117 23351 5120
rect 23293 5111 23351 5117
rect 13780 5052 16436 5080
rect 16485 5083 16543 5089
rect 13780 5040 13786 5052
rect 16485 5049 16497 5083
rect 16531 5080 16543 5083
rect 18598 5080 18604 5092
rect 16531 5052 18604 5080
rect 16531 5049 16543 5052
rect 16485 5043 16543 5049
rect 18598 5040 18604 5052
rect 18656 5040 18662 5092
rect 27448 5080 27476 5179
rect 43714 5176 43720 5228
rect 43772 5216 43778 5228
rect 46753 5219 46811 5225
rect 46753 5216 46765 5219
rect 43772 5188 46765 5216
rect 43772 5176 43778 5188
rect 46753 5185 46765 5188
rect 46799 5185 46811 5219
rect 46753 5179 46811 5185
rect 47121 5219 47179 5225
rect 47121 5185 47133 5219
rect 47167 5185 47179 5219
rect 47121 5179 47179 5185
rect 22066 5052 27476 5080
rect 12710 5012 12716 5024
rect 12268 4984 12716 5012
rect 12710 4972 12716 4984
rect 12768 4972 12774 5024
rect 12894 4972 12900 5024
rect 12952 4972 12958 5024
rect 13909 5015 13967 5021
rect 13909 4981 13921 5015
rect 13955 5012 13967 5015
rect 15378 5012 15384 5024
rect 13955 4984 15384 5012
rect 13955 4981 13967 4984
rect 13909 4975 13967 4981
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 15473 5015 15531 5021
rect 15473 4981 15485 5015
rect 15519 5012 15531 5015
rect 17126 5012 17132 5024
rect 15519 4984 17132 5012
rect 15519 4981 15531 4984
rect 15473 4975 15531 4981
rect 17126 4972 17132 4984
rect 17184 4972 17190 5024
rect 17218 4972 17224 5024
rect 17276 4972 17282 5024
rect 17862 4972 17868 5024
rect 17920 5012 17926 5024
rect 22066 5012 22094 5052
rect 27522 5040 27528 5092
rect 27580 5080 27586 5092
rect 42702 5080 42708 5092
rect 27580 5052 42708 5080
rect 27580 5040 27586 5052
rect 42702 5040 42708 5052
rect 42760 5040 42766 5092
rect 17920 4984 22094 5012
rect 17920 4972 17926 4984
rect 23198 4972 23204 5024
rect 23256 4972 23262 5024
rect 23474 4972 23480 5024
rect 23532 4972 23538 5024
rect 24121 5015 24179 5021
rect 24121 4981 24133 5015
rect 24167 5012 24179 5015
rect 26878 5012 26884 5024
rect 24167 4984 26884 5012
rect 24167 4981 24179 4984
rect 24121 4975 24179 4981
rect 26878 4972 26884 4984
rect 26936 4972 26942 5024
rect 27157 5015 27215 5021
rect 27157 4981 27169 5015
rect 27203 5012 27215 5015
rect 27430 5012 27436 5024
rect 27203 4984 27436 5012
rect 27203 4981 27215 4984
rect 27157 4975 27215 4981
rect 27430 4972 27436 4984
rect 27488 4972 27494 5024
rect 27617 5015 27675 5021
rect 27617 4981 27629 5015
rect 27663 5012 27675 5015
rect 29638 5012 29644 5024
rect 27663 4984 29644 5012
rect 27663 4981 27675 4984
rect 27617 4975 27675 4981
rect 29638 4972 29644 4984
rect 29696 4972 29702 5024
rect 46934 4972 46940 5024
rect 46992 4972 46998 5024
rect 47136 5012 47164 5179
rect 47136 4984 47900 5012
rect 1104 4922 47840 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 37950 4922
rect 38002 4870 38014 4922
rect 38066 4870 38078 4922
rect 38130 4870 38142 4922
rect 38194 4870 38206 4922
rect 38258 4870 43950 4922
rect 44002 4870 44014 4922
rect 44066 4870 44078 4922
rect 44130 4870 44142 4922
rect 44194 4870 44206 4922
rect 44258 4870 47840 4922
rect 1104 4848 47840 4870
rect 4157 4811 4215 4817
rect 4157 4777 4169 4811
rect 4203 4808 4215 4811
rect 7742 4808 7748 4820
rect 4203 4780 7748 4808
rect 4203 4777 4215 4780
rect 4157 4771 4215 4777
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 10410 4768 10416 4820
rect 10468 4808 10474 4820
rect 13722 4808 13728 4820
rect 10468 4780 13728 4808
rect 10468 4768 10474 4780
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 14734 4768 14740 4820
rect 14792 4808 14798 4820
rect 17862 4808 17868 4820
rect 14792 4780 17868 4808
rect 14792 4768 14798 4780
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 21634 4768 21640 4820
rect 21692 4808 21698 4820
rect 31754 4808 31760 4820
rect 21692 4780 31760 4808
rect 21692 4768 21698 4780
rect 31754 4768 31760 4780
rect 31812 4768 31818 4820
rect 42794 4808 42800 4820
rect 31864 4780 42800 4808
rect 2869 4743 2927 4749
rect 2869 4709 2881 4743
rect 2915 4740 2927 4743
rect 2915 4712 11836 4740
rect 2915 4709 2927 4712
rect 2869 4703 2927 4709
rect 4522 4672 4528 4684
rect 3988 4644 4528 4672
rect 2409 4607 2467 4613
rect 2409 4573 2421 4607
rect 2455 4604 2467 4607
rect 2590 4604 2596 4616
rect 2455 4576 2596 4604
rect 2455 4573 2467 4576
rect 2409 4567 2467 4573
rect 2590 4564 2596 4576
rect 2648 4564 2654 4616
rect 3988 4613 4016 4644
rect 4522 4632 4528 4644
rect 4580 4632 4586 4684
rect 6730 4632 6736 4684
rect 6788 4672 6794 4684
rect 11808 4672 11836 4712
rect 12342 4700 12348 4752
rect 12400 4740 12406 4752
rect 14826 4740 14832 4752
rect 12400 4712 14832 4740
rect 12400 4700 12406 4712
rect 14826 4700 14832 4712
rect 14884 4700 14890 4752
rect 17218 4700 17224 4752
rect 17276 4740 17282 4752
rect 25314 4740 25320 4752
rect 17276 4712 25320 4740
rect 17276 4700 17282 4712
rect 25314 4700 25320 4712
rect 25372 4700 25378 4752
rect 29638 4700 29644 4752
rect 29696 4740 29702 4752
rect 31864 4740 31892 4780
rect 42794 4768 42800 4780
rect 42852 4768 42858 4820
rect 29696 4712 31892 4740
rect 29696 4700 29702 4712
rect 40034 4700 40040 4752
rect 40092 4740 40098 4752
rect 40092 4712 47256 4740
rect 40092 4700 40098 4712
rect 16574 4672 16580 4684
rect 6788 4644 11652 4672
rect 11808 4644 16580 4672
rect 6788 4632 6794 4644
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4573 2743 4607
rect 2685 4567 2743 4573
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 4801 4607 4859 4613
rect 4801 4573 4813 4607
rect 4847 4604 4859 4607
rect 4847 4576 5212 4604
rect 4847 4573 4859 4576
rect 4801 4567 4859 4573
rect 2314 4496 2320 4548
rect 2372 4536 2378 4548
rect 2700 4536 2728 4567
rect 2372 4508 2728 4536
rect 4264 4536 4292 4567
rect 4890 4536 4896 4548
rect 4264 4508 4896 4536
rect 2372 4496 2378 4508
rect 4890 4496 4896 4508
rect 4948 4496 4954 4548
rect 5184 4536 5212 4576
rect 5258 4564 5264 4616
rect 5316 4604 5322 4616
rect 5537 4607 5595 4613
rect 5537 4604 5549 4607
rect 5316 4576 5549 4604
rect 5316 4564 5322 4576
rect 5537 4573 5549 4576
rect 5583 4573 5595 4607
rect 5537 4567 5595 4573
rect 6273 4607 6331 4613
rect 6273 4573 6285 4607
rect 6319 4604 6331 4607
rect 7466 4604 7472 4616
rect 6319 4576 7472 4604
rect 6319 4573 6331 4576
rect 6273 4567 6331 4573
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 5626 4536 5632 4548
rect 5184 4508 5632 4536
rect 5626 4496 5632 4508
rect 5684 4496 5690 4548
rect 8202 4536 8208 4548
rect 5736 4508 8208 4536
rect 2593 4471 2651 4477
rect 2593 4437 2605 4471
rect 2639 4468 2651 4471
rect 2774 4468 2780 4480
rect 2639 4440 2780 4468
rect 2639 4437 2651 4440
rect 2593 4431 2651 4437
rect 2774 4428 2780 4440
rect 2832 4428 2838 4480
rect 4430 4428 4436 4480
rect 4488 4428 4494 4480
rect 4985 4471 5043 4477
rect 4985 4437 4997 4471
rect 5031 4468 5043 4471
rect 5534 4468 5540 4480
rect 5031 4440 5540 4468
rect 5031 4437 5043 4440
rect 4985 4431 5043 4437
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 5736 4477 5764 4508
rect 8202 4496 8208 4508
rect 8260 4496 8266 4548
rect 5721 4471 5779 4477
rect 5721 4437 5733 4471
rect 5767 4437 5779 4471
rect 5721 4431 5779 4437
rect 6457 4471 6515 4477
rect 6457 4437 6469 4471
rect 6503 4468 6515 4471
rect 9582 4468 9588 4480
rect 6503 4440 9588 4468
rect 6503 4437 6515 4440
rect 6457 4431 6515 4437
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 11624 4468 11652 4644
rect 16574 4632 16580 4644
rect 16632 4632 16638 4684
rect 23198 4672 23204 4684
rect 17236 4644 23204 4672
rect 17236 4468 17264 4644
rect 23198 4632 23204 4644
rect 23256 4632 23262 4684
rect 27430 4632 27436 4684
rect 27488 4672 27494 4684
rect 41598 4672 41604 4684
rect 27488 4644 41604 4672
rect 27488 4632 27494 4644
rect 41598 4632 41604 4644
rect 41656 4632 41662 4684
rect 19242 4564 19248 4616
rect 19300 4564 19306 4616
rect 20898 4564 20904 4616
rect 20956 4604 20962 4616
rect 21177 4607 21235 4613
rect 21177 4604 21189 4607
rect 20956 4576 21189 4604
rect 20956 4564 20962 4576
rect 21177 4573 21189 4576
rect 21223 4573 21235 4607
rect 21177 4567 21235 4573
rect 26789 4607 26847 4613
rect 26789 4573 26801 4607
rect 26835 4604 26847 4607
rect 26881 4607 26939 4613
rect 26881 4604 26893 4607
rect 26835 4576 26893 4604
rect 26835 4573 26847 4576
rect 26789 4567 26847 4573
rect 26881 4573 26893 4576
rect 26927 4573 26939 4607
rect 26881 4567 26939 4573
rect 31754 4564 31760 4616
rect 31812 4604 31818 4616
rect 36998 4604 37004 4616
rect 31812 4576 37004 4604
rect 31812 4564 31818 4576
rect 36998 4564 37004 4576
rect 37056 4564 37062 4616
rect 37366 4564 37372 4616
rect 37424 4604 37430 4616
rect 47228 4613 47256 4712
rect 47394 4700 47400 4752
rect 47452 4700 47458 4752
rect 46845 4607 46903 4613
rect 46845 4604 46857 4607
rect 37424 4576 46857 4604
rect 37424 4564 37430 4576
rect 46845 4573 46857 4576
rect 46891 4573 46903 4607
rect 46845 4567 46903 4573
rect 47213 4607 47271 4613
rect 47213 4573 47225 4607
rect 47259 4573 47271 4607
rect 47213 4567 47271 4573
rect 19334 4496 19340 4548
rect 19392 4536 19398 4548
rect 47872 4536 47900 4984
rect 19392 4508 47900 4536
rect 19392 4496 19398 4508
rect 11624 4440 17264 4468
rect 19426 4428 19432 4480
rect 19484 4428 19490 4480
rect 21361 4471 21419 4477
rect 21361 4437 21373 4471
rect 21407 4468 21419 4471
rect 22002 4468 22008 4480
rect 21407 4440 22008 4468
rect 21407 4437 21419 4440
rect 21361 4431 21419 4437
rect 22002 4428 22008 4440
rect 22060 4428 22066 4480
rect 26694 4428 26700 4480
rect 26752 4428 26758 4480
rect 27065 4471 27123 4477
rect 27065 4437 27077 4471
rect 27111 4468 27123 4471
rect 37182 4468 37188 4480
rect 27111 4440 37188 4468
rect 27111 4437 27123 4440
rect 27065 4431 27123 4437
rect 37182 4428 37188 4440
rect 37240 4428 37246 4480
rect 47026 4428 47032 4480
rect 47084 4428 47090 4480
rect 1104 4378 47840 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 39010 4378
rect 39062 4326 39074 4378
rect 39126 4326 39138 4378
rect 39190 4326 39202 4378
rect 39254 4326 39266 4378
rect 39318 4326 45010 4378
rect 45062 4326 45074 4378
rect 45126 4326 45138 4378
rect 45190 4326 45202 4378
rect 45254 4326 45266 4378
rect 45318 4326 47840 4378
rect 1104 4304 47840 4326
rect 2774 4224 2780 4276
rect 2832 4264 2838 4276
rect 2832 4236 12388 4264
rect 2832 4224 2838 4236
rect 1118 4156 1124 4208
rect 1176 4196 1182 4208
rect 2225 4199 2283 4205
rect 2225 4196 2237 4199
rect 1176 4168 2237 4196
rect 1176 4156 1182 4168
rect 2225 4165 2237 4168
rect 2271 4165 2283 4199
rect 2225 4159 2283 4165
rect 4430 4156 4436 4208
rect 4488 4196 4494 4208
rect 5718 4196 5724 4208
rect 4488 4168 5724 4196
rect 4488 4156 4494 4168
rect 5718 4156 5724 4168
rect 5776 4156 5782 4208
rect 8202 4156 8208 4208
rect 8260 4196 8266 4208
rect 8260 4168 8892 4196
rect 8260 4156 8266 4168
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4128 7435 4131
rect 7834 4128 7840 4140
rect 7423 4100 7840 4128
rect 7423 4097 7435 4100
rect 7377 4091 7435 4097
rect 7834 4088 7840 4100
rect 7892 4088 7898 4140
rect 8481 4131 8539 4137
rect 8481 4097 8493 4131
rect 8527 4128 8539 4131
rect 8570 4128 8576 4140
rect 8527 4100 8576 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 8757 4131 8815 4137
rect 8757 4097 8769 4131
rect 8803 4097 8815 4131
rect 8864 4128 8892 4168
rect 11054 4156 11060 4208
rect 11112 4196 11118 4208
rect 12250 4196 12256 4208
rect 11112 4168 12256 4196
rect 11112 4156 11118 4168
rect 12250 4156 12256 4168
rect 12308 4156 12314 4208
rect 12360 4196 12388 4236
rect 16482 4224 16488 4276
rect 16540 4264 16546 4276
rect 26694 4264 26700 4276
rect 16540 4236 26700 4264
rect 16540 4224 16546 4236
rect 26694 4224 26700 4236
rect 26752 4224 26758 4276
rect 26786 4224 26792 4276
rect 26844 4264 26850 4276
rect 42426 4264 42432 4276
rect 26844 4236 42432 4264
rect 26844 4224 26850 4236
rect 42426 4224 42432 4236
rect 42484 4224 42490 4276
rect 15838 4196 15844 4208
rect 12360 4168 15844 4196
rect 15838 4156 15844 4168
rect 15896 4156 15902 4208
rect 16574 4156 16580 4208
rect 16632 4196 16638 4208
rect 16632 4168 18368 4196
rect 16632 4156 16638 4168
rect 18340 4128 18368 4168
rect 18414 4156 18420 4208
rect 18472 4196 18478 4208
rect 18693 4199 18751 4205
rect 18693 4196 18705 4199
rect 18472 4168 18705 4196
rect 18472 4156 18478 4168
rect 18693 4165 18705 4168
rect 18739 4165 18751 4199
rect 20622 4196 20628 4208
rect 18693 4159 18751 4165
rect 18800 4168 20628 4196
rect 18800 4128 18828 4168
rect 20622 4156 20628 4168
rect 20680 4156 20686 4208
rect 25866 4156 25872 4208
rect 25924 4196 25930 4208
rect 46014 4196 46020 4208
rect 25924 4168 46020 4196
rect 25924 4156 25930 4168
rect 46014 4156 46020 4168
rect 46072 4156 46078 4208
rect 8864 4100 17264 4128
rect 18340 4100 18828 4128
rect 18877 4131 18935 4137
rect 8757 4091 8815 4097
rect 2406 4020 2412 4072
rect 2464 4020 2470 4072
rect 8294 4020 8300 4072
rect 8352 4060 8358 4072
rect 8772 4060 8800 4091
rect 15746 4060 15752 4072
rect 8352 4032 8800 4060
rect 8864 4032 15752 4060
rect 8352 4020 8358 4032
rect 7558 3884 7564 3936
rect 7616 3884 7622 3936
rect 8665 3927 8723 3933
rect 8665 3893 8677 3927
rect 8711 3924 8723 3927
rect 8864 3924 8892 4032
rect 15746 4020 15752 4032
rect 15804 4020 15810 4072
rect 17236 4060 17264 4100
rect 18877 4097 18889 4131
rect 18923 4128 18935 4131
rect 20714 4128 20720 4140
rect 18923 4100 20720 4128
rect 18923 4097 18935 4100
rect 18877 4091 18935 4097
rect 20714 4088 20720 4100
rect 20772 4088 20778 4140
rect 40034 4088 40040 4140
rect 40092 4128 40098 4140
rect 40221 4131 40279 4137
rect 40221 4128 40233 4131
rect 40092 4100 40233 4128
rect 40092 4088 40098 4100
rect 40221 4097 40233 4100
rect 40267 4097 40279 4131
rect 40221 4091 40279 4097
rect 42426 4088 42432 4140
rect 42484 4128 42490 4140
rect 42705 4131 42763 4137
rect 42705 4128 42717 4131
rect 42484 4100 42717 4128
rect 42484 4088 42490 4100
rect 42705 4097 42717 4100
rect 42751 4097 42763 4131
rect 42705 4091 42763 4097
rect 46385 4131 46443 4137
rect 46385 4097 46397 4131
rect 46431 4128 46443 4131
rect 46477 4131 46535 4137
rect 46477 4128 46489 4131
rect 46431 4100 46489 4128
rect 46431 4097 46443 4100
rect 46385 4091 46443 4097
rect 46477 4097 46489 4100
rect 46523 4097 46535 4131
rect 46477 4091 46535 4097
rect 46753 4131 46811 4137
rect 46753 4097 46765 4131
rect 46799 4097 46811 4131
rect 46753 4091 46811 4097
rect 47121 4131 47179 4137
rect 47121 4097 47133 4131
rect 47167 4097 47179 4131
rect 47121 4091 47179 4097
rect 22462 4060 22468 4072
rect 17236 4032 22468 4060
rect 22462 4020 22468 4032
rect 22520 4020 22526 4072
rect 44358 4020 44364 4072
rect 44416 4060 44422 4072
rect 46768 4060 46796 4091
rect 44416 4032 46796 4060
rect 44416 4020 44422 4032
rect 23290 3952 23296 4004
rect 23348 3992 23354 4004
rect 30650 3992 30656 4004
rect 23348 3964 30656 3992
rect 23348 3952 23354 3964
rect 30650 3952 30656 3964
rect 30708 3952 30714 4004
rect 40405 3995 40463 4001
rect 40405 3961 40417 3995
rect 40451 3992 40463 3995
rect 47136 3992 47164 4091
rect 40451 3964 47164 3992
rect 40451 3961 40463 3964
rect 40405 3955 40463 3961
rect 47302 3952 47308 4004
rect 47360 3952 47366 4004
rect 8711 3896 8892 3924
rect 8941 3927 8999 3933
rect 8711 3893 8723 3896
rect 8665 3887 8723 3893
rect 8941 3893 8953 3927
rect 8987 3924 8999 3927
rect 15654 3924 15660 3936
rect 8987 3896 15660 3924
rect 8987 3893 8999 3896
rect 8941 3887 8999 3893
rect 15654 3884 15660 3896
rect 15712 3884 15718 3936
rect 18874 3884 18880 3936
rect 18932 3924 18938 3936
rect 28258 3924 28264 3936
rect 18932 3896 28264 3924
rect 18932 3884 18938 3896
rect 28258 3884 28264 3896
rect 28316 3884 28322 3936
rect 30834 3884 30840 3936
rect 30892 3924 30898 3936
rect 33502 3924 33508 3936
rect 30892 3896 33508 3924
rect 30892 3884 30898 3896
rect 33502 3884 33508 3896
rect 33560 3884 33566 3936
rect 42610 3884 42616 3936
rect 42668 3884 42674 3936
rect 46290 3884 46296 3936
rect 46348 3884 46354 3936
rect 46661 3927 46719 3933
rect 46661 3893 46673 3927
rect 46707 3924 46719 3927
rect 46842 3924 46848 3936
rect 46707 3896 46848 3924
rect 46707 3893 46719 3896
rect 46661 3887 46719 3893
rect 46842 3884 46848 3896
rect 46900 3884 46906 3936
rect 46934 3884 46940 3936
rect 46992 3884 46998 3936
rect 1104 3834 47840 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 37950 3834
rect 38002 3782 38014 3834
rect 38066 3782 38078 3834
rect 38130 3782 38142 3834
rect 38194 3782 38206 3834
rect 38258 3782 43950 3834
rect 44002 3782 44014 3834
rect 44066 3782 44078 3834
rect 44130 3782 44142 3834
rect 44194 3782 44206 3834
rect 44258 3782 47840 3834
rect 1104 3760 47840 3782
rect 15378 3680 15384 3732
rect 15436 3720 15442 3732
rect 38838 3720 38844 3732
rect 15436 3692 38844 3720
rect 15436 3680 15442 3692
rect 38838 3680 38844 3692
rect 38896 3680 38902 3732
rect 46014 3680 46020 3732
rect 46072 3680 46078 3732
rect 8478 3612 8484 3664
rect 8536 3652 8542 3664
rect 18874 3652 18880 3664
rect 8536 3624 18880 3652
rect 8536 3612 8542 3624
rect 18874 3612 18880 3624
rect 18932 3612 18938 3664
rect 23937 3655 23995 3661
rect 23937 3621 23949 3655
rect 23983 3652 23995 3655
rect 25038 3652 25044 3664
rect 23983 3624 25044 3652
rect 23983 3621 23995 3624
rect 23937 3615 23995 3621
rect 25038 3612 25044 3624
rect 25096 3612 25102 3664
rect 29822 3612 29828 3664
rect 29880 3612 29886 3664
rect 32953 3655 33011 3661
rect 32953 3652 32965 3655
rect 30668 3624 32965 3652
rect 16482 3584 16488 3596
rect 6886 3556 16488 3584
rect 1210 3476 1216 3528
rect 1268 3516 1274 3528
rect 6886 3516 6914 3556
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 20346 3544 20352 3596
rect 20404 3584 20410 3596
rect 30668 3584 30696 3624
rect 32953 3621 32965 3624
rect 32999 3621 33011 3655
rect 32953 3615 33011 3621
rect 46385 3655 46443 3661
rect 46385 3621 46397 3655
rect 46431 3652 46443 3655
rect 47026 3652 47032 3664
rect 46431 3624 47032 3652
rect 46431 3621 46443 3624
rect 46385 3615 46443 3621
rect 47026 3612 47032 3624
rect 47084 3612 47090 3664
rect 33962 3584 33968 3596
rect 20404 3556 30696 3584
rect 31726 3556 33968 3584
rect 20404 3544 20410 3556
rect 23753 3519 23811 3525
rect 23753 3516 23765 3519
rect 1268 3488 6914 3516
rect 9646 3488 23765 3516
rect 1268 3476 1274 3488
rect 6362 3408 6368 3460
rect 6420 3448 6426 3460
rect 9646 3448 9674 3488
rect 23753 3485 23765 3488
rect 23799 3485 23811 3519
rect 23753 3479 23811 3485
rect 24397 3519 24455 3525
rect 24397 3485 24409 3519
rect 24443 3485 24455 3519
rect 24397 3479 24455 3485
rect 28537 3519 28595 3525
rect 28537 3485 28549 3519
rect 28583 3516 28595 3519
rect 28629 3519 28687 3525
rect 28629 3516 28641 3519
rect 28583 3488 28641 3516
rect 28583 3485 28595 3488
rect 28537 3479 28595 3485
rect 28629 3485 28641 3488
rect 28675 3485 28687 3519
rect 28629 3479 28687 3485
rect 24412 3448 24440 3479
rect 28994 3476 29000 3528
rect 29052 3516 29058 3528
rect 29181 3519 29239 3525
rect 29181 3516 29193 3519
rect 29052 3488 29193 3516
rect 29052 3476 29058 3488
rect 29181 3485 29193 3488
rect 29227 3485 29239 3519
rect 29181 3479 29239 3485
rect 29638 3476 29644 3528
rect 29696 3476 29702 3528
rect 30098 3476 30104 3528
rect 30156 3476 30162 3528
rect 30561 3519 30619 3525
rect 30561 3485 30573 3519
rect 30607 3516 30619 3519
rect 30653 3519 30711 3525
rect 30653 3516 30665 3519
rect 30607 3488 30665 3516
rect 30607 3485 30619 3488
rect 30561 3479 30619 3485
rect 30653 3485 30665 3488
rect 30699 3485 30711 3519
rect 30653 3479 30711 3485
rect 31294 3476 31300 3528
rect 31352 3476 31358 3528
rect 28166 3448 28172 3460
rect 6420 3420 9674 3448
rect 22066 3420 24440 3448
rect 24596 3420 28172 3448
rect 6420 3408 6426 3420
rect 1302 3340 1308 3392
rect 1360 3380 1366 3392
rect 14734 3380 14740 3392
rect 1360 3352 14740 3380
rect 1360 3340 1366 3352
rect 14734 3340 14740 3352
rect 14792 3340 14798 3392
rect 17218 3340 17224 3392
rect 17276 3380 17282 3392
rect 22066 3380 22094 3420
rect 24596 3389 24624 3420
rect 28166 3408 28172 3420
rect 28224 3408 28230 3460
rect 29822 3408 29828 3460
rect 29880 3448 29886 3460
rect 30742 3448 30748 3460
rect 29880 3420 30748 3448
rect 29880 3408 29886 3420
rect 30742 3408 30748 3420
rect 30800 3408 30806 3460
rect 17276 3352 22094 3380
rect 24581 3383 24639 3389
rect 17276 3340 17282 3352
rect 24581 3349 24593 3383
rect 24627 3349 24639 3383
rect 24581 3343 24639 3349
rect 27522 3340 27528 3392
rect 27580 3380 27586 3392
rect 28445 3383 28503 3389
rect 28445 3380 28457 3383
rect 27580 3352 28457 3380
rect 27580 3340 27586 3352
rect 28445 3349 28457 3352
rect 28491 3349 28503 3383
rect 28445 3343 28503 3349
rect 28813 3383 28871 3389
rect 28813 3349 28825 3383
rect 28859 3380 28871 3383
rect 29270 3380 29276 3392
rect 28859 3352 29276 3380
rect 28859 3349 28871 3352
rect 28813 3343 28871 3349
rect 29270 3340 29276 3352
rect 29328 3340 29334 3392
rect 29362 3340 29368 3392
rect 29420 3340 29426 3392
rect 30285 3383 30343 3389
rect 30285 3349 30297 3383
rect 30331 3380 30343 3383
rect 30374 3380 30380 3392
rect 30331 3352 30380 3380
rect 30331 3349 30343 3352
rect 30285 3343 30343 3349
rect 30374 3340 30380 3352
rect 30432 3340 30438 3392
rect 30466 3340 30472 3392
rect 30524 3340 30530 3392
rect 30834 3340 30840 3392
rect 30892 3340 30898 3392
rect 31481 3383 31539 3389
rect 31481 3349 31493 3383
rect 31527 3380 31539 3383
rect 31726 3380 31754 3556
rect 33962 3544 33968 3556
rect 34020 3544 34026 3596
rect 42610 3544 42616 3596
rect 42668 3584 42674 3596
rect 42668 3556 46980 3584
rect 42668 3544 42674 3556
rect 31846 3476 31852 3528
rect 31904 3476 31910 3528
rect 32306 3476 32312 3528
rect 32364 3516 32370 3528
rect 32493 3519 32551 3525
rect 32493 3516 32505 3519
rect 32364 3488 32505 3516
rect 32364 3476 32370 3488
rect 32493 3485 32505 3488
rect 32539 3485 32551 3519
rect 32493 3479 32551 3485
rect 33045 3519 33103 3525
rect 33045 3485 33057 3519
rect 33091 3516 33103 3519
rect 33137 3519 33195 3525
rect 33137 3516 33149 3519
rect 33091 3488 33149 3516
rect 33091 3485 33103 3488
rect 33045 3479 33103 3485
rect 33137 3485 33149 3488
rect 33183 3485 33195 3519
rect 33137 3479 33195 3485
rect 46109 3519 46167 3525
rect 46109 3485 46121 3519
rect 46155 3516 46167 3519
rect 46201 3519 46259 3525
rect 46201 3516 46213 3519
rect 46155 3488 46213 3516
rect 46155 3485 46167 3488
rect 46109 3479 46167 3485
rect 46201 3485 46213 3488
rect 46247 3485 46259 3519
rect 46201 3479 46259 3485
rect 46474 3476 46480 3528
rect 46532 3516 46538 3528
rect 46952 3525 46980 3556
rect 46753 3519 46811 3525
rect 46753 3516 46765 3519
rect 46532 3488 46765 3516
rect 46532 3476 46538 3488
rect 46753 3485 46765 3488
rect 46799 3485 46811 3519
rect 46753 3479 46811 3485
rect 46937 3519 46995 3525
rect 46937 3485 46949 3519
rect 46983 3485 46995 3519
rect 46937 3479 46995 3485
rect 34698 3448 34704 3460
rect 32692 3420 34704 3448
rect 31527 3352 31754 3380
rect 31527 3349 31539 3352
rect 31481 3343 31539 3349
rect 32030 3340 32036 3392
rect 32088 3340 32094 3392
rect 32692 3389 32720 3420
rect 34698 3408 34704 3420
rect 34756 3408 34762 3460
rect 32677 3383 32735 3389
rect 32677 3349 32689 3383
rect 32723 3349 32735 3383
rect 32677 3343 32735 3349
rect 33321 3383 33379 3389
rect 33321 3349 33333 3383
rect 33367 3380 33379 3383
rect 35066 3380 35072 3392
rect 33367 3352 35072 3380
rect 33367 3349 33379 3352
rect 33321 3343 33379 3349
rect 35066 3340 35072 3352
rect 35124 3340 35130 3392
rect 46658 3340 46664 3392
rect 46716 3340 46722 3392
rect 47118 3340 47124 3392
rect 47176 3340 47182 3392
rect 1104 3290 47840 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 39010 3290
rect 39062 3238 39074 3290
rect 39126 3238 39138 3290
rect 39190 3238 39202 3290
rect 39254 3238 39266 3290
rect 39318 3238 45010 3290
rect 45062 3238 45074 3290
rect 45126 3238 45138 3290
rect 45190 3238 45202 3290
rect 45254 3238 45266 3290
rect 45318 3238 47840 3290
rect 1104 3216 47840 3238
rect 5994 3136 6000 3188
rect 6052 3176 6058 3188
rect 6052 3148 13768 3176
rect 6052 3136 6058 3148
rect 8662 3000 8668 3052
rect 8720 3040 8726 3052
rect 13740 3040 13768 3148
rect 13814 3136 13820 3188
rect 13872 3176 13878 3188
rect 14093 3179 14151 3185
rect 14093 3176 14105 3179
rect 13872 3148 14105 3176
rect 13872 3136 13878 3148
rect 14093 3145 14105 3148
rect 14139 3145 14151 3179
rect 14093 3139 14151 3145
rect 17770 3136 17776 3188
rect 17828 3136 17834 3188
rect 18141 3179 18199 3185
rect 18141 3145 18153 3179
rect 18187 3176 18199 3179
rect 45554 3176 45560 3188
rect 18187 3148 26188 3176
rect 18187 3145 18199 3148
rect 18141 3139 18199 3145
rect 14185 3111 14243 3117
rect 14185 3077 14197 3111
rect 14231 3108 14243 3111
rect 14369 3111 14427 3117
rect 14369 3108 14381 3111
rect 14231 3080 14381 3108
rect 14231 3077 14243 3080
rect 14185 3071 14243 3077
rect 14369 3077 14381 3080
rect 14415 3077 14427 3111
rect 14369 3071 14427 3077
rect 14550 3068 14556 3120
rect 14608 3068 14614 3120
rect 14734 3068 14740 3120
rect 14792 3108 14798 3120
rect 14792 3080 19748 3108
rect 14792 3068 14798 3080
rect 17218 3040 17224 3052
rect 8720 3012 12434 3040
rect 13740 3012 17224 3040
rect 8720 3000 8726 3012
rect 12406 2972 12434 3012
rect 17218 3000 17224 3012
rect 17276 3000 17282 3052
rect 17865 3043 17923 3049
rect 17865 3009 17877 3043
rect 17911 3040 17923 3043
rect 18049 3043 18107 3049
rect 18049 3040 18061 3043
rect 17911 3012 18061 3040
rect 17911 3009 17923 3012
rect 17865 3003 17923 3009
rect 18049 3009 18061 3012
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 19429 3043 19487 3049
rect 19429 3009 19441 3043
rect 19475 3040 19487 3043
rect 19613 3043 19671 3049
rect 19613 3040 19625 3043
rect 19475 3012 19625 3040
rect 19475 3009 19487 3012
rect 19429 3003 19487 3009
rect 19613 3009 19625 3012
rect 19659 3009 19671 3043
rect 19613 3003 19671 3009
rect 19337 2975 19395 2981
rect 19337 2972 19349 2975
rect 12406 2944 19349 2972
rect 19337 2941 19349 2944
rect 19383 2941 19395 2975
rect 19720 2972 19748 3080
rect 20806 3000 20812 3052
rect 20864 3040 20870 3052
rect 21913 3043 21971 3049
rect 21913 3040 21925 3043
rect 20864 3012 21925 3040
rect 20864 3000 20870 3012
rect 21913 3009 21925 3012
rect 21959 3009 21971 3043
rect 24765 3043 24823 3049
rect 24765 3040 24777 3043
rect 21913 3003 21971 3009
rect 22066 3012 24777 3040
rect 22066 2972 22094 3012
rect 24765 3009 24777 3012
rect 24811 3009 24823 3043
rect 24765 3003 24823 3009
rect 25961 3043 26019 3049
rect 25961 3009 25973 3043
rect 26007 3040 26019 3043
rect 26053 3043 26111 3049
rect 26053 3040 26065 3043
rect 26007 3012 26065 3040
rect 26007 3009 26019 3012
rect 25961 3003 26019 3009
rect 26053 3009 26065 3012
rect 26099 3009 26111 3043
rect 26160 3040 26188 3148
rect 26436 3148 45560 3176
rect 26436 3040 26464 3148
rect 45554 3136 45560 3148
rect 45612 3136 45618 3188
rect 47302 3136 47308 3188
rect 47360 3136 47366 3188
rect 27798 3068 27804 3120
rect 27856 3108 27862 3120
rect 27856 3080 28304 3108
rect 27856 3068 27862 3080
rect 26160 3012 26464 3040
rect 28077 3043 28135 3049
rect 26053 3003 26111 3009
rect 28077 3009 28089 3043
rect 28123 3040 28135 3043
rect 28169 3043 28227 3049
rect 28169 3040 28181 3043
rect 28123 3012 28181 3040
rect 28123 3009 28135 3012
rect 28077 3003 28135 3009
rect 28169 3009 28181 3012
rect 28215 3009 28227 3043
rect 28276 3040 28304 3080
rect 29362 3068 29368 3120
rect 29420 3108 29426 3120
rect 32674 3108 32680 3120
rect 29420 3080 32680 3108
rect 29420 3068 29426 3080
rect 32674 3068 32680 3080
rect 32732 3068 32738 3120
rect 43438 3108 43444 3120
rect 36556 3080 43444 3108
rect 29917 3043 29975 3049
rect 29917 3040 29929 3043
rect 28276 3012 29929 3040
rect 28169 3003 28227 3009
rect 29917 3009 29929 3012
rect 29963 3009 29975 3043
rect 29917 3003 29975 3009
rect 30650 3000 30656 3052
rect 30708 3000 30714 3052
rect 31110 3000 31116 3052
rect 31168 3000 31174 3052
rect 32030 3000 32036 3052
rect 32088 3040 32094 3052
rect 36556 3049 36584 3080
rect 43438 3068 43444 3080
rect 43496 3068 43502 3120
rect 33689 3043 33747 3049
rect 33689 3040 33701 3043
rect 32088 3012 33701 3040
rect 32088 3000 32094 3012
rect 33689 3009 33701 3012
rect 33735 3009 33747 3043
rect 33689 3003 33747 3009
rect 36541 3043 36599 3049
rect 36541 3009 36553 3043
rect 36587 3009 36599 3043
rect 36541 3003 36599 3009
rect 38838 3000 38844 3052
rect 38896 3000 38902 3052
rect 41598 3000 41604 3052
rect 41656 3040 41662 3052
rect 46385 3043 46443 3049
rect 46385 3040 46397 3043
rect 41656 3012 46397 3040
rect 41656 3000 41662 3012
rect 46385 3009 46397 3012
rect 46431 3009 46443 3043
rect 46385 3003 46443 3009
rect 46658 3000 46664 3052
rect 46716 3040 46722 3052
rect 46753 3043 46811 3049
rect 46753 3040 46765 3043
rect 46716 3012 46765 3040
rect 46716 3000 46722 3012
rect 46753 3009 46765 3012
rect 46799 3009 46811 3043
rect 46753 3003 46811 3009
rect 46842 3000 46848 3052
rect 46900 3040 46906 3052
rect 47121 3043 47179 3049
rect 47121 3040 47133 3043
rect 46900 3012 47133 3040
rect 46900 3000 46906 3012
rect 47121 3009 47133 3012
rect 47167 3009 47179 3043
rect 47121 3003 47179 3009
rect 19720 2944 22094 2972
rect 19337 2935 19395 2941
rect 24670 2932 24676 2984
rect 24728 2972 24734 2984
rect 25869 2975 25927 2981
rect 25869 2972 25881 2975
rect 24728 2944 25881 2972
rect 24728 2932 24734 2944
rect 25869 2941 25881 2944
rect 25915 2941 25927 2975
rect 25869 2935 25927 2941
rect 26160 2944 29868 2972
rect 7558 2864 7564 2916
rect 7616 2904 7622 2916
rect 19150 2904 19156 2916
rect 7616 2876 19156 2904
rect 7616 2864 7622 2876
rect 19150 2864 19156 2876
rect 19208 2864 19214 2916
rect 19797 2907 19855 2913
rect 19797 2873 19809 2907
rect 19843 2904 19855 2907
rect 26160 2904 26188 2944
rect 19843 2876 26188 2904
rect 26237 2907 26295 2913
rect 19843 2873 19855 2876
rect 19797 2867 19855 2873
rect 26237 2873 26249 2907
rect 26283 2904 26295 2907
rect 27798 2904 27804 2916
rect 26283 2876 27804 2904
rect 26283 2873 26295 2876
rect 26237 2867 26295 2873
rect 27798 2864 27804 2876
rect 27856 2864 27862 2916
rect 28353 2907 28411 2913
rect 27908 2876 28304 2904
rect 21818 2796 21824 2848
rect 21876 2836 21882 2848
rect 22097 2839 22155 2845
rect 22097 2836 22109 2839
rect 21876 2808 22109 2836
rect 21876 2796 21882 2808
rect 22097 2805 22109 2808
rect 22143 2805 22155 2839
rect 22097 2799 22155 2805
rect 24949 2839 25007 2845
rect 24949 2805 24961 2839
rect 24995 2836 25007 2839
rect 27908 2836 27936 2876
rect 24995 2808 27936 2836
rect 24995 2805 25007 2808
rect 24949 2799 25007 2805
rect 27982 2796 27988 2848
rect 28040 2796 28046 2848
rect 28276 2836 28304 2876
rect 28353 2873 28365 2907
rect 28399 2904 28411 2907
rect 29730 2904 29736 2916
rect 28399 2876 29736 2904
rect 28399 2873 28411 2876
rect 28353 2867 28411 2873
rect 29730 2864 29736 2876
rect 29788 2864 29794 2916
rect 29840 2904 29868 2944
rect 45646 2904 45652 2916
rect 29840 2876 45652 2904
rect 45646 2864 45652 2876
rect 45704 2864 45710 2916
rect 46569 2907 46627 2913
rect 46569 2873 46581 2907
rect 46615 2904 46627 2907
rect 47946 2904 47952 2916
rect 46615 2876 47952 2904
rect 46615 2873 46627 2876
rect 46569 2867 46627 2873
rect 47946 2864 47952 2876
rect 48004 2864 48010 2916
rect 28534 2836 28540 2848
rect 28276 2808 28540 2836
rect 28534 2796 28540 2808
rect 28592 2796 28598 2848
rect 29178 2796 29184 2848
rect 29236 2836 29242 2848
rect 30101 2839 30159 2845
rect 30101 2836 30113 2839
rect 29236 2808 30113 2836
rect 29236 2796 29242 2808
rect 30101 2805 30113 2808
rect 30147 2805 30159 2839
rect 30101 2799 30159 2805
rect 30282 2796 30288 2848
rect 30340 2836 30346 2848
rect 30837 2839 30895 2845
rect 30837 2836 30849 2839
rect 30340 2808 30849 2836
rect 30340 2796 30346 2808
rect 30837 2805 30849 2808
rect 30883 2805 30895 2839
rect 30837 2799 30895 2805
rect 31018 2796 31024 2848
rect 31076 2836 31082 2848
rect 31297 2839 31355 2845
rect 31297 2836 31309 2839
rect 31076 2808 31309 2836
rect 31076 2796 31082 2808
rect 31297 2805 31309 2808
rect 31343 2805 31355 2839
rect 31297 2799 31355 2805
rect 33594 2796 33600 2848
rect 33652 2836 33658 2848
rect 33873 2839 33931 2845
rect 33873 2836 33885 2839
rect 33652 2808 33885 2836
rect 33652 2796 33658 2808
rect 33873 2805 33885 2808
rect 33919 2805 33931 2839
rect 33873 2799 33931 2805
rect 36262 2796 36268 2848
rect 36320 2836 36326 2848
rect 36357 2839 36415 2845
rect 36357 2836 36369 2839
rect 36320 2808 36369 2836
rect 36320 2796 36326 2808
rect 36357 2805 36369 2808
rect 36403 2805 36415 2839
rect 36357 2799 36415 2805
rect 38746 2796 38752 2848
rect 38804 2836 38810 2848
rect 39025 2839 39083 2845
rect 39025 2836 39037 2839
rect 38804 2808 39037 2836
rect 38804 2796 38810 2808
rect 39025 2805 39037 2808
rect 39071 2805 39083 2839
rect 39025 2799 39083 2805
rect 46934 2796 46940 2848
rect 46992 2796 46998 2848
rect 1104 2746 47840 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 37950 2746
rect 38002 2694 38014 2746
rect 38066 2694 38078 2746
rect 38130 2694 38142 2746
rect 38194 2694 38206 2746
rect 38258 2694 43950 2746
rect 44002 2694 44014 2746
rect 44066 2694 44078 2746
rect 44130 2694 44142 2746
rect 44194 2694 44206 2746
rect 44258 2694 47840 2746
rect 1104 2672 47840 2694
rect 15838 2592 15844 2644
rect 15896 2632 15902 2644
rect 20622 2632 20628 2644
rect 15896 2604 20628 2632
rect 15896 2592 15902 2604
rect 20622 2592 20628 2604
rect 20680 2592 20686 2644
rect 25590 2632 25596 2644
rect 20732 2604 25596 2632
rect 15654 2524 15660 2576
rect 15712 2564 15718 2576
rect 20732 2564 20760 2604
rect 25590 2592 25596 2604
rect 25648 2592 25654 2644
rect 25700 2604 28304 2632
rect 15712 2536 20760 2564
rect 15712 2524 15718 2536
rect 22002 2524 22008 2576
rect 22060 2564 22066 2576
rect 25700 2564 25728 2604
rect 22060 2536 24532 2564
rect 22060 2524 22066 2536
rect 18984 2468 21404 2496
rect 16022 2388 16028 2440
rect 16080 2428 16086 2440
rect 18984 2428 19012 2468
rect 16080 2400 19012 2428
rect 16080 2388 16086 2400
rect 20622 2388 20628 2440
rect 20680 2388 20686 2440
rect 20714 2388 20720 2440
rect 20772 2428 20778 2440
rect 21376 2437 21404 2468
rect 23382 2456 23388 2508
rect 23440 2496 23446 2508
rect 23440 2468 23980 2496
rect 23440 2456 23446 2468
rect 20993 2431 21051 2437
rect 20993 2428 21005 2431
rect 20772 2400 21005 2428
rect 20772 2388 20778 2400
rect 20993 2397 21005 2400
rect 21039 2397 21051 2431
rect 20993 2391 21051 2397
rect 21361 2431 21419 2437
rect 21361 2397 21373 2431
rect 21407 2397 21419 2431
rect 21361 2391 21419 2397
rect 22094 2388 22100 2440
rect 22152 2388 22158 2440
rect 22462 2388 22468 2440
rect 22520 2388 22526 2440
rect 22830 2388 22836 2440
rect 22888 2388 22894 2440
rect 23198 2388 23204 2440
rect 23256 2388 23262 2440
rect 23566 2388 23572 2440
rect 23624 2388 23630 2440
rect 23952 2437 23980 2468
rect 24504 2437 24532 2536
rect 24596 2536 25728 2564
rect 23937 2431 23995 2437
rect 23937 2397 23949 2431
rect 23983 2397 23995 2431
rect 23937 2391 23995 2397
rect 24489 2431 24547 2437
rect 24489 2397 24501 2431
rect 24535 2397 24547 2431
rect 24489 2391 24547 2397
rect 10594 2320 10600 2372
rect 10652 2360 10658 2372
rect 24596 2360 24624 2536
rect 27890 2524 27896 2576
rect 27948 2524 27954 2576
rect 28166 2524 28172 2576
rect 28224 2524 28230 2576
rect 28276 2564 28304 2604
rect 28350 2592 28356 2644
rect 28408 2632 28414 2644
rect 28629 2635 28687 2641
rect 28629 2632 28641 2635
rect 28408 2604 28641 2632
rect 28408 2592 28414 2604
rect 28629 2601 28641 2604
rect 28675 2601 28687 2635
rect 29917 2635 29975 2641
rect 29917 2632 29929 2635
rect 28629 2595 28687 2601
rect 28736 2604 29929 2632
rect 28736 2564 28764 2604
rect 29917 2601 29929 2604
rect 29963 2601 29975 2635
rect 29917 2595 29975 2601
rect 30282 2592 30288 2644
rect 30340 2632 30346 2644
rect 31205 2635 31263 2641
rect 31205 2632 31217 2635
rect 30340 2604 31217 2632
rect 30340 2592 30346 2604
rect 31205 2601 31217 2604
rect 31251 2601 31263 2635
rect 31205 2595 31263 2601
rect 32858 2592 32864 2644
rect 32916 2632 32922 2644
rect 33781 2635 33839 2641
rect 33781 2632 33793 2635
rect 32916 2604 33793 2632
rect 32916 2592 32922 2604
rect 33781 2601 33793 2604
rect 33827 2601 33839 2635
rect 33781 2595 33839 2601
rect 35526 2592 35532 2644
rect 35584 2632 35590 2644
rect 36357 2635 36415 2641
rect 36357 2632 36369 2635
rect 35584 2604 36369 2632
rect 35584 2592 35590 2604
rect 36357 2601 36369 2604
rect 36403 2601 36415 2635
rect 36357 2595 36415 2601
rect 37642 2592 37648 2644
rect 37700 2632 37706 2644
rect 38565 2635 38623 2641
rect 38565 2632 38577 2635
rect 37700 2604 38577 2632
rect 37700 2592 37706 2604
rect 38565 2601 38577 2604
rect 38611 2601 38623 2635
rect 38565 2595 38623 2601
rect 47302 2592 47308 2644
rect 47360 2592 47366 2644
rect 28276 2536 28764 2564
rect 28810 2524 28816 2576
rect 28868 2564 28874 2576
rect 29641 2567 29699 2573
rect 29641 2564 29653 2567
rect 28868 2536 29653 2564
rect 28868 2524 28874 2536
rect 29641 2533 29653 2536
rect 29687 2533 29699 2567
rect 29641 2527 29699 2533
rect 29822 2524 29828 2576
rect 29880 2564 29886 2576
rect 30098 2564 30104 2576
rect 29880 2536 30104 2564
rect 29880 2524 29886 2536
rect 30098 2524 30104 2536
rect 30156 2524 30162 2576
rect 30374 2524 30380 2576
rect 30432 2564 30438 2576
rect 30432 2536 30604 2564
rect 30432 2524 30438 2536
rect 26878 2456 26884 2508
rect 26936 2496 26942 2508
rect 28184 2496 28212 2524
rect 26936 2468 27108 2496
rect 26936 2456 26942 2468
rect 24762 2388 24768 2440
rect 24820 2428 24826 2440
rect 24857 2431 24915 2437
rect 24857 2428 24869 2431
rect 24820 2400 24869 2428
rect 24820 2388 24826 2400
rect 24857 2397 24869 2400
rect 24903 2397 24915 2431
rect 24857 2391 24915 2397
rect 25038 2388 25044 2440
rect 25096 2388 25102 2440
rect 25222 2388 25228 2440
rect 25280 2388 25286 2440
rect 25590 2388 25596 2440
rect 25648 2388 25654 2440
rect 25958 2388 25964 2440
rect 26016 2388 26022 2440
rect 26326 2388 26332 2440
rect 26384 2388 26390 2440
rect 26602 2388 26608 2440
rect 26660 2428 26666 2440
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26660 2400 26985 2428
rect 26660 2388 26666 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 27080 2428 27108 2468
rect 28092 2468 28212 2496
rect 28092 2437 28120 2468
rect 28258 2456 28264 2508
rect 28316 2496 28322 2508
rect 30576 2496 30604 2536
rect 30650 2524 30656 2576
rect 30708 2564 30714 2576
rect 31481 2567 31539 2573
rect 31481 2564 31493 2567
rect 30708 2536 31493 2564
rect 30708 2524 30714 2536
rect 31481 2533 31493 2536
rect 31527 2533 31539 2567
rect 31481 2527 31539 2533
rect 32324 2536 32536 2564
rect 32324 2496 32352 2536
rect 28316 2468 30420 2496
rect 30576 2468 32352 2496
rect 32508 2496 32536 2536
rect 32582 2524 32588 2576
rect 32640 2564 32646 2576
rect 33413 2567 33471 2573
rect 33413 2564 33425 2567
rect 32640 2536 33425 2564
rect 32640 2524 32646 2536
rect 33413 2533 33425 2536
rect 33459 2533 33471 2567
rect 33413 2527 33471 2533
rect 34330 2524 34336 2576
rect 34388 2564 34394 2576
rect 35253 2567 35311 2573
rect 35253 2564 35265 2567
rect 34388 2536 35265 2564
rect 34388 2524 34394 2536
rect 35253 2533 35265 2536
rect 35299 2533 35311 2567
rect 35253 2527 35311 2533
rect 35802 2524 35808 2576
rect 35860 2564 35866 2576
rect 36633 2567 36691 2573
rect 36633 2564 36645 2567
rect 35860 2536 36645 2564
rect 35860 2524 35866 2536
rect 36633 2533 36645 2536
rect 36679 2533 36691 2567
rect 36633 2527 36691 2533
rect 36906 2524 36912 2576
rect 36964 2564 36970 2576
rect 37829 2567 37887 2573
rect 37829 2564 37841 2567
rect 36964 2536 37841 2564
rect 36964 2524 36970 2536
rect 37829 2533 37841 2536
rect 37875 2533 37887 2567
rect 37829 2527 37887 2533
rect 38378 2524 38384 2576
rect 38436 2564 38442 2576
rect 39301 2567 39359 2573
rect 39301 2564 39313 2567
rect 38436 2536 39313 2564
rect 38436 2524 38442 2536
rect 39301 2533 39313 2536
rect 39347 2533 39359 2567
rect 39301 2527 39359 2533
rect 39482 2524 39488 2576
rect 39540 2564 39546 2576
rect 40405 2567 40463 2573
rect 40405 2564 40417 2567
rect 39540 2536 40417 2564
rect 39540 2524 39546 2536
rect 40405 2533 40417 2536
rect 40451 2533 40463 2567
rect 40405 2527 40463 2533
rect 32508 2468 33272 2496
rect 28316 2456 28322 2468
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 27080 2400 27353 2428
rect 26973 2391 27031 2397
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 27341 2391 27399 2397
rect 27709 2431 27767 2437
rect 27709 2397 27721 2431
rect 27755 2397 27767 2431
rect 27709 2391 27767 2397
rect 28077 2431 28135 2437
rect 28077 2397 28089 2431
rect 28123 2397 28135 2431
rect 28077 2391 28135 2397
rect 28445 2431 28503 2437
rect 28445 2397 28457 2431
rect 28491 2428 28503 2431
rect 28534 2428 28540 2440
rect 28491 2400 28540 2428
rect 28491 2397 28503 2400
rect 28445 2391 28503 2397
rect 10652 2332 24624 2360
rect 25056 2360 25084 2388
rect 27724 2360 27752 2391
rect 28534 2388 28540 2400
rect 28592 2388 28598 2440
rect 28626 2388 28632 2440
rect 28684 2428 28690 2440
rect 28813 2431 28871 2437
rect 28813 2428 28825 2431
rect 28684 2400 28825 2428
rect 28684 2388 28690 2400
rect 28813 2397 28825 2400
rect 28859 2397 28871 2431
rect 28813 2391 28871 2397
rect 29825 2431 29883 2437
rect 29825 2397 29837 2431
rect 29871 2428 29883 2431
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29871 2400 29929 2428
rect 29871 2397 29883 2400
rect 29825 2391 29883 2397
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 30193 2431 30251 2437
rect 30193 2397 30205 2431
rect 30239 2428 30251 2431
rect 30285 2431 30343 2437
rect 30285 2428 30297 2431
rect 30239 2400 30297 2428
rect 30239 2397 30251 2400
rect 30193 2391 30251 2397
rect 30285 2397 30297 2400
rect 30331 2397 30343 2431
rect 30392 2428 30420 2468
rect 30837 2431 30895 2437
rect 30837 2428 30849 2431
rect 30392 2400 30849 2428
rect 30285 2391 30343 2397
rect 30837 2397 30849 2400
rect 30883 2428 30895 2431
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30883 2400 31033 2428
rect 30883 2397 30895 2400
rect 30837 2391 30895 2397
rect 31021 2397 31033 2400
rect 31067 2397 31079 2431
rect 31021 2391 31079 2397
rect 31665 2431 31723 2437
rect 31665 2397 31677 2431
rect 31711 2428 31723 2431
rect 31757 2431 31815 2437
rect 31757 2428 31769 2431
rect 31711 2400 31769 2428
rect 31711 2397 31723 2400
rect 31665 2391 31723 2397
rect 31757 2397 31769 2400
rect 31803 2397 31815 2431
rect 31757 2391 31815 2397
rect 32122 2388 32128 2440
rect 32180 2388 32186 2440
rect 32493 2431 32551 2437
rect 32493 2397 32505 2431
rect 32539 2428 32551 2431
rect 32674 2428 32680 2440
rect 32539 2400 32680 2428
rect 32539 2397 32551 2400
rect 32493 2391 32551 2397
rect 32674 2388 32680 2400
rect 32732 2388 32738 2440
rect 32766 2388 32772 2440
rect 32824 2428 32830 2440
rect 33244 2437 33272 2468
rect 36998 2456 37004 2508
rect 37056 2496 37062 2508
rect 40310 2496 40316 2508
rect 37056 2468 37872 2496
rect 37056 2456 37062 2468
rect 32861 2431 32919 2437
rect 32861 2428 32873 2431
rect 32824 2400 32873 2428
rect 32824 2388 32830 2400
rect 32861 2397 32873 2400
rect 32907 2397 32919 2431
rect 32861 2391 32919 2397
rect 33229 2431 33287 2437
rect 33229 2397 33241 2431
rect 33275 2397 33287 2431
rect 33229 2391 33287 2397
rect 33502 2388 33508 2440
rect 33560 2428 33566 2440
rect 33597 2431 33655 2437
rect 33597 2428 33609 2431
rect 33560 2400 33609 2428
rect 33560 2388 33566 2400
rect 33597 2397 33609 2400
rect 33643 2397 33655 2431
rect 33597 2391 33655 2397
rect 33962 2388 33968 2440
rect 34020 2388 34026 2440
rect 34698 2388 34704 2440
rect 34756 2388 34762 2440
rect 35066 2388 35072 2440
rect 35124 2388 35130 2440
rect 35434 2388 35440 2440
rect 35492 2388 35498 2440
rect 35618 2388 35624 2440
rect 35676 2428 35682 2440
rect 35805 2431 35863 2437
rect 35805 2428 35817 2431
rect 35676 2400 35817 2428
rect 35676 2388 35682 2400
rect 35805 2397 35817 2400
rect 35851 2397 35863 2431
rect 35805 2391 35863 2397
rect 36170 2388 36176 2440
rect 36228 2388 36234 2440
rect 36814 2388 36820 2440
rect 36872 2388 36878 2440
rect 37553 2431 37611 2437
rect 37553 2397 37565 2431
rect 37599 2397 37611 2431
rect 37553 2391 37611 2397
rect 37670 2431 37728 2437
rect 37670 2397 37682 2431
rect 37716 2428 37728 2431
rect 37844 2428 37872 2468
rect 37716 2400 37872 2428
rect 37936 2468 40316 2496
rect 37716 2397 37728 2400
rect 37670 2391 37728 2397
rect 25056 2332 27752 2360
rect 10652 2320 10658 2332
rect 29546 2320 29552 2372
rect 29604 2360 29610 2372
rect 29604 2332 30512 2360
rect 29604 2320 29610 2332
rect 20714 2252 20720 2304
rect 20772 2292 20778 2304
rect 20809 2295 20867 2301
rect 20809 2292 20821 2295
rect 20772 2264 20821 2292
rect 20772 2252 20778 2264
rect 20809 2261 20821 2264
rect 20855 2261 20867 2295
rect 20809 2255 20867 2261
rect 20898 2252 20904 2304
rect 20956 2292 20962 2304
rect 21177 2295 21235 2301
rect 21177 2292 21189 2295
rect 20956 2264 21189 2292
rect 20956 2252 20962 2264
rect 21177 2261 21189 2264
rect 21223 2261 21235 2295
rect 21177 2255 21235 2261
rect 21450 2252 21456 2304
rect 21508 2292 21514 2304
rect 21545 2295 21603 2301
rect 21545 2292 21557 2295
rect 21508 2264 21557 2292
rect 21508 2252 21514 2264
rect 21545 2261 21557 2264
rect 21591 2261 21603 2295
rect 21545 2255 21603 2261
rect 22186 2252 22192 2304
rect 22244 2292 22250 2304
rect 22281 2295 22339 2301
rect 22281 2292 22293 2295
rect 22244 2264 22293 2292
rect 22244 2252 22250 2264
rect 22281 2261 22293 2264
rect 22327 2261 22339 2295
rect 22281 2255 22339 2261
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22649 2295 22707 2301
rect 22649 2292 22661 2295
rect 22612 2264 22661 2292
rect 22612 2252 22618 2264
rect 22649 2261 22661 2264
rect 22695 2261 22707 2295
rect 22649 2255 22707 2261
rect 22922 2252 22928 2304
rect 22980 2292 22986 2304
rect 23017 2295 23075 2301
rect 23017 2292 23029 2295
rect 22980 2264 23029 2292
rect 22980 2252 22986 2264
rect 23017 2261 23029 2264
rect 23063 2261 23075 2295
rect 23017 2255 23075 2261
rect 23290 2252 23296 2304
rect 23348 2292 23354 2304
rect 23385 2295 23443 2301
rect 23385 2292 23397 2295
rect 23348 2264 23397 2292
rect 23348 2252 23354 2264
rect 23385 2261 23397 2264
rect 23431 2261 23443 2295
rect 23385 2255 23443 2261
rect 23658 2252 23664 2304
rect 23716 2292 23722 2304
rect 23753 2295 23811 2301
rect 23753 2292 23765 2295
rect 23716 2264 23765 2292
rect 23716 2252 23722 2264
rect 23753 2261 23765 2264
rect 23799 2261 23811 2295
rect 23753 2255 23811 2261
rect 24026 2252 24032 2304
rect 24084 2292 24090 2304
rect 24121 2295 24179 2301
rect 24121 2292 24133 2295
rect 24084 2264 24133 2292
rect 24084 2252 24090 2264
rect 24121 2261 24133 2264
rect 24167 2261 24179 2295
rect 24121 2255 24179 2261
rect 24394 2252 24400 2304
rect 24452 2292 24458 2304
rect 24673 2295 24731 2301
rect 24673 2292 24685 2295
rect 24452 2264 24685 2292
rect 24452 2252 24458 2264
rect 24673 2261 24685 2264
rect 24719 2261 24731 2295
rect 24673 2255 24731 2261
rect 25038 2252 25044 2304
rect 25096 2252 25102 2304
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 25409 2295 25467 2301
rect 25409 2292 25421 2295
rect 25188 2264 25421 2292
rect 25188 2252 25194 2264
rect 25409 2261 25421 2264
rect 25455 2261 25467 2295
rect 25409 2255 25467 2261
rect 25498 2252 25504 2304
rect 25556 2292 25562 2304
rect 25777 2295 25835 2301
rect 25777 2292 25789 2295
rect 25556 2264 25789 2292
rect 25556 2252 25562 2264
rect 25777 2261 25789 2264
rect 25823 2261 25835 2295
rect 25777 2255 25835 2261
rect 25866 2252 25872 2304
rect 25924 2292 25930 2304
rect 26145 2295 26203 2301
rect 26145 2292 26157 2295
rect 25924 2264 26157 2292
rect 25924 2252 25930 2264
rect 26145 2261 26157 2264
rect 26191 2261 26203 2295
rect 26145 2255 26203 2261
rect 26234 2252 26240 2304
rect 26292 2292 26298 2304
rect 26513 2295 26571 2301
rect 26513 2292 26525 2295
rect 26292 2264 26525 2292
rect 26292 2252 26298 2264
rect 26513 2261 26525 2264
rect 26559 2261 26571 2295
rect 26513 2255 26571 2261
rect 26602 2252 26608 2304
rect 26660 2292 26666 2304
rect 27157 2295 27215 2301
rect 27157 2292 27169 2295
rect 26660 2264 27169 2292
rect 26660 2252 26666 2264
rect 27157 2261 27169 2264
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 27338 2252 27344 2304
rect 27396 2292 27402 2304
rect 27525 2295 27583 2301
rect 27525 2292 27537 2295
rect 27396 2264 27537 2292
rect 27396 2252 27402 2264
rect 27525 2261 27537 2264
rect 27571 2261 27583 2295
rect 27525 2255 27583 2261
rect 27706 2252 27712 2304
rect 27764 2292 27770 2304
rect 28261 2295 28319 2301
rect 28261 2292 28273 2295
rect 27764 2264 28273 2292
rect 27764 2252 27770 2264
rect 28261 2261 28273 2264
rect 28307 2261 28319 2295
rect 28261 2255 28319 2261
rect 28902 2252 28908 2304
rect 28960 2292 28966 2304
rect 28997 2295 29055 2301
rect 28997 2292 29009 2295
rect 28960 2264 29009 2292
rect 28960 2252 28966 2264
rect 28997 2261 29009 2264
rect 29043 2261 29055 2295
rect 28997 2255 29055 2261
rect 30098 2252 30104 2304
rect 30156 2252 30162 2304
rect 30484 2301 30512 2332
rect 31386 2320 31392 2372
rect 31444 2360 31450 2372
rect 31444 2332 32352 2360
rect 31444 2320 31450 2332
rect 30469 2295 30527 2301
rect 30469 2261 30481 2295
rect 30515 2261 30527 2295
rect 30469 2255 30527 2261
rect 30558 2252 30564 2304
rect 30616 2292 30622 2304
rect 32324 2301 32352 2332
rect 32398 2320 32404 2372
rect 32456 2360 32462 2372
rect 32456 2332 33088 2360
rect 32456 2320 32462 2332
rect 31757 2295 31815 2301
rect 31757 2292 31769 2295
rect 30616 2264 31769 2292
rect 30616 2252 30622 2264
rect 31757 2261 31769 2264
rect 31803 2261 31815 2295
rect 31757 2255 31815 2261
rect 32309 2295 32367 2301
rect 32309 2261 32321 2295
rect 32355 2261 32367 2295
rect 32309 2255 32367 2261
rect 32674 2252 32680 2304
rect 32732 2252 32738 2304
rect 33060 2301 33088 2332
rect 35158 2320 35164 2372
rect 35216 2360 35222 2372
rect 37568 2360 37596 2391
rect 37936 2360 37964 2468
rect 40310 2456 40316 2468
rect 40368 2456 40374 2508
rect 40494 2456 40500 2508
rect 40552 2496 40558 2508
rect 40552 2468 41414 2496
rect 40552 2456 40558 2468
rect 38010 2388 38016 2440
rect 38068 2388 38074 2440
rect 38102 2388 38108 2440
rect 38160 2428 38166 2440
rect 38381 2431 38439 2437
rect 38381 2428 38393 2431
rect 38160 2400 38393 2428
rect 38160 2388 38166 2400
rect 38381 2397 38393 2400
rect 38427 2397 38439 2431
rect 38381 2391 38439 2397
rect 38470 2388 38476 2440
rect 38528 2428 38534 2440
rect 38749 2431 38807 2437
rect 38749 2428 38761 2431
rect 38528 2400 38761 2428
rect 38528 2388 38534 2400
rect 38749 2397 38761 2400
rect 38795 2397 38807 2431
rect 38749 2391 38807 2397
rect 38838 2388 38844 2440
rect 38896 2428 38902 2440
rect 39117 2431 39175 2437
rect 39117 2428 39129 2431
rect 38896 2400 39129 2428
rect 38896 2388 38902 2400
rect 39117 2397 39129 2400
rect 39163 2397 39175 2431
rect 39117 2391 39175 2397
rect 39206 2388 39212 2440
rect 39264 2428 39270 2440
rect 39853 2431 39911 2437
rect 39853 2428 39865 2431
rect 39264 2400 39865 2428
rect 39264 2388 39270 2400
rect 39853 2397 39865 2400
rect 39899 2397 39911 2431
rect 39853 2391 39911 2397
rect 40034 2388 40040 2440
rect 40092 2428 40098 2440
rect 40221 2431 40279 2437
rect 40221 2428 40233 2431
rect 40092 2400 40233 2428
rect 40092 2388 40098 2400
rect 40221 2397 40233 2400
rect 40267 2397 40279 2431
rect 41386 2428 41414 2468
rect 42794 2456 42800 2508
rect 42852 2496 42858 2508
rect 42852 2468 46060 2496
rect 42852 2456 42858 2468
rect 46032 2437 46060 2468
rect 46198 2456 46204 2508
rect 46256 2496 46262 2508
rect 46256 2468 46796 2496
rect 46256 2456 46262 2468
rect 45649 2431 45707 2437
rect 45649 2428 45661 2431
rect 41386 2400 45661 2428
rect 40221 2391 40279 2397
rect 45649 2397 45661 2400
rect 45695 2397 45707 2431
rect 45649 2391 45707 2397
rect 46017 2431 46075 2437
rect 46017 2397 46029 2431
rect 46063 2397 46075 2431
rect 46017 2391 46075 2397
rect 46382 2388 46388 2440
rect 46440 2388 46446 2440
rect 46768 2437 46796 2468
rect 46753 2431 46811 2437
rect 46753 2397 46765 2431
rect 46799 2397 46811 2431
rect 46753 2391 46811 2397
rect 47026 2388 47032 2440
rect 47084 2428 47090 2440
rect 47121 2431 47179 2437
rect 47121 2428 47133 2431
rect 47084 2400 47133 2428
rect 47084 2388 47090 2400
rect 47121 2397 47133 2400
rect 47167 2397 47179 2431
rect 47121 2391 47179 2397
rect 35216 2332 36032 2360
rect 37568 2332 37964 2360
rect 35216 2320 35222 2332
rect 33045 2295 33103 2301
rect 33045 2261 33057 2295
rect 33091 2261 33103 2295
rect 33045 2255 33103 2261
rect 33502 2252 33508 2304
rect 33560 2292 33566 2304
rect 34149 2295 34207 2301
rect 34149 2292 34161 2295
rect 33560 2264 34161 2292
rect 33560 2252 33566 2264
rect 34149 2261 34161 2264
rect 34195 2261 34207 2295
rect 34149 2255 34207 2261
rect 34238 2252 34244 2304
rect 34296 2292 34302 2304
rect 34885 2295 34943 2301
rect 34885 2292 34897 2295
rect 34296 2264 34897 2292
rect 34296 2252 34302 2264
rect 34885 2261 34897 2264
rect 34931 2261 34943 2295
rect 34885 2255 34943 2261
rect 34974 2252 34980 2304
rect 35032 2292 35038 2304
rect 36004 2301 36032 2332
rect 35621 2295 35679 2301
rect 35621 2292 35633 2295
rect 35032 2264 35633 2292
rect 35032 2252 35038 2264
rect 35621 2261 35633 2264
rect 35667 2261 35679 2295
rect 35621 2255 35679 2261
rect 35989 2295 36047 2301
rect 35989 2261 36001 2295
rect 36035 2261 36047 2295
rect 35989 2255 36047 2261
rect 36722 2252 36728 2304
rect 36780 2292 36786 2304
rect 37369 2295 37427 2301
rect 37369 2292 37381 2295
rect 36780 2264 37381 2292
rect 36780 2252 36786 2264
rect 37369 2261 37381 2264
rect 37415 2261 37427 2295
rect 37369 2255 37427 2261
rect 38194 2252 38200 2304
rect 38252 2252 38258 2304
rect 38562 2252 38568 2304
rect 38620 2292 38626 2304
rect 38933 2295 38991 2301
rect 38933 2292 38945 2295
rect 38620 2264 38945 2292
rect 38620 2252 38626 2264
rect 38933 2261 38945 2264
rect 38979 2261 38991 2295
rect 38933 2255 38991 2261
rect 39390 2252 39396 2304
rect 39448 2292 39454 2304
rect 40037 2295 40095 2301
rect 40037 2292 40049 2295
rect 39448 2264 40049 2292
rect 39448 2252 39454 2264
rect 40037 2261 40049 2264
rect 40083 2261 40095 2295
rect 40037 2255 40095 2261
rect 45830 2252 45836 2304
rect 45888 2252 45894 2304
rect 46198 2252 46204 2304
rect 46256 2252 46262 2304
rect 46566 2252 46572 2304
rect 46624 2252 46630 2304
rect 46934 2252 46940 2304
rect 46992 2252 46998 2304
rect 1104 2202 47840 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 39010 2202
rect 39062 2150 39074 2202
rect 39126 2150 39138 2202
rect 39190 2150 39202 2202
rect 39254 2150 39266 2202
rect 39318 2150 45010 2202
rect 45062 2150 45074 2202
rect 45126 2150 45138 2202
rect 45190 2150 45202 2202
rect 45254 2150 45266 2202
rect 45318 2150 47840 2202
rect 1104 2128 47840 2150
rect 19150 2048 19156 2100
rect 19208 2088 19214 2100
rect 19208 2060 24716 2088
rect 19208 2048 19214 2060
rect 10502 1980 10508 2032
rect 10560 2020 10566 2032
rect 24118 2020 24124 2032
rect 10560 1992 24124 2020
rect 10560 1980 10566 1992
rect 24118 1980 24124 1992
rect 24176 1980 24182 2032
rect 24688 2020 24716 2060
rect 27430 2048 27436 2100
rect 27488 2088 27494 2100
rect 27890 2088 27896 2100
rect 27488 2060 27896 2088
rect 27488 2048 27494 2060
rect 27890 2048 27896 2060
rect 27948 2048 27954 2100
rect 29270 2048 29276 2100
rect 29328 2088 29334 2100
rect 29328 2060 30696 2088
rect 29328 2048 29334 2060
rect 25958 2020 25964 2032
rect 24688 1992 25964 2020
rect 25958 1980 25964 1992
rect 26016 1980 26022 2032
rect 30668 2020 30696 2060
rect 30742 2048 30748 2100
rect 30800 2088 30806 2100
rect 32766 2088 32772 2100
rect 30800 2060 32772 2088
rect 30800 2048 30806 2060
rect 32766 2048 32772 2060
rect 32824 2048 32830 2100
rect 32122 2020 32128 2032
rect 30668 1992 32128 2020
rect 32122 1980 32128 1992
rect 32180 1980 32186 2032
rect 37182 1980 37188 2032
rect 37240 2020 37246 2032
rect 40494 2020 40500 2032
rect 37240 1992 40500 2020
rect 37240 1980 37246 1992
rect 40494 1980 40500 1992
rect 40552 1980 40558 2032
rect 11422 1912 11428 1964
rect 11480 1952 11486 1964
rect 24486 1952 24492 1964
rect 11480 1924 24492 1952
rect 11480 1912 11486 1924
rect 24486 1912 24492 1924
rect 24544 1912 24550 1964
rect 25222 1952 25228 1964
rect 24596 1924 25228 1952
rect 15746 1844 15752 1896
rect 15804 1884 15810 1896
rect 24596 1884 24624 1924
rect 25222 1912 25228 1924
rect 25280 1912 25286 1964
rect 36538 1912 36544 1964
rect 36596 1952 36602 1964
rect 43530 1952 43536 1964
rect 36596 1924 43536 1952
rect 36596 1912 36602 1924
rect 43530 1912 43536 1924
rect 43588 1912 43594 1964
rect 15804 1856 24624 1884
rect 15804 1844 15810 1856
rect 30006 1844 30012 1896
rect 30064 1884 30070 1896
rect 46382 1884 46388 1896
rect 30064 1856 46388 1884
rect 30064 1844 30070 1856
rect 46382 1844 46388 1856
rect 46440 1844 46446 1896
rect 9582 1776 9588 1828
rect 9640 1816 9646 1828
rect 26326 1816 26332 1828
rect 9640 1788 26332 1816
rect 9640 1776 9646 1788
rect 26326 1776 26332 1788
rect 26384 1776 26390 1828
rect 30098 1816 30104 1828
rect 28966 1788 30104 1816
rect 7742 1708 7748 1760
rect 7800 1748 7806 1760
rect 23198 1748 23204 1760
rect 7800 1720 23204 1748
rect 7800 1708 7806 1720
rect 23198 1708 23204 1720
rect 23256 1708 23262 1760
rect 24118 1708 24124 1760
rect 24176 1748 24182 1760
rect 28966 1748 28994 1788
rect 30098 1776 30104 1788
rect 30156 1776 30162 1828
rect 24176 1720 28994 1748
rect 24176 1708 24182 1720
rect 11330 1640 11336 1692
rect 11388 1680 11394 1692
rect 28626 1680 28632 1692
rect 11388 1652 28632 1680
rect 11388 1640 11394 1652
rect 28626 1640 28632 1652
rect 28684 1640 28690 1692
rect 28718 1640 28724 1692
rect 28776 1680 28782 1692
rect 28902 1680 28908 1692
rect 28776 1652 28908 1680
rect 28776 1640 28782 1652
rect 28902 1640 28908 1652
rect 28960 1640 28966 1692
rect 26418 1572 26424 1624
rect 26476 1612 26482 1624
rect 36538 1612 36544 1624
rect 26476 1584 36544 1612
rect 26476 1572 26482 1584
rect 36538 1572 36544 1584
rect 36596 1572 36602 1624
rect 19426 1504 19432 1556
rect 19484 1544 19490 1556
rect 35618 1544 35624 1556
rect 19484 1516 35624 1544
rect 19484 1504 19490 1516
rect 35618 1504 35624 1516
rect 35676 1504 35682 1556
rect 25314 1436 25320 1488
rect 25372 1476 25378 1488
rect 38010 1476 38016 1488
rect 25372 1448 38016 1476
rect 25372 1436 25378 1448
rect 38010 1436 38016 1448
rect 38068 1436 38074 1488
rect 38102 1436 38108 1488
rect 38160 1476 38166 1488
rect 38562 1476 38568 1488
rect 38160 1448 38568 1476
rect 38160 1436 38166 1448
rect 38562 1436 38568 1448
rect 38620 1436 38626 1488
rect 24486 1368 24492 1420
rect 24544 1408 24550 1420
rect 30558 1408 30564 1420
rect 24544 1380 30564 1408
rect 24544 1368 24550 1380
rect 30558 1368 30564 1380
rect 30616 1368 30622 1420
rect 31754 1368 31760 1420
rect 31812 1408 31818 1420
rect 32674 1408 32680 1420
rect 31812 1380 32680 1408
rect 31812 1368 31818 1380
rect 32674 1368 32680 1380
rect 32732 1368 32738 1420
rect 37274 1368 37280 1420
rect 37332 1408 37338 1420
rect 38194 1408 38200 1420
rect 37332 1380 38200 1408
rect 37332 1368 37338 1380
rect 38194 1368 38200 1380
rect 38252 1368 38258 1420
rect 39574 1368 39580 1420
rect 39632 1408 39638 1420
rect 41322 1408 41328 1420
rect 39632 1380 41328 1408
rect 39632 1368 39638 1380
rect 41322 1368 41328 1380
rect 41380 1368 41386 1420
rect 5718 1300 5724 1352
rect 5776 1340 5782 1352
rect 22830 1340 22836 1352
rect 5776 1312 22836 1340
rect 5776 1300 5782 1312
rect 22830 1300 22836 1312
rect 22888 1300 22894 1352
rect 32490 1300 32496 1352
rect 32548 1340 32554 1352
rect 32950 1340 32956 1352
rect 32548 1312 32956 1340
rect 32548 1300 32554 1312
rect 32950 1300 32956 1312
rect 33008 1300 33014 1352
rect 5534 1232 5540 1284
rect 5592 1272 5598 1284
rect 22094 1272 22100 1284
rect 5592 1244 22100 1272
rect 5592 1232 5598 1244
rect 22094 1232 22100 1244
rect 22152 1232 22158 1284
rect 13354 620 13360 672
rect 13412 660 13418 672
rect 24670 660 24676 672
rect 13412 632 24676 660
rect 13412 620 13418 632
rect 24670 620 24676 632
rect 24728 620 24734 672
rect 20346 552 20352 604
rect 20404 592 20410 604
rect 32306 592 32312 604
rect 20404 564 32312 592
rect 20404 552 20410 564
rect 32306 552 32312 564
rect 32364 552 32370 604
rect 7098 484 7104 536
rect 7156 524 7162 536
rect 23474 524 23480 536
rect 7156 496 23480 524
rect 7156 484 7162 496
rect 23474 484 23480 496
rect 23532 484 23538 536
rect 3418 416 3424 468
rect 3476 456 3482 468
rect 20806 456 20812 468
rect 3476 428 20812 456
rect 3476 416 3482 428
rect 20806 416 20812 428
rect 20864 416 20870 468
rect 10778 348 10784 400
rect 10836 388 10842 400
rect 28994 388 29000 400
rect 10836 360 29000 388
rect 10836 348 10842 360
rect 28994 348 29000 360
rect 29052 348 29058 400
rect 10410 280 10416 332
rect 10468 320 10474 332
rect 29638 320 29644 332
rect 10468 292 29644 320
rect 10468 280 10474 292
rect 29638 280 29644 292
rect 29696 280 29702 332
rect 32950 280 32956 332
rect 33008 320 33014 332
rect 41690 320 41696 332
rect 33008 292 41696 320
rect 33008 280 33014 292
rect 41690 280 41696 292
rect 41748 280 41754 332
rect 10042 212 10048 264
rect 10100 252 10106 264
rect 29822 252 29828 264
rect 10100 224 29828 252
rect 10100 212 10106 224
rect 29822 212 29828 224
rect 29880 212 29886 264
rect 30926 212 30932 264
rect 30984 252 30990 264
rect 42426 252 42432 264
rect 30984 224 42432 252
rect 30984 212 30990 224
rect 42426 212 42432 224
rect 42484 212 42490 264
rect 8938 144 8944 196
rect 8996 144 9002 196
rect 9674 144 9680 196
rect 9732 184 9738 196
rect 30466 184 30472 196
rect 9732 156 30472 184
rect 9732 144 9738 156
rect 30466 144 30472 156
rect 30524 144 30530 196
rect 31202 144 31208 196
rect 31260 184 31266 196
rect 42794 184 42800 196
rect 31260 156 42800 184
rect 31260 144 31266 156
rect 42794 144 42800 156
rect 42852 144 42858 196
rect 8956 116 8984 144
rect 31846 116 31852 128
rect 8956 88 31852 116
rect 31846 76 31852 88
rect 31904 76 31910 128
rect 33778 76 33784 128
rect 33836 116 33842 128
rect 41966 116 41972 128
rect 33836 88 41972 116
rect 33836 76 33842 88
rect 41966 76 41972 88
rect 42024 76 42030 128
rect 18230 8 18236 60
rect 18288 48 18294 60
rect 44818 48 44824 60
rect 18288 20 44824 48
rect 18288 8 18294 20
rect 44818 8 44824 20
rect 44876 8 44882 60
<< via1 >>
rect 33876 9188 33928 9240
rect 38568 9188 38620 9240
rect 19524 9120 19576 9172
rect 46020 9120 46072 9172
rect 33968 9052 34020 9104
rect 40408 9052 40460 9104
rect 37280 8984 37332 9036
rect 6644 8916 6696 8968
rect 38752 8916 38804 8968
rect 23940 8848 23992 8900
rect 46388 8848 46440 8900
rect 4068 8780 4120 8832
rect 26516 8780 26568 8832
rect 41236 8780 41288 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 39010 8678 39062 8730
rect 39074 8678 39126 8730
rect 39138 8678 39190 8730
rect 39202 8678 39254 8730
rect 39266 8678 39318 8730
rect 45010 8678 45062 8730
rect 45074 8678 45126 8730
rect 45138 8678 45190 8730
rect 45202 8678 45254 8730
rect 45266 8678 45318 8730
rect 1400 8576 1452 8628
rect 3700 8576 3752 8628
rect 4068 8576 4120 8628
rect 6000 8576 6052 8628
rect 8300 8576 8352 8628
rect 10600 8576 10652 8628
rect 12900 8576 12952 8628
rect 15384 8576 15436 8628
rect 17500 8576 17552 8628
rect 19800 8576 19852 8628
rect 22100 8576 22152 8628
rect 24400 8576 24452 8628
rect 26700 8576 26752 8628
rect 29000 8576 29052 8628
rect 31300 8576 31352 8628
rect 33600 8576 33652 8628
rect 34060 8576 34112 8628
rect 35900 8576 35952 8628
rect 38200 8576 38252 8628
rect 40500 8576 40552 8628
rect 42800 8576 42852 8628
rect 45376 8576 45428 8628
rect 45836 8619 45888 8628
rect 45836 8585 45845 8619
rect 45845 8585 45879 8619
rect 45879 8585 45888 8619
rect 45836 8576 45888 8585
rect 46204 8619 46256 8628
rect 46204 8585 46213 8619
rect 46213 8585 46247 8619
rect 46247 8585 46256 8619
rect 46204 8576 46256 8585
rect 47400 8576 47452 8628
rect 22192 8508 22244 8560
rect 34244 8508 34296 8560
rect 6644 8483 6696 8492
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 6644 8440 6696 8449
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 10692 8483 10744 8492
rect 10692 8449 10701 8483
rect 10701 8449 10735 8483
rect 10735 8449 10744 8483
rect 10692 8440 10744 8449
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 15384 8440 15436 8492
rect 17868 8483 17920 8492
rect 17868 8449 17877 8483
rect 17877 8449 17911 8483
rect 17911 8449 17920 8483
rect 17868 8440 17920 8449
rect 20628 8440 20680 8492
rect 23480 8440 23532 8492
rect 25872 8440 25924 8492
rect 29276 8440 29328 8492
rect 29368 8483 29420 8492
rect 29368 8449 29377 8483
rect 29377 8449 29411 8483
rect 29411 8449 29420 8483
rect 29368 8440 29420 8449
rect 33876 8440 33928 8492
rect 33968 8483 34020 8492
rect 33968 8449 33977 8483
rect 33977 8449 34011 8483
rect 34011 8449 34020 8483
rect 33968 8440 34020 8449
rect 37188 8440 37240 8492
rect 39580 8440 39632 8492
rect 40868 8483 40920 8492
rect 40868 8449 40877 8483
rect 40877 8449 40911 8483
rect 40911 8449 40920 8483
rect 40868 8440 40920 8449
rect 43168 8483 43220 8492
rect 43168 8449 43177 8483
rect 43177 8449 43211 8483
rect 43211 8449 43220 8483
rect 43168 8440 43220 8449
rect 45468 8483 45520 8492
rect 45468 8449 45477 8483
rect 45477 8449 45511 8483
rect 45511 8449 45520 8483
rect 45468 8440 45520 8449
rect 46020 8483 46072 8492
rect 46020 8449 46029 8483
rect 46029 8449 46063 8483
rect 46063 8449 46072 8483
rect 46020 8440 46072 8449
rect 46388 8483 46440 8492
rect 46388 8449 46397 8483
rect 46397 8449 46431 8483
rect 46431 8449 46440 8483
rect 46388 8440 46440 8449
rect 46756 8483 46808 8492
rect 46756 8449 46765 8483
rect 46765 8449 46799 8483
rect 46799 8449 46808 8483
rect 46756 8440 46808 8449
rect 37832 8372 37884 8424
rect 41236 8372 41288 8424
rect 29276 8236 29328 8288
rect 39948 8304 40000 8356
rect 47216 8304 47268 8356
rect 47308 8347 47360 8356
rect 47308 8313 47317 8347
rect 47317 8313 47351 8347
rect 47351 8313 47360 8347
rect 47308 8304 47360 8313
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 37950 8134 38002 8186
rect 38014 8134 38066 8186
rect 38078 8134 38130 8186
rect 38142 8134 38194 8186
rect 38206 8134 38258 8186
rect 43950 8134 44002 8186
rect 44014 8134 44066 8186
rect 44078 8134 44130 8186
rect 44142 8134 44194 8186
rect 44206 8134 44258 8186
rect 8392 8032 8444 8084
rect 10692 8032 10744 8084
rect 19524 8075 19576 8084
rect 19524 8041 19533 8075
rect 19533 8041 19567 8075
rect 19567 8041 19576 8075
rect 19524 8032 19576 8041
rect 20536 8075 20588 8084
rect 20536 8041 20545 8075
rect 20545 8041 20579 8075
rect 20579 8041 20588 8075
rect 20536 8032 20588 8041
rect 20628 8075 20680 8084
rect 20628 8041 20637 8075
rect 20637 8041 20671 8075
rect 20671 8041 20680 8075
rect 20628 8032 20680 8041
rect 21732 8075 21784 8084
rect 21732 8041 21741 8075
rect 21741 8041 21775 8075
rect 21775 8041 21784 8075
rect 21732 8032 21784 8041
rect 22192 8032 22244 8084
rect 23480 8075 23532 8084
rect 23480 8041 23489 8075
rect 23489 8041 23523 8075
rect 23523 8041 23532 8075
rect 23480 8032 23532 8041
rect 23940 8075 23992 8084
rect 23940 8041 23949 8075
rect 23949 8041 23983 8075
rect 23983 8041 23992 8075
rect 23940 8032 23992 8041
rect 25872 8032 25924 8084
rect 26516 8075 26568 8084
rect 26516 8041 26525 8075
rect 26525 8041 26559 8075
rect 26559 8041 26568 8075
rect 26516 8032 26568 8041
rect 29368 8032 29420 8084
rect 37832 8075 37884 8084
rect 37832 8041 37841 8075
rect 37841 8041 37875 8075
rect 37875 8041 37884 8075
rect 37832 8032 37884 8041
rect 43812 8032 43864 8084
rect 7564 7964 7616 8016
rect 11612 7964 11664 8016
rect 11796 7964 11848 8016
rect 46664 8075 46716 8084
rect 46664 8041 46673 8075
rect 46673 8041 46707 8075
rect 46707 8041 46716 8075
rect 46664 8032 46716 8041
rect 1032 7828 1084 7880
rect 10048 7871 10100 7880
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 10140 7828 10192 7880
rect 14188 7828 14240 7880
rect 19340 7871 19392 7880
rect 19340 7837 19349 7871
rect 19349 7837 19383 7871
rect 19383 7837 19392 7871
rect 19340 7828 19392 7837
rect 20352 7871 20404 7880
rect 20352 7837 20361 7871
rect 20361 7837 20395 7871
rect 20395 7837 20404 7871
rect 20352 7828 20404 7837
rect 20812 7871 20864 7880
rect 20812 7837 20821 7871
rect 20821 7837 20855 7871
rect 20855 7837 20864 7871
rect 20812 7828 20864 7837
rect 3792 7760 3844 7812
rect 11888 7692 11940 7744
rect 16028 7692 16080 7744
rect 20720 7692 20772 7744
rect 23388 7760 23440 7812
rect 23756 7871 23808 7880
rect 23756 7837 23765 7871
rect 23765 7837 23799 7871
rect 23799 7837 23808 7871
rect 23756 7828 23808 7837
rect 25596 7871 25648 7880
rect 25596 7837 25605 7871
rect 25605 7837 25639 7871
rect 25639 7837 25648 7871
rect 25596 7828 25648 7837
rect 26240 7871 26292 7880
rect 26240 7837 26249 7871
rect 26249 7837 26283 7871
rect 26283 7837 26292 7871
rect 26240 7828 26292 7837
rect 26332 7871 26384 7880
rect 26332 7837 26341 7871
rect 26341 7837 26375 7871
rect 26375 7837 26384 7871
rect 26332 7828 26384 7837
rect 26516 7828 26568 7880
rect 29920 7828 29972 7880
rect 24952 7760 25004 7812
rect 24676 7692 24728 7744
rect 36544 7760 36596 7812
rect 39672 7828 39724 7880
rect 39856 7760 39908 7812
rect 46020 7871 46072 7880
rect 46020 7837 46029 7871
rect 46029 7837 46063 7871
rect 46063 7837 46072 7871
rect 46020 7828 46072 7837
rect 46112 7871 46164 7880
rect 46112 7837 46121 7871
rect 46121 7837 46155 7871
rect 46155 7837 46164 7871
rect 46112 7828 46164 7837
rect 47216 7871 47268 7880
rect 47216 7837 47225 7871
rect 47225 7837 47259 7871
rect 47259 7837 47268 7871
rect 47216 7828 47268 7837
rect 46572 7760 46624 7812
rect 29736 7735 29788 7744
rect 29736 7701 29745 7735
rect 29745 7701 29779 7735
rect 29779 7701 29788 7735
rect 29736 7692 29788 7701
rect 30472 7692 30524 7744
rect 36176 7692 36228 7744
rect 36820 7692 36872 7744
rect 40132 7692 40184 7744
rect 40316 7692 40368 7744
rect 44824 7692 44876 7744
rect 45376 7692 45428 7744
rect 45928 7692 45980 7744
rect 46296 7735 46348 7744
rect 46296 7701 46305 7735
rect 46305 7701 46339 7735
rect 46339 7701 46348 7735
rect 46296 7692 46348 7701
rect 47032 7735 47084 7744
rect 47032 7701 47041 7735
rect 47041 7701 47075 7735
rect 47075 7701 47084 7735
rect 47032 7692 47084 7701
rect 47400 7735 47452 7744
rect 47400 7701 47409 7735
rect 47409 7701 47443 7735
rect 47443 7701 47452 7735
rect 47400 7692 47452 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 39010 7590 39062 7642
rect 39074 7590 39126 7642
rect 39138 7590 39190 7642
rect 39202 7590 39254 7642
rect 39266 7590 39318 7642
rect 45010 7590 45062 7642
rect 45074 7590 45126 7642
rect 45138 7590 45190 7642
rect 45202 7590 45254 7642
rect 45266 7590 45318 7642
rect 4160 7488 4212 7540
rect 1584 7420 1636 7472
rect 10048 7352 10100 7404
rect 1860 7284 1912 7336
rect 10140 7284 10192 7336
rect 11612 7463 11664 7472
rect 11612 7429 11621 7463
rect 11621 7429 11655 7463
rect 11655 7429 11664 7463
rect 11612 7420 11664 7429
rect 12992 7488 13044 7540
rect 15384 7488 15436 7540
rect 17868 7531 17920 7540
rect 17868 7497 17877 7531
rect 17877 7497 17911 7531
rect 17911 7497 17920 7531
rect 17868 7488 17920 7497
rect 20536 7488 20588 7540
rect 23572 7488 23624 7540
rect 29736 7488 29788 7540
rect 36452 7488 36504 7540
rect 37280 7488 37332 7540
rect 38752 7531 38804 7540
rect 38752 7497 38761 7531
rect 38761 7497 38795 7531
rect 38795 7497 38804 7531
rect 38752 7488 38804 7497
rect 39580 7531 39632 7540
rect 39580 7497 39589 7531
rect 39589 7497 39623 7531
rect 39623 7497 39632 7531
rect 39580 7488 39632 7497
rect 40868 7488 40920 7540
rect 43444 7488 43496 7540
rect 45376 7488 45428 7540
rect 46756 7488 46808 7540
rect 46940 7531 46992 7540
rect 46940 7497 46949 7531
rect 46949 7497 46983 7531
rect 46983 7497 46992 7531
rect 46940 7488 46992 7497
rect 20352 7420 20404 7472
rect 20812 7420 20864 7472
rect 31208 7420 31260 7472
rect 36544 7420 36596 7472
rect 11796 7395 11848 7404
rect 11796 7361 11805 7395
rect 11805 7361 11839 7395
rect 11839 7361 11848 7395
rect 11796 7352 11848 7361
rect 14188 7284 14240 7336
rect 18052 7395 18104 7404
rect 18052 7361 18061 7395
rect 18061 7361 18095 7395
rect 18095 7361 18104 7395
rect 18052 7352 18104 7361
rect 33784 7284 33836 7336
rect 38936 7284 38988 7336
rect 39580 7284 39632 7336
rect 45928 7352 45980 7404
rect 45744 7284 45796 7336
rect 46572 7352 46624 7404
rect 47492 7284 47544 7336
rect 11980 7191 12032 7200
rect 11980 7157 11989 7191
rect 11989 7157 12023 7191
rect 12023 7157 12032 7191
rect 11980 7148 12032 7157
rect 22928 7191 22980 7200
rect 22928 7157 22937 7191
rect 22937 7157 22971 7191
rect 22971 7157 22980 7191
rect 22928 7148 22980 7157
rect 23296 7191 23348 7200
rect 23296 7157 23305 7191
rect 23305 7157 23339 7191
rect 23339 7157 23348 7191
rect 23296 7148 23348 7157
rect 27620 7148 27672 7200
rect 37372 7148 37424 7200
rect 38660 7148 38712 7200
rect 40592 7216 40644 7268
rect 40224 7148 40276 7200
rect 47308 7191 47360 7200
rect 47308 7157 47317 7191
rect 47317 7157 47351 7191
rect 47351 7157 47360 7191
rect 47308 7148 47360 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 37950 7046 38002 7098
rect 38014 7046 38066 7098
rect 38078 7046 38130 7098
rect 38142 7046 38194 7098
rect 38206 7046 38258 7098
rect 43950 7046 44002 7098
rect 44014 7046 44066 7098
rect 44078 7046 44130 7098
rect 44142 7046 44194 7098
rect 44206 7046 44258 7098
rect 23296 6944 23348 6996
rect 43720 6944 43772 6996
rect 46020 6944 46072 6996
rect 12348 6808 12400 6860
rect 1308 6740 1360 6792
rect 36452 6876 36504 6928
rect 44364 6876 44416 6928
rect 43812 6808 43864 6860
rect 12256 6672 12308 6724
rect 36544 6672 36596 6724
rect 38568 6672 38620 6724
rect 18972 6604 19024 6656
rect 25872 6604 25924 6656
rect 26332 6647 26384 6656
rect 26332 6613 26341 6647
rect 26341 6613 26375 6647
rect 26375 6613 26384 6647
rect 26332 6604 26384 6613
rect 39948 6604 40000 6656
rect 44640 6740 44692 6792
rect 46296 6808 46348 6860
rect 46020 6783 46072 6792
rect 46020 6749 46029 6783
rect 46029 6749 46063 6783
rect 46063 6749 46072 6783
rect 46020 6740 46072 6749
rect 46664 6783 46716 6792
rect 46664 6749 46673 6783
rect 46673 6749 46707 6783
rect 46707 6749 46716 6783
rect 46664 6740 46716 6749
rect 42708 6672 42760 6724
rect 47124 6740 47176 6792
rect 42800 6604 42852 6656
rect 43168 6604 43220 6656
rect 45468 6604 45520 6656
rect 47032 6647 47084 6656
rect 47032 6613 47041 6647
rect 47041 6613 47075 6647
rect 47075 6613 47084 6647
rect 47032 6604 47084 6613
rect 47400 6647 47452 6656
rect 47400 6613 47409 6647
rect 47409 6613 47443 6647
rect 47443 6613 47452 6647
rect 47400 6604 47452 6613
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 39010 6502 39062 6554
rect 39074 6502 39126 6554
rect 39138 6502 39190 6554
rect 39202 6502 39254 6554
rect 39266 6502 39318 6554
rect 45010 6502 45062 6554
rect 45074 6502 45126 6554
rect 45138 6502 45190 6554
rect 45202 6502 45254 6554
rect 45266 6502 45318 6554
rect 8668 6400 8720 6452
rect 23296 6400 23348 6452
rect 26332 6400 26384 6452
rect 40040 6400 40092 6452
rect 40408 6400 40460 6452
rect 47308 6443 47360 6452
rect 47308 6409 47317 6443
rect 47317 6409 47351 6443
rect 47351 6409 47360 6443
rect 47308 6400 47360 6409
rect 18052 6332 18104 6384
rect 30932 6332 30984 6384
rect 36544 6332 36596 6384
rect 47216 6332 47268 6384
rect 3424 6264 3476 6316
rect 30380 6264 30432 6316
rect 1308 6196 1360 6248
rect 26516 6196 26568 6248
rect 45376 6264 45428 6316
rect 46572 6307 46624 6316
rect 46572 6273 46581 6307
rect 46581 6273 46615 6307
rect 46615 6273 46624 6307
rect 46572 6264 46624 6273
rect 44916 6196 44968 6248
rect 480 6128 532 6180
rect 27620 6128 27672 6180
rect 37188 6128 37240 6180
rect 24768 6060 24820 6112
rect 35440 6060 35492 6112
rect 46756 6103 46808 6112
rect 46756 6069 46765 6103
rect 46765 6069 46799 6103
rect 46799 6069 46808 6103
rect 46756 6060 46808 6069
rect 46940 6103 46992 6112
rect 46940 6069 46949 6103
rect 46949 6069 46983 6103
rect 46983 6069 46992 6103
rect 46940 6060 46992 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 37950 5958 38002 6010
rect 38014 5958 38066 6010
rect 38078 5958 38130 6010
rect 38142 5958 38194 6010
rect 38206 5958 38258 6010
rect 43950 5958 44002 6010
rect 44014 5958 44066 6010
rect 44078 5958 44130 6010
rect 44142 5958 44194 6010
rect 44206 5958 44258 6010
rect 8668 5899 8720 5908
rect 8668 5865 8677 5899
rect 8677 5865 8711 5899
rect 8711 5865 8720 5899
rect 8668 5856 8720 5865
rect 12164 5856 12216 5908
rect 19248 5856 19300 5908
rect 20720 5856 20772 5908
rect 24676 5788 24728 5840
rect 42800 5856 42852 5908
rect 43812 5856 43864 5908
rect 46940 5788 46992 5840
rect 47400 5831 47452 5840
rect 47400 5797 47409 5831
rect 47409 5797 47443 5831
rect 47443 5797 47452 5831
rect 47400 5788 47452 5797
rect 18972 5720 19024 5772
rect 46112 5720 46164 5772
rect 12624 5652 12676 5704
rect 15936 5652 15988 5704
rect 22008 5652 22060 5704
rect 27528 5652 27580 5704
rect 32772 5695 32824 5704
rect 32772 5661 32781 5695
rect 32781 5661 32815 5695
rect 32815 5661 32824 5695
rect 32772 5652 32824 5661
rect 45560 5652 45612 5704
rect 47216 5695 47268 5704
rect 47216 5661 47225 5695
rect 47225 5661 47259 5695
rect 47259 5661 47268 5695
rect 47216 5652 47268 5661
rect 18972 5584 19024 5636
rect 30472 5584 30524 5636
rect 14924 5516 14976 5568
rect 47124 5584 47176 5636
rect 46204 5516 46256 5568
rect 47032 5559 47084 5568
rect 47032 5525 47041 5559
rect 47041 5525 47075 5559
rect 47075 5525 47084 5559
rect 47032 5516 47084 5525
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 39010 5414 39062 5466
rect 39074 5414 39126 5466
rect 39138 5414 39190 5466
rect 39202 5414 39254 5466
rect 39266 5414 39318 5466
rect 45010 5414 45062 5466
rect 45074 5414 45126 5466
rect 45138 5414 45190 5466
rect 45202 5414 45254 5466
rect 45266 5414 45318 5466
rect 11428 5312 11480 5364
rect 11520 5312 11572 5364
rect 11060 5244 11112 5296
rect 10416 5219 10468 5228
rect 10416 5185 10425 5219
rect 10425 5185 10459 5219
rect 10459 5185 10468 5219
rect 10416 5176 10468 5185
rect 12348 5219 12400 5228
rect 12348 5185 12357 5219
rect 12357 5185 12391 5219
rect 12391 5185 12400 5219
rect 12348 5176 12400 5185
rect 15476 5244 15528 5296
rect 11888 5040 11940 5092
rect 8484 4972 8536 5024
rect 10508 4972 10560 5024
rect 10600 5015 10652 5024
rect 10600 4981 10609 5015
rect 10609 4981 10643 5015
rect 10643 4981 10652 5015
rect 10600 4972 10652 4981
rect 11336 5015 11388 5024
rect 11336 4981 11345 5015
rect 11345 4981 11379 5015
rect 11379 4981 11388 5015
rect 11336 4972 11388 4981
rect 14280 5108 14332 5160
rect 16212 5176 16264 5228
rect 16672 5176 16724 5228
rect 17040 5219 17092 5228
rect 17040 5185 17049 5219
rect 17049 5185 17083 5219
rect 17083 5185 17092 5219
rect 17040 5176 17092 5185
rect 17408 5176 17460 5228
rect 22008 5355 22060 5364
rect 22008 5321 22017 5355
rect 22017 5321 22051 5355
rect 22051 5321 22060 5355
rect 22008 5312 22060 5321
rect 21640 5244 21692 5296
rect 46572 5312 46624 5364
rect 47308 5355 47360 5364
rect 47308 5321 47317 5355
rect 47317 5321 47351 5355
rect 47351 5321 47360 5355
rect 47308 5312 47360 5321
rect 26608 5244 26660 5296
rect 45652 5244 45704 5296
rect 47216 5244 47268 5296
rect 21732 5176 21784 5228
rect 15568 5108 15620 5160
rect 12532 5083 12584 5092
rect 12532 5049 12541 5083
rect 12541 5049 12575 5083
rect 12575 5049 12584 5083
rect 12532 5040 12584 5049
rect 13728 5040 13780 5092
rect 24032 5176 24084 5228
rect 26976 5219 27028 5228
rect 26976 5185 26985 5219
rect 26985 5185 27019 5219
rect 27019 5185 27028 5219
rect 26976 5176 27028 5185
rect 18604 5040 18656 5092
rect 43720 5176 43772 5228
rect 12716 4972 12768 5024
rect 12900 5015 12952 5024
rect 12900 4981 12909 5015
rect 12909 4981 12943 5015
rect 12943 4981 12952 5015
rect 12900 4972 12952 4981
rect 15384 4972 15436 5024
rect 17132 4972 17184 5024
rect 17224 5015 17276 5024
rect 17224 4981 17233 5015
rect 17233 4981 17267 5015
rect 17267 4981 17276 5015
rect 17224 4972 17276 4981
rect 17868 4972 17920 5024
rect 27528 5040 27580 5092
rect 42708 5040 42760 5092
rect 23204 5015 23256 5024
rect 23204 4981 23213 5015
rect 23213 4981 23247 5015
rect 23247 4981 23256 5015
rect 23204 4972 23256 4981
rect 23480 5015 23532 5024
rect 23480 4981 23489 5015
rect 23489 4981 23523 5015
rect 23523 4981 23532 5015
rect 23480 4972 23532 4981
rect 26884 4972 26936 5024
rect 27436 4972 27488 5024
rect 29644 4972 29696 5024
rect 46940 5015 46992 5024
rect 46940 4981 46949 5015
rect 46949 4981 46983 5015
rect 46983 4981 46992 5015
rect 46940 4972 46992 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 37950 4870 38002 4922
rect 38014 4870 38066 4922
rect 38078 4870 38130 4922
rect 38142 4870 38194 4922
rect 38206 4870 38258 4922
rect 43950 4870 44002 4922
rect 44014 4870 44066 4922
rect 44078 4870 44130 4922
rect 44142 4870 44194 4922
rect 44206 4870 44258 4922
rect 7748 4768 7800 4820
rect 10416 4768 10468 4820
rect 13728 4768 13780 4820
rect 14740 4768 14792 4820
rect 17868 4768 17920 4820
rect 21640 4768 21692 4820
rect 31760 4768 31812 4820
rect 2596 4564 2648 4616
rect 4528 4632 4580 4684
rect 6736 4632 6788 4684
rect 12348 4700 12400 4752
rect 14832 4700 14884 4752
rect 17224 4700 17276 4752
rect 25320 4700 25372 4752
rect 29644 4700 29696 4752
rect 42800 4768 42852 4820
rect 40040 4700 40092 4752
rect 2320 4496 2372 4548
rect 4896 4496 4948 4548
rect 5264 4564 5316 4616
rect 7472 4564 7524 4616
rect 5632 4496 5684 4548
rect 2780 4428 2832 4480
rect 4436 4471 4488 4480
rect 4436 4437 4445 4471
rect 4445 4437 4479 4471
rect 4479 4437 4488 4471
rect 4436 4428 4488 4437
rect 5540 4428 5592 4480
rect 8208 4496 8260 4548
rect 9588 4428 9640 4480
rect 16580 4632 16632 4684
rect 23204 4632 23256 4684
rect 27436 4632 27488 4684
rect 41604 4632 41656 4684
rect 19248 4607 19300 4616
rect 19248 4573 19257 4607
rect 19257 4573 19291 4607
rect 19291 4573 19300 4607
rect 19248 4564 19300 4573
rect 20904 4564 20956 4616
rect 31760 4564 31812 4616
rect 37004 4564 37056 4616
rect 37372 4564 37424 4616
rect 47400 4743 47452 4752
rect 47400 4709 47409 4743
rect 47409 4709 47443 4743
rect 47443 4709 47452 4743
rect 47400 4700 47452 4709
rect 19340 4496 19392 4548
rect 19432 4471 19484 4480
rect 19432 4437 19441 4471
rect 19441 4437 19475 4471
rect 19475 4437 19484 4471
rect 19432 4428 19484 4437
rect 22008 4428 22060 4480
rect 26700 4471 26752 4480
rect 26700 4437 26709 4471
rect 26709 4437 26743 4471
rect 26743 4437 26752 4471
rect 26700 4428 26752 4437
rect 37188 4428 37240 4480
rect 47032 4471 47084 4480
rect 47032 4437 47041 4471
rect 47041 4437 47075 4471
rect 47075 4437 47084 4471
rect 47032 4428 47084 4437
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 39010 4326 39062 4378
rect 39074 4326 39126 4378
rect 39138 4326 39190 4378
rect 39202 4326 39254 4378
rect 39266 4326 39318 4378
rect 45010 4326 45062 4378
rect 45074 4326 45126 4378
rect 45138 4326 45190 4378
rect 45202 4326 45254 4378
rect 45266 4326 45318 4378
rect 2780 4224 2832 4276
rect 1124 4156 1176 4208
rect 4436 4156 4488 4208
rect 5724 4156 5776 4208
rect 8208 4156 8260 4208
rect 7840 4088 7892 4140
rect 8576 4088 8628 4140
rect 11060 4156 11112 4208
rect 12256 4156 12308 4208
rect 16488 4224 16540 4276
rect 26700 4224 26752 4276
rect 26792 4224 26844 4276
rect 42432 4224 42484 4276
rect 15844 4156 15896 4208
rect 16580 4156 16632 4208
rect 18420 4199 18472 4208
rect 18420 4165 18429 4199
rect 18429 4165 18463 4199
rect 18463 4165 18472 4199
rect 18420 4156 18472 4165
rect 20628 4156 20680 4208
rect 25872 4156 25924 4208
rect 46020 4156 46072 4208
rect 2412 4063 2464 4072
rect 2412 4029 2421 4063
rect 2421 4029 2455 4063
rect 2455 4029 2464 4063
rect 2412 4020 2464 4029
rect 8300 4020 8352 4072
rect 7564 3927 7616 3936
rect 7564 3893 7573 3927
rect 7573 3893 7607 3927
rect 7607 3893 7616 3927
rect 7564 3884 7616 3893
rect 15752 4020 15804 4072
rect 20720 4088 20772 4140
rect 40040 4131 40092 4140
rect 40040 4097 40049 4131
rect 40049 4097 40083 4131
rect 40083 4097 40092 4131
rect 40040 4088 40092 4097
rect 42432 4131 42484 4140
rect 42432 4097 42441 4131
rect 42441 4097 42475 4131
rect 42475 4097 42484 4131
rect 42432 4088 42484 4097
rect 22468 4020 22520 4072
rect 44364 4020 44416 4072
rect 23296 3952 23348 4004
rect 30656 3952 30708 4004
rect 47308 3995 47360 4004
rect 47308 3961 47317 3995
rect 47317 3961 47351 3995
rect 47351 3961 47360 3995
rect 47308 3952 47360 3961
rect 15660 3884 15712 3936
rect 18880 3884 18932 3936
rect 28264 3884 28316 3936
rect 30840 3884 30892 3936
rect 33508 3884 33560 3936
rect 42616 3927 42668 3936
rect 42616 3893 42625 3927
rect 42625 3893 42659 3927
rect 42659 3893 42668 3927
rect 42616 3884 42668 3893
rect 46296 3927 46348 3936
rect 46296 3893 46305 3927
rect 46305 3893 46339 3927
rect 46339 3893 46348 3927
rect 46296 3884 46348 3893
rect 46848 3884 46900 3936
rect 46940 3927 46992 3936
rect 46940 3893 46949 3927
rect 46949 3893 46983 3927
rect 46983 3893 46992 3927
rect 46940 3884 46992 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 37950 3782 38002 3834
rect 38014 3782 38066 3834
rect 38078 3782 38130 3834
rect 38142 3782 38194 3834
rect 38206 3782 38258 3834
rect 43950 3782 44002 3834
rect 44014 3782 44066 3834
rect 44078 3782 44130 3834
rect 44142 3782 44194 3834
rect 44206 3782 44258 3834
rect 15384 3680 15436 3732
rect 38844 3680 38896 3732
rect 46020 3723 46072 3732
rect 46020 3689 46029 3723
rect 46029 3689 46063 3723
rect 46063 3689 46072 3723
rect 46020 3680 46072 3689
rect 8484 3612 8536 3664
rect 18880 3612 18932 3664
rect 25044 3612 25096 3664
rect 29828 3655 29880 3664
rect 29828 3621 29837 3655
rect 29837 3621 29871 3655
rect 29871 3621 29880 3655
rect 29828 3612 29880 3621
rect 1216 3476 1268 3528
rect 16488 3544 16540 3596
rect 20352 3544 20404 3596
rect 47032 3612 47084 3664
rect 6368 3408 6420 3460
rect 29000 3476 29052 3528
rect 29644 3519 29696 3528
rect 29644 3485 29653 3519
rect 29653 3485 29687 3519
rect 29687 3485 29696 3519
rect 29644 3476 29696 3485
rect 30104 3519 30156 3528
rect 30104 3485 30113 3519
rect 30113 3485 30147 3519
rect 30147 3485 30156 3519
rect 30104 3476 30156 3485
rect 31300 3519 31352 3528
rect 31300 3485 31309 3519
rect 31309 3485 31343 3519
rect 31343 3485 31352 3519
rect 31300 3476 31352 3485
rect 1308 3340 1360 3392
rect 14740 3340 14792 3392
rect 17224 3340 17276 3392
rect 28172 3408 28224 3460
rect 29828 3408 29880 3460
rect 30748 3408 30800 3460
rect 27528 3340 27580 3392
rect 29276 3340 29328 3392
rect 29368 3383 29420 3392
rect 29368 3349 29377 3383
rect 29377 3349 29411 3383
rect 29411 3349 29420 3383
rect 29368 3340 29420 3349
rect 30380 3340 30432 3392
rect 30472 3383 30524 3392
rect 30472 3349 30481 3383
rect 30481 3349 30515 3383
rect 30515 3349 30524 3383
rect 30472 3340 30524 3349
rect 30840 3383 30892 3392
rect 30840 3349 30849 3383
rect 30849 3349 30883 3383
rect 30883 3349 30892 3383
rect 30840 3340 30892 3349
rect 33968 3544 34020 3596
rect 42616 3544 42668 3596
rect 31852 3519 31904 3528
rect 31852 3485 31861 3519
rect 31861 3485 31895 3519
rect 31895 3485 31904 3519
rect 31852 3476 31904 3485
rect 32312 3476 32364 3528
rect 46480 3519 46532 3528
rect 46480 3485 46489 3519
rect 46489 3485 46523 3519
rect 46523 3485 46532 3519
rect 46480 3476 46532 3485
rect 32036 3383 32088 3392
rect 32036 3349 32045 3383
rect 32045 3349 32079 3383
rect 32079 3349 32088 3383
rect 32036 3340 32088 3349
rect 34704 3408 34756 3460
rect 35072 3340 35124 3392
rect 46664 3383 46716 3392
rect 46664 3349 46673 3383
rect 46673 3349 46707 3383
rect 46707 3349 46716 3383
rect 46664 3340 46716 3349
rect 47124 3383 47176 3392
rect 47124 3349 47133 3383
rect 47133 3349 47167 3383
rect 47167 3349 47176 3383
rect 47124 3340 47176 3349
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 39010 3238 39062 3290
rect 39074 3238 39126 3290
rect 39138 3238 39190 3290
rect 39202 3238 39254 3290
rect 39266 3238 39318 3290
rect 45010 3238 45062 3290
rect 45074 3238 45126 3290
rect 45138 3238 45190 3290
rect 45202 3238 45254 3290
rect 45266 3238 45318 3290
rect 6000 3136 6052 3188
rect 8668 3000 8720 3052
rect 13820 3136 13872 3188
rect 17776 3179 17828 3188
rect 17776 3145 17785 3179
rect 17785 3145 17819 3179
rect 17819 3145 17828 3179
rect 17776 3136 17828 3145
rect 14556 3111 14608 3120
rect 14556 3077 14565 3111
rect 14565 3077 14599 3111
rect 14599 3077 14608 3111
rect 14556 3068 14608 3077
rect 14740 3068 14792 3120
rect 17224 3000 17276 3052
rect 20812 3000 20864 3052
rect 45560 3136 45612 3188
rect 47308 3179 47360 3188
rect 47308 3145 47317 3179
rect 47317 3145 47351 3179
rect 47351 3145 47360 3179
rect 47308 3136 47360 3145
rect 27804 3068 27856 3120
rect 29368 3068 29420 3120
rect 32680 3068 32732 3120
rect 30656 3043 30708 3052
rect 30656 3009 30665 3043
rect 30665 3009 30699 3043
rect 30699 3009 30708 3043
rect 30656 3000 30708 3009
rect 31116 3043 31168 3052
rect 31116 3009 31125 3043
rect 31125 3009 31159 3043
rect 31159 3009 31168 3043
rect 31116 3000 31168 3009
rect 32036 3000 32088 3052
rect 43444 3068 43496 3120
rect 38844 3043 38896 3052
rect 38844 3009 38853 3043
rect 38853 3009 38887 3043
rect 38887 3009 38896 3043
rect 38844 3000 38896 3009
rect 41604 3000 41656 3052
rect 46664 3000 46716 3052
rect 46848 3000 46900 3052
rect 24676 2932 24728 2984
rect 7564 2864 7616 2916
rect 19156 2864 19208 2916
rect 27804 2864 27856 2916
rect 21824 2796 21876 2848
rect 27988 2839 28040 2848
rect 27988 2805 27997 2839
rect 27997 2805 28031 2839
rect 28031 2805 28040 2839
rect 27988 2796 28040 2805
rect 29736 2864 29788 2916
rect 45652 2864 45704 2916
rect 47952 2864 48004 2916
rect 28540 2796 28592 2848
rect 29184 2796 29236 2848
rect 30288 2796 30340 2848
rect 31024 2796 31076 2848
rect 33600 2796 33652 2848
rect 36268 2796 36320 2848
rect 38752 2796 38804 2848
rect 46940 2839 46992 2848
rect 46940 2805 46949 2839
rect 46949 2805 46983 2839
rect 46983 2805 46992 2839
rect 46940 2796 46992 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 37950 2694 38002 2746
rect 38014 2694 38066 2746
rect 38078 2694 38130 2746
rect 38142 2694 38194 2746
rect 38206 2694 38258 2746
rect 43950 2694 44002 2746
rect 44014 2694 44066 2746
rect 44078 2694 44130 2746
rect 44142 2694 44194 2746
rect 44206 2694 44258 2746
rect 15844 2592 15896 2644
rect 20628 2592 20680 2644
rect 15660 2524 15712 2576
rect 25596 2592 25648 2644
rect 22008 2524 22060 2576
rect 16028 2388 16080 2440
rect 20628 2431 20680 2440
rect 20628 2397 20637 2431
rect 20637 2397 20671 2431
rect 20671 2397 20680 2431
rect 20628 2388 20680 2397
rect 20720 2388 20772 2440
rect 23388 2456 23440 2508
rect 22100 2431 22152 2440
rect 22100 2397 22109 2431
rect 22109 2397 22143 2431
rect 22143 2397 22152 2431
rect 22100 2388 22152 2397
rect 22468 2431 22520 2440
rect 22468 2397 22477 2431
rect 22477 2397 22511 2431
rect 22511 2397 22520 2431
rect 22468 2388 22520 2397
rect 22836 2431 22888 2440
rect 22836 2397 22845 2431
rect 22845 2397 22879 2431
rect 22879 2397 22888 2431
rect 22836 2388 22888 2397
rect 23204 2431 23256 2440
rect 23204 2397 23213 2431
rect 23213 2397 23247 2431
rect 23247 2397 23256 2431
rect 23204 2388 23256 2397
rect 23572 2431 23624 2440
rect 23572 2397 23581 2431
rect 23581 2397 23615 2431
rect 23615 2397 23624 2431
rect 23572 2388 23624 2397
rect 10600 2320 10652 2372
rect 27896 2567 27948 2576
rect 27896 2533 27905 2567
rect 27905 2533 27939 2567
rect 27939 2533 27948 2567
rect 27896 2524 27948 2533
rect 28172 2524 28224 2576
rect 28356 2592 28408 2644
rect 30288 2592 30340 2644
rect 32864 2592 32916 2644
rect 35532 2592 35584 2644
rect 37648 2592 37700 2644
rect 47308 2635 47360 2644
rect 47308 2601 47317 2635
rect 47317 2601 47351 2635
rect 47351 2601 47360 2635
rect 47308 2592 47360 2601
rect 28816 2524 28868 2576
rect 29828 2524 29880 2576
rect 30104 2524 30156 2576
rect 30380 2524 30432 2576
rect 26884 2456 26936 2508
rect 24768 2388 24820 2440
rect 25044 2388 25096 2440
rect 25228 2431 25280 2440
rect 25228 2397 25237 2431
rect 25237 2397 25271 2431
rect 25271 2397 25280 2431
rect 25228 2388 25280 2397
rect 25596 2431 25648 2440
rect 25596 2397 25605 2431
rect 25605 2397 25639 2431
rect 25639 2397 25648 2431
rect 25596 2388 25648 2397
rect 25964 2431 26016 2440
rect 25964 2397 25973 2431
rect 25973 2397 26007 2431
rect 26007 2397 26016 2431
rect 25964 2388 26016 2397
rect 26332 2431 26384 2440
rect 26332 2397 26341 2431
rect 26341 2397 26375 2431
rect 26375 2397 26384 2431
rect 26332 2388 26384 2397
rect 26608 2388 26660 2440
rect 28264 2456 28316 2508
rect 30656 2524 30708 2576
rect 32588 2524 32640 2576
rect 34336 2524 34388 2576
rect 35808 2524 35860 2576
rect 36912 2524 36964 2576
rect 38384 2524 38436 2576
rect 39488 2524 39540 2576
rect 28540 2388 28592 2440
rect 28632 2388 28684 2440
rect 32128 2431 32180 2440
rect 32128 2397 32137 2431
rect 32137 2397 32171 2431
rect 32171 2397 32180 2431
rect 32128 2388 32180 2397
rect 32680 2388 32732 2440
rect 32772 2388 32824 2440
rect 37004 2456 37056 2508
rect 33508 2388 33560 2440
rect 33968 2431 34020 2440
rect 33968 2397 33977 2431
rect 33977 2397 34011 2431
rect 34011 2397 34020 2431
rect 33968 2388 34020 2397
rect 34704 2431 34756 2440
rect 34704 2397 34713 2431
rect 34713 2397 34747 2431
rect 34747 2397 34756 2431
rect 34704 2388 34756 2397
rect 35072 2431 35124 2440
rect 35072 2397 35081 2431
rect 35081 2397 35115 2431
rect 35115 2397 35124 2431
rect 35072 2388 35124 2397
rect 35440 2431 35492 2440
rect 35440 2397 35449 2431
rect 35449 2397 35483 2431
rect 35483 2397 35492 2431
rect 35440 2388 35492 2397
rect 35624 2388 35676 2440
rect 36176 2431 36228 2440
rect 36176 2397 36185 2431
rect 36185 2397 36219 2431
rect 36219 2397 36228 2431
rect 36176 2388 36228 2397
rect 36820 2431 36872 2440
rect 36820 2397 36829 2431
rect 36829 2397 36863 2431
rect 36863 2397 36872 2431
rect 36820 2388 36872 2397
rect 29552 2320 29604 2372
rect 20720 2252 20772 2304
rect 20904 2252 20956 2304
rect 21456 2252 21508 2304
rect 22192 2252 22244 2304
rect 22560 2252 22612 2304
rect 22928 2252 22980 2304
rect 23296 2252 23348 2304
rect 23664 2252 23716 2304
rect 24032 2252 24084 2304
rect 24400 2252 24452 2304
rect 25044 2295 25096 2304
rect 25044 2261 25053 2295
rect 25053 2261 25087 2295
rect 25087 2261 25096 2295
rect 25044 2252 25096 2261
rect 25136 2252 25188 2304
rect 25504 2252 25556 2304
rect 25872 2252 25924 2304
rect 26240 2252 26292 2304
rect 26608 2252 26660 2304
rect 27344 2252 27396 2304
rect 27712 2252 27764 2304
rect 28908 2252 28960 2304
rect 30104 2295 30156 2304
rect 30104 2261 30113 2295
rect 30113 2261 30147 2295
rect 30147 2261 30156 2295
rect 30104 2252 30156 2261
rect 31392 2320 31444 2372
rect 30564 2252 30616 2304
rect 32404 2320 32456 2372
rect 32680 2295 32732 2304
rect 32680 2261 32689 2295
rect 32689 2261 32723 2295
rect 32723 2261 32732 2295
rect 32680 2252 32732 2261
rect 35164 2320 35216 2372
rect 40316 2456 40368 2508
rect 40500 2456 40552 2508
rect 38016 2431 38068 2440
rect 38016 2397 38025 2431
rect 38025 2397 38059 2431
rect 38059 2397 38068 2431
rect 38016 2388 38068 2397
rect 38108 2388 38160 2440
rect 38476 2388 38528 2440
rect 38844 2388 38896 2440
rect 39212 2388 39264 2440
rect 40040 2388 40092 2440
rect 42800 2456 42852 2508
rect 46204 2456 46256 2508
rect 46388 2431 46440 2440
rect 46388 2397 46397 2431
rect 46397 2397 46431 2431
rect 46431 2397 46440 2431
rect 46388 2388 46440 2397
rect 47032 2388 47084 2440
rect 33508 2252 33560 2304
rect 34244 2252 34296 2304
rect 34980 2252 35032 2304
rect 36728 2252 36780 2304
rect 38200 2295 38252 2304
rect 38200 2261 38209 2295
rect 38209 2261 38243 2295
rect 38243 2261 38252 2295
rect 38200 2252 38252 2261
rect 38568 2252 38620 2304
rect 39396 2252 39448 2304
rect 45836 2295 45888 2304
rect 45836 2261 45845 2295
rect 45845 2261 45879 2295
rect 45879 2261 45888 2295
rect 45836 2252 45888 2261
rect 46204 2295 46256 2304
rect 46204 2261 46213 2295
rect 46213 2261 46247 2295
rect 46247 2261 46256 2295
rect 46204 2252 46256 2261
rect 46572 2295 46624 2304
rect 46572 2261 46581 2295
rect 46581 2261 46615 2295
rect 46615 2261 46624 2295
rect 46572 2252 46624 2261
rect 46940 2295 46992 2304
rect 46940 2261 46949 2295
rect 46949 2261 46983 2295
rect 46983 2261 46992 2295
rect 46940 2252 46992 2261
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 39010 2150 39062 2202
rect 39074 2150 39126 2202
rect 39138 2150 39190 2202
rect 39202 2150 39254 2202
rect 39266 2150 39318 2202
rect 45010 2150 45062 2202
rect 45074 2150 45126 2202
rect 45138 2150 45190 2202
rect 45202 2150 45254 2202
rect 45266 2150 45318 2202
rect 19156 2048 19208 2100
rect 10508 1980 10560 2032
rect 24124 1980 24176 2032
rect 27436 2048 27488 2100
rect 27896 2048 27948 2100
rect 29276 2048 29328 2100
rect 25964 1980 26016 2032
rect 30748 2048 30800 2100
rect 32772 2048 32824 2100
rect 32128 1980 32180 2032
rect 37188 1980 37240 2032
rect 40500 1980 40552 2032
rect 11428 1912 11480 1964
rect 24492 1912 24544 1964
rect 15752 1844 15804 1896
rect 25228 1912 25280 1964
rect 36544 1912 36596 1964
rect 43536 1912 43588 1964
rect 30012 1844 30064 1896
rect 46388 1844 46440 1896
rect 9588 1776 9640 1828
rect 26332 1776 26384 1828
rect 7748 1708 7800 1760
rect 23204 1708 23256 1760
rect 24124 1708 24176 1760
rect 30104 1776 30156 1828
rect 11336 1640 11388 1692
rect 28632 1640 28684 1692
rect 28724 1640 28776 1692
rect 28908 1640 28960 1692
rect 26424 1572 26476 1624
rect 36544 1572 36596 1624
rect 19432 1504 19484 1556
rect 35624 1504 35676 1556
rect 25320 1436 25372 1488
rect 38016 1436 38068 1488
rect 38108 1436 38160 1488
rect 38568 1436 38620 1488
rect 24492 1368 24544 1420
rect 30564 1368 30616 1420
rect 31760 1368 31812 1420
rect 32680 1368 32732 1420
rect 37280 1368 37332 1420
rect 38200 1368 38252 1420
rect 39580 1368 39632 1420
rect 41328 1368 41380 1420
rect 5724 1300 5776 1352
rect 22836 1300 22888 1352
rect 32496 1300 32548 1352
rect 32956 1300 33008 1352
rect 5540 1232 5592 1284
rect 22100 1232 22152 1284
rect 13360 620 13412 672
rect 24676 620 24728 672
rect 20352 552 20404 604
rect 32312 552 32364 604
rect 7104 484 7156 536
rect 23480 484 23532 536
rect 3424 416 3476 468
rect 20812 416 20864 468
rect 10784 348 10836 400
rect 29000 348 29052 400
rect 10416 280 10468 332
rect 29644 280 29696 332
rect 32956 280 33008 332
rect 41696 280 41748 332
rect 10048 212 10100 264
rect 29828 212 29880 264
rect 30932 212 30984 264
rect 42432 212 42484 264
rect 8944 144 8996 196
rect 9680 144 9732 196
rect 30472 144 30524 196
rect 31208 144 31260 196
rect 42800 144 42852 196
rect 31852 76 31904 128
rect 33784 76 33836 128
rect 41972 76 42024 128
rect 18236 8 18288 60
rect 44824 8 44876 60
<< metal2 >>
rect 1398 11194 1454 11250
rect 3698 11194 3754 11250
rect 5998 11194 6054 11250
rect 8298 11194 8354 11250
rect 10598 11194 10654 11250
rect 12898 11194 12954 11250
rect 15198 11194 15254 11250
rect 17498 11194 17554 11250
rect 19798 11194 19854 11250
rect 22098 11194 22154 11250
rect 24398 11194 24454 11250
rect 26698 11194 26754 11250
rect 28998 11194 29054 11250
rect 31298 11194 31354 11250
rect 33598 11194 33654 11250
rect 35898 11194 35954 11250
rect 38198 11194 38254 11250
rect 40498 11194 40554 11250
rect 42798 11194 42854 11250
rect 45098 11194 45154 11250
rect 45204 11206 45416 11234
rect 202 9888 258 9897
rect 202 9823 258 9832
rect 216 6497 244 9823
rect 1030 9344 1086 9353
rect 1030 9279 1086 9288
rect 1044 7886 1072 9279
rect 1412 8634 1440 11194
rect 2870 8800 2926 8809
rect 2870 8735 2926 8744
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 2884 8401 2912 8735
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 3712 8634 3740 11194
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 4080 8634 4108 8774
rect 6012 8634 6040 11194
rect 7562 9072 7618 9081
rect 7562 9007 7618 9016
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6656 8498 6684 8910
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 2870 8392 2926 8401
rect 2870 8327 2926 8336
rect 1766 8256 1822 8265
rect 1766 8191 1822 8200
rect 1032 7880 1084 7886
rect 1780 7857 1808 8191
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 7576 8022 7604 9007
rect 8312 8634 8340 11194
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 10612 8634 10640 11194
rect 12254 9616 12310 9625
rect 12254 9551 12310 9560
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 8404 8090 8432 8434
rect 10704 8090 10732 8434
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 7564 8016 7616 8022
rect 7564 7958 7616 7964
rect 11612 8016 11664 8022
rect 11612 7958 11664 7964
rect 11796 8016 11848 8022
rect 11796 7958 11848 7964
rect 10048 7880 10100 7886
rect 1032 7822 1084 7828
rect 1766 7848 1822 7857
rect 10048 7822 10100 7828
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 1766 7783 1822 7792
rect 3792 7812 3844 7818
rect 3792 7754 3844 7760
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 1584 7472 1636 7478
rect 1306 7440 1362 7449
rect 1584 7414 1636 7420
rect 1306 7375 1362 7384
rect 1320 6798 1348 7375
rect 1308 6792 1360 6798
rect 1308 6734 1360 6740
rect 202 6488 258 6497
rect 202 6423 258 6432
rect 1308 6248 1360 6254
rect 1308 6190 1360 6196
rect 480 6180 532 6186
rect 480 6122 532 6128
rect 492 4457 520 6122
rect 478 4448 534 4457
rect 478 4383 534 4392
rect 1124 4208 1176 4214
rect 1124 4150 1176 4156
rect 1136 1465 1164 4150
rect 1320 3913 1348 6190
rect 1306 3904 1362 3913
rect 1306 3839 1362 3848
rect 1216 3528 1268 3534
rect 1216 3470 1268 3476
rect 1228 2009 1256 3470
rect 1308 3392 1360 3398
rect 1308 3334 1360 3340
rect 1214 2000 1270 2009
rect 1214 1935 1270 1944
rect 1320 1737 1348 3334
rect 1306 1728 1362 1737
rect 1306 1663 1362 1672
rect 1122 1456 1178 1465
rect 1122 1391 1178 1400
rect 1596 56 1624 7414
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1766 4992 1822 5001
rect 1766 4927 1822 4936
rect 1780 4593 1808 4927
rect 1766 4584 1822 4593
rect 1766 4519 1822 4528
rect 1872 2530 1900 7278
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 2410 6488 2466 6497
rect 3010 6491 3318 6500
rect 2410 6423 2466 6432
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2424 5953 2452 6423
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 2410 5944 2466 5953
rect 2410 5879 2466 5888
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2320 4548 2372 4554
rect 2320 4490 2372 4496
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 1872 2502 1992 2530
rect 1964 56 1992 2502
rect 2332 56 2360 4490
rect 2412 4072 2464 4078
rect 2410 4040 2412 4049
rect 2464 4040 2466 4049
rect 2410 3975 2466 3984
rect 2608 82 2636 4558
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2792 4282 2820 4422
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 3436 626 3464 6258
rect 3344 598 3464 626
rect 2608 56 2728 82
rect 3068 56 3188 82
rect 1582 0 1638 56
rect 1950 0 2006 56
rect 2318 0 2374 56
rect 2608 54 2742 56
rect 2686 0 2742 54
rect 3054 54 3188 56
rect 3054 0 3110 54
rect 3160 42 3188 54
rect 3344 42 3372 598
rect 3424 468 3476 474
rect 3424 410 3476 416
rect 3436 56 3464 410
rect 3804 56 3832 7754
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4172 56 4200 7482
rect 10060 7410 10088 7822
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 10152 7342 10180 7822
rect 11624 7478 11652 7958
rect 11612 7472 11664 7478
rect 11612 7414 11664 7420
rect 11808 7410 11836 7958
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 7746 6760 7802 6769
rect 7746 6695 7802 6704
rect 5814 6488 5870 6497
rect 5814 6423 5870 6432
rect 4528 4684 4580 4690
rect 4528 4626 4580 4632
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4448 4214 4476 4422
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4540 56 4568 4626
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 4896 4548 4948 4554
rect 4896 4490 4948 4496
rect 4908 56 4936 4490
rect 5276 56 5304 4558
rect 5632 4548 5684 4554
rect 5632 4490 5684 4496
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5552 1290 5580 4422
rect 5540 1284 5592 1290
rect 5540 1226 5592 1232
rect 5644 56 5672 4490
rect 5724 4208 5776 4214
rect 5724 4150 5776 4156
rect 5736 1358 5764 4150
rect 5828 2417 5856 6423
rect 7760 5953 7788 6695
rect 8758 6624 8814 6633
rect 8758 6559 8814 6568
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7746 5944 7802 5953
rect 7950 5947 8258 5956
rect 8680 5914 8708 6394
rect 8772 6089 8800 6559
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 8850 6488 8906 6497
rect 9010 6491 9318 6500
rect 8850 6423 8906 6432
rect 8758 6080 8814 6089
rect 8758 6015 8814 6024
rect 7746 5879 7802 5888
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8864 5817 8892 6423
rect 11900 6361 11928 7686
rect 12162 7304 12218 7313
rect 12162 7239 12218 7248
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11886 6352 11942 6361
rect 11886 6287 11942 6296
rect 11518 6216 11574 6225
rect 11518 6151 11574 6160
rect 8666 5808 8722 5817
rect 8666 5743 8722 5752
rect 8850 5808 8906 5817
rect 8850 5743 8906 5752
rect 7654 5672 7710 5681
rect 7654 5607 7710 5616
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 5814 2408 5870 2417
rect 5814 2343 5870 2352
rect 5724 1352 5776 1358
rect 5724 1294 5776 1300
rect 6012 56 6040 3130
rect 6380 56 6408 3402
rect 6748 56 6776 4626
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7104 536 7156 542
rect 7104 478 7156 484
rect 7116 56 7144 478
rect 7484 56 7512 4558
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7576 2922 7604 3878
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7668 2553 7696 5607
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7654 2544 7710 2553
rect 7654 2479 7710 2488
rect 7760 1766 7788 4762
rect 8208 4548 8260 4554
rect 8208 4490 8260 4496
rect 8220 4214 8248 4490
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 7748 1760 7800 1766
rect 7748 1702 7800 1708
rect 7852 56 7880 4082
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 8312 3618 8340 4014
rect 8496 3670 8524 4966
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8220 3590 8340 3618
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8220 2938 8248 3590
rect 8220 2910 8340 2938
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 8312 2530 8340 2910
rect 8220 2502 8340 2530
rect 8220 56 8248 2502
rect 8588 56 8616 4082
rect 8680 3058 8708 5743
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 11532 5370 11560 6151
rect 11992 5681 12020 7142
rect 12176 5914 12204 7239
rect 12268 6730 12296 9551
rect 12912 8634 12940 11194
rect 15212 8922 15240 11194
rect 15212 8894 15424 8922
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 15396 8634 15424 8894
rect 17512 8634 17540 11194
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 19338 8528 19394 8537
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 17868 8492 17920 8498
rect 19338 8463 19394 8472
rect 17868 8434 17920 8440
rect 13004 7546 13032 8434
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 12346 7440 12402 7449
rect 12346 7375 12402 7384
rect 12360 6866 12388 7375
rect 14200 7342 14228 7822
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 15396 7546 15424 8434
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 12714 6488 12770 6497
rect 15010 6491 15318 6500
rect 12714 6423 12770 6432
rect 12728 6225 12756 6423
rect 12714 6216 12770 6225
rect 12714 6151 12770 6160
rect 13726 6080 13782 6089
rect 13726 6015 13782 6024
rect 12164 5908 12216 5914
rect 12164 5850 12216 5856
rect 12624 5704 12676 5710
rect 11978 5672 12034 5681
rect 12624 5646 12676 5652
rect 11978 5607 12034 5616
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 10428 4826 10456 5170
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 9600 1834 9628 4422
rect 10520 2038 10548 4966
rect 10612 2378 10640 4966
rect 11072 4214 11100 5238
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 10600 2372 10652 2378
rect 10600 2314 10652 2320
rect 10508 2032 10560 2038
rect 10508 1974 10560 1980
rect 9588 1828 9640 1834
rect 9588 1770 9640 1776
rect 11348 1698 11376 4966
rect 11440 1970 11468 5306
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 11888 5092 11940 5098
rect 11888 5034 11940 5040
rect 11428 1964 11480 1970
rect 11428 1906 11480 1912
rect 11518 1864 11574 1873
rect 11518 1799 11574 1808
rect 11336 1692 11388 1698
rect 11336 1634 11388 1640
rect 11150 504 11206 513
rect 11150 439 11206 448
rect 10784 400 10836 406
rect 10784 342 10836 348
rect 10416 332 10468 338
rect 10416 274 10468 280
rect 10048 264 10100 270
rect 9310 232 9366 241
rect 8944 196 8996 202
rect 10048 206 10100 212
rect 9310 167 9366 176
rect 9680 196 9732 202
rect 8944 138 8996 144
rect 8956 56 8984 138
rect 9324 56 9352 167
rect 9680 138 9732 144
rect 9692 56 9720 138
rect 10060 56 10088 206
rect 10428 56 10456 274
rect 10796 56 10824 342
rect 11164 56 11192 439
rect 11532 56 11560 1799
rect 11900 56 11928 5034
rect 12360 4758 12388 5170
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 12348 4752 12400 4758
rect 12348 4694 12400 4700
rect 12256 4208 12308 4214
rect 12256 4150 12308 4156
rect 12268 56 12296 4150
rect 12544 2553 12572 5034
rect 12530 2544 12586 2553
rect 12530 2479 12586 2488
rect 12636 56 12664 5646
rect 13740 5098 13768 6015
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 14280 5160 14332 5166
rect 13818 5128 13874 5137
rect 13728 5092 13780 5098
rect 14280 5102 14332 5108
rect 13818 5063 13874 5072
rect 13728 5034 13780 5040
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 3160 14 3372 42
rect 3422 0 3478 56
rect 3790 0 3846 56
rect 4158 0 4214 56
rect 4526 0 4582 56
rect 4894 0 4950 56
rect 5262 0 5318 56
rect 5630 0 5686 56
rect 5998 0 6054 56
rect 6366 0 6422 56
rect 6734 0 6790 56
rect 7102 0 7158 56
rect 7470 0 7526 56
rect 7838 0 7894 56
rect 8206 0 8262 56
rect 8574 0 8630 56
rect 8942 0 8998 56
rect 9310 0 9366 56
rect 9678 0 9734 56
rect 10046 0 10102 56
rect 10414 0 10470 56
rect 10782 0 10838 56
rect 11150 0 11206 56
rect 11518 0 11574 56
rect 11886 0 11942 56
rect 12254 0 12310 56
rect 12622 0 12678 56
rect 12728 42 12756 4966
rect 12912 2417 12940 4966
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 12898 2408 12954 2417
rect 12898 2343 12954 2352
rect 13360 672 13412 678
rect 13360 614 13412 620
rect 12912 56 13032 82
rect 13372 56 13400 614
rect 13740 56 13768 4762
rect 13832 3194 13860 5063
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 14292 3074 14320 5102
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14554 3768 14610 3777
rect 14554 3703 14610 3712
rect 14568 3126 14596 3703
rect 14752 3398 14780 4762
rect 14832 4752 14884 4758
rect 14832 4694 14884 4700
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 13832 3046 14320 3074
rect 14556 3120 14608 3126
rect 14556 3062 14608 3068
rect 14740 3120 14792 3126
rect 14740 3062 14792 3068
rect 12912 54 13046 56
rect 12912 42 12940 54
rect 12728 14 12940 42
rect 12990 0 13046 54
rect 13358 0 13414 56
rect 13726 0 13782 56
rect 13832 42 13860 3046
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 14016 56 14136 82
rect 14476 56 14596 82
rect 14016 54 14150 56
rect 14016 42 14044 54
rect 13832 14 14044 42
rect 14094 0 14150 54
rect 14462 54 14596 56
rect 14462 0 14518 54
rect 14568 42 14596 54
rect 14752 42 14780 3062
rect 14844 56 14872 4694
rect 14936 1737 14964 5510
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 15476 5296 15528 5302
rect 15476 5238 15528 5244
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 15396 3738 15424 4966
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 15010 3227 15318 3236
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 14922 1728 14978 1737
rect 14922 1663 14978 1672
rect 15212 56 15332 82
rect 14568 14 14780 42
rect 14830 0 14886 56
rect 15198 54 15332 56
rect 15198 0 15254 54
rect 15304 42 15332 54
rect 15488 42 15516 5238
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 15580 56 15608 5102
rect 15844 4208 15896 4214
rect 15844 4150 15896 4156
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15672 2582 15700 3878
rect 15660 2576 15712 2582
rect 15660 2518 15712 2524
rect 15764 1902 15792 4014
rect 15856 2650 15884 4150
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 15752 1896 15804 1902
rect 15752 1838 15804 1844
rect 15948 56 15976 5646
rect 16040 2446 16068 7686
rect 17880 7546 17908 8434
rect 19352 7886 19380 8463
rect 19536 8090 19564 9114
rect 19812 8634 19840 11194
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 22112 8634 22140 11194
rect 23940 8900 23992 8906
rect 23940 8842 23992 8848
rect 19800 8628 19852 8634
rect 19800 8570 19852 8576
rect 22100 8628 22152 8634
rect 22100 8570 22152 8576
rect 22192 8560 22244 8566
rect 22192 8502 22244 8508
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 19950 8188 20258 8197
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 20640 8090 20668 8434
rect 21730 8392 21786 8401
rect 21730 8327 21786 8336
rect 21744 8090 21772 8327
rect 22204 8090 22232 8502
rect 23480 8492 23532 8498
rect 23480 8434 23532 8440
rect 23492 8090 23520 8434
rect 23952 8090 23980 8842
rect 24412 8634 24440 11194
rect 26516 8832 26568 8838
rect 26516 8774 26568 8780
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 25872 8492 25924 8498
rect 25872 8434 25924 8440
rect 25884 8090 25912 8434
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 26528 8090 26556 8774
rect 26712 8634 26740 11194
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 29012 8634 29040 11194
rect 31312 8634 31340 11194
rect 33010 8732 33318 8741
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 33010 8667 33318 8676
rect 33612 8634 33640 11194
rect 33876 9240 33928 9246
rect 33876 9182 33928 9188
rect 26700 8628 26752 8634
rect 26700 8570 26752 8576
rect 29000 8628 29052 8634
rect 29000 8570 29052 8576
rect 31300 8628 31352 8634
rect 31300 8570 31352 8576
rect 33600 8628 33652 8634
rect 33600 8570 33652 8576
rect 33888 8498 33916 9182
rect 33968 9104 34020 9110
rect 33968 9046 34020 9052
rect 33980 8498 34008 9046
rect 35912 8634 35940 11194
rect 37280 9036 37332 9042
rect 37280 8978 37332 8984
rect 34060 8628 34112 8634
rect 34060 8570 34112 8576
rect 35900 8628 35952 8634
rect 35900 8570 35952 8576
rect 34072 8514 34100 8570
rect 34244 8560 34296 8566
rect 34072 8508 34244 8514
rect 34072 8502 34296 8508
rect 29276 8492 29328 8498
rect 29276 8434 29328 8440
rect 29368 8492 29420 8498
rect 29368 8434 29420 8440
rect 33876 8492 33928 8498
rect 33876 8434 33928 8440
rect 33968 8492 34020 8498
rect 34072 8486 34284 8502
rect 37188 8492 37240 8498
rect 33968 8434 34020 8440
rect 37188 8434 37240 8440
rect 29288 8294 29316 8434
rect 29276 8288 29328 8294
rect 29276 8230 29328 8236
rect 29380 8090 29408 8434
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 20536 8084 20588 8090
rect 20536 8026 20588 8032
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 21732 8084 21784 8090
rect 21732 8026 21784 8032
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 23940 8084 23992 8090
rect 23940 8026 23992 8032
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 26516 8084 26568 8090
rect 26516 8026 26568 8032
rect 29368 8084 29420 8090
rect 29368 8026 29420 8032
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 20364 7478 20392 7822
rect 20548 7546 20576 8026
rect 25594 7984 25650 7993
rect 25594 7919 25650 7928
rect 26330 7984 26386 7993
rect 26330 7919 26386 7928
rect 25608 7886 25636 7919
rect 26344 7886 26372 7919
rect 20812 7880 20864 7886
rect 23756 7880 23808 7886
rect 20812 7822 20864 7828
rect 23754 7848 23756 7857
rect 25596 7880 25648 7886
rect 23808 7848 23810 7857
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20352 7472 20404 7478
rect 20352 7414 20404 7420
rect 18052 7404 18104 7410
rect 18052 7346 18104 7352
rect 18064 6390 18092 7346
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 19246 6896 19302 6905
rect 19246 6831 19302 6840
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 18052 6384 18104 6390
rect 18052 6326 18104 6332
rect 18418 6352 18474 6361
rect 18418 6287 18474 6296
rect 17958 5264 18014 5273
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 17408 5228 17460 5234
rect 17958 5199 18014 5208
rect 17408 5170 17460 5176
rect 16224 2774 16252 5170
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 16488 4276 16540 4282
rect 16488 4218 16540 4224
rect 16500 3602 16528 4218
rect 16592 4214 16620 4626
rect 16580 4208 16632 4214
rect 16580 4150 16632 4156
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16224 2746 16344 2774
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 16316 56 16344 2746
rect 16684 56 16712 5170
rect 17052 56 17080 5170
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17144 1601 17172 4966
rect 17236 4758 17264 4966
rect 17224 4752 17276 4758
rect 17224 4694 17276 4700
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17236 3058 17264 3334
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17130 1592 17186 1601
rect 17130 1527 17186 1536
rect 17420 56 17448 5170
rect 17868 5024 17920 5030
rect 17774 4992 17830 5001
rect 17868 4966 17920 4972
rect 17774 4927 17830 4936
rect 17788 3194 17816 4927
rect 17880 4826 17908 4966
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17972 2961 18000 5199
rect 18432 4214 18460 6287
rect 18984 5778 19012 6598
rect 19260 5914 19288 6831
rect 19614 6352 19670 6361
rect 19614 6287 19670 6296
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 18972 5772 19024 5778
rect 18972 5714 19024 5720
rect 18972 5636 19024 5642
rect 18972 5578 19024 5584
rect 18604 5092 18656 5098
rect 18604 5034 18656 5040
rect 18420 4208 18472 4214
rect 18420 4150 18472 4156
rect 17958 2952 18014 2961
rect 17958 2887 18014 2896
rect 18616 2009 18644 5034
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18892 3670 18920 3878
rect 18880 3664 18932 3670
rect 18880 3606 18932 3612
rect 18984 2774 19012 5578
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19156 2916 19208 2922
rect 19156 2858 19208 2864
rect 18892 2746 19012 2774
rect 18602 2000 18658 2009
rect 18602 1935 18658 1944
rect 18510 368 18566 377
rect 18510 303 18566 312
rect 17774 96 17830 105
rect 15304 14 15516 42
rect 15566 0 15622 56
rect 15934 0 15990 56
rect 16302 0 16358 56
rect 16670 0 16726 56
rect 17038 0 17094 56
rect 17406 0 17462 56
rect 18156 66 18276 82
rect 18156 60 18288 66
rect 18156 56 18236 60
rect 17774 0 17830 40
rect 18142 54 18236 56
rect 18142 0 18198 54
rect 18524 56 18552 303
rect 18892 56 18920 2746
rect 19168 2106 19196 2858
rect 19156 2100 19208 2106
rect 19156 2042 19208 2048
rect 19260 56 19288 4558
rect 19340 4548 19392 4554
rect 19340 4490 19392 4496
rect 19352 3777 19380 4490
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19338 3768 19394 3777
rect 19338 3703 19394 3712
rect 19444 1562 19472 4422
rect 19432 1556 19484 1562
rect 19432 1498 19484 1504
rect 19628 56 19656 6287
rect 20732 6066 20760 7686
rect 20824 7478 20852 7822
rect 23388 7812 23440 7818
rect 25596 7822 25648 7828
rect 26240 7880 26292 7886
rect 26240 7822 26292 7828
rect 26332 7880 26384 7886
rect 26332 7822 26384 7828
rect 26516 7880 26568 7886
rect 26516 7822 26568 7828
rect 29920 7880 29972 7886
rect 29920 7822 29972 7828
rect 23754 7783 23810 7792
rect 24952 7812 25004 7818
rect 23388 7754 23440 7760
rect 24952 7754 25004 7760
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 20812 7472 20864 7478
rect 20812 7414 20864 7420
rect 22928 7200 22980 7206
rect 22928 7142 22980 7148
rect 23296 7200 23348 7206
rect 23296 7142 23348 7148
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 20732 6038 20852 6066
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 20628 4208 20680 4214
rect 20628 4150 20680 4156
rect 20640 4026 20668 4150
rect 20732 4146 20760 5850
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 20640 3998 20760 4026
rect 19950 3836 20258 3845
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 20352 3596 20404 3602
rect 20352 3538 20404 3544
rect 19950 2748 20258 2757
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 20364 762 20392 3538
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 20640 2446 20668 2586
rect 20732 2446 20760 3998
rect 20824 3058 20852 6038
rect 22008 5704 22060 5710
rect 22008 5646 22060 5652
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 21730 5400 21786 5409
rect 22020 5370 22048 5646
rect 21730 5335 21786 5344
rect 22008 5364 22060 5370
rect 21640 5296 21692 5302
rect 21640 5238 21692 5244
rect 21652 4826 21680 5238
rect 21744 5234 21772 5335
rect 22008 5306 22060 5312
rect 21732 5228 21784 5234
rect 21732 5170 21784 5176
rect 21640 4820 21692 4826
rect 21640 4762 21692 4768
rect 20904 4616 20956 4622
rect 22940 4593 22968 7142
rect 23308 7002 23336 7142
rect 23296 6996 23348 7002
rect 23296 6938 23348 6944
rect 23296 6452 23348 6458
rect 23296 6394 23348 6400
rect 23204 5024 23256 5030
rect 23204 4966 23256 4972
rect 23216 4690 23244 4966
rect 23204 4684 23256 4690
rect 23204 4626 23256 4632
rect 20904 4558 20956 4564
rect 22926 4584 22982 4593
rect 20812 3052 20864 3058
rect 20812 2994 20864 3000
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 20720 2440 20772 2446
rect 20916 2394 20944 4558
rect 22926 4519 22982 4528
rect 22008 4480 22060 4486
rect 22008 4422 22060 4428
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 21824 2848 21876 2854
rect 21824 2790 21876 2796
rect 20720 2382 20772 2388
rect 20824 2366 20944 2394
rect 20720 2304 20772 2310
rect 20720 2246 20772 2252
rect 20272 734 20392 762
rect 19996 56 20116 82
rect 18236 2 18288 8
rect 18510 0 18566 56
rect 18878 0 18934 56
rect 19246 0 19302 56
rect 19614 0 19670 56
rect 19982 54 20116 56
rect 19982 0 20038 54
rect 20088 42 20116 54
rect 20272 42 20300 734
rect 20352 604 20404 610
rect 20352 546 20404 552
rect 20364 56 20392 546
rect 20732 56 20760 2246
rect 20824 474 20852 2366
rect 20904 2304 20956 2310
rect 20904 2246 20956 2252
rect 21456 2304 21508 2310
rect 21456 2246 21508 2252
rect 20812 468 20864 474
rect 20812 410 20864 416
rect 20088 14 20300 42
rect 20350 0 20406 56
rect 20718 0 20774 56
rect 20916 42 20944 2246
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 21008 56 21128 82
rect 21468 56 21496 2246
rect 21836 56 21864 2790
rect 22020 2582 22048 4422
rect 22468 4072 22520 4078
rect 22468 4014 22520 4020
rect 22008 2576 22060 2582
rect 22008 2518 22060 2524
rect 22480 2446 22508 4014
rect 23308 4010 23336 6394
rect 23296 4004 23348 4010
rect 23296 3946 23348 3952
rect 23400 2514 23428 7754
rect 24676 7744 24728 7750
rect 24676 7686 24728 7692
rect 23572 7540 23624 7546
rect 23572 7482 23624 7488
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 23388 2508 23440 2514
rect 23388 2450 23440 2456
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 22468 2440 22520 2446
rect 22468 2382 22520 2388
rect 22836 2440 22888 2446
rect 22836 2382 22888 2388
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 22112 1290 22140 2382
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 22100 1284 22152 1290
rect 22100 1226 22152 1232
rect 22204 56 22232 2246
rect 22572 56 22600 2246
rect 22848 1358 22876 2382
rect 22928 2304 22980 2310
rect 22928 2246 22980 2252
rect 22836 1352 22888 1358
rect 22836 1294 22888 1300
rect 22940 56 22968 2246
rect 23216 1766 23244 2382
rect 23296 2304 23348 2310
rect 23296 2246 23348 2252
rect 23204 1760 23256 1766
rect 23204 1702 23256 1708
rect 23308 56 23336 2246
rect 23492 542 23520 4966
rect 23584 2446 23612 7482
rect 24688 5846 24716 7686
rect 24768 6112 24820 6118
rect 24768 6054 24820 6060
rect 24676 5840 24728 5846
rect 24676 5782 24728 5788
rect 24030 5400 24086 5409
rect 24030 5335 24086 5344
rect 24044 5234 24072 5335
rect 24032 5228 24084 5234
rect 24032 5170 24084 5176
rect 24676 2984 24728 2990
rect 24676 2926 24728 2932
rect 23572 2440 23624 2446
rect 23572 2382 23624 2388
rect 23664 2304 23716 2310
rect 23664 2246 23716 2252
rect 24032 2304 24084 2310
rect 24032 2246 24084 2252
rect 24400 2304 24452 2310
rect 24400 2246 24452 2252
rect 23480 536 23532 542
rect 23480 478 23532 484
rect 23676 56 23704 2246
rect 24044 56 24072 2246
rect 24124 2032 24176 2038
rect 24124 1974 24176 1980
rect 24136 1766 24164 1974
rect 24124 1760 24176 1766
rect 24124 1702 24176 1708
rect 24412 56 24440 2246
rect 24492 1964 24544 1970
rect 24492 1906 24544 1912
rect 24504 1426 24532 1906
rect 24492 1420 24544 1426
rect 24492 1362 24544 1368
rect 24688 678 24716 2926
rect 24780 2446 24808 6054
rect 24964 2961 24992 7754
rect 26252 7426 26280 7822
rect 26252 7398 26464 7426
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 25872 6656 25924 6662
rect 25872 6598 25924 6604
rect 26332 6656 26384 6662
rect 26332 6598 26384 6604
rect 25320 4752 25372 4758
rect 25884 4729 25912 6598
rect 26344 6458 26372 6598
rect 26332 6452 26384 6458
rect 26332 6394 26384 6400
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 25320 4694 25372 4700
rect 25870 4720 25926 4729
rect 25044 3664 25096 3670
rect 25044 3606 25096 3612
rect 24950 2952 25006 2961
rect 24950 2887 25006 2896
rect 25056 2446 25084 3606
rect 24768 2440 24820 2446
rect 24768 2382 24820 2388
rect 25044 2440 25096 2446
rect 25044 2382 25096 2388
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 25044 2304 25096 2310
rect 24780 2252 25044 2258
rect 24780 2246 25096 2252
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 24780 2230 25084 2246
rect 24676 672 24728 678
rect 24676 614 24728 620
rect 24780 56 24808 2230
rect 25148 56 25176 2246
rect 25240 1970 25268 2382
rect 25228 1964 25280 1970
rect 25228 1906 25280 1912
rect 25332 1494 25360 4694
rect 25870 4655 25926 4664
rect 25872 4208 25924 4214
rect 25872 4150 25924 4156
rect 25884 3097 25912 4150
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 25870 3088 25926 3097
rect 25870 3023 25926 3032
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 25596 2644 25648 2650
rect 25596 2586 25648 2592
rect 25608 2446 25636 2586
rect 25596 2440 25648 2446
rect 25596 2382 25648 2388
rect 25964 2440 26016 2446
rect 25964 2382 26016 2388
rect 26332 2440 26384 2446
rect 26332 2382 26384 2388
rect 25504 2304 25556 2310
rect 25504 2246 25556 2252
rect 25872 2304 25924 2310
rect 25872 2246 25924 2252
rect 25320 1488 25372 1494
rect 25320 1430 25372 1436
rect 25516 56 25544 2246
rect 25884 56 25912 2246
rect 25976 2038 26004 2382
rect 26240 2304 26292 2310
rect 26240 2246 26292 2252
rect 25964 2032 26016 2038
rect 25964 1974 26016 1980
rect 26252 56 26280 2246
rect 26344 1834 26372 2382
rect 26332 1828 26384 1834
rect 26332 1770 26384 1776
rect 26436 1630 26464 7398
rect 26528 6254 26556 7822
rect 29736 7744 29788 7750
rect 29736 7686 29788 7692
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 29748 7546 29776 7686
rect 29736 7540 29788 7546
rect 29736 7482 29788 7488
rect 27620 7200 27672 7206
rect 27620 7142 27672 7148
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 26516 6248 26568 6254
rect 26516 6190 26568 6196
rect 27632 6186 27660 7142
rect 27620 6180 27672 6186
rect 27620 6122 27672 6128
rect 27528 5704 27580 5710
rect 27528 5646 27580 5652
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 26608 5296 26660 5302
rect 26608 5238 26660 5244
rect 26620 2446 26648 5238
rect 26976 5228 27028 5234
rect 26976 5170 27028 5176
rect 26988 5137 27016 5170
rect 26974 5128 27030 5137
rect 27540 5098 27568 5646
rect 26974 5063 27030 5072
rect 27528 5092 27580 5098
rect 27528 5034 27580 5040
rect 26884 5024 26936 5030
rect 26884 4966 26936 4972
rect 27436 5024 27488 5030
rect 27436 4966 27488 4972
rect 29644 5024 29696 5030
rect 29644 4966 29696 4972
rect 26700 4480 26752 4486
rect 26700 4422 26752 4428
rect 26712 4282 26740 4422
rect 26700 4276 26752 4282
rect 26700 4218 26752 4224
rect 26792 4276 26844 4282
rect 26792 4218 26844 4224
rect 26804 3505 26832 4218
rect 26790 3496 26846 3505
rect 26790 3431 26846 3440
rect 26896 2514 26924 4966
rect 27448 4690 27476 4966
rect 29656 4758 29684 4966
rect 29644 4752 29696 4758
rect 29644 4694 29696 4700
rect 27436 4684 27488 4690
rect 27436 4626 27488 4632
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 28264 3936 28316 3942
rect 28264 3878 28316 3884
rect 28172 3460 28224 3466
rect 28172 3402 28224 3408
rect 27528 3392 27580 3398
rect 27528 3334 27580 3340
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 26884 2508 26936 2514
rect 26884 2450 26936 2456
rect 26608 2440 26660 2446
rect 26608 2382 26660 2388
rect 26608 2304 26660 2310
rect 26608 2246 26660 2252
rect 27344 2304 27396 2310
rect 27344 2246 27396 2252
rect 26424 1624 26476 1630
rect 26424 1566 26476 1572
rect 26620 56 26648 2246
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 27356 354 27384 2246
rect 27436 2100 27488 2106
rect 27436 2042 27488 2048
rect 27264 326 27384 354
rect 26988 56 27108 82
rect 21008 54 21142 56
rect 21008 42 21036 54
rect 20916 14 21036 42
rect 21086 0 21142 54
rect 21454 0 21510 56
rect 21822 0 21878 56
rect 22190 0 22246 56
rect 22558 0 22614 56
rect 22926 0 22982 56
rect 23294 0 23350 56
rect 23662 0 23718 56
rect 24030 0 24086 56
rect 24398 0 24454 56
rect 24766 0 24822 56
rect 25134 0 25190 56
rect 25502 0 25558 56
rect 25870 0 25926 56
rect 26238 0 26294 56
rect 26606 0 26662 56
rect 26974 54 27108 56
rect 26974 0 27030 54
rect 27080 42 27108 54
rect 27264 42 27292 326
rect 27448 218 27476 2042
rect 27540 513 27568 3334
rect 27804 3120 27856 3126
rect 27804 3062 27856 3068
rect 27816 2922 27844 3062
rect 27804 2916 27856 2922
rect 27804 2858 27856 2864
rect 27988 2848 28040 2854
rect 27988 2790 28040 2796
rect 27896 2576 27948 2582
rect 27896 2518 27948 2524
rect 27712 2304 27764 2310
rect 27712 2246 27764 2252
rect 27526 504 27582 513
rect 27526 439 27582 448
rect 27356 190 27476 218
rect 27356 56 27384 190
rect 27724 56 27752 2246
rect 27908 2106 27936 2518
rect 27896 2100 27948 2106
rect 27896 2042 27948 2048
rect 28000 1873 28028 2790
rect 28184 2582 28212 3402
rect 28172 2576 28224 2582
rect 28172 2518 28224 2524
rect 28276 2514 28304 3878
rect 29828 3664 29880 3670
rect 29828 3606 29880 3612
rect 29000 3528 29052 3534
rect 29000 3470 29052 3476
rect 29644 3528 29696 3534
rect 29644 3470 29696 3476
rect 28540 2848 28592 2854
rect 28540 2790 28592 2796
rect 28356 2644 28408 2650
rect 28356 2586 28408 2592
rect 28264 2508 28316 2514
rect 28264 2450 28316 2456
rect 27986 1864 28042 1873
rect 27986 1799 28042 1808
rect 28092 56 28212 82
rect 27080 14 27292 42
rect 27342 0 27398 56
rect 27710 0 27766 56
rect 28078 54 28212 56
rect 28078 0 28134 54
rect 28184 42 28212 54
rect 28368 42 28396 2586
rect 28552 2446 28580 2790
rect 28816 2576 28868 2582
rect 28816 2518 28868 2524
rect 28540 2440 28592 2446
rect 28540 2382 28592 2388
rect 28632 2440 28684 2446
rect 28632 2382 28684 2388
rect 28644 1698 28672 2382
rect 28632 1692 28684 1698
rect 28632 1634 28684 1640
rect 28724 1692 28776 1698
rect 28724 1634 28776 1640
rect 28460 56 28580 82
rect 28184 14 28396 42
rect 28446 54 28580 56
rect 28446 0 28502 54
rect 28552 42 28580 54
rect 28736 42 28764 1634
rect 28828 56 28856 2518
rect 28908 2304 28960 2310
rect 28908 2246 28960 2252
rect 28920 1698 28948 2246
rect 28908 1692 28960 1698
rect 28908 1634 28960 1640
rect 29012 406 29040 3470
rect 29276 3392 29328 3398
rect 29276 3334 29328 3340
rect 29368 3392 29420 3398
rect 29368 3334 29420 3340
rect 29184 2848 29236 2854
rect 29184 2790 29236 2796
rect 29000 400 29052 406
rect 29000 342 29052 348
rect 29196 56 29224 2790
rect 29288 2106 29316 3334
rect 29380 3126 29408 3334
rect 29368 3120 29420 3126
rect 29368 3062 29420 3068
rect 29552 2372 29604 2378
rect 29552 2314 29604 2320
rect 29276 2100 29328 2106
rect 29276 2042 29328 2048
rect 29564 56 29592 2314
rect 29656 338 29684 3470
rect 29840 3466 29868 3606
rect 29828 3460 29880 3466
rect 29828 3402 29880 3408
rect 29734 3088 29790 3097
rect 29734 3023 29790 3032
rect 29748 2922 29776 3023
rect 29736 2916 29788 2922
rect 29736 2858 29788 2864
rect 29828 2576 29880 2582
rect 29828 2518 29880 2524
rect 29644 332 29696 338
rect 29644 274 29696 280
rect 29840 270 29868 2518
rect 29932 513 29960 7822
rect 36544 7812 36596 7818
rect 36544 7754 36596 7760
rect 30472 7744 30524 7750
rect 30472 7686 30524 7692
rect 36176 7744 36228 7750
rect 36176 7686 36228 7692
rect 30378 6352 30434 6361
rect 30378 6287 30380 6296
rect 30432 6287 30434 6296
rect 30380 6258 30432 6264
rect 30484 5642 30512 7686
rect 33010 7644 33318 7653
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 31208 7472 31260 7478
rect 31208 7414 31260 7420
rect 30932 6384 30984 6390
rect 30932 6326 30984 6332
rect 30472 5636 30524 5642
rect 30472 5578 30524 5584
rect 30010 4040 30066 4049
rect 30010 3975 30066 3984
rect 30656 4004 30708 4010
rect 30024 1902 30052 3975
rect 30656 3946 30708 3952
rect 30104 3528 30156 3534
rect 30104 3470 30156 3476
rect 30116 2582 30144 3470
rect 30380 3392 30432 3398
rect 30380 3334 30432 3340
rect 30472 3392 30524 3398
rect 30472 3334 30524 3340
rect 30288 2848 30340 2854
rect 30208 2808 30288 2836
rect 30104 2576 30156 2582
rect 30104 2518 30156 2524
rect 30104 2304 30156 2310
rect 30104 2246 30156 2252
rect 30012 1896 30064 1902
rect 30012 1838 30064 1844
rect 30116 1834 30144 2246
rect 30104 1828 30156 1834
rect 30104 1770 30156 1776
rect 29918 504 29974 513
rect 29918 439 29974 448
rect 29828 264 29880 270
rect 29828 206 29880 212
rect 29932 56 30052 82
rect 28552 14 28764 42
rect 28814 0 28870 56
rect 29182 0 29238 56
rect 29550 0 29606 56
rect 29918 54 30052 56
rect 29918 0 29974 54
rect 30024 42 30052 54
rect 30208 42 30236 2808
rect 30288 2790 30340 2796
rect 30288 2644 30340 2650
rect 30288 2586 30340 2592
rect 30300 56 30328 2586
rect 30392 2582 30420 3334
rect 30380 2576 30432 2582
rect 30380 2518 30432 2524
rect 30484 202 30512 3334
rect 30668 3058 30696 3946
rect 30840 3936 30892 3942
rect 30840 3878 30892 3884
rect 30748 3460 30800 3466
rect 30748 3402 30800 3408
rect 30656 3052 30708 3058
rect 30656 2994 30708 3000
rect 30656 2576 30708 2582
rect 30656 2518 30708 2524
rect 30564 2304 30616 2310
rect 30564 2246 30616 2252
rect 30576 1426 30604 2246
rect 30564 1420 30616 1426
rect 30564 1362 30616 1368
rect 30472 196 30524 202
rect 30472 138 30524 144
rect 30668 56 30696 2518
rect 30760 2106 30788 3402
rect 30852 3398 30880 3878
rect 30840 3392 30892 3398
rect 30840 3334 30892 3340
rect 30748 2100 30800 2106
rect 30748 2042 30800 2048
rect 30944 270 30972 6326
rect 31114 3088 31170 3097
rect 31114 3023 31116 3032
rect 31168 3023 31170 3032
rect 31116 2994 31168 3000
rect 31024 2848 31076 2854
rect 31024 2790 31076 2796
rect 30932 264 30984 270
rect 30932 206 30984 212
rect 31036 56 31064 2790
rect 31220 202 31248 7414
rect 33784 7336 33836 7342
rect 33784 7278 33836 7284
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 33010 6556 33318 6565
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 32770 5808 32826 5817
rect 32770 5743 32826 5752
rect 32784 5710 32812 5743
rect 32772 5704 32824 5710
rect 32494 5672 32550 5681
rect 32772 5646 32824 5652
rect 32494 5607 32550 5616
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 31760 4820 31812 4826
rect 31760 4762 31812 4768
rect 31772 4622 31800 4762
rect 31760 4616 31812 4622
rect 31760 4558 31812 4564
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 31300 3528 31352 3534
rect 31300 3470 31352 3476
rect 31852 3528 31904 3534
rect 31852 3470 31904 3476
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 31312 241 31340 3470
rect 31392 2372 31444 2378
rect 31392 2314 31444 2320
rect 31298 232 31354 241
rect 31208 196 31260 202
rect 31298 167 31354 176
rect 31208 138 31260 144
rect 31404 56 31432 2314
rect 31760 1420 31812 1426
rect 31760 1362 31812 1368
rect 31772 56 31800 1362
rect 31864 134 31892 3470
rect 32036 3392 32088 3398
rect 32036 3334 32088 3340
rect 32048 3058 32076 3334
rect 32036 3052 32088 3058
rect 32036 2994 32088 3000
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 32128 2440 32180 2446
rect 32128 2382 32180 2388
rect 32140 2038 32168 2382
rect 32128 2032 32180 2038
rect 32128 1974 32180 1980
rect 32324 610 32352 3470
rect 32404 2372 32456 2378
rect 32404 2314 32456 2320
rect 32312 604 32364 610
rect 32312 546 32364 552
rect 31852 128 31904 134
rect 31852 70 31904 76
rect 32140 56 32260 82
rect 30024 14 30236 42
rect 30286 0 30342 56
rect 30654 0 30710 56
rect 31022 0 31078 56
rect 31390 0 31446 56
rect 31758 0 31814 56
rect 32126 54 32260 56
rect 32126 0 32182 54
rect 32232 42 32260 54
rect 32416 42 32444 2314
rect 32508 1358 32536 5607
rect 33010 5468 33318 5477
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 33010 5403 33318 5412
rect 33010 4380 33318 4389
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 33508 3936 33560 3942
rect 33508 3878 33560 3884
rect 33010 3292 33318 3301
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 32680 3120 32732 3126
rect 32680 3062 32732 3068
rect 32588 2576 32640 2582
rect 32588 2518 32640 2524
rect 32496 1352 32548 1358
rect 32496 1294 32548 1300
rect 32600 1170 32628 2518
rect 32692 2446 32720 3062
rect 32864 2644 32916 2650
rect 32864 2586 32916 2592
rect 32680 2440 32732 2446
rect 32680 2382 32732 2388
rect 32772 2440 32824 2446
rect 32772 2382 32824 2388
rect 32680 2304 32732 2310
rect 32680 2246 32732 2252
rect 32692 1426 32720 2246
rect 32784 2106 32812 2382
rect 32772 2100 32824 2106
rect 32772 2042 32824 2048
rect 32680 1420 32732 1426
rect 32680 1362 32732 1368
rect 32508 1142 32628 1170
rect 32508 56 32536 1142
rect 32876 56 32904 2586
rect 33520 2446 33548 3878
rect 33600 2848 33652 2854
rect 33600 2790 33652 2796
rect 33508 2440 33560 2446
rect 33508 2382 33560 2388
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 33010 2204 33318 2213
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 32956 1352 33008 1358
rect 32956 1294 33008 1300
rect 32968 338 32996 1294
rect 32956 332 33008 338
rect 32956 274 33008 280
rect 33244 56 33364 82
rect 32232 14 32444 42
rect 32494 0 32550 56
rect 32862 0 32918 56
rect 33230 54 33364 56
rect 33230 0 33286 54
rect 33336 42 33364 54
rect 33520 42 33548 2246
rect 33612 56 33640 2790
rect 33796 134 33824 7278
rect 35440 6112 35492 6118
rect 35440 6054 35492 6060
rect 33968 3596 34020 3602
rect 33968 3538 34020 3544
rect 33980 2446 34008 3538
rect 34704 3460 34756 3466
rect 34704 3402 34756 3408
rect 34336 2576 34388 2582
rect 34336 2518 34388 2524
rect 33968 2440 34020 2446
rect 33968 2382 34020 2388
rect 34244 2304 34296 2310
rect 34244 2246 34296 2252
rect 33784 128 33836 134
rect 33784 70 33836 76
rect 33980 56 34100 82
rect 33336 14 33548 42
rect 33598 0 33654 56
rect 33966 54 34100 56
rect 33966 0 34022 54
rect 34072 42 34100 54
rect 34256 42 34284 2246
rect 34348 56 34376 2518
rect 34716 2446 34744 3402
rect 35072 3392 35124 3398
rect 35072 3334 35124 3340
rect 35084 2446 35112 3334
rect 35452 2446 35480 6054
rect 35532 2644 35584 2650
rect 35532 2586 35584 2592
rect 34704 2440 34756 2446
rect 34704 2382 34756 2388
rect 35072 2440 35124 2446
rect 35072 2382 35124 2388
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 35164 2372 35216 2378
rect 35164 2314 35216 2320
rect 34980 2304 35032 2310
rect 34980 2246 35032 2252
rect 34716 56 34836 82
rect 34072 14 34284 42
rect 34334 0 34390 56
rect 34702 54 34836 56
rect 34702 0 34758 54
rect 34808 42 34836 54
rect 34992 42 35020 2246
rect 35176 1170 35204 2314
rect 35544 1170 35572 2586
rect 35808 2576 35860 2582
rect 35808 2518 35860 2524
rect 35624 2440 35676 2446
rect 35624 2382 35676 2388
rect 35636 1562 35664 2382
rect 35624 1556 35676 1562
rect 35624 1498 35676 1504
rect 35084 1142 35204 1170
rect 35452 1142 35572 1170
rect 35084 56 35112 1142
rect 35452 56 35480 1142
rect 35820 56 35848 2518
rect 36188 2446 36216 7686
rect 36452 7540 36504 7546
rect 36452 7482 36504 7488
rect 36464 6934 36492 7482
rect 36556 7478 36584 7754
rect 36820 7744 36872 7750
rect 36820 7686 36872 7692
rect 36544 7472 36596 7478
rect 36544 7414 36596 7420
rect 36452 6928 36504 6934
rect 36452 6870 36504 6876
rect 36544 6724 36596 6730
rect 36544 6666 36596 6672
rect 36556 6390 36584 6666
rect 36544 6384 36596 6390
rect 36544 6326 36596 6332
rect 36268 2848 36320 2854
rect 36268 2790 36320 2796
rect 36176 2440 36228 2446
rect 36176 2382 36228 2388
rect 36280 1442 36308 2790
rect 36832 2446 36860 7686
rect 37200 6186 37228 8434
rect 37292 7546 37320 8978
rect 38212 8634 38240 11194
rect 38568 9240 38620 9246
rect 38568 9182 38620 9188
rect 38200 8628 38252 8634
rect 38200 8570 38252 8576
rect 37832 8424 37884 8430
rect 37832 8366 37884 8372
rect 37844 8090 37872 8366
rect 37950 8188 38258 8197
rect 37950 8186 37956 8188
rect 38012 8186 38036 8188
rect 38092 8186 38116 8188
rect 38172 8186 38196 8188
rect 38252 8186 38258 8188
rect 38012 8134 38014 8186
rect 38194 8134 38196 8186
rect 37950 8132 37956 8134
rect 38012 8132 38036 8134
rect 38092 8132 38116 8134
rect 38172 8132 38196 8134
rect 38252 8132 38258 8134
rect 37950 8123 38258 8132
rect 37832 8084 37884 8090
rect 37832 8026 37884 8032
rect 37280 7540 37332 7546
rect 37280 7482 37332 7488
rect 37372 7200 37424 7206
rect 37372 7142 37424 7148
rect 37188 6180 37240 6186
rect 37188 6122 37240 6128
rect 37384 4622 37412 7142
rect 37950 7100 38258 7109
rect 37950 7098 37956 7100
rect 38012 7098 38036 7100
rect 38092 7098 38116 7100
rect 38172 7098 38196 7100
rect 38252 7098 38258 7100
rect 38012 7046 38014 7098
rect 38194 7046 38196 7098
rect 37950 7044 37956 7046
rect 38012 7044 38036 7046
rect 38092 7044 38116 7046
rect 38172 7044 38196 7046
rect 38252 7044 38258 7046
rect 37950 7035 38258 7044
rect 38580 6730 38608 9182
rect 40408 9104 40460 9110
rect 40408 9046 40460 9052
rect 38752 8968 38804 8974
rect 38752 8910 38804 8916
rect 38764 7546 38792 8910
rect 39010 8732 39318 8741
rect 39010 8730 39016 8732
rect 39072 8730 39096 8732
rect 39152 8730 39176 8732
rect 39232 8730 39256 8732
rect 39312 8730 39318 8732
rect 39072 8678 39074 8730
rect 39254 8678 39256 8730
rect 39010 8676 39016 8678
rect 39072 8676 39096 8678
rect 39152 8676 39176 8678
rect 39232 8676 39256 8678
rect 39312 8676 39318 8678
rect 39010 8667 39318 8676
rect 39580 8492 39632 8498
rect 39580 8434 39632 8440
rect 39010 7644 39318 7653
rect 39010 7642 39016 7644
rect 39072 7642 39096 7644
rect 39152 7642 39176 7644
rect 39232 7642 39256 7644
rect 39312 7642 39318 7644
rect 39072 7590 39074 7642
rect 39254 7590 39256 7642
rect 39010 7588 39016 7590
rect 39072 7588 39096 7590
rect 39152 7588 39176 7590
rect 39232 7588 39256 7590
rect 39312 7588 39318 7590
rect 39010 7579 39318 7588
rect 39592 7546 39620 8434
rect 39948 8356 40000 8362
rect 39948 8298 40000 8304
rect 39672 7880 39724 7886
rect 39672 7822 39724 7828
rect 38752 7540 38804 7546
rect 38752 7482 38804 7488
rect 39580 7540 39632 7546
rect 39580 7482 39632 7488
rect 38936 7336 38988 7342
rect 38672 7284 38936 7290
rect 38672 7278 38988 7284
rect 39580 7336 39632 7342
rect 39580 7278 39632 7284
rect 38672 7262 38976 7278
rect 38672 7206 38700 7262
rect 38660 7200 38712 7206
rect 38660 7142 38712 7148
rect 38568 6724 38620 6730
rect 38568 6666 38620 6672
rect 39010 6556 39318 6565
rect 39010 6554 39016 6556
rect 39072 6554 39096 6556
rect 39152 6554 39176 6556
rect 39232 6554 39256 6556
rect 39312 6554 39318 6556
rect 39072 6502 39074 6554
rect 39254 6502 39256 6554
rect 39010 6500 39016 6502
rect 39072 6500 39096 6502
rect 39152 6500 39176 6502
rect 39232 6500 39256 6502
rect 39312 6500 39318 6502
rect 39010 6491 39318 6500
rect 37950 6012 38258 6021
rect 37950 6010 37956 6012
rect 38012 6010 38036 6012
rect 38092 6010 38116 6012
rect 38172 6010 38196 6012
rect 38252 6010 38258 6012
rect 38012 5958 38014 6010
rect 38194 5958 38196 6010
rect 37950 5956 37956 5958
rect 38012 5956 38036 5958
rect 38092 5956 38116 5958
rect 38172 5956 38196 5958
rect 38252 5956 38258 5958
rect 37950 5947 38258 5956
rect 39010 5468 39318 5477
rect 39010 5466 39016 5468
rect 39072 5466 39096 5468
rect 39152 5466 39176 5468
rect 39232 5466 39256 5468
rect 39312 5466 39318 5468
rect 39072 5414 39074 5466
rect 39254 5414 39256 5466
rect 39010 5412 39016 5414
rect 39072 5412 39096 5414
rect 39152 5412 39176 5414
rect 39232 5412 39256 5414
rect 39312 5412 39318 5414
rect 39010 5403 39318 5412
rect 37950 4924 38258 4933
rect 37950 4922 37956 4924
rect 38012 4922 38036 4924
rect 38092 4922 38116 4924
rect 38172 4922 38196 4924
rect 38252 4922 38258 4924
rect 38012 4870 38014 4922
rect 38194 4870 38196 4922
rect 37950 4868 37956 4870
rect 38012 4868 38036 4870
rect 38092 4868 38116 4870
rect 38172 4868 38196 4870
rect 38252 4868 38258 4870
rect 37950 4859 38258 4868
rect 37004 4616 37056 4622
rect 37004 4558 37056 4564
rect 37372 4616 37424 4622
rect 37372 4558 37424 4564
rect 36912 2576 36964 2582
rect 36912 2518 36964 2524
rect 36820 2440 36872 2446
rect 36820 2382 36872 2388
rect 36728 2304 36780 2310
rect 36728 2246 36780 2252
rect 36544 1964 36596 1970
rect 36544 1906 36596 1912
rect 36556 1630 36584 1906
rect 36544 1624 36596 1630
rect 36544 1566 36596 1572
rect 36188 1414 36308 1442
rect 36188 56 36216 1414
rect 36556 56 36676 82
rect 34808 14 35020 42
rect 35070 0 35126 56
rect 35438 0 35494 56
rect 35806 0 35862 56
rect 36174 0 36230 56
rect 36542 54 36676 56
rect 36542 0 36598 54
rect 36648 42 36676 54
rect 36740 42 36768 2246
rect 36924 56 36952 2518
rect 37016 2514 37044 4558
rect 37188 4480 37240 4486
rect 37188 4422 37240 4428
rect 37004 2508 37056 2514
rect 37004 2450 37056 2456
rect 37200 2038 37228 4422
rect 39010 4380 39318 4389
rect 39010 4378 39016 4380
rect 39072 4378 39096 4380
rect 39152 4378 39176 4380
rect 39232 4378 39256 4380
rect 39312 4378 39318 4380
rect 39072 4326 39074 4378
rect 39254 4326 39256 4378
rect 39010 4324 39016 4326
rect 39072 4324 39096 4326
rect 39152 4324 39176 4326
rect 39232 4324 39256 4326
rect 39312 4324 39318 4326
rect 39010 4315 39318 4324
rect 37950 3836 38258 3845
rect 37950 3834 37956 3836
rect 38012 3834 38036 3836
rect 38092 3834 38116 3836
rect 38172 3834 38196 3836
rect 38252 3834 38258 3836
rect 38012 3782 38014 3834
rect 38194 3782 38196 3834
rect 37950 3780 37956 3782
rect 38012 3780 38036 3782
rect 38092 3780 38116 3782
rect 38172 3780 38196 3782
rect 38252 3780 38258 3782
rect 37950 3771 38258 3780
rect 38844 3732 38896 3738
rect 38844 3674 38896 3680
rect 38856 3058 38884 3674
rect 39010 3292 39318 3301
rect 39010 3290 39016 3292
rect 39072 3290 39096 3292
rect 39152 3290 39176 3292
rect 39232 3290 39256 3292
rect 39312 3290 39318 3292
rect 39072 3238 39074 3290
rect 39254 3238 39256 3290
rect 39010 3236 39016 3238
rect 39072 3236 39096 3238
rect 39152 3236 39176 3238
rect 39232 3236 39256 3238
rect 39312 3236 39318 3238
rect 39010 3227 39318 3236
rect 38844 3052 38896 3058
rect 38844 2994 38896 3000
rect 38752 2848 38804 2854
rect 38752 2790 38804 2796
rect 37950 2748 38258 2757
rect 37950 2746 37956 2748
rect 38012 2746 38036 2748
rect 38092 2746 38116 2748
rect 38172 2746 38196 2748
rect 38252 2746 38258 2748
rect 38012 2694 38014 2746
rect 38194 2694 38196 2746
rect 37950 2692 37956 2694
rect 38012 2692 38036 2694
rect 38092 2692 38116 2694
rect 38172 2692 38196 2694
rect 38252 2692 38258 2694
rect 37950 2683 38258 2692
rect 37648 2644 37700 2650
rect 37648 2586 37700 2592
rect 37188 2032 37240 2038
rect 37188 1974 37240 1980
rect 37280 1420 37332 1426
rect 37280 1362 37332 1368
rect 37292 56 37320 1362
rect 37660 56 37688 2586
rect 38384 2576 38436 2582
rect 38384 2518 38436 2524
rect 38016 2440 38068 2446
rect 38016 2382 38068 2388
rect 38108 2440 38160 2446
rect 38108 2382 38160 2388
rect 38028 1494 38056 2382
rect 38120 2009 38148 2382
rect 38200 2304 38252 2310
rect 38200 2246 38252 2252
rect 38106 2000 38162 2009
rect 38106 1935 38162 1944
rect 38016 1488 38068 1494
rect 38016 1430 38068 1436
rect 38108 1488 38160 1494
rect 38108 1430 38160 1436
rect 38120 1170 38148 1430
rect 38212 1426 38240 2246
rect 38200 1420 38252 1426
rect 38200 1362 38252 1368
rect 38028 1142 38148 1170
rect 38028 56 38056 1142
rect 38396 56 38424 2518
rect 38476 2440 38528 2446
rect 38476 2382 38528 2388
rect 38488 1601 38516 2382
rect 38568 2304 38620 2310
rect 38568 2246 38620 2252
rect 38474 1592 38530 1601
rect 38474 1527 38530 1536
rect 38580 1494 38608 2246
rect 38568 1488 38620 1494
rect 38568 1430 38620 1436
rect 38764 56 38792 2790
rect 39488 2576 39540 2582
rect 39488 2518 39540 2524
rect 38844 2440 38896 2446
rect 39212 2440 39264 2446
rect 38844 2382 38896 2388
rect 39210 2408 39212 2417
rect 39264 2408 39266 2417
rect 38856 1737 38884 2382
rect 39210 2343 39266 2352
rect 39396 2304 39448 2310
rect 39396 2246 39448 2252
rect 39010 2204 39318 2213
rect 39010 2202 39016 2204
rect 39072 2202 39096 2204
rect 39152 2202 39176 2204
rect 39232 2202 39256 2204
rect 39312 2202 39318 2204
rect 39072 2150 39074 2202
rect 39254 2150 39256 2202
rect 39010 2148 39016 2150
rect 39072 2148 39096 2150
rect 39152 2148 39176 2150
rect 39232 2148 39256 2150
rect 39312 2148 39318 2150
rect 39010 2139 39318 2148
rect 38842 1728 38898 1737
rect 38842 1663 38898 1672
rect 39132 56 39252 82
rect 36648 14 36768 42
rect 36910 0 36966 56
rect 37278 0 37334 56
rect 37646 0 37702 56
rect 38014 0 38070 56
rect 38382 0 38438 56
rect 38750 0 38806 56
rect 39118 54 39252 56
rect 39118 0 39174 54
rect 39224 42 39252 54
rect 39408 42 39436 2246
rect 39500 56 39528 2518
rect 39592 1426 39620 7278
rect 39580 1420 39632 1426
rect 39580 1362 39632 1368
rect 39684 377 39712 7822
rect 39856 7812 39908 7818
rect 39856 7754 39908 7760
rect 39670 368 39726 377
rect 39670 303 39726 312
rect 39868 56 39896 7754
rect 39960 6662 39988 8298
rect 40132 7744 40184 7750
rect 40132 7686 40184 7692
rect 40316 7744 40368 7750
rect 40316 7686 40368 7692
rect 39948 6656 40000 6662
rect 39948 6598 40000 6604
rect 40040 6452 40092 6458
rect 40040 6394 40092 6400
rect 40052 4758 40080 6394
rect 40040 4752 40092 4758
rect 40040 4694 40092 4700
rect 40038 4176 40094 4185
rect 40038 4111 40040 4120
rect 40092 4111 40094 4120
rect 40040 4082 40092 4088
rect 40038 2544 40094 2553
rect 40038 2479 40094 2488
rect 40052 2446 40080 2479
rect 40040 2440 40092 2446
rect 40040 2382 40092 2388
rect 40144 105 40172 7686
rect 40224 7200 40276 7206
rect 40224 7142 40276 7148
rect 40130 96 40186 105
rect 39224 14 39436 42
rect 39486 0 39542 56
rect 39854 0 39910 56
rect 40236 56 40264 7142
rect 40328 2514 40356 7686
rect 40420 6458 40448 9046
rect 40512 8634 40540 11194
rect 41236 8832 41288 8838
rect 41236 8774 41288 8780
rect 40500 8628 40552 8634
rect 40500 8570 40552 8576
rect 40868 8492 40920 8498
rect 40868 8434 40920 8440
rect 40880 7546 40908 8434
rect 41248 8430 41276 8774
rect 42812 8634 42840 11194
rect 45112 11098 45140 11194
rect 45204 11098 45232 11206
rect 45112 11070 45232 11098
rect 45010 8732 45318 8741
rect 45010 8730 45016 8732
rect 45072 8730 45096 8732
rect 45152 8730 45176 8732
rect 45232 8730 45256 8732
rect 45312 8730 45318 8732
rect 45072 8678 45074 8730
rect 45254 8678 45256 8730
rect 45010 8676 45016 8678
rect 45072 8676 45096 8678
rect 45152 8676 45176 8678
rect 45232 8676 45256 8678
rect 45312 8676 45318 8678
rect 45010 8667 45318 8676
rect 45388 8634 45416 11206
rect 47398 11194 47454 11250
rect 45926 9888 45982 9897
rect 45926 9823 45982 9832
rect 45834 8800 45890 8809
rect 45834 8735 45890 8744
rect 45848 8634 45876 8735
rect 42800 8628 42852 8634
rect 42800 8570 42852 8576
rect 45376 8628 45428 8634
rect 45376 8570 45428 8576
rect 45836 8628 45888 8634
rect 45836 8570 45888 8576
rect 43168 8492 43220 8498
rect 43168 8434 43220 8440
rect 45468 8492 45520 8498
rect 45468 8434 45520 8440
rect 41236 8424 41288 8430
rect 41236 8366 41288 8372
rect 40868 7540 40920 7546
rect 40868 7482 40920 7488
rect 40592 7268 40644 7274
rect 40592 7210 40644 7216
rect 40408 6452 40460 6458
rect 40408 6394 40460 6400
rect 40316 2508 40368 2514
rect 40316 2450 40368 2456
rect 40500 2508 40552 2514
rect 40500 2450 40552 2456
rect 40512 2038 40540 2450
rect 40500 2032 40552 2038
rect 40500 1974 40552 1980
rect 40604 56 40632 7210
rect 42708 6724 42760 6730
rect 42708 6666 42760 6672
rect 40958 6216 41014 6225
rect 40958 6151 41014 6160
rect 40972 56 41000 6151
rect 42720 5098 42748 6666
rect 43180 6662 43208 8434
rect 43950 8188 44258 8197
rect 43950 8186 43956 8188
rect 44012 8186 44036 8188
rect 44092 8186 44116 8188
rect 44172 8186 44196 8188
rect 44252 8186 44258 8188
rect 44012 8134 44014 8186
rect 44194 8134 44196 8186
rect 43950 8132 43956 8134
rect 44012 8132 44036 8134
rect 44092 8132 44116 8134
rect 44172 8132 44196 8134
rect 44252 8132 44258 8134
rect 43950 8123 44258 8132
rect 43812 8084 43864 8090
rect 43812 8026 43864 8032
rect 43444 7540 43496 7546
rect 43444 7482 43496 7488
rect 42800 6656 42852 6662
rect 42800 6598 42852 6604
rect 43168 6656 43220 6662
rect 43168 6598 43220 6604
rect 42812 5914 42840 6598
rect 42800 5908 42852 5914
rect 42800 5850 42852 5856
rect 42708 5092 42760 5098
rect 42708 5034 42760 5040
rect 42800 4820 42852 4826
rect 42800 4762 42852 4768
rect 41604 4684 41656 4690
rect 41604 4626 41656 4632
rect 41616 3058 41644 4626
rect 42432 4276 42484 4282
rect 42432 4218 42484 4224
rect 42444 4146 42472 4218
rect 42432 4140 42484 4146
rect 42432 4082 42484 4088
rect 42616 3936 42668 3942
rect 42616 3878 42668 3884
rect 42628 3602 42656 3878
rect 42616 3596 42668 3602
rect 42616 3538 42668 3544
rect 41604 3052 41656 3058
rect 41604 2994 41656 3000
rect 42812 2514 42840 4762
rect 43456 3126 43484 7482
rect 43720 6996 43772 7002
rect 43720 6938 43772 6944
rect 43732 5234 43760 6938
rect 43824 6866 43852 8026
rect 44824 7744 44876 7750
rect 44824 7686 44876 7692
rect 45376 7744 45428 7750
rect 45376 7686 45428 7692
rect 43950 7100 44258 7109
rect 43950 7098 43956 7100
rect 44012 7098 44036 7100
rect 44092 7098 44116 7100
rect 44172 7098 44196 7100
rect 44252 7098 44258 7100
rect 44012 7046 44014 7098
rect 44194 7046 44196 7098
rect 43950 7044 43956 7046
rect 44012 7044 44036 7046
rect 44092 7044 44116 7046
rect 44172 7044 44196 7046
rect 44252 7044 44258 7046
rect 43950 7035 44258 7044
rect 44364 6928 44416 6934
rect 44364 6870 44416 6876
rect 43812 6860 43864 6866
rect 43812 6802 43864 6808
rect 43950 6012 44258 6021
rect 43950 6010 43956 6012
rect 44012 6010 44036 6012
rect 44092 6010 44116 6012
rect 44172 6010 44196 6012
rect 44252 6010 44258 6012
rect 44012 5958 44014 6010
rect 44194 5958 44196 6010
rect 43950 5956 43956 5958
rect 44012 5956 44036 5958
rect 44092 5956 44116 5958
rect 44172 5956 44196 5958
rect 44252 5956 44258 5958
rect 43950 5947 44258 5956
rect 43812 5908 43864 5914
rect 43812 5850 43864 5856
rect 43720 5228 43772 5234
rect 43720 5170 43772 5176
rect 43444 3120 43496 3126
rect 43444 3062 43496 3068
rect 43166 2952 43222 2961
rect 43166 2887 43222 2896
rect 42800 2508 42852 2514
rect 42800 2450 42852 2456
rect 41328 1420 41380 1426
rect 41328 1362 41380 1368
rect 41340 56 41368 1362
rect 41696 332 41748 338
rect 41696 274 41748 280
rect 41708 56 41736 274
rect 42432 264 42484 270
rect 42432 206 42484 212
rect 41972 128 42024 134
rect 42024 76 42104 82
rect 41972 70 42104 76
rect 41984 56 42104 70
rect 42444 56 42472 206
rect 42800 196 42852 202
rect 42800 138 42852 144
rect 42812 56 42840 138
rect 43180 56 43208 2887
rect 43536 1964 43588 1970
rect 43536 1906 43588 1912
rect 43548 56 43576 1906
rect 43824 1408 43852 5850
rect 43950 4924 44258 4933
rect 43950 4922 43956 4924
rect 44012 4922 44036 4924
rect 44092 4922 44116 4924
rect 44172 4922 44196 4924
rect 44252 4922 44258 4924
rect 44012 4870 44014 4922
rect 44194 4870 44196 4922
rect 43950 4868 43956 4870
rect 44012 4868 44036 4870
rect 44092 4868 44116 4870
rect 44172 4868 44196 4870
rect 44252 4868 44258 4870
rect 43950 4859 44258 4868
rect 44376 4078 44404 6870
rect 44640 6792 44692 6798
rect 44640 6734 44692 6740
rect 44364 4072 44416 4078
rect 44364 4014 44416 4020
rect 43950 3836 44258 3845
rect 43950 3834 43956 3836
rect 44012 3834 44036 3836
rect 44092 3834 44116 3836
rect 44172 3834 44196 3836
rect 44252 3834 44258 3836
rect 44012 3782 44014 3834
rect 44194 3782 44196 3834
rect 43950 3780 43956 3782
rect 44012 3780 44036 3782
rect 44092 3780 44116 3782
rect 44172 3780 44196 3782
rect 44252 3780 44258 3782
rect 43950 3771 44258 3780
rect 43950 2748 44258 2757
rect 43950 2746 43956 2748
rect 44012 2746 44036 2748
rect 44092 2746 44116 2748
rect 44172 2746 44196 2748
rect 44252 2746 44258 2748
rect 44012 2694 44014 2746
rect 44194 2694 44196 2746
rect 43950 2692 43956 2694
rect 44012 2692 44036 2694
rect 44092 2692 44116 2694
rect 44172 2692 44196 2694
rect 44252 2692 44258 2694
rect 43950 2683 44258 2692
rect 43824 1380 43944 1408
rect 43916 56 43944 1380
rect 44270 504 44326 513
rect 44270 439 44326 448
rect 44284 56 44312 439
rect 44652 56 44680 6734
rect 44836 66 44864 7686
rect 45010 7644 45318 7653
rect 45010 7642 45016 7644
rect 45072 7642 45096 7644
rect 45152 7642 45176 7644
rect 45232 7642 45256 7644
rect 45312 7642 45318 7644
rect 45072 7590 45074 7642
rect 45254 7590 45256 7642
rect 45010 7588 45016 7590
rect 45072 7588 45096 7590
rect 45152 7588 45176 7590
rect 45232 7588 45256 7590
rect 45312 7588 45318 7590
rect 45010 7579 45318 7588
rect 45388 7546 45416 7686
rect 45376 7540 45428 7546
rect 45376 7482 45428 7488
rect 45480 6662 45508 8434
rect 45940 7750 45968 9823
rect 46294 9616 46350 9625
rect 46294 9551 46350 9560
rect 46020 9172 46072 9178
rect 46020 9114 46072 9120
rect 46032 8498 46060 9114
rect 46204 8628 46256 8634
rect 46204 8570 46256 8576
rect 46216 8537 46244 8570
rect 46202 8528 46258 8537
rect 46020 8492 46072 8498
rect 46202 8463 46258 8472
rect 46020 8434 46072 8440
rect 46020 7880 46072 7886
rect 46020 7822 46072 7828
rect 46112 7880 46164 7886
rect 46112 7822 46164 7828
rect 45928 7744 45980 7750
rect 45928 7686 45980 7692
rect 45928 7404 45980 7410
rect 45928 7346 45980 7352
rect 45744 7336 45796 7342
rect 45744 7278 45796 7284
rect 45468 6656 45520 6662
rect 45468 6598 45520 6604
rect 45010 6556 45318 6565
rect 45010 6554 45016 6556
rect 45072 6554 45096 6556
rect 45152 6554 45176 6556
rect 45232 6554 45256 6556
rect 45312 6554 45318 6556
rect 45072 6502 45074 6554
rect 45254 6502 45256 6554
rect 45010 6500 45016 6502
rect 45072 6500 45096 6502
rect 45152 6500 45176 6502
rect 45232 6500 45256 6502
rect 45312 6500 45318 6502
rect 45010 6491 45318 6500
rect 45376 6316 45428 6322
rect 45376 6258 45428 6264
rect 44916 6248 44968 6254
rect 44916 6190 44968 6196
rect 44928 1408 44956 6190
rect 45010 5468 45318 5477
rect 45010 5466 45016 5468
rect 45072 5466 45096 5468
rect 45152 5466 45176 5468
rect 45232 5466 45256 5468
rect 45312 5466 45318 5468
rect 45072 5414 45074 5466
rect 45254 5414 45256 5466
rect 45010 5412 45016 5414
rect 45072 5412 45096 5414
rect 45152 5412 45176 5414
rect 45232 5412 45256 5414
rect 45312 5412 45318 5414
rect 45010 5403 45318 5412
rect 45010 4380 45318 4389
rect 45010 4378 45016 4380
rect 45072 4378 45096 4380
rect 45152 4378 45176 4380
rect 45232 4378 45256 4380
rect 45312 4378 45318 4380
rect 45072 4326 45074 4378
rect 45254 4326 45256 4378
rect 45010 4324 45016 4326
rect 45072 4324 45096 4326
rect 45152 4324 45176 4326
rect 45232 4324 45256 4326
rect 45312 4324 45318 4326
rect 45010 4315 45318 4324
rect 45010 3292 45318 3301
rect 45010 3290 45016 3292
rect 45072 3290 45096 3292
rect 45152 3290 45176 3292
rect 45232 3290 45256 3292
rect 45312 3290 45318 3292
rect 45072 3238 45074 3290
rect 45254 3238 45256 3290
rect 45010 3236 45016 3238
rect 45072 3236 45096 3238
rect 45152 3236 45176 3238
rect 45232 3236 45256 3238
rect 45312 3236 45318 3238
rect 45010 3227 45318 3236
rect 45010 2204 45318 2213
rect 45010 2202 45016 2204
rect 45072 2202 45096 2204
rect 45152 2202 45176 2204
rect 45232 2202 45256 2204
rect 45312 2202 45318 2204
rect 45072 2150 45074 2202
rect 45254 2150 45256 2202
rect 45010 2148 45016 2150
rect 45072 2148 45096 2150
rect 45152 2148 45176 2150
rect 45232 2148 45256 2150
rect 45312 2148 45318 2150
rect 45010 2139 45318 2148
rect 44928 1380 45048 1408
rect 44824 60 44876 66
rect 40130 31 40186 40
rect 40222 0 40278 56
rect 40590 0 40646 56
rect 40958 0 41014 56
rect 41326 0 41382 56
rect 41694 0 41750 56
rect 41984 54 42118 56
rect 42062 0 42118 54
rect 42430 0 42486 56
rect 42798 0 42854 56
rect 43166 0 43222 56
rect 43534 0 43590 56
rect 43902 0 43958 56
rect 44270 0 44326 56
rect 44638 0 44694 56
rect 45020 56 45048 1380
rect 45388 56 45416 6258
rect 45560 5704 45612 5710
rect 45560 5646 45612 5652
rect 45572 3194 45600 5646
rect 45652 5296 45704 5302
rect 45652 5238 45704 5244
rect 45560 3188 45612 3194
rect 45560 3130 45612 3136
rect 45664 2922 45692 5238
rect 45652 2916 45704 2922
rect 45652 2858 45704 2864
rect 45756 56 45784 7278
rect 45940 2774 45968 7346
rect 46032 7002 46060 7822
rect 46020 6996 46072 7002
rect 46020 6938 46072 6944
rect 46020 6792 46072 6798
rect 46018 6760 46020 6769
rect 46072 6760 46074 6769
rect 46018 6695 46074 6704
rect 46124 5778 46152 7822
rect 46308 7750 46336 9551
rect 46938 9344 46994 9353
rect 46938 9279 46994 9288
rect 46662 9072 46718 9081
rect 46662 9007 46718 9016
rect 46388 8900 46440 8906
rect 46388 8842 46440 8848
rect 46400 8498 46428 8842
rect 46388 8492 46440 8498
rect 46388 8434 46440 8440
rect 46676 8090 46704 9007
rect 46756 8492 46808 8498
rect 46756 8434 46808 8440
rect 46664 8084 46716 8090
rect 46664 8026 46716 8032
rect 46572 7812 46624 7818
rect 46572 7754 46624 7760
rect 46296 7744 46348 7750
rect 46296 7686 46348 7692
rect 46584 7410 46612 7754
rect 46768 7546 46796 8434
rect 46952 7546 46980 9279
rect 47412 8634 47440 11194
rect 47400 8628 47452 8634
rect 47400 8570 47452 8576
rect 47216 8356 47268 8362
rect 47216 8298 47268 8304
rect 47308 8356 47360 8362
rect 47308 8298 47360 8304
rect 47228 8265 47256 8298
rect 47214 8256 47270 8265
rect 47214 8191 47270 8200
rect 47320 7993 47348 8298
rect 47306 7984 47362 7993
rect 47306 7919 47362 7928
rect 47216 7880 47268 7886
rect 47216 7822 47268 7828
rect 47032 7744 47084 7750
rect 47032 7686 47084 7692
rect 46756 7540 46808 7546
rect 46756 7482 46808 7488
rect 46940 7540 46992 7546
rect 46940 7482 46992 7488
rect 47044 7449 47072 7686
rect 47030 7440 47086 7449
rect 46572 7404 46624 7410
rect 47030 7375 47086 7384
rect 46572 7346 46624 7352
rect 46296 6860 46348 6866
rect 46296 6802 46348 6808
rect 46112 5772 46164 5778
rect 46112 5714 46164 5720
rect 46204 5568 46256 5574
rect 46204 5510 46256 5516
rect 46020 4208 46072 4214
rect 46020 4150 46072 4156
rect 46032 3738 46060 4150
rect 46020 3732 46072 3738
rect 46020 3674 46072 3680
rect 45940 2746 46152 2774
rect 45836 2304 45888 2310
rect 45836 2246 45888 2252
rect 45848 2009 45876 2246
rect 45834 2000 45890 2009
rect 45834 1935 45890 1944
rect 46124 56 46152 2746
rect 46216 2514 46244 5510
rect 46308 4026 46336 6802
rect 46664 6792 46716 6798
rect 46664 6734 46716 6740
rect 47124 6792 47176 6798
rect 47124 6734 47176 6740
rect 46572 6316 46624 6322
rect 46572 6258 46624 6264
rect 46584 5370 46612 6258
rect 46572 5364 46624 5370
rect 46572 5306 46624 5312
rect 46478 4584 46534 4593
rect 46478 4519 46534 4528
rect 46308 3998 46428 4026
rect 46296 3936 46348 3942
rect 46296 3878 46348 3884
rect 46308 3641 46336 3878
rect 46294 3632 46350 3641
rect 46294 3567 46350 3576
rect 46400 2774 46428 3998
rect 46492 3534 46520 4519
rect 46480 3528 46532 3534
rect 46480 3470 46532 3476
rect 46676 3482 46704 6734
rect 47032 6656 47084 6662
rect 47030 6624 47032 6633
rect 47084 6624 47086 6633
rect 47030 6559 47086 6568
rect 46756 6112 46808 6118
rect 46754 6080 46756 6089
rect 46940 6112 46992 6118
rect 46808 6080 46810 6089
rect 46940 6054 46992 6060
rect 46754 6015 46810 6024
rect 46952 5846 46980 6054
rect 46940 5840 46992 5846
rect 46940 5782 46992 5788
rect 47136 5642 47164 6734
rect 47228 6390 47256 7822
rect 47400 7744 47452 7750
rect 47398 7712 47400 7721
rect 47452 7712 47454 7721
rect 47398 7647 47454 7656
rect 47492 7336 47544 7342
rect 47492 7278 47544 7284
rect 47308 7200 47360 7206
rect 47306 7168 47308 7177
rect 47360 7168 47362 7177
rect 47306 7103 47362 7112
rect 47398 6896 47454 6905
rect 47398 6831 47454 6840
rect 47412 6662 47440 6831
rect 47400 6656 47452 6662
rect 47400 6598 47452 6604
rect 47308 6452 47360 6458
rect 47308 6394 47360 6400
rect 47216 6384 47268 6390
rect 47320 6361 47348 6394
rect 47216 6326 47268 6332
rect 47306 6352 47362 6361
rect 47306 6287 47362 6296
rect 47400 5840 47452 5846
rect 47398 5808 47400 5817
rect 47452 5808 47454 5817
rect 47398 5743 47454 5752
rect 47216 5704 47268 5710
rect 47216 5646 47268 5652
rect 47124 5636 47176 5642
rect 47124 5578 47176 5584
rect 47032 5568 47084 5574
rect 47030 5536 47032 5545
rect 47084 5536 47086 5545
rect 47030 5471 47086 5480
rect 47228 5302 47256 5646
rect 47308 5364 47360 5370
rect 47308 5306 47360 5312
rect 47216 5296 47268 5302
rect 47320 5273 47348 5306
rect 47216 5238 47268 5244
rect 47306 5264 47362 5273
rect 47306 5199 47362 5208
rect 47504 5114 47532 7278
rect 47228 5086 47532 5114
rect 46940 5024 46992 5030
rect 46938 4992 46940 5001
rect 46992 4992 46994 5001
rect 46938 4927 46994 4936
rect 47032 4480 47084 4486
rect 47030 4448 47032 4457
rect 47084 4448 47086 4457
rect 47030 4383 47086 4392
rect 46848 3936 46900 3942
rect 46940 3936 46992 3942
rect 46848 3878 46900 3884
rect 46938 3904 46940 3913
rect 46992 3904 46994 3913
rect 46676 3454 46796 3482
rect 46664 3392 46716 3398
rect 46664 3334 46716 3340
rect 46676 3058 46704 3334
rect 46664 3052 46716 3058
rect 46664 2994 46716 3000
rect 46768 2774 46796 3454
rect 46860 3058 46888 3878
rect 46938 3839 46994 3848
rect 47032 3664 47084 3670
rect 47032 3606 47084 3612
rect 46848 3052 46900 3058
rect 46848 2994 46900 3000
rect 46940 2848 46992 2854
rect 46938 2816 46940 2825
rect 46992 2816 46994 2825
rect 46400 2746 46520 2774
rect 46768 2746 46888 2774
rect 46938 2751 46994 2760
rect 46204 2508 46256 2514
rect 46204 2450 46256 2456
rect 46388 2440 46440 2446
rect 46388 2382 46440 2388
rect 46204 2304 46256 2310
rect 46204 2246 46256 2252
rect 46216 1737 46244 2246
rect 46400 1902 46428 2382
rect 46388 1896 46440 1902
rect 46388 1838 46440 1844
rect 46202 1728 46258 1737
rect 46202 1663 46258 1672
rect 46492 56 46520 2746
rect 46572 2304 46624 2310
rect 46572 2246 46624 2252
rect 46584 1465 46612 2246
rect 46570 1456 46626 1465
rect 46570 1391 46626 1400
rect 46860 56 46888 2746
rect 47044 2446 47072 3606
rect 47124 3392 47176 3398
rect 47122 3360 47124 3369
rect 47176 3360 47178 3369
rect 47122 3295 47178 3304
rect 47032 2440 47084 2446
rect 47032 2382 47084 2388
rect 46940 2304 46992 2310
rect 46938 2272 46940 2281
rect 46992 2272 46994 2281
rect 46938 2207 46994 2216
rect 47228 56 47256 5086
rect 47400 4752 47452 4758
rect 47398 4720 47400 4729
rect 47452 4720 47454 4729
rect 47398 4655 47454 4664
rect 47306 4176 47362 4185
rect 47306 4111 47362 4120
rect 47320 4010 47348 4111
rect 47308 4004 47360 4010
rect 47308 3946 47360 3952
rect 47306 3632 47362 3641
rect 47306 3567 47362 3576
rect 47320 3194 47348 3567
rect 47308 3188 47360 3194
rect 47308 3130 47360 3136
rect 47306 3088 47362 3097
rect 47306 3023 47362 3032
rect 47320 2650 47348 3023
rect 47952 2916 48004 2922
rect 47952 2858 48004 2864
rect 47308 2644 47360 2650
rect 47308 2586 47360 2592
rect 47964 2553 47992 2858
rect 47950 2544 48006 2553
rect 47950 2479 48006 2488
rect 44824 2 44876 8
rect 45006 0 45062 56
rect 45374 0 45430 56
rect 45742 0 45798 56
rect 46110 0 46166 56
rect 46478 0 46534 56
rect 46846 0 46902 56
rect 47214 0 47270 56
<< via2 >>
rect 202 9832 258 9888
rect 1030 9288 1086 9344
rect 2870 8744 2926 8800
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 7562 9016 7618 9072
rect 2870 8336 2926 8392
rect 1766 8200 1822 8256
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 12254 9560 12310 9616
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 1766 7792 1822 7848
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 1306 7384 1362 7440
rect 202 6432 258 6488
rect 478 4392 534 4448
rect 1306 3848 1362 3904
rect 1214 1944 1270 2000
rect 1306 1672 1362 1728
rect 1122 1400 1178 1456
rect 1766 4936 1822 4992
rect 1766 4528 1822 4584
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 2410 6432 2466 6488
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 2410 5888 2466 5944
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 2410 4020 2412 4040
rect 2412 4020 2464 4040
rect 2464 4020 2466 4040
rect 2410 3984 2466 4020
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 7746 6704 7802 6760
rect 5814 6432 5870 6488
rect 8758 6568 8814 6624
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 7746 5888 7802 5944
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 8850 6432 8906 6488
rect 8758 6024 8814 6080
rect 12162 7248 12218 7304
rect 11886 6296 11942 6352
rect 11518 6160 11574 6216
rect 8666 5752 8722 5808
rect 8850 5752 8906 5808
rect 7654 5616 7710 5672
rect 5814 2352 5870 2408
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 7654 2488 7710 2544
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 19338 8472 19394 8528
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 12346 7384 12402 7440
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 12714 6432 12770 6488
rect 12714 6160 12770 6216
rect 13726 6024 13782 6080
rect 11978 5616 12034 5672
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 11518 1808 11574 1864
rect 11150 448 11206 504
rect 9310 176 9366 232
rect 12530 2488 12586 2544
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 13818 5072 13874 5128
rect 12898 2352 12954 2408
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 14554 3712 14610 3768
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 14922 1672 14978 1728
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 21730 8336 21786 8392
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 25594 7928 25650 7984
rect 26330 7928 26386 7984
rect 23754 7828 23756 7848
rect 23756 7828 23808 7848
rect 23808 7828 23810 7848
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 19246 6840 19302 6896
rect 18418 6296 18474 6352
rect 17958 5208 18014 5264
rect 17130 1536 17186 1592
rect 17774 4936 17830 4992
rect 19614 6296 19670 6352
rect 17958 2896 18014 2952
rect 18602 1944 18658 2000
rect 18510 312 18566 368
rect 17774 40 17830 96
rect 19338 3712 19394 3768
rect 23754 7792 23810 7828
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 21730 5344 21786 5400
rect 22926 4528 22982 4584
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 24030 5344 24086 5400
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 24950 2896 25006 2952
rect 25870 4664 25926 4720
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 25870 3032 25926 3088
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 26974 5072 27030 5128
rect 26790 3440 26846 3496
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 27526 448 27582 504
rect 27986 1808 28042 1864
rect 29734 3032 29790 3088
rect 30378 6316 30434 6352
rect 30378 6296 30380 6316
rect 30380 6296 30432 6316
rect 30432 6296 30434 6316
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 30010 3984 30066 4040
rect 29918 448 29974 504
rect 31114 3052 31170 3088
rect 31114 3032 31116 3052
rect 31116 3032 31168 3052
rect 31168 3032 31170 3052
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 32770 5752 32826 5808
rect 32494 5616 32550 5672
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 31298 176 31354 232
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
rect 37956 8186 38012 8188
rect 38036 8186 38092 8188
rect 38116 8186 38172 8188
rect 38196 8186 38252 8188
rect 37956 8134 38002 8186
rect 38002 8134 38012 8186
rect 38036 8134 38066 8186
rect 38066 8134 38078 8186
rect 38078 8134 38092 8186
rect 38116 8134 38130 8186
rect 38130 8134 38142 8186
rect 38142 8134 38172 8186
rect 38196 8134 38206 8186
rect 38206 8134 38252 8186
rect 37956 8132 38012 8134
rect 38036 8132 38092 8134
rect 38116 8132 38172 8134
rect 38196 8132 38252 8134
rect 37956 7098 38012 7100
rect 38036 7098 38092 7100
rect 38116 7098 38172 7100
rect 38196 7098 38252 7100
rect 37956 7046 38002 7098
rect 38002 7046 38012 7098
rect 38036 7046 38066 7098
rect 38066 7046 38078 7098
rect 38078 7046 38092 7098
rect 38116 7046 38130 7098
rect 38130 7046 38142 7098
rect 38142 7046 38172 7098
rect 38196 7046 38206 7098
rect 38206 7046 38252 7098
rect 37956 7044 38012 7046
rect 38036 7044 38092 7046
rect 38116 7044 38172 7046
rect 38196 7044 38252 7046
rect 39016 8730 39072 8732
rect 39096 8730 39152 8732
rect 39176 8730 39232 8732
rect 39256 8730 39312 8732
rect 39016 8678 39062 8730
rect 39062 8678 39072 8730
rect 39096 8678 39126 8730
rect 39126 8678 39138 8730
rect 39138 8678 39152 8730
rect 39176 8678 39190 8730
rect 39190 8678 39202 8730
rect 39202 8678 39232 8730
rect 39256 8678 39266 8730
rect 39266 8678 39312 8730
rect 39016 8676 39072 8678
rect 39096 8676 39152 8678
rect 39176 8676 39232 8678
rect 39256 8676 39312 8678
rect 39016 7642 39072 7644
rect 39096 7642 39152 7644
rect 39176 7642 39232 7644
rect 39256 7642 39312 7644
rect 39016 7590 39062 7642
rect 39062 7590 39072 7642
rect 39096 7590 39126 7642
rect 39126 7590 39138 7642
rect 39138 7590 39152 7642
rect 39176 7590 39190 7642
rect 39190 7590 39202 7642
rect 39202 7590 39232 7642
rect 39256 7590 39266 7642
rect 39266 7590 39312 7642
rect 39016 7588 39072 7590
rect 39096 7588 39152 7590
rect 39176 7588 39232 7590
rect 39256 7588 39312 7590
rect 39016 6554 39072 6556
rect 39096 6554 39152 6556
rect 39176 6554 39232 6556
rect 39256 6554 39312 6556
rect 39016 6502 39062 6554
rect 39062 6502 39072 6554
rect 39096 6502 39126 6554
rect 39126 6502 39138 6554
rect 39138 6502 39152 6554
rect 39176 6502 39190 6554
rect 39190 6502 39202 6554
rect 39202 6502 39232 6554
rect 39256 6502 39266 6554
rect 39266 6502 39312 6554
rect 39016 6500 39072 6502
rect 39096 6500 39152 6502
rect 39176 6500 39232 6502
rect 39256 6500 39312 6502
rect 37956 6010 38012 6012
rect 38036 6010 38092 6012
rect 38116 6010 38172 6012
rect 38196 6010 38252 6012
rect 37956 5958 38002 6010
rect 38002 5958 38012 6010
rect 38036 5958 38066 6010
rect 38066 5958 38078 6010
rect 38078 5958 38092 6010
rect 38116 5958 38130 6010
rect 38130 5958 38142 6010
rect 38142 5958 38172 6010
rect 38196 5958 38206 6010
rect 38206 5958 38252 6010
rect 37956 5956 38012 5958
rect 38036 5956 38092 5958
rect 38116 5956 38172 5958
rect 38196 5956 38252 5958
rect 39016 5466 39072 5468
rect 39096 5466 39152 5468
rect 39176 5466 39232 5468
rect 39256 5466 39312 5468
rect 39016 5414 39062 5466
rect 39062 5414 39072 5466
rect 39096 5414 39126 5466
rect 39126 5414 39138 5466
rect 39138 5414 39152 5466
rect 39176 5414 39190 5466
rect 39190 5414 39202 5466
rect 39202 5414 39232 5466
rect 39256 5414 39266 5466
rect 39266 5414 39312 5466
rect 39016 5412 39072 5414
rect 39096 5412 39152 5414
rect 39176 5412 39232 5414
rect 39256 5412 39312 5414
rect 37956 4922 38012 4924
rect 38036 4922 38092 4924
rect 38116 4922 38172 4924
rect 38196 4922 38252 4924
rect 37956 4870 38002 4922
rect 38002 4870 38012 4922
rect 38036 4870 38066 4922
rect 38066 4870 38078 4922
rect 38078 4870 38092 4922
rect 38116 4870 38130 4922
rect 38130 4870 38142 4922
rect 38142 4870 38172 4922
rect 38196 4870 38206 4922
rect 38206 4870 38252 4922
rect 37956 4868 38012 4870
rect 38036 4868 38092 4870
rect 38116 4868 38172 4870
rect 38196 4868 38252 4870
rect 39016 4378 39072 4380
rect 39096 4378 39152 4380
rect 39176 4378 39232 4380
rect 39256 4378 39312 4380
rect 39016 4326 39062 4378
rect 39062 4326 39072 4378
rect 39096 4326 39126 4378
rect 39126 4326 39138 4378
rect 39138 4326 39152 4378
rect 39176 4326 39190 4378
rect 39190 4326 39202 4378
rect 39202 4326 39232 4378
rect 39256 4326 39266 4378
rect 39266 4326 39312 4378
rect 39016 4324 39072 4326
rect 39096 4324 39152 4326
rect 39176 4324 39232 4326
rect 39256 4324 39312 4326
rect 37956 3834 38012 3836
rect 38036 3834 38092 3836
rect 38116 3834 38172 3836
rect 38196 3834 38252 3836
rect 37956 3782 38002 3834
rect 38002 3782 38012 3834
rect 38036 3782 38066 3834
rect 38066 3782 38078 3834
rect 38078 3782 38092 3834
rect 38116 3782 38130 3834
rect 38130 3782 38142 3834
rect 38142 3782 38172 3834
rect 38196 3782 38206 3834
rect 38206 3782 38252 3834
rect 37956 3780 38012 3782
rect 38036 3780 38092 3782
rect 38116 3780 38172 3782
rect 38196 3780 38252 3782
rect 39016 3290 39072 3292
rect 39096 3290 39152 3292
rect 39176 3290 39232 3292
rect 39256 3290 39312 3292
rect 39016 3238 39062 3290
rect 39062 3238 39072 3290
rect 39096 3238 39126 3290
rect 39126 3238 39138 3290
rect 39138 3238 39152 3290
rect 39176 3238 39190 3290
rect 39190 3238 39202 3290
rect 39202 3238 39232 3290
rect 39256 3238 39266 3290
rect 39266 3238 39312 3290
rect 39016 3236 39072 3238
rect 39096 3236 39152 3238
rect 39176 3236 39232 3238
rect 39256 3236 39312 3238
rect 37956 2746 38012 2748
rect 38036 2746 38092 2748
rect 38116 2746 38172 2748
rect 38196 2746 38252 2748
rect 37956 2694 38002 2746
rect 38002 2694 38012 2746
rect 38036 2694 38066 2746
rect 38066 2694 38078 2746
rect 38078 2694 38092 2746
rect 38116 2694 38130 2746
rect 38130 2694 38142 2746
rect 38142 2694 38172 2746
rect 38196 2694 38206 2746
rect 38206 2694 38252 2746
rect 37956 2692 38012 2694
rect 38036 2692 38092 2694
rect 38116 2692 38172 2694
rect 38196 2692 38252 2694
rect 38106 1944 38162 2000
rect 38474 1536 38530 1592
rect 39210 2388 39212 2408
rect 39212 2388 39264 2408
rect 39264 2388 39266 2408
rect 39210 2352 39266 2388
rect 39016 2202 39072 2204
rect 39096 2202 39152 2204
rect 39176 2202 39232 2204
rect 39256 2202 39312 2204
rect 39016 2150 39062 2202
rect 39062 2150 39072 2202
rect 39096 2150 39126 2202
rect 39126 2150 39138 2202
rect 39138 2150 39152 2202
rect 39176 2150 39190 2202
rect 39190 2150 39202 2202
rect 39202 2150 39232 2202
rect 39256 2150 39266 2202
rect 39266 2150 39312 2202
rect 39016 2148 39072 2150
rect 39096 2148 39152 2150
rect 39176 2148 39232 2150
rect 39256 2148 39312 2150
rect 38842 1672 38898 1728
rect 39670 312 39726 368
rect 40038 4140 40094 4176
rect 40038 4120 40040 4140
rect 40040 4120 40092 4140
rect 40092 4120 40094 4140
rect 40038 2488 40094 2544
rect 40130 40 40186 96
rect 45016 8730 45072 8732
rect 45096 8730 45152 8732
rect 45176 8730 45232 8732
rect 45256 8730 45312 8732
rect 45016 8678 45062 8730
rect 45062 8678 45072 8730
rect 45096 8678 45126 8730
rect 45126 8678 45138 8730
rect 45138 8678 45152 8730
rect 45176 8678 45190 8730
rect 45190 8678 45202 8730
rect 45202 8678 45232 8730
rect 45256 8678 45266 8730
rect 45266 8678 45312 8730
rect 45016 8676 45072 8678
rect 45096 8676 45152 8678
rect 45176 8676 45232 8678
rect 45256 8676 45312 8678
rect 45926 9832 45982 9888
rect 45834 8744 45890 8800
rect 40958 6160 41014 6216
rect 43956 8186 44012 8188
rect 44036 8186 44092 8188
rect 44116 8186 44172 8188
rect 44196 8186 44252 8188
rect 43956 8134 44002 8186
rect 44002 8134 44012 8186
rect 44036 8134 44066 8186
rect 44066 8134 44078 8186
rect 44078 8134 44092 8186
rect 44116 8134 44130 8186
rect 44130 8134 44142 8186
rect 44142 8134 44172 8186
rect 44196 8134 44206 8186
rect 44206 8134 44252 8186
rect 43956 8132 44012 8134
rect 44036 8132 44092 8134
rect 44116 8132 44172 8134
rect 44196 8132 44252 8134
rect 43956 7098 44012 7100
rect 44036 7098 44092 7100
rect 44116 7098 44172 7100
rect 44196 7098 44252 7100
rect 43956 7046 44002 7098
rect 44002 7046 44012 7098
rect 44036 7046 44066 7098
rect 44066 7046 44078 7098
rect 44078 7046 44092 7098
rect 44116 7046 44130 7098
rect 44130 7046 44142 7098
rect 44142 7046 44172 7098
rect 44196 7046 44206 7098
rect 44206 7046 44252 7098
rect 43956 7044 44012 7046
rect 44036 7044 44092 7046
rect 44116 7044 44172 7046
rect 44196 7044 44252 7046
rect 43956 6010 44012 6012
rect 44036 6010 44092 6012
rect 44116 6010 44172 6012
rect 44196 6010 44252 6012
rect 43956 5958 44002 6010
rect 44002 5958 44012 6010
rect 44036 5958 44066 6010
rect 44066 5958 44078 6010
rect 44078 5958 44092 6010
rect 44116 5958 44130 6010
rect 44130 5958 44142 6010
rect 44142 5958 44172 6010
rect 44196 5958 44206 6010
rect 44206 5958 44252 6010
rect 43956 5956 44012 5958
rect 44036 5956 44092 5958
rect 44116 5956 44172 5958
rect 44196 5956 44252 5958
rect 43166 2896 43222 2952
rect 43956 4922 44012 4924
rect 44036 4922 44092 4924
rect 44116 4922 44172 4924
rect 44196 4922 44252 4924
rect 43956 4870 44002 4922
rect 44002 4870 44012 4922
rect 44036 4870 44066 4922
rect 44066 4870 44078 4922
rect 44078 4870 44092 4922
rect 44116 4870 44130 4922
rect 44130 4870 44142 4922
rect 44142 4870 44172 4922
rect 44196 4870 44206 4922
rect 44206 4870 44252 4922
rect 43956 4868 44012 4870
rect 44036 4868 44092 4870
rect 44116 4868 44172 4870
rect 44196 4868 44252 4870
rect 43956 3834 44012 3836
rect 44036 3834 44092 3836
rect 44116 3834 44172 3836
rect 44196 3834 44252 3836
rect 43956 3782 44002 3834
rect 44002 3782 44012 3834
rect 44036 3782 44066 3834
rect 44066 3782 44078 3834
rect 44078 3782 44092 3834
rect 44116 3782 44130 3834
rect 44130 3782 44142 3834
rect 44142 3782 44172 3834
rect 44196 3782 44206 3834
rect 44206 3782 44252 3834
rect 43956 3780 44012 3782
rect 44036 3780 44092 3782
rect 44116 3780 44172 3782
rect 44196 3780 44252 3782
rect 43956 2746 44012 2748
rect 44036 2746 44092 2748
rect 44116 2746 44172 2748
rect 44196 2746 44252 2748
rect 43956 2694 44002 2746
rect 44002 2694 44012 2746
rect 44036 2694 44066 2746
rect 44066 2694 44078 2746
rect 44078 2694 44092 2746
rect 44116 2694 44130 2746
rect 44130 2694 44142 2746
rect 44142 2694 44172 2746
rect 44196 2694 44206 2746
rect 44206 2694 44252 2746
rect 43956 2692 44012 2694
rect 44036 2692 44092 2694
rect 44116 2692 44172 2694
rect 44196 2692 44252 2694
rect 44270 448 44326 504
rect 45016 7642 45072 7644
rect 45096 7642 45152 7644
rect 45176 7642 45232 7644
rect 45256 7642 45312 7644
rect 45016 7590 45062 7642
rect 45062 7590 45072 7642
rect 45096 7590 45126 7642
rect 45126 7590 45138 7642
rect 45138 7590 45152 7642
rect 45176 7590 45190 7642
rect 45190 7590 45202 7642
rect 45202 7590 45232 7642
rect 45256 7590 45266 7642
rect 45266 7590 45312 7642
rect 45016 7588 45072 7590
rect 45096 7588 45152 7590
rect 45176 7588 45232 7590
rect 45256 7588 45312 7590
rect 46294 9560 46350 9616
rect 46202 8472 46258 8528
rect 45016 6554 45072 6556
rect 45096 6554 45152 6556
rect 45176 6554 45232 6556
rect 45256 6554 45312 6556
rect 45016 6502 45062 6554
rect 45062 6502 45072 6554
rect 45096 6502 45126 6554
rect 45126 6502 45138 6554
rect 45138 6502 45152 6554
rect 45176 6502 45190 6554
rect 45190 6502 45202 6554
rect 45202 6502 45232 6554
rect 45256 6502 45266 6554
rect 45266 6502 45312 6554
rect 45016 6500 45072 6502
rect 45096 6500 45152 6502
rect 45176 6500 45232 6502
rect 45256 6500 45312 6502
rect 45016 5466 45072 5468
rect 45096 5466 45152 5468
rect 45176 5466 45232 5468
rect 45256 5466 45312 5468
rect 45016 5414 45062 5466
rect 45062 5414 45072 5466
rect 45096 5414 45126 5466
rect 45126 5414 45138 5466
rect 45138 5414 45152 5466
rect 45176 5414 45190 5466
rect 45190 5414 45202 5466
rect 45202 5414 45232 5466
rect 45256 5414 45266 5466
rect 45266 5414 45312 5466
rect 45016 5412 45072 5414
rect 45096 5412 45152 5414
rect 45176 5412 45232 5414
rect 45256 5412 45312 5414
rect 45016 4378 45072 4380
rect 45096 4378 45152 4380
rect 45176 4378 45232 4380
rect 45256 4378 45312 4380
rect 45016 4326 45062 4378
rect 45062 4326 45072 4378
rect 45096 4326 45126 4378
rect 45126 4326 45138 4378
rect 45138 4326 45152 4378
rect 45176 4326 45190 4378
rect 45190 4326 45202 4378
rect 45202 4326 45232 4378
rect 45256 4326 45266 4378
rect 45266 4326 45312 4378
rect 45016 4324 45072 4326
rect 45096 4324 45152 4326
rect 45176 4324 45232 4326
rect 45256 4324 45312 4326
rect 45016 3290 45072 3292
rect 45096 3290 45152 3292
rect 45176 3290 45232 3292
rect 45256 3290 45312 3292
rect 45016 3238 45062 3290
rect 45062 3238 45072 3290
rect 45096 3238 45126 3290
rect 45126 3238 45138 3290
rect 45138 3238 45152 3290
rect 45176 3238 45190 3290
rect 45190 3238 45202 3290
rect 45202 3238 45232 3290
rect 45256 3238 45266 3290
rect 45266 3238 45312 3290
rect 45016 3236 45072 3238
rect 45096 3236 45152 3238
rect 45176 3236 45232 3238
rect 45256 3236 45312 3238
rect 45016 2202 45072 2204
rect 45096 2202 45152 2204
rect 45176 2202 45232 2204
rect 45256 2202 45312 2204
rect 45016 2150 45062 2202
rect 45062 2150 45072 2202
rect 45096 2150 45126 2202
rect 45126 2150 45138 2202
rect 45138 2150 45152 2202
rect 45176 2150 45190 2202
rect 45190 2150 45202 2202
rect 45202 2150 45232 2202
rect 45256 2150 45266 2202
rect 45266 2150 45312 2202
rect 45016 2148 45072 2150
rect 45096 2148 45152 2150
rect 45176 2148 45232 2150
rect 45256 2148 45312 2150
rect 46018 6740 46020 6760
rect 46020 6740 46072 6760
rect 46072 6740 46074 6760
rect 46018 6704 46074 6740
rect 46938 9288 46994 9344
rect 46662 9016 46718 9072
rect 47214 8200 47270 8256
rect 47306 7928 47362 7984
rect 47030 7384 47086 7440
rect 45834 1944 45890 2000
rect 46478 4528 46534 4584
rect 46294 3576 46350 3632
rect 47030 6604 47032 6624
rect 47032 6604 47084 6624
rect 47084 6604 47086 6624
rect 47030 6568 47086 6604
rect 46754 6060 46756 6080
rect 46756 6060 46808 6080
rect 46808 6060 46810 6080
rect 46754 6024 46810 6060
rect 47398 7692 47400 7712
rect 47400 7692 47452 7712
rect 47452 7692 47454 7712
rect 47398 7656 47454 7692
rect 47306 7148 47308 7168
rect 47308 7148 47360 7168
rect 47360 7148 47362 7168
rect 47306 7112 47362 7148
rect 47398 6840 47454 6896
rect 47306 6296 47362 6352
rect 47398 5788 47400 5808
rect 47400 5788 47452 5808
rect 47452 5788 47454 5808
rect 47398 5752 47454 5788
rect 47030 5516 47032 5536
rect 47032 5516 47084 5536
rect 47084 5516 47086 5536
rect 47030 5480 47086 5516
rect 47306 5208 47362 5264
rect 46938 4972 46940 4992
rect 46940 4972 46992 4992
rect 46992 4972 46994 4992
rect 46938 4936 46994 4972
rect 47030 4428 47032 4448
rect 47032 4428 47084 4448
rect 47084 4428 47086 4448
rect 47030 4392 47086 4428
rect 46938 3884 46940 3904
rect 46940 3884 46992 3904
rect 46992 3884 46994 3904
rect 46938 3848 46994 3884
rect 46938 2796 46940 2816
rect 46940 2796 46992 2816
rect 46992 2796 46994 2816
rect 46938 2760 46994 2796
rect 46202 1672 46258 1728
rect 46570 1400 46626 1456
rect 47122 3340 47124 3360
rect 47124 3340 47176 3360
rect 47176 3340 47178 3360
rect 47122 3304 47178 3340
rect 46938 2252 46940 2272
rect 46940 2252 46992 2272
rect 46992 2252 46994 2272
rect 46938 2216 46994 2252
rect 47398 4700 47400 4720
rect 47400 4700 47452 4720
rect 47452 4700 47454 4720
rect 47398 4664 47454 4700
rect 47306 4120 47362 4176
rect 47306 3576 47362 3632
rect 47306 3032 47362 3088
rect 47950 2488 48006 2544
<< metal3 >>
rect 0 9890 120 9920
rect 197 9890 263 9893
rect 0 9888 263 9890
rect 0 9832 202 9888
rect 258 9832 263 9888
rect 0 9830 263 9832
rect 0 9800 120 9830
rect 197 9827 263 9830
rect 45921 9890 45987 9893
rect 48880 9890 49000 9920
rect 45921 9888 49000 9890
rect 45921 9832 45926 9888
rect 45982 9832 49000 9888
rect 45921 9830 49000 9832
rect 45921 9827 45987 9830
rect 48880 9800 49000 9830
rect 0 9618 120 9648
rect 12249 9618 12315 9621
rect 0 9616 12315 9618
rect 0 9560 12254 9616
rect 12310 9560 12315 9616
rect 0 9558 12315 9560
rect 0 9528 120 9558
rect 12249 9555 12315 9558
rect 46289 9618 46355 9621
rect 48880 9618 49000 9648
rect 46289 9616 49000 9618
rect 46289 9560 46294 9616
rect 46350 9560 49000 9616
rect 46289 9558 49000 9560
rect 46289 9555 46355 9558
rect 48880 9528 49000 9558
rect 0 9346 120 9376
rect 1025 9346 1091 9349
rect 0 9344 1091 9346
rect 0 9288 1030 9344
rect 1086 9288 1091 9344
rect 0 9286 1091 9288
rect 0 9256 120 9286
rect 1025 9283 1091 9286
rect 46933 9346 46999 9349
rect 48880 9346 49000 9376
rect 46933 9344 49000 9346
rect 46933 9288 46938 9344
rect 46994 9288 49000 9344
rect 46933 9286 49000 9288
rect 46933 9283 46999 9286
rect 48880 9256 49000 9286
rect 0 9074 120 9104
rect 7557 9074 7623 9077
rect 0 9072 7623 9074
rect 0 9016 7562 9072
rect 7618 9016 7623 9072
rect 0 9014 7623 9016
rect 0 8984 120 9014
rect 7557 9011 7623 9014
rect 46657 9074 46723 9077
rect 48880 9074 49000 9104
rect 46657 9072 49000 9074
rect 46657 9016 46662 9072
rect 46718 9016 49000 9072
rect 46657 9014 49000 9016
rect 46657 9011 46723 9014
rect 48880 8984 49000 9014
rect 0 8802 120 8832
rect 2865 8802 2931 8805
rect 0 8800 2931 8802
rect 0 8744 2870 8800
rect 2926 8744 2931 8800
rect 0 8742 2931 8744
rect 0 8712 120 8742
rect 2865 8739 2931 8742
rect 45829 8802 45895 8805
rect 48880 8802 49000 8832
rect 45829 8800 49000 8802
rect 45829 8744 45834 8800
rect 45890 8744 49000 8800
rect 45829 8742 49000 8744
rect 45829 8739 45895 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 33006 8671 33322 8672
rect 39006 8736 39322 8737
rect 39006 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39322 8736
rect 39006 8671 39322 8672
rect 45006 8736 45322 8737
rect 45006 8672 45012 8736
rect 45076 8672 45092 8736
rect 45156 8672 45172 8736
rect 45236 8672 45252 8736
rect 45316 8672 45322 8736
rect 48880 8712 49000 8742
rect 45006 8671 45322 8672
rect 0 8530 120 8560
rect 19333 8530 19399 8533
rect 0 8528 19399 8530
rect 0 8472 19338 8528
rect 19394 8472 19399 8528
rect 0 8470 19399 8472
rect 0 8440 120 8470
rect 19333 8467 19399 8470
rect 46197 8530 46263 8533
rect 48880 8530 49000 8560
rect 46197 8528 49000 8530
rect 46197 8472 46202 8528
rect 46258 8472 49000 8528
rect 46197 8470 49000 8472
rect 46197 8467 46263 8470
rect 48880 8440 49000 8470
rect 2865 8394 2931 8397
rect 21725 8394 21791 8397
rect 2865 8392 21791 8394
rect 2865 8336 2870 8392
rect 2926 8336 21730 8392
rect 21786 8336 21791 8392
rect 2865 8334 21791 8336
rect 2865 8331 2931 8334
rect 21725 8331 21791 8334
rect 0 8258 120 8288
rect 1761 8258 1827 8261
rect 0 8256 1827 8258
rect 0 8200 1766 8256
rect 1822 8200 1827 8256
rect 0 8198 1827 8200
rect 0 8168 120 8198
rect 1761 8195 1827 8198
rect 47209 8258 47275 8261
rect 48880 8258 49000 8288
rect 47209 8256 49000 8258
rect 47209 8200 47214 8256
rect 47270 8200 49000 8256
rect 47209 8198 49000 8200
rect 47209 8195 47275 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 37946 8192 38262 8193
rect 37946 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38262 8192
rect 37946 8127 38262 8128
rect 43946 8192 44262 8193
rect 43946 8128 43952 8192
rect 44016 8128 44032 8192
rect 44096 8128 44112 8192
rect 44176 8128 44192 8192
rect 44256 8128 44262 8192
rect 48880 8168 49000 8198
rect 43946 8127 44262 8128
rect 0 7986 120 8016
rect 25589 7986 25655 7989
rect 26325 7986 26391 7989
rect 0 7984 26391 7986
rect 0 7928 25594 7984
rect 25650 7928 26330 7984
rect 26386 7928 26391 7984
rect 0 7926 26391 7928
rect 0 7896 120 7926
rect 25589 7923 25655 7926
rect 26325 7923 26391 7926
rect 47301 7986 47367 7989
rect 48880 7986 49000 8016
rect 47301 7984 49000 7986
rect 47301 7928 47306 7984
rect 47362 7928 49000 7984
rect 47301 7926 49000 7928
rect 47301 7923 47367 7926
rect 48880 7896 49000 7926
rect 1761 7850 1827 7853
rect 23749 7850 23815 7853
rect 1761 7848 23815 7850
rect 1761 7792 1766 7848
rect 1822 7792 23754 7848
rect 23810 7792 23815 7848
rect 1761 7790 23815 7792
rect 1761 7787 1827 7790
rect 23749 7787 23815 7790
rect 0 7714 120 7744
rect 47393 7714 47459 7717
rect 48880 7714 49000 7744
rect 0 7654 2882 7714
rect 0 7624 120 7654
rect 0 7442 120 7472
rect 1301 7442 1367 7445
rect 0 7440 1367 7442
rect 0 7384 1306 7440
rect 1362 7384 1367 7440
rect 0 7382 1367 7384
rect 2822 7442 2882 7654
rect 47393 7712 49000 7714
rect 47393 7656 47398 7712
rect 47454 7656 49000 7712
rect 47393 7654 49000 7656
rect 47393 7651 47459 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 33006 7583 33322 7584
rect 39006 7648 39322 7649
rect 39006 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39322 7648
rect 39006 7583 39322 7584
rect 45006 7648 45322 7649
rect 45006 7584 45012 7648
rect 45076 7584 45092 7648
rect 45156 7584 45172 7648
rect 45236 7584 45252 7648
rect 45316 7584 45322 7648
rect 48880 7624 49000 7654
rect 45006 7583 45322 7584
rect 12341 7442 12407 7445
rect 2822 7440 12407 7442
rect 2822 7384 12346 7440
rect 12402 7384 12407 7440
rect 2822 7382 12407 7384
rect 0 7352 120 7382
rect 1301 7379 1367 7382
rect 12341 7379 12407 7382
rect 47025 7442 47091 7445
rect 48880 7442 49000 7472
rect 47025 7440 49000 7442
rect 47025 7384 47030 7440
rect 47086 7384 49000 7440
rect 47025 7382 49000 7384
rect 47025 7379 47091 7382
rect 48880 7352 49000 7382
rect 12157 7306 12223 7309
rect 1718 7304 12223 7306
rect 1718 7248 12162 7304
rect 12218 7248 12223 7304
rect 1718 7246 12223 7248
rect 0 7170 120 7200
rect 1718 7170 1778 7246
rect 12157 7243 12223 7246
rect 0 7110 1778 7170
rect 47301 7170 47367 7173
rect 48880 7170 49000 7200
rect 47301 7168 49000 7170
rect 47301 7112 47306 7168
rect 47362 7112 49000 7168
rect 47301 7110 49000 7112
rect 0 7080 120 7110
rect 47301 7107 47367 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 37946 7104 38262 7105
rect 37946 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38262 7104
rect 37946 7039 38262 7040
rect 43946 7104 44262 7105
rect 43946 7040 43952 7104
rect 44016 7040 44032 7104
rect 44096 7040 44112 7104
rect 44176 7040 44192 7104
rect 44256 7040 44262 7104
rect 48880 7080 49000 7110
rect 43946 7039 44262 7040
rect 0 6898 120 6928
rect 19241 6898 19307 6901
rect 0 6896 19307 6898
rect 0 6840 19246 6896
rect 19302 6840 19307 6896
rect 0 6838 19307 6840
rect 0 6808 120 6838
rect 19241 6835 19307 6838
rect 47393 6898 47459 6901
rect 48880 6898 49000 6928
rect 47393 6896 49000 6898
rect 47393 6840 47398 6896
rect 47454 6840 49000 6896
rect 47393 6838 49000 6840
rect 47393 6835 47459 6838
rect 48880 6808 49000 6838
rect 7741 6762 7807 6765
rect 46013 6762 46079 6765
rect 2822 6702 6930 6762
rect 0 6626 120 6656
rect 2822 6626 2882 6702
rect 0 6566 2882 6626
rect 6870 6626 6930 6702
rect 7741 6760 46079 6762
rect 7741 6704 7746 6760
rect 7802 6704 46018 6760
rect 46074 6704 46079 6760
rect 7741 6702 46079 6704
rect 7741 6699 7807 6702
rect 46013 6699 46079 6702
rect 8753 6626 8819 6629
rect 6870 6624 8819 6626
rect 6870 6568 8758 6624
rect 8814 6568 8819 6624
rect 6870 6566 8819 6568
rect 0 6536 120 6566
rect 8753 6563 8819 6566
rect 47025 6626 47091 6629
rect 48880 6626 49000 6656
rect 47025 6624 49000 6626
rect 47025 6568 47030 6624
rect 47086 6568 49000 6624
rect 47025 6566 49000 6568
rect 47025 6563 47091 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 33006 6495 33322 6496
rect 39006 6560 39322 6561
rect 39006 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39322 6560
rect 39006 6495 39322 6496
rect 45006 6560 45322 6561
rect 45006 6496 45012 6560
rect 45076 6496 45092 6560
rect 45156 6496 45172 6560
rect 45236 6496 45252 6560
rect 45316 6496 45322 6560
rect 48880 6536 49000 6566
rect 45006 6495 45322 6496
rect 197 6490 263 6493
rect 2405 6490 2471 6493
rect 197 6488 2471 6490
rect 197 6432 202 6488
rect 258 6432 2410 6488
rect 2466 6432 2471 6488
rect 197 6430 2471 6432
rect 197 6427 263 6430
rect 2405 6427 2471 6430
rect 5809 6490 5875 6493
rect 8845 6490 8911 6493
rect 5809 6488 8911 6490
rect 5809 6432 5814 6488
rect 5870 6432 8850 6488
rect 8906 6432 8911 6488
rect 5809 6430 8911 6432
rect 5809 6427 5875 6430
rect 8845 6427 8911 6430
rect 12709 6490 12775 6493
rect 12709 6488 14842 6490
rect 12709 6432 12714 6488
rect 12770 6432 14842 6488
rect 12709 6430 14842 6432
rect 12709 6427 12775 6430
rect 0 6354 120 6384
rect 11881 6354 11947 6357
rect 14782 6354 14842 6430
rect 18413 6354 18479 6357
rect 0 6294 11714 6354
rect 0 6264 120 6294
rect 11513 6218 11579 6221
rect 1718 6216 11579 6218
rect 1718 6160 11518 6216
rect 11574 6160 11579 6216
rect 1718 6158 11579 6160
rect 11654 6218 11714 6294
rect 11881 6352 12956 6354
rect 11881 6296 11886 6352
rect 11942 6296 12956 6352
rect 11881 6294 12956 6296
rect 14782 6352 18479 6354
rect 14782 6296 18418 6352
rect 18474 6296 18479 6352
rect 14782 6294 18479 6296
rect 11881 6291 11947 6294
rect 12709 6218 12775 6221
rect 11654 6216 12775 6218
rect 11654 6160 12714 6216
rect 12770 6160 12775 6216
rect 11654 6158 12775 6160
rect 12896 6218 12956 6294
rect 18413 6291 18479 6294
rect 19609 6354 19675 6357
rect 30373 6354 30439 6357
rect 19609 6352 30439 6354
rect 19609 6296 19614 6352
rect 19670 6296 30378 6352
rect 30434 6296 30439 6352
rect 19609 6294 30439 6296
rect 19609 6291 19675 6294
rect 30373 6291 30439 6294
rect 47301 6354 47367 6357
rect 48880 6354 49000 6384
rect 47301 6352 49000 6354
rect 47301 6296 47306 6352
rect 47362 6296 49000 6352
rect 47301 6294 49000 6296
rect 47301 6291 47367 6294
rect 48880 6264 49000 6294
rect 40953 6218 41019 6221
rect 12896 6216 41019 6218
rect 12896 6160 40958 6216
rect 41014 6160 41019 6216
rect 12896 6158 41019 6160
rect 0 6082 120 6112
rect 1718 6082 1778 6158
rect 11513 6155 11579 6158
rect 12709 6155 12775 6158
rect 40953 6155 41019 6158
rect 0 6022 1778 6082
rect 8753 6082 8819 6085
rect 13721 6082 13787 6085
rect 8753 6080 13787 6082
rect 8753 6024 8758 6080
rect 8814 6024 13726 6080
rect 13782 6024 13787 6080
rect 8753 6022 13787 6024
rect 0 5992 120 6022
rect 8753 6019 8819 6022
rect 13721 6019 13787 6022
rect 46749 6082 46815 6085
rect 48880 6082 49000 6112
rect 46749 6080 49000 6082
rect 46749 6024 46754 6080
rect 46810 6024 49000 6080
rect 46749 6022 49000 6024
rect 46749 6019 46815 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 37946 6016 38262 6017
rect 37946 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38262 6016
rect 37946 5951 38262 5952
rect 43946 6016 44262 6017
rect 43946 5952 43952 6016
rect 44016 5952 44032 6016
rect 44096 5952 44112 6016
rect 44176 5952 44192 6016
rect 44256 5952 44262 6016
rect 48880 5992 49000 6022
rect 43946 5951 44262 5952
rect 2405 5946 2471 5949
rect 7741 5946 7807 5949
rect 2405 5944 7807 5946
rect 2405 5888 2410 5944
rect 2466 5888 7746 5944
rect 7802 5888 7807 5944
rect 2405 5886 7807 5888
rect 2405 5883 2471 5886
rect 7741 5883 7807 5886
rect 0 5810 120 5840
rect 8661 5810 8727 5813
rect 0 5750 3802 5810
rect 0 5720 120 5750
rect 3742 5674 3802 5750
rect 6870 5808 8727 5810
rect 6870 5752 8666 5808
rect 8722 5752 8727 5808
rect 6870 5750 8727 5752
rect 6870 5674 6930 5750
rect 8661 5747 8727 5750
rect 8845 5810 8911 5813
rect 32765 5810 32831 5813
rect 8845 5808 32831 5810
rect 8845 5752 8850 5808
rect 8906 5752 32770 5808
rect 32826 5752 32831 5808
rect 8845 5750 32831 5752
rect 8845 5747 8911 5750
rect 32765 5747 32831 5750
rect 47393 5810 47459 5813
rect 48880 5810 49000 5840
rect 47393 5808 49000 5810
rect 47393 5752 47398 5808
rect 47454 5752 49000 5808
rect 47393 5750 49000 5752
rect 47393 5747 47459 5750
rect 48880 5720 49000 5750
rect 2822 5614 3618 5674
rect 3742 5614 6930 5674
rect 7649 5674 7715 5677
rect 11973 5674 12039 5677
rect 32489 5674 32555 5677
rect 7649 5672 9506 5674
rect 7649 5616 7654 5672
rect 7710 5616 9506 5672
rect 7649 5614 9506 5616
rect 0 5538 120 5568
rect 2822 5538 2882 5614
rect 0 5478 2882 5538
rect 3558 5538 3618 5614
rect 7649 5611 7715 5614
rect 9446 5538 9506 5614
rect 11973 5672 32555 5674
rect 11973 5616 11978 5672
rect 12034 5616 32494 5672
rect 32550 5616 32555 5672
rect 11973 5614 32555 5616
rect 11973 5611 12039 5614
rect 32489 5611 32555 5614
rect 47025 5538 47091 5541
rect 48880 5538 49000 5568
rect 3558 5478 8770 5538
rect 9446 5478 14842 5538
rect 0 5448 120 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 0 5266 120 5296
rect 8710 5266 8770 5478
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 0 5206 6930 5266
rect 8710 5206 14658 5266
rect 0 5176 120 5206
rect 6870 5130 6930 5206
rect 13813 5130 13879 5133
rect 6870 5128 13879 5130
rect 6870 5072 13818 5128
rect 13874 5072 13879 5128
rect 6870 5070 13879 5072
rect 13813 5067 13879 5070
rect 0 4994 120 5024
rect 1761 4994 1827 4997
rect 0 4992 1827 4994
rect 0 4936 1766 4992
rect 1822 4936 1827 4992
rect 0 4934 1827 4936
rect 14598 4994 14658 5206
rect 14782 5130 14842 5478
rect 47025 5536 49000 5538
rect 47025 5480 47030 5536
rect 47086 5480 49000 5536
rect 47025 5478 49000 5480
rect 47025 5475 47091 5478
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 33006 5407 33322 5408
rect 39006 5472 39322 5473
rect 39006 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39322 5472
rect 39006 5407 39322 5408
rect 45006 5472 45322 5473
rect 45006 5408 45012 5472
rect 45076 5408 45092 5472
rect 45156 5408 45172 5472
rect 45236 5408 45252 5472
rect 45316 5408 45322 5472
rect 48880 5448 49000 5478
rect 45006 5407 45322 5408
rect 21725 5402 21791 5405
rect 24025 5402 24091 5405
rect 21725 5400 24091 5402
rect 21725 5344 21730 5400
rect 21786 5344 24030 5400
rect 24086 5344 24091 5400
rect 21725 5342 24091 5344
rect 21725 5339 21791 5342
rect 24025 5339 24091 5342
rect 17953 5266 18019 5269
rect 47301 5266 47367 5269
rect 48880 5266 49000 5296
rect 17953 5264 31770 5266
rect 17953 5208 17958 5264
rect 18014 5208 31770 5264
rect 17953 5206 31770 5208
rect 17953 5203 18019 5206
rect 26969 5130 27035 5133
rect 14782 5128 27035 5130
rect 14782 5072 26974 5128
rect 27030 5072 27035 5128
rect 14782 5070 27035 5072
rect 26969 5067 27035 5070
rect 17769 4994 17835 4997
rect 14598 4992 17835 4994
rect 14598 4936 17774 4992
rect 17830 4936 17835 4992
rect 14598 4934 17835 4936
rect 0 4904 120 4934
rect 1761 4931 1827 4934
rect 17769 4931 17835 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 0 4722 120 4752
rect 25865 4722 25931 4725
rect 0 4720 25931 4722
rect 0 4664 25870 4720
rect 25926 4664 25931 4720
rect 0 4662 25931 4664
rect 0 4632 120 4662
rect 25865 4659 25931 4662
rect 1761 4586 1827 4589
rect 22921 4586 22987 4589
rect 1761 4584 22987 4586
rect 1761 4528 1766 4584
rect 1822 4528 22926 4584
rect 22982 4528 22987 4584
rect 1761 4526 22987 4528
rect 31710 4586 31770 5206
rect 47301 5264 49000 5266
rect 47301 5208 47306 5264
rect 47362 5208 49000 5264
rect 47301 5206 49000 5208
rect 47301 5203 47367 5206
rect 48880 5176 49000 5206
rect 46933 4994 46999 4997
rect 48880 4994 49000 5024
rect 46933 4992 49000 4994
rect 46933 4936 46938 4992
rect 46994 4936 49000 4992
rect 46933 4934 49000 4936
rect 46933 4931 46999 4934
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 37946 4928 38262 4929
rect 37946 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38262 4928
rect 37946 4863 38262 4864
rect 43946 4928 44262 4929
rect 43946 4864 43952 4928
rect 44016 4864 44032 4928
rect 44096 4864 44112 4928
rect 44176 4864 44192 4928
rect 44256 4864 44262 4928
rect 48880 4904 49000 4934
rect 43946 4863 44262 4864
rect 47393 4722 47459 4725
rect 48880 4722 49000 4752
rect 47393 4720 49000 4722
rect 47393 4664 47398 4720
rect 47454 4664 49000 4720
rect 47393 4662 49000 4664
rect 47393 4659 47459 4662
rect 48880 4632 49000 4662
rect 46473 4586 46539 4589
rect 31710 4584 46539 4586
rect 31710 4528 46478 4584
rect 46534 4528 46539 4584
rect 31710 4526 46539 4528
rect 1761 4523 1827 4526
rect 22921 4523 22987 4526
rect 46473 4523 46539 4526
rect 0 4450 120 4480
rect 473 4450 539 4453
rect 0 4448 539 4450
rect 0 4392 478 4448
rect 534 4392 539 4448
rect 0 4390 539 4392
rect 0 4360 120 4390
rect 473 4387 539 4390
rect 47025 4450 47091 4453
rect 48880 4450 49000 4480
rect 47025 4448 49000 4450
rect 47025 4392 47030 4448
rect 47086 4392 49000 4448
rect 47025 4390 49000 4392
rect 47025 4387 47091 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 33006 4319 33322 4320
rect 39006 4384 39322 4385
rect 39006 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39322 4384
rect 39006 4319 39322 4320
rect 45006 4384 45322 4385
rect 45006 4320 45012 4384
rect 45076 4320 45092 4384
rect 45156 4320 45172 4384
rect 45236 4320 45252 4384
rect 45316 4320 45322 4384
rect 48880 4360 49000 4390
rect 45006 4319 45322 4320
rect 0 4178 120 4208
rect 40033 4178 40099 4181
rect 0 4176 40099 4178
rect 0 4120 40038 4176
rect 40094 4120 40099 4176
rect 0 4118 40099 4120
rect 0 4088 120 4118
rect 40033 4115 40099 4118
rect 47301 4178 47367 4181
rect 48880 4178 49000 4208
rect 47301 4176 49000 4178
rect 47301 4120 47306 4176
rect 47362 4120 49000 4176
rect 47301 4118 49000 4120
rect 47301 4115 47367 4118
rect 48880 4088 49000 4118
rect 2405 4042 2471 4045
rect 30005 4042 30071 4045
rect 2405 4040 30071 4042
rect 2405 3984 2410 4040
rect 2466 3984 30010 4040
rect 30066 3984 30071 4040
rect 2405 3982 30071 3984
rect 2405 3979 2471 3982
rect 30005 3979 30071 3982
rect 0 3906 120 3936
rect 1301 3906 1367 3909
rect 0 3904 1367 3906
rect 0 3848 1306 3904
rect 1362 3848 1367 3904
rect 0 3846 1367 3848
rect 0 3816 120 3846
rect 1301 3843 1367 3846
rect 46933 3906 46999 3909
rect 48880 3906 49000 3936
rect 46933 3904 49000 3906
rect 46933 3848 46938 3904
rect 46994 3848 49000 3904
rect 46933 3846 49000 3848
rect 46933 3843 46999 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 37946 3840 38262 3841
rect 37946 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38262 3840
rect 37946 3775 38262 3776
rect 43946 3840 44262 3841
rect 43946 3776 43952 3840
rect 44016 3776 44032 3840
rect 44096 3776 44112 3840
rect 44176 3776 44192 3840
rect 44256 3776 44262 3840
rect 48880 3816 49000 3846
rect 43946 3775 44262 3776
rect 14549 3770 14615 3773
rect 19333 3770 19399 3773
rect 14549 3768 19399 3770
rect 14549 3712 14554 3768
rect 14610 3712 19338 3768
rect 19394 3712 19399 3768
rect 14549 3710 19399 3712
rect 14549 3707 14615 3710
rect 19333 3707 19399 3710
rect 0 3634 120 3664
rect 46289 3634 46355 3637
rect 0 3632 46355 3634
rect 0 3576 46294 3632
rect 46350 3576 46355 3632
rect 0 3574 46355 3576
rect 0 3544 120 3574
rect 46289 3571 46355 3574
rect 47301 3634 47367 3637
rect 48880 3634 49000 3664
rect 47301 3632 49000 3634
rect 47301 3576 47306 3632
rect 47362 3576 49000 3632
rect 47301 3574 49000 3576
rect 47301 3571 47367 3574
rect 48880 3544 49000 3574
rect 26785 3498 26851 3501
rect 2822 3496 26851 3498
rect 2822 3440 26790 3496
rect 26846 3440 26851 3496
rect 2822 3438 26851 3440
rect 0 3362 120 3392
rect 2822 3362 2882 3438
rect 26785 3435 26851 3438
rect 0 3302 2882 3362
rect 47117 3362 47183 3365
rect 48880 3362 49000 3392
rect 47117 3360 49000 3362
rect 47117 3304 47122 3360
rect 47178 3304 49000 3360
rect 47117 3302 49000 3304
rect 0 3272 120 3302
rect 47117 3299 47183 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 33006 3231 33322 3232
rect 39006 3296 39322 3297
rect 39006 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39322 3296
rect 39006 3231 39322 3232
rect 45006 3296 45322 3297
rect 45006 3232 45012 3296
rect 45076 3232 45092 3296
rect 45156 3232 45172 3296
rect 45236 3232 45252 3296
rect 45316 3232 45322 3296
rect 48880 3272 49000 3302
rect 45006 3231 45322 3232
rect 0 3090 120 3120
rect 25865 3090 25931 3093
rect 0 3088 25931 3090
rect 0 3032 25870 3088
rect 25926 3032 25931 3088
rect 0 3030 25931 3032
rect 0 3000 120 3030
rect 25865 3027 25931 3030
rect 29729 3090 29795 3093
rect 31109 3090 31175 3093
rect 29729 3088 31175 3090
rect 29729 3032 29734 3088
rect 29790 3032 31114 3088
rect 31170 3032 31175 3088
rect 29729 3030 31175 3032
rect 29729 3027 29795 3030
rect 31109 3027 31175 3030
rect 47301 3090 47367 3093
rect 48880 3090 49000 3120
rect 47301 3088 49000 3090
rect 47301 3032 47306 3088
rect 47362 3032 49000 3088
rect 47301 3030 49000 3032
rect 47301 3027 47367 3030
rect 48880 3000 49000 3030
rect 17953 2954 18019 2957
rect 1718 2952 18019 2954
rect 1718 2896 17958 2952
rect 18014 2896 18019 2952
rect 1718 2894 18019 2896
rect 0 2818 120 2848
rect 1718 2818 1778 2894
rect 17953 2891 18019 2894
rect 24945 2954 25011 2957
rect 43161 2954 43227 2957
rect 24945 2952 43227 2954
rect 24945 2896 24950 2952
rect 25006 2896 43166 2952
rect 43222 2896 43227 2952
rect 24945 2894 43227 2896
rect 24945 2891 25011 2894
rect 43161 2891 43227 2894
rect 0 2758 1778 2818
rect 46933 2818 46999 2821
rect 48880 2818 49000 2848
rect 46933 2816 49000 2818
rect 46933 2760 46938 2816
rect 46994 2760 49000 2816
rect 46933 2758 49000 2760
rect 0 2728 120 2758
rect 46933 2755 46999 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 37946 2752 38262 2753
rect 37946 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38262 2752
rect 37946 2687 38262 2688
rect 43946 2752 44262 2753
rect 43946 2688 43952 2752
rect 44016 2688 44032 2752
rect 44096 2688 44112 2752
rect 44176 2688 44192 2752
rect 44256 2688 44262 2752
rect 48880 2728 49000 2758
rect 43946 2687 44262 2688
rect 0 2546 120 2576
rect 7649 2546 7715 2549
rect 0 2544 7715 2546
rect 0 2488 7654 2544
rect 7710 2488 7715 2544
rect 0 2486 7715 2488
rect 0 2456 120 2486
rect 7649 2483 7715 2486
rect 12525 2546 12591 2549
rect 40033 2546 40099 2549
rect 12525 2544 40099 2546
rect 12525 2488 12530 2544
rect 12586 2488 40038 2544
rect 40094 2488 40099 2544
rect 12525 2486 40099 2488
rect 12525 2483 12591 2486
rect 40033 2483 40099 2486
rect 47945 2546 48011 2549
rect 48880 2546 49000 2576
rect 47945 2544 49000 2546
rect 47945 2488 47950 2544
rect 48006 2488 49000 2544
rect 47945 2486 49000 2488
rect 47945 2483 48011 2486
rect 48880 2456 49000 2486
rect 5809 2410 5875 2413
rect 2822 2408 5875 2410
rect 2822 2352 5814 2408
rect 5870 2352 5875 2408
rect 2822 2350 5875 2352
rect 0 2274 120 2304
rect 2822 2274 2882 2350
rect 5809 2347 5875 2350
rect 12893 2410 12959 2413
rect 39205 2410 39271 2413
rect 12893 2408 39271 2410
rect 12893 2352 12898 2408
rect 12954 2352 39210 2408
rect 39266 2352 39271 2408
rect 12893 2350 39271 2352
rect 12893 2347 12959 2350
rect 39205 2347 39271 2350
rect 0 2214 2882 2274
rect 46933 2274 46999 2277
rect 48880 2274 49000 2304
rect 46933 2272 49000 2274
rect 46933 2216 46938 2272
rect 46994 2216 49000 2272
rect 46933 2214 49000 2216
rect 0 2184 120 2214
rect 46933 2211 46999 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 33006 2143 33322 2144
rect 39006 2208 39322 2209
rect 39006 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39322 2208
rect 39006 2143 39322 2144
rect 45006 2208 45322 2209
rect 45006 2144 45012 2208
rect 45076 2144 45092 2208
rect 45156 2144 45172 2208
rect 45236 2144 45252 2208
rect 45316 2144 45322 2208
rect 48880 2184 49000 2214
rect 45006 2143 45322 2144
rect 0 2002 120 2032
rect 1209 2002 1275 2005
rect 0 2000 1275 2002
rect 0 1944 1214 2000
rect 1270 1944 1275 2000
rect 0 1942 1275 1944
rect 0 1912 120 1942
rect 1209 1939 1275 1942
rect 18597 2002 18663 2005
rect 38101 2002 38167 2005
rect 18597 2000 38167 2002
rect 18597 1944 18602 2000
rect 18658 1944 38106 2000
rect 38162 1944 38167 2000
rect 18597 1942 38167 1944
rect 18597 1939 18663 1942
rect 38101 1939 38167 1942
rect 45829 2002 45895 2005
rect 48880 2002 49000 2032
rect 45829 2000 49000 2002
rect 45829 1944 45834 2000
rect 45890 1944 49000 2000
rect 45829 1942 49000 1944
rect 45829 1939 45895 1942
rect 48880 1912 49000 1942
rect 11513 1866 11579 1869
rect 27981 1866 28047 1869
rect 11513 1864 28047 1866
rect 11513 1808 11518 1864
rect 11574 1808 27986 1864
rect 28042 1808 28047 1864
rect 11513 1806 28047 1808
rect 11513 1803 11579 1806
rect 27981 1803 28047 1806
rect 0 1730 120 1760
rect 1301 1730 1367 1733
rect 0 1728 1367 1730
rect 0 1672 1306 1728
rect 1362 1672 1367 1728
rect 0 1670 1367 1672
rect 0 1640 120 1670
rect 1301 1667 1367 1670
rect 14917 1730 14983 1733
rect 38837 1730 38903 1733
rect 14917 1728 38903 1730
rect 14917 1672 14922 1728
rect 14978 1672 38842 1728
rect 38898 1672 38903 1728
rect 14917 1670 38903 1672
rect 14917 1667 14983 1670
rect 38837 1667 38903 1670
rect 46197 1730 46263 1733
rect 48880 1730 49000 1760
rect 46197 1728 49000 1730
rect 46197 1672 46202 1728
rect 46258 1672 49000 1728
rect 46197 1670 49000 1672
rect 46197 1667 46263 1670
rect 48880 1640 49000 1670
rect 17125 1594 17191 1597
rect 38469 1594 38535 1597
rect 17125 1592 38535 1594
rect 17125 1536 17130 1592
rect 17186 1536 38474 1592
rect 38530 1536 38535 1592
rect 17125 1534 38535 1536
rect 17125 1531 17191 1534
rect 38469 1531 38535 1534
rect 0 1458 120 1488
rect 1117 1458 1183 1461
rect 0 1456 1183 1458
rect 0 1400 1122 1456
rect 1178 1400 1183 1456
rect 0 1398 1183 1400
rect 0 1368 120 1398
rect 1117 1395 1183 1398
rect 46565 1458 46631 1461
rect 48880 1458 49000 1488
rect 46565 1456 49000 1458
rect 46565 1400 46570 1456
rect 46626 1400 49000 1456
rect 46565 1398 49000 1400
rect 46565 1395 46631 1398
rect 48880 1368 49000 1398
rect 11145 506 11211 509
rect 27521 506 27587 509
rect 11145 504 27587 506
rect 11145 448 11150 504
rect 11206 448 27526 504
rect 27582 448 27587 504
rect 11145 446 27587 448
rect 11145 443 11211 446
rect 27521 443 27587 446
rect 29913 506 29979 509
rect 44265 506 44331 509
rect 29913 504 44331 506
rect 29913 448 29918 504
rect 29974 448 44270 504
rect 44326 448 44331 504
rect 29913 446 44331 448
rect 29913 443 29979 446
rect 44265 443 44331 446
rect 18505 370 18571 373
rect 39665 370 39731 373
rect 18505 368 39731 370
rect 18505 312 18510 368
rect 18566 312 39670 368
rect 39726 312 39731 368
rect 18505 310 39731 312
rect 18505 307 18571 310
rect 39665 307 39731 310
rect 9305 234 9371 237
rect 31293 234 31359 237
rect 9305 232 31359 234
rect 9305 176 9310 232
rect 9366 176 31298 232
rect 31354 176 31359 232
rect 9305 174 31359 176
rect 9305 171 9371 174
rect 31293 171 31359 174
rect 17769 98 17835 101
rect 40125 98 40191 101
rect 17769 96 40191 98
rect 17769 40 17774 96
rect 17830 40 40130 96
rect 40186 40 40191 96
rect 17769 38 40191 40
rect 17769 35 17835 38
rect 40125 35 40191 38
<< via3 >>
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 39012 8732 39076 8736
rect 39012 8676 39016 8732
rect 39016 8676 39072 8732
rect 39072 8676 39076 8732
rect 39012 8672 39076 8676
rect 39092 8732 39156 8736
rect 39092 8676 39096 8732
rect 39096 8676 39152 8732
rect 39152 8676 39156 8732
rect 39092 8672 39156 8676
rect 39172 8732 39236 8736
rect 39172 8676 39176 8732
rect 39176 8676 39232 8732
rect 39232 8676 39236 8732
rect 39172 8672 39236 8676
rect 39252 8732 39316 8736
rect 39252 8676 39256 8732
rect 39256 8676 39312 8732
rect 39312 8676 39316 8732
rect 39252 8672 39316 8676
rect 45012 8732 45076 8736
rect 45012 8676 45016 8732
rect 45016 8676 45072 8732
rect 45072 8676 45076 8732
rect 45012 8672 45076 8676
rect 45092 8732 45156 8736
rect 45092 8676 45096 8732
rect 45096 8676 45152 8732
rect 45152 8676 45156 8732
rect 45092 8672 45156 8676
rect 45172 8732 45236 8736
rect 45172 8676 45176 8732
rect 45176 8676 45232 8732
rect 45232 8676 45236 8732
rect 45172 8672 45236 8676
rect 45252 8732 45316 8736
rect 45252 8676 45256 8732
rect 45256 8676 45312 8732
rect 45312 8676 45316 8732
rect 45252 8672 45316 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 37952 8188 38016 8192
rect 37952 8132 37956 8188
rect 37956 8132 38012 8188
rect 38012 8132 38016 8188
rect 37952 8128 38016 8132
rect 38032 8188 38096 8192
rect 38032 8132 38036 8188
rect 38036 8132 38092 8188
rect 38092 8132 38096 8188
rect 38032 8128 38096 8132
rect 38112 8188 38176 8192
rect 38112 8132 38116 8188
rect 38116 8132 38172 8188
rect 38172 8132 38176 8188
rect 38112 8128 38176 8132
rect 38192 8188 38256 8192
rect 38192 8132 38196 8188
rect 38196 8132 38252 8188
rect 38252 8132 38256 8188
rect 38192 8128 38256 8132
rect 43952 8188 44016 8192
rect 43952 8132 43956 8188
rect 43956 8132 44012 8188
rect 44012 8132 44016 8188
rect 43952 8128 44016 8132
rect 44032 8188 44096 8192
rect 44032 8132 44036 8188
rect 44036 8132 44092 8188
rect 44092 8132 44096 8188
rect 44032 8128 44096 8132
rect 44112 8188 44176 8192
rect 44112 8132 44116 8188
rect 44116 8132 44172 8188
rect 44172 8132 44176 8188
rect 44112 8128 44176 8132
rect 44192 8188 44256 8192
rect 44192 8132 44196 8188
rect 44196 8132 44252 8188
rect 44252 8132 44256 8188
rect 44192 8128 44256 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 39012 7644 39076 7648
rect 39012 7588 39016 7644
rect 39016 7588 39072 7644
rect 39072 7588 39076 7644
rect 39012 7584 39076 7588
rect 39092 7644 39156 7648
rect 39092 7588 39096 7644
rect 39096 7588 39152 7644
rect 39152 7588 39156 7644
rect 39092 7584 39156 7588
rect 39172 7644 39236 7648
rect 39172 7588 39176 7644
rect 39176 7588 39232 7644
rect 39232 7588 39236 7644
rect 39172 7584 39236 7588
rect 39252 7644 39316 7648
rect 39252 7588 39256 7644
rect 39256 7588 39312 7644
rect 39312 7588 39316 7644
rect 39252 7584 39316 7588
rect 45012 7644 45076 7648
rect 45012 7588 45016 7644
rect 45016 7588 45072 7644
rect 45072 7588 45076 7644
rect 45012 7584 45076 7588
rect 45092 7644 45156 7648
rect 45092 7588 45096 7644
rect 45096 7588 45152 7644
rect 45152 7588 45156 7644
rect 45092 7584 45156 7588
rect 45172 7644 45236 7648
rect 45172 7588 45176 7644
rect 45176 7588 45232 7644
rect 45232 7588 45236 7644
rect 45172 7584 45236 7588
rect 45252 7644 45316 7648
rect 45252 7588 45256 7644
rect 45256 7588 45312 7644
rect 45312 7588 45316 7644
rect 45252 7584 45316 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 37952 7100 38016 7104
rect 37952 7044 37956 7100
rect 37956 7044 38012 7100
rect 38012 7044 38016 7100
rect 37952 7040 38016 7044
rect 38032 7100 38096 7104
rect 38032 7044 38036 7100
rect 38036 7044 38092 7100
rect 38092 7044 38096 7100
rect 38032 7040 38096 7044
rect 38112 7100 38176 7104
rect 38112 7044 38116 7100
rect 38116 7044 38172 7100
rect 38172 7044 38176 7100
rect 38112 7040 38176 7044
rect 38192 7100 38256 7104
rect 38192 7044 38196 7100
rect 38196 7044 38252 7100
rect 38252 7044 38256 7100
rect 38192 7040 38256 7044
rect 43952 7100 44016 7104
rect 43952 7044 43956 7100
rect 43956 7044 44012 7100
rect 44012 7044 44016 7100
rect 43952 7040 44016 7044
rect 44032 7100 44096 7104
rect 44032 7044 44036 7100
rect 44036 7044 44092 7100
rect 44092 7044 44096 7100
rect 44032 7040 44096 7044
rect 44112 7100 44176 7104
rect 44112 7044 44116 7100
rect 44116 7044 44172 7100
rect 44172 7044 44176 7100
rect 44112 7040 44176 7044
rect 44192 7100 44256 7104
rect 44192 7044 44196 7100
rect 44196 7044 44252 7100
rect 44252 7044 44256 7100
rect 44192 7040 44256 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 39012 6556 39076 6560
rect 39012 6500 39016 6556
rect 39016 6500 39072 6556
rect 39072 6500 39076 6556
rect 39012 6496 39076 6500
rect 39092 6556 39156 6560
rect 39092 6500 39096 6556
rect 39096 6500 39152 6556
rect 39152 6500 39156 6556
rect 39092 6496 39156 6500
rect 39172 6556 39236 6560
rect 39172 6500 39176 6556
rect 39176 6500 39232 6556
rect 39232 6500 39236 6556
rect 39172 6496 39236 6500
rect 39252 6556 39316 6560
rect 39252 6500 39256 6556
rect 39256 6500 39312 6556
rect 39312 6500 39316 6556
rect 39252 6496 39316 6500
rect 45012 6556 45076 6560
rect 45012 6500 45016 6556
rect 45016 6500 45072 6556
rect 45072 6500 45076 6556
rect 45012 6496 45076 6500
rect 45092 6556 45156 6560
rect 45092 6500 45096 6556
rect 45096 6500 45152 6556
rect 45152 6500 45156 6556
rect 45092 6496 45156 6500
rect 45172 6556 45236 6560
rect 45172 6500 45176 6556
rect 45176 6500 45232 6556
rect 45232 6500 45236 6556
rect 45172 6496 45236 6500
rect 45252 6556 45316 6560
rect 45252 6500 45256 6556
rect 45256 6500 45312 6556
rect 45312 6500 45316 6556
rect 45252 6496 45316 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 37952 6012 38016 6016
rect 37952 5956 37956 6012
rect 37956 5956 38012 6012
rect 38012 5956 38016 6012
rect 37952 5952 38016 5956
rect 38032 6012 38096 6016
rect 38032 5956 38036 6012
rect 38036 5956 38092 6012
rect 38092 5956 38096 6012
rect 38032 5952 38096 5956
rect 38112 6012 38176 6016
rect 38112 5956 38116 6012
rect 38116 5956 38172 6012
rect 38172 5956 38176 6012
rect 38112 5952 38176 5956
rect 38192 6012 38256 6016
rect 38192 5956 38196 6012
rect 38196 5956 38252 6012
rect 38252 5956 38256 6012
rect 38192 5952 38256 5956
rect 43952 6012 44016 6016
rect 43952 5956 43956 6012
rect 43956 5956 44012 6012
rect 44012 5956 44016 6012
rect 43952 5952 44016 5956
rect 44032 6012 44096 6016
rect 44032 5956 44036 6012
rect 44036 5956 44092 6012
rect 44092 5956 44096 6012
rect 44032 5952 44096 5956
rect 44112 6012 44176 6016
rect 44112 5956 44116 6012
rect 44116 5956 44172 6012
rect 44172 5956 44176 6012
rect 44112 5952 44176 5956
rect 44192 6012 44256 6016
rect 44192 5956 44196 6012
rect 44196 5956 44252 6012
rect 44252 5956 44256 6012
rect 44192 5952 44256 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 39012 5468 39076 5472
rect 39012 5412 39016 5468
rect 39016 5412 39072 5468
rect 39072 5412 39076 5468
rect 39012 5408 39076 5412
rect 39092 5468 39156 5472
rect 39092 5412 39096 5468
rect 39096 5412 39152 5468
rect 39152 5412 39156 5468
rect 39092 5408 39156 5412
rect 39172 5468 39236 5472
rect 39172 5412 39176 5468
rect 39176 5412 39232 5468
rect 39232 5412 39236 5468
rect 39172 5408 39236 5412
rect 39252 5468 39316 5472
rect 39252 5412 39256 5468
rect 39256 5412 39312 5468
rect 39312 5412 39316 5468
rect 39252 5408 39316 5412
rect 45012 5468 45076 5472
rect 45012 5412 45016 5468
rect 45016 5412 45072 5468
rect 45072 5412 45076 5468
rect 45012 5408 45076 5412
rect 45092 5468 45156 5472
rect 45092 5412 45096 5468
rect 45096 5412 45152 5468
rect 45152 5412 45156 5468
rect 45092 5408 45156 5412
rect 45172 5468 45236 5472
rect 45172 5412 45176 5468
rect 45176 5412 45232 5468
rect 45232 5412 45236 5468
rect 45172 5408 45236 5412
rect 45252 5468 45316 5472
rect 45252 5412 45256 5468
rect 45256 5412 45312 5468
rect 45312 5412 45316 5468
rect 45252 5408 45316 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 37952 4924 38016 4928
rect 37952 4868 37956 4924
rect 37956 4868 38012 4924
rect 38012 4868 38016 4924
rect 37952 4864 38016 4868
rect 38032 4924 38096 4928
rect 38032 4868 38036 4924
rect 38036 4868 38092 4924
rect 38092 4868 38096 4924
rect 38032 4864 38096 4868
rect 38112 4924 38176 4928
rect 38112 4868 38116 4924
rect 38116 4868 38172 4924
rect 38172 4868 38176 4924
rect 38112 4864 38176 4868
rect 38192 4924 38256 4928
rect 38192 4868 38196 4924
rect 38196 4868 38252 4924
rect 38252 4868 38256 4924
rect 38192 4864 38256 4868
rect 43952 4924 44016 4928
rect 43952 4868 43956 4924
rect 43956 4868 44012 4924
rect 44012 4868 44016 4924
rect 43952 4864 44016 4868
rect 44032 4924 44096 4928
rect 44032 4868 44036 4924
rect 44036 4868 44092 4924
rect 44092 4868 44096 4924
rect 44032 4864 44096 4868
rect 44112 4924 44176 4928
rect 44112 4868 44116 4924
rect 44116 4868 44172 4924
rect 44172 4868 44176 4924
rect 44112 4864 44176 4868
rect 44192 4924 44256 4928
rect 44192 4868 44196 4924
rect 44196 4868 44252 4924
rect 44252 4868 44256 4924
rect 44192 4864 44256 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 39012 4380 39076 4384
rect 39012 4324 39016 4380
rect 39016 4324 39072 4380
rect 39072 4324 39076 4380
rect 39012 4320 39076 4324
rect 39092 4380 39156 4384
rect 39092 4324 39096 4380
rect 39096 4324 39152 4380
rect 39152 4324 39156 4380
rect 39092 4320 39156 4324
rect 39172 4380 39236 4384
rect 39172 4324 39176 4380
rect 39176 4324 39232 4380
rect 39232 4324 39236 4380
rect 39172 4320 39236 4324
rect 39252 4380 39316 4384
rect 39252 4324 39256 4380
rect 39256 4324 39312 4380
rect 39312 4324 39316 4380
rect 39252 4320 39316 4324
rect 45012 4380 45076 4384
rect 45012 4324 45016 4380
rect 45016 4324 45072 4380
rect 45072 4324 45076 4380
rect 45012 4320 45076 4324
rect 45092 4380 45156 4384
rect 45092 4324 45096 4380
rect 45096 4324 45152 4380
rect 45152 4324 45156 4380
rect 45092 4320 45156 4324
rect 45172 4380 45236 4384
rect 45172 4324 45176 4380
rect 45176 4324 45232 4380
rect 45232 4324 45236 4380
rect 45172 4320 45236 4324
rect 45252 4380 45316 4384
rect 45252 4324 45256 4380
rect 45256 4324 45312 4380
rect 45312 4324 45316 4380
rect 45252 4320 45316 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 37952 3836 38016 3840
rect 37952 3780 37956 3836
rect 37956 3780 38012 3836
rect 38012 3780 38016 3836
rect 37952 3776 38016 3780
rect 38032 3836 38096 3840
rect 38032 3780 38036 3836
rect 38036 3780 38092 3836
rect 38092 3780 38096 3836
rect 38032 3776 38096 3780
rect 38112 3836 38176 3840
rect 38112 3780 38116 3836
rect 38116 3780 38172 3836
rect 38172 3780 38176 3836
rect 38112 3776 38176 3780
rect 38192 3836 38256 3840
rect 38192 3780 38196 3836
rect 38196 3780 38252 3836
rect 38252 3780 38256 3836
rect 38192 3776 38256 3780
rect 43952 3836 44016 3840
rect 43952 3780 43956 3836
rect 43956 3780 44012 3836
rect 44012 3780 44016 3836
rect 43952 3776 44016 3780
rect 44032 3836 44096 3840
rect 44032 3780 44036 3836
rect 44036 3780 44092 3836
rect 44092 3780 44096 3836
rect 44032 3776 44096 3780
rect 44112 3836 44176 3840
rect 44112 3780 44116 3836
rect 44116 3780 44172 3836
rect 44172 3780 44176 3836
rect 44112 3776 44176 3780
rect 44192 3836 44256 3840
rect 44192 3780 44196 3836
rect 44196 3780 44252 3836
rect 44252 3780 44256 3836
rect 44192 3776 44256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 39012 3292 39076 3296
rect 39012 3236 39016 3292
rect 39016 3236 39072 3292
rect 39072 3236 39076 3292
rect 39012 3232 39076 3236
rect 39092 3292 39156 3296
rect 39092 3236 39096 3292
rect 39096 3236 39152 3292
rect 39152 3236 39156 3292
rect 39092 3232 39156 3236
rect 39172 3292 39236 3296
rect 39172 3236 39176 3292
rect 39176 3236 39232 3292
rect 39232 3236 39236 3292
rect 39172 3232 39236 3236
rect 39252 3292 39316 3296
rect 39252 3236 39256 3292
rect 39256 3236 39312 3292
rect 39312 3236 39316 3292
rect 39252 3232 39316 3236
rect 45012 3292 45076 3296
rect 45012 3236 45016 3292
rect 45016 3236 45072 3292
rect 45072 3236 45076 3292
rect 45012 3232 45076 3236
rect 45092 3292 45156 3296
rect 45092 3236 45096 3292
rect 45096 3236 45152 3292
rect 45152 3236 45156 3292
rect 45092 3232 45156 3236
rect 45172 3292 45236 3296
rect 45172 3236 45176 3292
rect 45176 3236 45232 3292
rect 45232 3236 45236 3292
rect 45172 3232 45236 3236
rect 45252 3292 45316 3296
rect 45252 3236 45256 3292
rect 45256 3236 45312 3292
rect 45312 3236 45316 3292
rect 45252 3232 45316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 37952 2748 38016 2752
rect 37952 2692 37956 2748
rect 37956 2692 38012 2748
rect 38012 2692 38016 2748
rect 37952 2688 38016 2692
rect 38032 2748 38096 2752
rect 38032 2692 38036 2748
rect 38036 2692 38092 2748
rect 38092 2692 38096 2748
rect 38032 2688 38096 2692
rect 38112 2748 38176 2752
rect 38112 2692 38116 2748
rect 38116 2692 38172 2748
rect 38172 2692 38176 2748
rect 38112 2688 38176 2692
rect 38192 2748 38256 2752
rect 38192 2692 38196 2748
rect 38196 2692 38252 2748
rect 38252 2692 38256 2748
rect 38192 2688 38256 2692
rect 43952 2748 44016 2752
rect 43952 2692 43956 2748
rect 43956 2692 44012 2748
rect 44012 2692 44016 2748
rect 43952 2688 44016 2692
rect 44032 2748 44096 2752
rect 44032 2692 44036 2748
rect 44036 2692 44092 2748
rect 44092 2692 44096 2748
rect 44032 2688 44096 2692
rect 44112 2748 44176 2752
rect 44112 2692 44116 2748
rect 44116 2692 44172 2748
rect 44172 2692 44176 2748
rect 44112 2688 44176 2692
rect 44192 2748 44256 2752
rect 44192 2692 44196 2748
rect 44196 2692 44252 2748
rect 44252 2692 44256 2748
rect 44192 2688 44256 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
rect 39012 2204 39076 2208
rect 39012 2148 39016 2204
rect 39016 2148 39072 2204
rect 39072 2148 39076 2204
rect 39012 2144 39076 2148
rect 39092 2204 39156 2208
rect 39092 2148 39096 2204
rect 39096 2148 39152 2204
rect 39152 2148 39156 2204
rect 39092 2144 39156 2148
rect 39172 2204 39236 2208
rect 39172 2148 39176 2204
rect 39176 2148 39232 2204
rect 39232 2148 39236 2204
rect 39172 2144 39236 2148
rect 39252 2204 39316 2208
rect 39252 2148 39256 2204
rect 39256 2148 39312 2204
rect 39312 2148 39316 2204
rect 39252 2144 39316 2148
rect 45012 2204 45076 2208
rect 45012 2148 45016 2204
rect 45016 2148 45072 2204
rect 45072 2148 45076 2204
rect 45012 2144 45076 2148
rect 45092 2204 45156 2208
rect 45092 2148 45096 2204
rect 45096 2148 45152 2204
rect 45152 2148 45156 2204
rect 45092 2144 45156 2148
rect 45172 2204 45236 2208
rect 45172 2148 45176 2204
rect 45176 2148 45232 2204
rect 45232 2148 45236 2204
rect 45172 2144 45236 2148
rect 45252 2204 45316 2208
rect 45252 2148 45256 2204
rect 45256 2148 45312 2204
rect 45312 2148 45316 2204
rect 45252 2144 45316 2148
<< metal4 >>
rect 1944 8192 2264 11250
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 8736 3324 11250
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11250
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 8736 9324 11250
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 8192 14264 11250
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13944 0 14264 2688
rect 15004 8736 15324 11250
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 8192 20264 11250
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19944 0 20264 2688
rect 21004 8736 21324 11250
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 21004 6560 21324 7584
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25944 8192 26264 11250
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25944 0 26264 2688
rect 27004 8736 27324 11250
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 31944 8192 32264 11250
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 0 32264 2688
rect 33004 8736 33324 11250
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
rect 37944 8192 38264 11250
rect 37944 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38264 8192
rect 37944 7104 38264 8128
rect 37944 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38264 7104
rect 37944 6016 38264 7040
rect 37944 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38264 6016
rect 37944 4928 38264 5952
rect 37944 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38264 4928
rect 37944 3840 38264 4864
rect 37944 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38264 3840
rect 37944 2752 38264 3776
rect 37944 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38264 2752
rect 37944 0 38264 2688
rect 39004 8736 39324 11250
rect 39004 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39324 8736
rect 39004 7648 39324 8672
rect 39004 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39324 7648
rect 39004 6560 39324 7584
rect 39004 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39324 6560
rect 39004 5472 39324 6496
rect 39004 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39324 5472
rect 39004 4384 39324 5408
rect 39004 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39324 4384
rect 39004 3296 39324 4320
rect 39004 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39324 3296
rect 39004 2208 39324 3232
rect 39004 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39324 2208
rect 39004 0 39324 2144
rect 43944 8192 44264 11250
rect 43944 8128 43952 8192
rect 44016 8128 44032 8192
rect 44096 8128 44112 8192
rect 44176 8128 44192 8192
rect 44256 8128 44264 8192
rect 43944 7104 44264 8128
rect 43944 7040 43952 7104
rect 44016 7040 44032 7104
rect 44096 7040 44112 7104
rect 44176 7040 44192 7104
rect 44256 7040 44264 7104
rect 43944 6016 44264 7040
rect 43944 5952 43952 6016
rect 44016 5952 44032 6016
rect 44096 5952 44112 6016
rect 44176 5952 44192 6016
rect 44256 5952 44264 6016
rect 43944 4928 44264 5952
rect 43944 4864 43952 4928
rect 44016 4864 44032 4928
rect 44096 4864 44112 4928
rect 44176 4864 44192 4928
rect 44256 4864 44264 4928
rect 43944 3840 44264 4864
rect 43944 3776 43952 3840
rect 44016 3776 44032 3840
rect 44096 3776 44112 3840
rect 44176 3776 44192 3840
rect 44256 3776 44264 3840
rect 43944 2752 44264 3776
rect 43944 2688 43952 2752
rect 44016 2688 44032 2752
rect 44096 2688 44112 2752
rect 44176 2688 44192 2752
rect 44256 2688 44264 2752
rect 43944 0 44264 2688
rect 45004 8736 45324 11250
rect 45004 8672 45012 8736
rect 45076 8672 45092 8736
rect 45156 8672 45172 8736
rect 45236 8672 45252 8736
rect 45316 8672 45324 8736
rect 45004 7648 45324 8672
rect 45004 7584 45012 7648
rect 45076 7584 45092 7648
rect 45156 7584 45172 7648
rect 45236 7584 45252 7648
rect 45316 7584 45324 7648
rect 45004 6560 45324 7584
rect 45004 6496 45012 6560
rect 45076 6496 45092 6560
rect 45156 6496 45172 6560
rect 45236 6496 45252 6560
rect 45316 6496 45324 6560
rect 45004 5472 45324 6496
rect 45004 5408 45012 5472
rect 45076 5408 45092 5472
rect 45156 5408 45172 5472
rect 45236 5408 45252 5472
rect 45316 5408 45324 5472
rect 45004 4384 45324 5408
rect 45004 4320 45012 4384
rect 45076 4320 45092 4384
rect 45156 4320 45172 4384
rect 45236 4320 45252 4384
rect 45316 4320 45324 4384
rect 45004 3296 45324 4320
rect 45004 3232 45012 3296
rect 45076 3232 45092 3296
rect 45156 3232 45172 3296
rect 45236 3232 45252 3296
rect 45316 3232 45324 3296
rect 45004 2208 45324 3232
rect 45004 2144 45012 2208
rect 45076 2144 45092 2208
rect 45156 2144 45172 2208
rect 45236 2144 45252 2208
rect 45316 2144 45324 2208
rect 45004 0 45324 2144
use sky130_fd_sc_hd__clkbuf_2  _000_
timestamp -3599
transform 1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _001_
timestamp -3599
transform 1 0 27416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _002_
timestamp -3599
transform 1 0 26864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _003_
timestamp -3599
transform 1 0 32936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _004_
timestamp -3599
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _005_
timestamp -3599
transform -1 0 46736 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _006_
timestamp -3599
transform -1 0 46460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _007_
timestamp -3599
transform -1 0 42688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _008_
timestamp -3599
transform -1 0 46736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _009_
timestamp -3599
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _010_
timestamp -3599
transform -1 0 40480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _011_
timestamp -3599
transform 1 0 33212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _012_
timestamp -3599
transform 1 0 26128 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _013_
timestamp -3599
transform 1 0 23092 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _014_
timestamp -3599
transform 1 0 14260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _015_
timestamp -3599
transform 1 0 17940 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _016_
timestamp -3599
transform 1 0 19504 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _017_
timestamp -3599
transform 1 0 24932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _018_
timestamp -3599
transform 1 0 18584 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _019_
timestamp -3599
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _020_
timestamp -3599
transform 1 0 19688 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _021_
timestamp -3599
transform 1 0 18124 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _022_
timestamp -3599
transform 1 0 26864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _023_
timestamp -3599
transform 1 0 18584 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _024_
timestamp -3599
transform 1 0 26312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _025_
timestamp -3599
transform -1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _026_
timestamp -3599
transform 1 0 19320 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _027_
timestamp -3599
transform 1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _028_
timestamp -3599
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _029_
timestamp -3599
transform 1 0 1932 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _030_
timestamp -3599
transform 1 0 15732 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _031_
timestamp -3599
transform 1 0 46184 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _032_
timestamp -3599
transform -1 0 38364 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _033_
timestamp -3599
transform -1 0 39008 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _034_
timestamp -3599
transform -1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _035_
timestamp -3599
transform -1 0 10304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _036_
timestamp -3599
transform -1 0 12328 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp -3599
transform -1 0 15088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _038_
timestamp -3599
transform 1 0 17848 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _039_
timestamp -3599
transform 1 0 20608 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp -3599
transform 1 0 23460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp -3599
transform 1 0 26036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _042_
timestamp -3599
transform -1 0 40296 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp -3599
transform 1 0 29808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _044_
timestamp -3599
transform -1 0 41584 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp -3599
transform 1 0 42412 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp -3599
transform 1 0 43332 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp -3599
transform 1 0 39560 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp -3599
transform 1 0 40756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp -3599
transform 1 0 44528 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp -3599
transform 1 0 46460 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp -3599
transform -1 0 46736 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _052_
timestamp -3599
transform 1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _053_
timestamp -3599
transform 1 0 2668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _054_
timestamp -3599
transform 1 0 11960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _055_
timestamp -3599
transform -1 0 16192 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _056_
timestamp -3599
transform 1 0 4784 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _057_
timestamp -3599
transform 1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _058_
timestamp -3599
transform 1 0 4232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _059_
timestamp -3599
transform 1 0 3956 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp -3599
transform -1 0 20608 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp -3599
transform -1 0 21160 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp -3599
transform -1 0 21436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp -3599
transform -1 0 22264 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _064_
timestamp -3599
transform 1 0 8464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _065_
timestamp -3599
transform 1 0 8740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _066_
timestamp -3599
transform 1 0 7360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _067_
timestamp -3599
transform 1 0 6256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp -3599
transform -1 0 23920 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp -3599
transform -1 0 24196 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp -3599
transform -1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp -3599
transform -1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp -3599
transform -1 0 25024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _073_
timestamp -3599
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _074_
timestamp -3599
transform 1 0 10396 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp -3599
transform -1 0 26312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _076_
timestamp -3599
transform 1 0 9200 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp -3599
transform -1 0 8740 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _078_
timestamp -3599
transform 1 0 8096 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _079_
timestamp -3599
transform 1 0 8372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp -3599
transform -1 0 28428 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp -3599
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp -3599
transform -1 0 29440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp -3599
transform -1 0 29900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp -3599
transform -1 0 30360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp -3599
transform -1 0 30912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp -3599
transform -1 0 31556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp -3599
transform -1 0 32108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp -3599
transform -1 0 32752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp -3599
transform -1 0 33396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp -3599
transform -1 0 34040 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _091_
timestamp -3599
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp -3599
transform -1 0 35604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp -3599
transform 1 0 39376 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _094_
timestamp -3599
transform -1 0 45724 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp -3599
transform 1 0 40388 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _096_
timestamp -3599
transform 1 0 17480 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _097_
timestamp -3599
transform 1 0 17020 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp -3599
transform -1 0 16560 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _099_
timestamp -3599
transform 1 0 15272 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _100_
timestamp -3599
transform 1 0 14536 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _101_
timestamp -3599
transform 1 0 13708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _102_
timestamp -3599
transform 1 0 12696 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _103_
timestamp -3599
transform 1 0 12236 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp -3599
transform -1 0 38088 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform -1 0 40204 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform 1 0 33028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform -1 0 26128 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform 1 0 22908 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform -1 0 14260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform -1 0 17940 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 19504 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform -1 0 18584 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform -1 0 22264 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform 1 0 19504 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform 1 0 17940 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform 1 0 26680 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform 1 0 25576 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform -1 0 24196 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform -1 0 19780 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp -3599
transform 1 0 21712 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp -3599
transform -1 0 26864 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp -3599
transform 1 0 15548 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp -3599
transform 1 0 46000 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp -3599
transform -1 0 32936 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp -3599
transform -1 0 27416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp -3599
transform -1 0 46920 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp -3599
transform -1 0 46184 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp -3599
transform -1 0 42872 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp -3599
transform 1 0 46276 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp -3599
transform 1 0 46920 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp -3599
transform -1 0 8096 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp -3599
transform -1 0 12052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp -3599
transform -1 0 23460 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp -3599
transform 1 0 23184 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp -3599
transform -1 0 30636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp -3599
transform -1 0 28612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp -3599
transform 1 0 27968 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp -3599
transform -1 0 35328 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp -3599
transform 1 0 33580 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp -3599
transform -1 0 33120 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp -3599
transform -1 0 40388 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp -3599
transform -1 0 45448 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp -3599
transform -1 0 30084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp -3599
transform 1 0 30084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp -3599
transform 1 0 30820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp -3599
transform -1 0 31924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp -3599
transform -1 0 26036 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_45
timestamp -3599
transform 1 0 23460 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_46
timestamp -3599
transform 1 0 25852 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636964856
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636964856
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636964856
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636964856
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636964856
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636964856
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636964856
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636964856
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -3599
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636964856
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636964856
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -3599
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636964856
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636964856
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -3599
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636964856
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636964856
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp -3599
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636964856
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_209
timestamp -3599
transform 1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_225
timestamp -3599
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_253
timestamp -3599
transform 1 0 24380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp -3599
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -3599
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_321
timestamp -3599
transform 1 0 30636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp -3599
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp -3599
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp -3599
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp -3599
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_429
timestamp 1636964856
transform 1 0 40572 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_441
timestamp -3599
transform 1 0 41676 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp -3599
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1636964856
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1636964856
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp -3599
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_477
timestamp -3599
transform 1 0 44988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_483
timestamp -3599
transform 1 0 45540 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636964856
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636964856
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636964856
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636964856
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp -3599
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -3599
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636964856
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636964856
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636964856
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636964856
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp -3599
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -3599
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636964856
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636964856
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_137
timestamp -3599
transform 1 0 13708 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_147
timestamp 1636964856
transform 1 0 14628 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp -3599
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -3599
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636964856
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_187
timestamp -3599
transform 1 0 18308 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_195
timestamp -3599
transform 1 0 19044 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_204
timestamp 1636964856
transform 1 0 19872 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_216
timestamp -3599
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_225
timestamp -3599
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_230
timestamp 1636964856
transform 1 0 22264 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_242
timestamp 1636964856
transform 1 0 23368 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_254
timestamp -3599
transform 1 0 24472 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_260
timestamp -3599
transform 1 0 25024 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_268
timestamp -3599
transform 1 0 25760 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_274
timestamp -3599
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_281
timestamp -3599
transform 1 0 26956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_289
timestamp -3599
transform 1 0 27692 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_297
timestamp 1636964856
transform 1 0 28428 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_309
timestamp -3599
transform 1 0 29532 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_317
timestamp -3599
transform 1 0 30268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_325
timestamp -3599
transform 1 0 31004 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_330
timestamp -3599
transform 1 0 31464 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636964856
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_349
timestamp -3599
transform 1 0 33212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_353
timestamp -3599
transform 1 0 33580 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_358
timestamp 1636964856
transform 1 0 34040 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_370
timestamp 1636964856
transform 1 0 35144 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_386
timestamp -3599
transform 1 0 36616 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636964856
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_405
timestamp -3599
transform 1 0 38364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_409
timestamp -3599
transform 1 0 38732 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_414
timestamp 1636964856
transform 1 0 39192 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_426
timestamp 1636964856
transform 1 0 40296 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_438
timestamp -3599
transform 1 0 41400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp -3599
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1636964856
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1636964856
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1636964856
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_485
timestamp -3599
transform 1 0 45724 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_491
timestamp -3599
transform 1 0 46276 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636964856
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636964856
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636964856
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636964856
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636964856
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636964856
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636964856
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636964856
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636964856
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636964856
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp -3599
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp -3599
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636964856
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636964856
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636964856
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636964856
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp -3599
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp -3599
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636964856
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636964856
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636964856
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636964856
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_245
timestamp -3599
transform 1 0 23644 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp -3599
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_256
timestamp 1636964856
transform 1 0 24656 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_268
timestamp 1636964856
transform 1 0 25760 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_280
timestamp 1636964856
transform 1 0 26864 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_292
timestamp -3599
transform 1 0 27968 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_296
timestamp -3599
transform 1 0 28336 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_302
timestamp -3599
transform 1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_309
timestamp -3599
transform 1 0 29532 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_313
timestamp -3599
transform 1 0 29900 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_318
timestamp -3599
transform 1 0 30360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_324
timestamp -3599
transform 1 0 30912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_331
timestamp -3599
transform 1 0 31556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_337
timestamp -3599
transform 1 0 32108 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_344
timestamp -3599
transform 1 0 32752 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_351
timestamp 1636964856
transform 1 0 33396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp -3599
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636964856
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636964856
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636964856
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1636964856
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp -3599
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp -3599
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636964856
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636964856
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1636964856
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1636964856
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp -3599
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp -3599
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_477
timestamp -3599
transform 1 0 44988 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_485
timestamp -3599
transform 1 0 45724 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_502
timestamp -3599
transform 1 0 47288 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636964856
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636964856
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636964856
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp -3599
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -3599
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp -3599
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_65
timestamp -3599
transform 1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_71
timestamp -3599
transform 1 0 7636 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_79
timestamp -3599
transform 1 0 8372 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_86
timestamp 1636964856
transform 1 0 9016 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_98
timestamp 1636964856
transform 1 0 10120 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp -3599
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636964856
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636964856
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636964856
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636964856
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp -3599
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -3599
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636964856
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_181
timestamp -3599
transform 1 0 17756 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_187
timestamp -3599
transform 1 0 18308 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_194
timestamp 1636964856
transform 1 0 18952 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_206
timestamp 1636964856
transform 1 0 20056 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_218
timestamp -3599
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636964856
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636964856
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636964856
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636964856
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp -3599
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp -3599
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636964856
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636964856
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636964856
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636964856
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp -3599
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp -3599
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636964856
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636964856
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636964856
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636964856
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp -3599
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp -3599
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636964856
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636964856
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_417
timestamp -3599
transform 1 0 39468 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_428
timestamp 1636964856
transform 1 0 40480 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_440
timestamp -3599
transform 1 0 41584 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_454
timestamp 1636964856
transform 1 0 42872 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_466
timestamp 1636964856
transform 1 0 43976 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_478
timestamp 1636964856
transform 1 0 45080 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_490
timestamp -3599
transform 1 0 46184 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_11
timestamp -3599
transform 1 0 2116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp -3599
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp -3599
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_37
timestamp -3599
transform 1 0 4508 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_43
timestamp -3599
transform 1 0 5060 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_47
timestamp -3599
transform 1 0 5428 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_51
timestamp -3599
transform 1 0 5796 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_55
timestamp -3599
transform 1 0 6164 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_59
timestamp 1636964856
transform 1 0 6532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_71
timestamp 1636964856
transform 1 0 7636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -3599
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636964856
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636964856
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636964856
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636964856
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp -3599
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp -3599
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636964856
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636964856
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636964856
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636964856
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp -3599
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp -3599
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_200
timestamp 1636964856
transform 1 0 19504 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_212
timestamp -3599
transform 1 0 20608 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636964856
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636964856
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp -3599
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp -3599
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636964856
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636964856
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_277
timestamp -3599
transform 1 0 26588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_283
timestamp 1636964856
transform 1 0 27140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_295
timestamp 1636964856
transform 1 0 28244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp -3599
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636964856
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636964856
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1636964856
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1636964856
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp -3599
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp -3599
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636964856
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636964856
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1636964856
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1636964856
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp -3599
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp -3599
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636964856
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636964856
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1636964856
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1636964856
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp -3599
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp -3599
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1636964856
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_489
timestamp -3599
transform 1 0 46092 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636964856
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636964856
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636964856
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636964856
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp -3599
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp -3599
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636964856
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_69
timestamp -3599
transform 1 0 7452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_75
timestamp -3599
transform 1 0 8004 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_82
timestamp -3599
transform 1 0 8648 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_91
timestamp -3599
transform 1 0 9476 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_99
timestamp -3599
transform 1 0 10212 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_104
timestamp -3599
transform 1 0 10672 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_108
timestamp -3599
transform 1 0 11040 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp -3599
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_125
timestamp -3599
transform 1 0 12604 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_129
timestamp -3599
transform 1 0 12972 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_140
timestamp 1636964856
transform 1 0 13984 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_152
timestamp -3599
transform 1 0 15088 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_157
timestamp -3599
transform 1 0 15548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_176
timestamp -3599
transform 1 0 17296 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636964856
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636964856
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636964856
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp -3599
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp -3599
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_230
timestamp -3599
transform 1 0 22264 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_238
timestamp -3599
transform 1 0 23000 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_242
timestamp -3599
transform 1 0 23368 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_251
timestamp -3599
transform 1 0 24196 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_262
timestamp 1636964856
transform 1 0 25208 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp -3599
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_289
timestamp 1636964856
transform 1 0 27692 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_301
timestamp 1636964856
transform 1 0 28796 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_313
timestamp 1636964856
transform 1 0 29900 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_325
timestamp -3599
transform 1 0 31004 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_333
timestamp -3599
transform 1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636964856
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636964856
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636964856
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636964856
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp -3599
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp -3599
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636964856
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1636964856
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1636964856
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1636964856
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp -3599
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp -3599
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1636964856
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1636964856
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1636964856
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_485
timestamp -3599
transform 1 0 45724 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_493
timestamp -3599
transform 1 0 46460 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636964856
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636964856
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636964856
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636964856
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636964856
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636964856
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_77
timestamp -3599
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp -3599
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636964856
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636964856
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636964856
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1636964856
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp -3599
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp -3599
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp -3599
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_145
timestamp -3599
transform 1 0 14444 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_149
timestamp 1636964856
transform 1 0 14812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_161
timestamp 1636964856
transform 1 0 15916 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_173
timestamp -3599
transform 1 0 17020 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_181
timestamp -3599
transform 1 0 17756 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp -3599
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp -3599
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_197
timestamp -3599
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_205
timestamp 1636964856
transform 1 0 19964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_217
timestamp 1636964856
transform 1 0 21068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_229
timestamp 1636964856
transform 1 0 22172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_241
timestamp -3599
transform 1 0 23276 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp -3599
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636964856
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636964856
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1636964856
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1636964856
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp -3599
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp -3599
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636964856
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1636964856
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_333
timestamp -3599
transform 1 0 31740 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_341
timestamp -3599
transform 1 0 32476 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_349
timestamp 1636964856
transform 1 0 33212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_361
timestamp -3599
transform 1 0 34316 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636964856
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1636964856
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1636964856
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1636964856
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp -3599
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp -3599
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1636964856
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1636964856
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1636964856
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1636964856
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp -3599
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp -3599
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1636964856
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_489
timestamp -3599
transform 1 0 46092 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636964856
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636964856
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636964856
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636964856
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp -3599
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -3599
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636964856
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636964856
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636964856
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1636964856
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp -3599
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp -3599
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636964856
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636964856
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1636964856
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1636964856
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp -3599
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp -3599
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636964856
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636964856
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1636964856
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1636964856
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp -3599
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp -3599
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp -3599
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_230
timestamp 1636964856
transform 1 0 22264 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_242
timestamp 1636964856
transform 1 0 23368 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_254
timestamp 1636964856
transform 1 0 24472 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_266
timestamp 1636964856
transform 1 0 25576 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp -3599
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636964856
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1636964856
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1636964856
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1636964856
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp -3599
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp -3599
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1636964856
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_349
timestamp -3599
transform 1 0 33212 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_358
timestamp 1636964856
transform 1 0 34040 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_370
timestamp 1636964856
transform 1 0 35144 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_382
timestamp -3599
transform 1 0 36248 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_390
timestamp -3599
transform 1 0 36984 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1636964856
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1636964856
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1636964856
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1636964856
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp -3599
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp -3599
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_452
timestamp -3599
transform 1 0 42688 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_458
timestamp -3599
transform 1 0 43240 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_462
timestamp 1636964856
transform 1 0 43608 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_474
timestamp 1636964856
transform 1 0 44712 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_486
timestamp -3599
transform 1 0 45816 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636964856
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636964856
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -3599
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636964856
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636964856
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636964856
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636964856
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp -3599
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp -3599
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636964856
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1636964856
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1636964856
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1636964856
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp -3599
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp -3599
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636964856
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_153
timestamp -3599
transform 1 0 15180 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_163
timestamp 1636964856
transform 1 0 16100 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_175
timestamp 1636964856
transform 1 0 17204 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_187
timestamp -3599
transform 1 0 18308 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp -3599
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636964856
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636964856
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1636964856
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1636964856
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp -3599
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp -3599
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636964856
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_265
timestamp -3599
transform 1 0 25484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_269
timestamp -3599
transform 1 0 25852 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_275
timestamp -3599
transform 1 0 26404 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_283
timestamp 1636964856
transform 1 0 27140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_295
timestamp 1636964856
transform 1 0 28244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp -3599
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1636964856
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1636964856
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1636964856
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1636964856
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp -3599
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp -3599
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1636964856
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1636964856
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1636964856
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1636964856
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp -3599
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp -3599
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_421
timestamp -3599
transform 1 0 39836 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_426
timestamp -3599
transform 1 0 40296 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_434
timestamp -3599
transform 1 0 41032 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_440
timestamp 1636964856
transform 1 0 41584 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_452
timestamp 1636964856
transform 1 0 42688 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_464
timestamp -3599
transform 1 0 43792 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp -3599
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_477
timestamp -3599
transform 1 0 44988 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_485
timestamp -3599
transform 1 0 45724 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_496
timestamp -3599
transform 1 0 46736 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636964856
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636964856
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636964856
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1636964856
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp -3599
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -3599
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636964856
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636964856
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1636964856
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1636964856
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp -3599
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp -3599
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_122
timestamp 1636964856
transform 1 0 12328 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_134
timestamp 1636964856
transform 1 0 13432 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_146
timestamp -3599
transform 1 0 14536 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_152
timestamp 1636964856
transform 1 0 15088 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp -3599
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636964856
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_181
timestamp -3599
transform 1 0 17756 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_185
timestamp 1636964856
transform 1 0 18124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_197
timestamp 1636964856
transform 1 0 19228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_209
timestamp 1636964856
transform 1 0 20332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp -3599
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1636964856
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_242
timestamp 1636964856
transform 1 0 23368 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_254
timestamp 1636964856
transform 1 0 24472 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_266
timestamp 1636964856
transform 1 0 25576 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp -3599
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636964856
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1636964856
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1636964856
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1636964856
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp -3599
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp -3599
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_337
timestamp -3599
transform 1 0 32108 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_345
timestamp -3599
transform 1 0 32844 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_352
timestamp 1636964856
transform 1 0 33488 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_364
timestamp 1636964856
transform 1 0 34592 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_376
timestamp 1636964856
transform 1 0 35696 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_388
timestamp -3599
transform 1 0 36800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_393
timestamp -3599
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_405
timestamp -3599
transform 1 0 38364 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_412
timestamp -3599
transform 1 0 39008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_421
timestamp -3599
transform 1 0 39836 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_429
timestamp -3599
transform 1 0 40572 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_434
timestamp 1636964856
transform 1 0 41032 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_446
timestamp -3599
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1636964856
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1636964856
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1636964856
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_485
timestamp -3599
transform 1 0 45724 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_13
timestamp 1636964856
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp -3599
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636964856
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636964856
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1636964856
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_65
timestamp -3599
transform 1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_73
timestamp -3599
transform 1 0 7820 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_79
timestamp -3599
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp -3599
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636964856
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_100
timestamp 1636964856
transform 1 0 10304 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_112
timestamp -3599
transform 1 0 11408 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1636964856
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp -3599
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp -3599
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1636964856
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_153
timestamp -3599
transform 1 0 15180 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_164
timestamp 1636964856
transform 1 0 16192 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_176
timestamp 1636964856
transform 1 0 17296 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_188
timestamp -3599
transform 1 0 18400 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_197
timestamp -3599
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_203
timestamp -3599
transform 1 0 19780 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_218
timestamp -3599
transform 1 0 21160 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_229
timestamp 1636964856
transform 1 0 22172 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp -3599
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1636964856
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_265
timestamp -3599
transform 1 0 25484 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_268
timestamp -3599
transform 1 0 25760 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1636964856
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1636964856
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp -3599
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp -3599
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_315
timestamp 1636964856
transform 1 0 30084 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_327
timestamp 1636964856
transform 1 0 31188 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_339
timestamp 1636964856
transform 1 0 32292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_351
timestamp 1636964856
transform 1 0 33396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp -3599
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_365
timestamp -3599
transform 1 0 34684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_369
timestamp -3599
transform 1 0 35052 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_375
timestamp 1636964856
transform 1 0 35604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_387
timestamp -3599
transform 1 0 36708 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_395
timestamp -3599
transform 1 0 37444 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_402
timestamp 1636964856
transform 1 0 38088 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_414
timestamp -3599
transform 1 0 39192 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp -3599
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_421
timestamp -3599
transform 1 0 39836 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_430
timestamp 1636964856
transform 1 0 40664 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_442
timestamp 1636964856
transform 1 0 41768 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_454
timestamp 1636964856
transform 1 0 42872 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_466
timestamp -3599
transform 1 0 43976 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_474
timestamp -3599
transform 1 0 44712 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_477
timestamp -3599
transform 1 0 44988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_7
timestamp 1636964856
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_19
timestamp -3599
transform 1 0 2852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_27
timestamp -3599
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_33
timestamp 1636964856
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_45
timestamp -3599
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp -3599
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_61
timestamp 1636964856
transform 1 0 6716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_73
timestamp -3599
transform 1 0 7820 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_83
timestamp -3599
transform 1 0 8740 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_85
timestamp 1636964856
transform 1 0 8924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_97
timestamp -3599
transform 1 0 10028 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_103
timestamp -3599
transform 1 0 10580 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp -3599
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1636964856
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_125
timestamp -3599
transform 1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_133
timestamp -3599
transform 1 0 13340 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_139
timestamp -3599
transform 1 0 13892 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_141
timestamp 1636964856
transform 1 0 14076 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_153
timestamp -3599
transform 1 0 15180 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_158
timestamp -3599
transform 1 0 15640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp -3599
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_169
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_177
timestamp -3599
transform 1 0 17388 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_183
timestamp 1636964856
transform 1 0 17940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_195
timestamp -3599
transform 1 0 19044 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_197
timestamp -3599
transform 1 0 19228 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_203
timestamp -3599
transform 1 0 19780 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_208
timestamp 1636964856
transform 1 0 20240 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp -3599
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_225
timestamp -3599
transform 1 0 21804 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_233
timestamp 1636964856
transform 1 0 22540 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_245
timestamp -3599
transform 1 0 23644 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_251
timestamp -3599
transform 1 0 24196 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_253
timestamp -3599
transform 1 0 24380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_258
timestamp 1636964856
transform 1 0 24840 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_270
timestamp -3599
transform 1 0 25944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp -3599
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_285
timestamp 1636964856
transform 1 0 27324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_297
timestamp -3599
transform 1 0 28428 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_303
timestamp -3599
transform 1 0 28980 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_309
timestamp 1636964856
transform 1 0 29532 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_321
timestamp -3599
transform 1 0 30636 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp -3599
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1636964856
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_349
timestamp -3599
transform 1 0 33212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_353
timestamp -3599
transform 1 0 33580 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_358
timestamp -3599
transform 1 0 34040 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_365
timestamp 1636964856
transform 1 0 34684 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_377
timestamp -3599
transform 1 0 35788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_383
timestamp -3599
transform 1 0 36340 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp -3599
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_393
timestamp -3599
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_401
timestamp -3599
transform 1 0 37996 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_408
timestamp 1636964856
transform 1 0 38640 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_421
timestamp -3599
transform 1 0 39836 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_433
timestamp 1636964856
transform 1 0 40940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_445
timestamp -3599
transform 1 0 42044 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_449
timestamp -3599
transform 1 0 42412 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_453
timestamp -3599
transform 1 0 42780 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_458
timestamp 1636964856
transform 1 0 43240 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_470
timestamp -3599
transform 1 0 44344 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_477
timestamp -3599
transform 1 0 44988 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_483
timestamp -3599
transform 1 0 45540 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output1
timestamp -3599
transform 1 0 46368 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform 1 0 46828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform 1 0 47196 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform 1 0 46736 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 46828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform 1 0 47196 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 46552 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -3599
transform 1 0 47104 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -3599
transform 1 0 46828 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -3599
transform 1 0 46000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp -3599
transform 1 0 47196 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp -3599
transform 1 0 47104 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp -3599
transform 1 0 46828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp -3599
transform 1 0 47196 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp -3599
transform 1 0 47104 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -3599
transform 1 0 46368 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp -3599
transform 1 0 46000 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp -3599
transform 1 0 45632 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp -3599
transform 1 0 46460 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp -3599
transform 1 0 46736 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp -3599
transform 1 0 45632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp -3599
transform 1 0 46092 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp -3599
transform -1 0 46092 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp -3599
transform 1 0 46736 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp -3599
transform 1 0 46368 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp -3599
transform 1 0 46736 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp -3599
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp -3599
transform 1 0 46920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp -3599
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp -3599
transform 1 0 46736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp -3599
transform -1 0 4140 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp -3599
transform -1 0 27324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp -3599
transform -1 0 29440 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp -3599
transform -1 0 31740 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp -3599
transform -1 0 34040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp -3599
transform -1 0 36340 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp -3599
transform -1 0 38640 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp -3599
transform -1 0 40940 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp -3599
transform -1 0 43240 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp -3599
transform -1 0 45540 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp -3599
transform 1 0 46736 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp -3599
transform -1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp -3599
transform 1 0 8372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp -3599
transform 1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp -3599
transform 1 0 12972 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp -3599
transform 1 0 15272 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp -3599
transform -1 0 17940 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp -3599
transform -1 0 20240 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp -3599
transform -1 0 22540 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp -3599
transform -1 0 24840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp -3599
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp -3599
transform 1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp -3599
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp -3599
transform 1 0 21896 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp -3599
transform 1 0 22080 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp -3599
transform 1 0 22448 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp -3599
transform 1 0 22816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp -3599
transform 1 0 23184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp -3599
transform 1 0 23552 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp -3599
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp -3599
transform 1 0 24472 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp -3599
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp -3599
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp -3599
transform 1 0 25576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp -3599
transform 1 0 25944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp -3599
transform 1 0 26312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp -3599
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp -3599
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp -3599
transform 1 0 27692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp -3599
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp -3599
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp -3599
transform 1 0 32476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp -3599
transform 1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp -3599
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform 1 0 33948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform 1 0 33672 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform 1 0 28796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform -1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform 1 0 29900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform 1 0 30268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform 1 0 30636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform -1 0 31740 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform 1 0 31096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform 1 0 38732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform 1 0 39100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform 1 0 39836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform 1 0 40204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform 1 0 35052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform 1 0 35420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform -1 0 36892 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform -1 0 36616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform -1 0 37628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform 1 0 37628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform 1 0 37996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output105
timestamp -3599
transform -1 0 1748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 47840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 47840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 47840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 47840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 47840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 47840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 47840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 47840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 47840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 47840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 47840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 47840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_38
timestamp -3599
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_39
timestamp -3599
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_40
timestamp -3599
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_41
timestamp -3599
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_45
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_46
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_47
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_48
timestamp -3599
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_49
timestamp -3599
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_50
timestamp -3599
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_52
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_53
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_54
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_55
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_56
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_57
timestamp -3599
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_58
timestamp -3599
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_59
timestamp -3599
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_60
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_61
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_62
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_63
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_64
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_65
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_66
timestamp -3599
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_67
timestamp -3599
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_68
timestamp -3599
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_69
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_70
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_71
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_72
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_73
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_74
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_75
timestamp -3599
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_76
timestamp -3599
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_77
timestamp -3599
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_78
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_79
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_80
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_81
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_82
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_83
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_84
timestamp -3599
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_85
timestamp -3599
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_86
timestamp -3599
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_87
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_88
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_89
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_90
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_91
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_92
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_93
timestamp -3599
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_94
timestamp -3599
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_95
timestamp -3599
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_96
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_97
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_98
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_99
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_100
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_101
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_102
timestamp -3599
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_103
timestamp -3599
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_104
timestamp -3599
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_105
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_106
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_107
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_108
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_109
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_110
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_111
timestamp -3599
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_112
timestamp -3599
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_113
timestamp -3599
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_114
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_115
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_116
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_117
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_118
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_119
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_120
timestamp -3599
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_121
timestamp -3599
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_122
timestamp -3599
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_123
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_124
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_125
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_126
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_127
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp -3599
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp -3599
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp -3599
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_132
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_133
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_136
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_137
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_138
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_139
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_140
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_141
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_142
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_143
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_144
timestamp -3599
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_145
timestamp -3599
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_146
timestamp -3599
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_147
timestamp -3599
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_148
timestamp -3599
transform 1 0 44896 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_149
timestamp -3599
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 9800 120 9920 0 FreeSans 480 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 48880 1368 49000 1488 0 FreeSans 480 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 48880 4088 49000 4208 0 FreeSans 480 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 48880 4360 49000 4480 0 FreeSans 480 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 48880 4632 49000 4752 0 FreeSans 480 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 48880 4904 49000 5024 0 FreeSans 480 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 48880 5176 49000 5296 0 FreeSans 480 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 48880 5448 49000 5568 0 FreeSans 480 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 48880 5720 49000 5840 0 FreeSans 480 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 48880 5992 49000 6112 0 FreeSans 480 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 48880 6264 49000 6384 0 FreeSans 480 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 48880 6536 49000 6656 0 FreeSans 480 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 48880 1640 49000 1760 0 FreeSans 480 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 48880 6808 49000 6928 0 FreeSans 480 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 48880 7080 49000 7200 0 FreeSans 480 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 48880 7352 49000 7472 0 FreeSans 480 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 48880 7624 49000 7744 0 FreeSans 480 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 48880 7896 49000 8016 0 FreeSans 480 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 48880 8168 49000 8288 0 FreeSans 480 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 48880 8440 49000 8560 0 FreeSans 480 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 48880 8712 49000 8832 0 FreeSans 480 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 48880 8984 49000 9104 0 FreeSans 480 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 48880 9256 49000 9376 0 FreeSans 480 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 48880 1912 49000 2032 0 FreeSans 480 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 48880 9528 49000 9648 0 FreeSans 480 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 48880 9800 49000 9920 0 FreeSans 480 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 48880 2184 49000 2304 0 FreeSans 480 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 48880 2456 49000 2576 0 FreeSans 480 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 48880 2728 49000 2848 0 FreeSans 480 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 48880 3000 49000 3120 0 FreeSans 480 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 48880 3272 49000 3392 0 FreeSans 480 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 48880 3544 49000 3664 0 FreeSans 480 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 48880 3816 49000 3936 0 FreeSans 480 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 40222 0 40278 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 43902 0 43958 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 44270 0 44326 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 44638 0 44694 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 45006 0 45062 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 45374 0 45430 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 45742 0 45798 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 46110 0 46166 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 46478 0 46534 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 46846 0 46902 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 47214 0 47270 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 40590 0 40646 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 40958 0 41014 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 41326 0 41382 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 41694 0 41750 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 42062 0 42118 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 42430 0 42486 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 42798 0 42854 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 43166 0 43222 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 43534 0 43590 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 3698 11194 3754 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 26698 11194 26754 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 28998 11194 29054 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 31298 11194 31354 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 33598 11194 33654 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 35898 11194 35954 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 38198 11194 38254 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 40498 11194 40554 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 42798 11194 42854 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 45098 11194 45154 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 47398 11194 47454 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 5998 11194 6054 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 8298 11194 8354 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 10598 11194 10654 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 12898 11194 12954 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 15198 11194 15254 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 17498 11194 17554 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 19798 11194 19854 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 22098 11194 22154 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 24398 11194 24454 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 1582 0 1638 56 0 FreeSans 224 0 0 0 N1END[0]
port 104 nsew signal input
flabel metal2 s 1950 0 2006 56 0 FreeSans 224 0 0 0 N1END[1]
port 105 nsew signal input
flabel metal2 s 2318 0 2374 56 0 FreeSans 224 0 0 0 N1END[2]
port 106 nsew signal input
flabel metal2 s 2686 0 2742 56 0 FreeSans 224 0 0 0 N1END[3]
port 107 nsew signal input
flabel metal2 s 5998 0 6054 56 0 FreeSans 224 0 0 0 N2END[0]
port 108 nsew signal input
flabel metal2 s 6366 0 6422 56 0 FreeSans 224 0 0 0 N2END[1]
port 109 nsew signal input
flabel metal2 s 6734 0 6790 56 0 FreeSans 224 0 0 0 N2END[2]
port 110 nsew signal input
flabel metal2 s 7102 0 7158 56 0 FreeSans 224 0 0 0 N2END[3]
port 111 nsew signal input
flabel metal2 s 7470 0 7526 56 0 FreeSans 224 0 0 0 N2END[4]
port 112 nsew signal input
flabel metal2 s 7838 0 7894 56 0 FreeSans 224 0 0 0 N2END[5]
port 113 nsew signal input
flabel metal2 s 8206 0 8262 56 0 FreeSans 224 0 0 0 N2END[6]
port 114 nsew signal input
flabel metal2 s 8574 0 8630 56 0 FreeSans 224 0 0 0 N2END[7]
port 115 nsew signal input
flabel metal2 s 3054 0 3110 56 0 FreeSans 224 0 0 0 N2MID[0]
port 116 nsew signal input
flabel metal2 s 3422 0 3478 56 0 FreeSans 224 0 0 0 N2MID[1]
port 117 nsew signal input
flabel metal2 s 3790 0 3846 56 0 FreeSans 224 0 0 0 N2MID[2]
port 118 nsew signal input
flabel metal2 s 4158 0 4214 56 0 FreeSans 224 0 0 0 N2MID[3]
port 119 nsew signal input
flabel metal2 s 4526 0 4582 56 0 FreeSans 224 0 0 0 N2MID[4]
port 120 nsew signal input
flabel metal2 s 4894 0 4950 56 0 FreeSans 224 0 0 0 N2MID[5]
port 121 nsew signal input
flabel metal2 s 5262 0 5318 56 0 FreeSans 224 0 0 0 N2MID[6]
port 122 nsew signal input
flabel metal2 s 5630 0 5686 56 0 FreeSans 224 0 0 0 N2MID[7]
port 123 nsew signal input
flabel metal2 s 8942 0 8998 56 0 FreeSans 224 0 0 0 N4END[0]
port 124 nsew signal input
flabel metal2 s 12622 0 12678 56 0 FreeSans 224 0 0 0 N4END[10]
port 125 nsew signal input
flabel metal2 s 12990 0 13046 56 0 FreeSans 224 0 0 0 N4END[11]
port 126 nsew signal input
flabel metal2 s 13358 0 13414 56 0 FreeSans 224 0 0 0 N4END[12]
port 127 nsew signal input
flabel metal2 s 13726 0 13782 56 0 FreeSans 224 0 0 0 N4END[13]
port 128 nsew signal input
flabel metal2 s 14094 0 14150 56 0 FreeSans 224 0 0 0 N4END[14]
port 129 nsew signal input
flabel metal2 s 14462 0 14518 56 0 FreeSans 224 0 0 0 N4END[15]
port 130 nsew signal input
flabel metal2 s 9310 0 9366 56 0 FreeSans 224 0 0 0 N4END[1]
port 131 nsew signal input
flabel metal2 s 9678 0 9734 56 0 FreeSans 224 0 0 0 N4END[2]
port 132 nsew signal input
flabel metal2 s 10046 0 10102 56 0 FreeSans 224 0 0 0 N4END[3]
port 133 nsew signal input
flabel metal2 s 10414 0 10470 56 0 FreeSans 224 0 0 0 N4END[4]
port 134 nsew signal input
flabel metal2 s 10782 0 10838 56 0 FreeSans 224 0 0 0 N4END[5]
port 135 nsew signal input
flabel metal2 s 11150 0 11206 56 0 FreeSans 224 0 0 0 N4END[6]
port 136 nsew signal input
flabel metal2 s 11518 0 11574 56 0 FreeSans 224 0 0 0 N4END[7]
port 137 nsew signal input
flabel metal2 s 11886 0 11942 56 0 FreeSans 224 0 0 0 N4END[8]
port 138 nsew signal input
flabel metal2 s 12254 0 12310 56 0 FreeSans 224 0 0 0 N4END[9]
port 139 nsew signal input
flabel metal2 s 14830 0 14886 56 0 FreeSans 224 0 0 0 NN4END[0]
port 140 nsew signal input
flabel metal2 s 18510 0 18566 56 0 FreeSans 224 0 0 0 NN4END[10]
port 141 nsew signal input
flabel metal2 s 18878 0 18934 56 0 FreeSans 224 0 0 0 NN4END[11]
port 142 nsew signal input
flabel metal2 s 19246 0 19302 56 0 FreeSans 224 0 0 0 NN4END[12]
port 143 nsew signal input
flabel metal2 s 19614 0 19670 56 0 FreeSans 224 0 0 0 NN4END[13]
port 144 nsew signal input
flabel metal2 s 19982 0 20038 56 0 FreeSans 224 0 0 0 NN4END[14]
port 145 nsew signal input
flabel metal2 s 20350 0 20406 56 0 FreeSans 224 0 0 0 NN4END[15]
port 146 nsew signal input
flabel metal2 s 15198 0 15254 56 0 FreeSans 224 0 0 0 NN4END[1]
port 147 nsew signal input
flabel metal2 s 15566 0 15622 56 0 FreeSans 224 0 0 0 NN4END[2]
port 148 nsew signal input
flabel metal2 s 15934 0 15990 56 0 FreeSans 224 0 0 0 NN4END[3]
port 149 nsew signal input
flabel metal2 s 16302 0 16358 56 0 FreeSans 224 0 0 0 NN4END[4]
port 150 nsew signal input
flabel metal2 s 16670 0 16726 56 0 FreeSans 224 0 0 0 NN4END[5]
port 151 nsew signal input
flabel metal2 s 17038 0 17094 56 0 FreeSans 224 0 0 0 NN4END[6]
port 152 nsew signal input
flabel metal2 s 17406 0 17462 56 0 FreeSans 224 0 0 0 NN4END[7]
port 153 nsew signal input
flabel metal2 s 17774 0 17830 56 0 FreeSans 224 0 0 0 NN4END[8]
port 154 nsew signal input
flabel metal2 s 18142 0 18198 56 0 FreeSans 224 0 0 0 NN4END[9]
port 155 nsew signal input
flabel metal2 s 20718 0 20774 56 0 FreeSans 224 0 0 0 S1BEG[0]
port 156 nsew signal output
flabel metal2 s 21086 0 21142 56 0 FreeSans 224 0 0 0 S1BEG[1]
port 157 nsew signal output
flabel metal2 s 21454 0 21510 56 0 FreeSans 224 0 0 0 S1BEG[2]
port 158 nsew signal output
flabel metal2 s 21822 0 21878 56 0 FreeSans 224 0 0 0 S1BEG[3]
port 159 nsew signal output
flabel metal2 s 22190 0 22246 56 0 FreeSans 224 0 0 0 S2BEG[0]
port 160 nsew signal output
flabel metal2 s 22558 0 22614 56 0 FreeSans 224 0 0 0 S2BEG[1]
port 161 nsew signal output
flabel metal2 s 22926 0 22982 56 0 FreeSans 224 0 0 0 S2BEG[2]
port 162 nsew signal output
flabel metal2 s 23294 0 23350 56 0 FreeSans 224 0 0 0 S2BEG[3]
port 163 nsew signal output
flabel metal2 s 23662 0 23718 56 0 FreeSans 224 0 0 0 S2BEG[4]
port 164 nsew signal output
flabel metal2 s 24030 0 24086 56 0 FreeSans 224 0 0 0 S2BEG[5]
port 165 nsew signal output
flabel metal2 s 24398 0 24454 56 0 FreeSans 224 0 0 0 S2BEG[6]
port 166 nsew signal output
flabel metal2 s 24766 0 24822 56 0 FreeSans 224 0 0 0 S2BEG[7]
port 167 nsew signal output
flabel metal2 s 25134 0 25190 56 0 FreeSans 224 0 0 0 S2BEGb[0]
port 168 nsew signal output
flabel metal2 s 25502 0 25558 56 0 FreeSans 224 0 0 0 S2BEGb[1]
port 169 nsew signal output
flabel metal2 s 25870 0 25926 56 0 FreeSans 224 0 0 0 S2BEGb[2]
port 170 nsew signal output
flabel metal2 s 26238 0 26294 56 0 FreeSans 224 0 0 0 S2BEGb[3]
port 171 nsew signal output
flabel metal2 s 26606 0 26662 56 0 FreeSans 224 0 0 0 S2BEGb[4]
port 172 nsew signal output
flabel metal2 s 26974 0 27030 56 0 FreeSans 224 0 0 0 S2BEGb[5]
port 173 nsew signal output
flabel metal2 s 27342 0 27398 56 0 FreeSans 224 0 0 0 S2BEGb[6]
port 174 nsew signal output
flabel metal2 s 27710 0 27766 56 0 FreeSans 224 0 0 0 S2BEGb[7]
port 175 nsew signal output
flabel metal2 s 28078 0 28134 56 0 FreeSans 224 0 0 0 S4BEG[0]
port 176 nsew signal output
flabel metal2 s 31758 0 31814 56 0 FreeSans 224 0 0 0 S4BEG[10]
port 177 nsew signal output
flabel metal2 s 32126 0 32182 56 0 FreeSans 224 0 0 0 S4BEG[11]
port 178 nsew signal output
flabel metal2 s 32494 0 32550 56 0 FreeSans 224 0 0 0 S4BEG[12]
port 179 nsew signal output
flabel metal2 s 32862 0 32918 56 0 FreeSans 224 0 0 0 S4BEG[13]
port 180 nsew signal output
flabel metal2 s 33230 0 33286 56 0 FreeSans 224 0 0 0 S4BEG[14]
port 181 nsew signal output
flabel metal2 s 33598 0 33654 56 0 FreeSans 224 0 0 0 S4BEG[15]
port 182 nsew signal output
flabel metal2 s 28446 0 28502 56 0 FreeSans 224 0 0 0 S4BEG[1]
port 183 nsew signal output
flabel metal2 s 28814 0 28870 56 0 FreeSans 224 0 0 0 S4BEG[2]
port 184 nsew signal output
flabel metal2 s 29182 0 29238 56 0 FreeSans 224 0 0 0 S4BEG[3]
port 185 nsew signal output
flabel metal2 s 29550 0 29606 56 0 FreeSans 224 0 0 0 S4BEG[4]
port 186 nsew signal output
flabel metal2 s 29918 0 29974 56 0 FreeSans 224 0 0 0 S4BEG[5]
port 187 nsew signal output
flabel metal2 s 30286 0 30342 56 0 FreeSans 224 0 0 0 S4BEG[6]
port 188 nsew signal output
flabel metal2 s 30654 0 30710 56 0 FreeSans 224 0 0 0 S4BEG[7]
port 189 nsew signal output
flabel metal2 s 31022 0 31078 56 0 FreeSans 224 0 0 0 S4BEG[8]
port 190 nsew signal output
flabel metal2 s 31390 0 31446 56 0 FreeSans 224 0 0 0 S4BEG[9]
port 191 nsew signal output
flabel metal2 s 33966 0 34022 56 0 FreeSans 224 0 0 0 SS4BEG[0]
port 192 nsew signal output
flabel metal2 s 37646 0 37702 56 0 FreeSans 224 0 0 0 SS4BEG[10]
port 193 nsew signal output
flabel metal2 s 38014 0 38070 56 0 FreeSans 224 0 0 0 SS4BEG[11]
port 194 nsew signal output
flabel metal2 s 38382 0 38438 56 0 FreeSans 224 0 0 0 SS4BEG[12]
port 195 nsew signal output
flabel metal2 s 38750 0 38806 56 0 FreeSans 224 0 0 0 SS4BEG[13]
port 196 nsew signal output
flabel metal2 s 39118 0 39174 56 0 FreeSans 224 0 0 0 SS4BEG[14]
port 197 nsew signal output
flabel metal2 s 39486 0 39542 56 0 FreeSans 224 0 0 0 SS4BEG[15]
port 198 nsew signal output
flabel metal2 s 34334 0 34390 56 0 FreeSans 224 0 0 0 SS4BEG[1]
port 199 nsew signal output
flabel metal2 s 34702 0 34758 56 0 FreeSans 224 0 0 0 SS4BEG[2]
port 200 nsew signal output
flabel metal2 s 35070 0 35126 56 0 FreeSans 224 0 0 0 SS4BEG[3]
port 201 nsew signal output
flabel metal2 s 35438 0 35494 56 0 FreeSans 224 0 0 0 SS4BEG[4]
port 202 nsew signal output
flabel metal2 s 35806 0 35862 56 0 FreeSans 224 0 0 0 SS4BEG[5]
port 203 nsew signal output
flabel metal2 s 36174 0 36230 56 0 FreeSans 224 0 0 0 SS4BEG[6]
port 204 nsew signal output
flabel metal2 s 36542 0 36598 56 0 FreeSans 224 0 0 0 SS4BEG[7]
port 205 nsew signal output
flabel metal2 s 36910 0 36966 56 0 FreeSans 224 0 0 0 SS4BEG[8]
port 206 nsew signal output
flabel metal2 s 37278 0 37334 56 0 FreeSans 224 0 0 0 SS4BEG[9]
port 207 nsew signal output
flabel metal2 s 39854 0 39910 56 0 FreeSans 224 0 0 0 UserCLK
port 208 nsew signal input
flabel metal2 s 1398 11194 1454 11250 0 FreeSans 224 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal4 s 3004 0 3324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 3004 11190 3324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 11190 9324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 11190 15324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 11190 21324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 11190 27324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 11190 33324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 0 39324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 0 39324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 11190 39324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 45004 0 45324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 45004 0 45324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 45004 11190 45324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 1944 11190 2264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 0 8264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 11190 8264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 0 14264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 11190 14264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 0 20264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 11190 20264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 0 26264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 11190 26264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 0 32264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 11190 32264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 0 38264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 0 38264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 11190 38264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 43944 0 44264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 43944 0 44264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 43944 11190 44264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
rlabel metal1 24472 8704 24472 8704 0 VGND
rlabel metal1 24472 8160 24472 8160 0 VPWR
rlabel metal3 620 1428 620 1428 0 FrameData[0]
rlabel via2 40066 4131 40066 4131 0 FrameData[10]
rlabel metal3 298 4420 298 4420 0 FrameData[11]
rlabel metal1 25944 6630 25944 6630 0 FrameData[12]
rlabel metal3 942 4964 942 4964 0 FrameData[13]
rlabel metal3 3495 5236 3495 5236 0 FrameData[14]
rlabel metal3 1471 5508 1471 5508 0 FrameData[15]
rlabel metal3 1931 5780 1931 5780 0 FrameData[16]
rlabel metal3 919 6052 919 6052 0 FrameData[17]
rlabel metal3 11684 6256 11684 6256 0 FrameData[18]
rlabel metal3 1471 6596 1471 6596 0 FrameData[19]
rlabel metal3 712 1700 712 1700 0 FrameData[1]
rlabel metal1 19412 5882 19412 5882 0 FrameData[20]
rlabel metal3 919 7140 919 7140 0 FrameData[21]
rlabel metal3 712 7412 712 7412 0 FrameData[22]
rlabel metal3 1471 7684 1471 7684 0 FrameData[23]
rlabel metal2 25622 7905 25622 7905 0 FrameData[24]
rlabel metal3 942 8228 942 8228 0 FrameData[25]
rlabel metal2 19366 8177 19366 8177 0 FrameData[26]
rlabel metal3 1494 8772 1494 8772 0 FrameData[27]
rlabel metal2 7590 8517 7590 8517 0 FrameData[28]
rlabel metal3 574 9316 574 9316 0 FrameData[29]
rlabel metal3 666 1972 666 1972 0 FrameData[2]
rlabel metal3 6186 9588 6186 9588 0 FrameData[30]
rlabel metal3 1334 6460 1334 6460 0 FrameData[31]
rlabel metal3 1471 2244 1471 2244 0 FrameData[3]
rlabel metal2 7682 4080 7682 4080 0 FrameData[4]
rlabel metal3 919 2788 919 2788 0 FrameData[5]
rlabel metal2 25898 3621 25898 3621 0 FrameData[6]
rlabel metal3 1471 3332 1471 3332 0 FrameData[7]
rlabel metal2 46322 3757 46322 3757 0 FrameData[8]
rlabel metal3 712 3876 712 3876 0 FrameData[9]
rlabel metal3 47754 1428 47754 1428 0 FrameData_O[0]
rlabel metal3 48122 4148 48122 4148 0 FrameData_O[10]
rlabel metal3 47984 4420 47984 4420 0 FrameData_O[11]
rlabel metal3 48168 4692 48168 4692 0 FrameData_O[12]
rlabel metal3 47938 4964 47938 4964 0 FrameData_O[13]
rlabel metal3 48122 5236 48122 5236 0 FrameData_O[14]
rlabel metal3 47984 5508 47984 5508 0 FrameData_O[15]
rlabel metal3 48168 5780 48168 5780 0 FrameData_O[16]
rlabel metal3 47846 6052 47846 6052 0 FrameData_O[17]
rlabel metal3 48122 6324 48122 6324 0 FrameData_O[18]
rlabel metal3 47984 6596 47984 6596 0 FrameData_O[19]
rlabel metal3 47570 1700 47570 1700 0 FrameData_O[1]
rlabel metal3 48168 6868 48168 6868 0 FrameData_O[20]
rlabel metal3 48122 7140 48122 7140 0 FrameData_O[21]
rlabel metal3 47984 7412 47984 7412 0 FrameData_O[22]
rlabel metal3 48168 7684 48168 7684 0 FrameData_O[23]
rlabel metal3 48122 7956 48122 7956 0 FrameData_O[24]
rlabel metal3 48076 8228 48076 8228 0 FrameData_O[25]
rlabel metal3 47570 8500 47570 8500 0 FrameData_O[26]
rlabel metal2 45862 8687 45862 8687 0 FrameData_O[27]
rlabel metal2 46690 8551 46690 8551 0 FrameData_O[28]
rlabel metal2 46966 8415 46966 8415 0 FrameData_O[29]
rlabel metal3 47386 1972 47386 1972 0 FrameData_O[2]
rlabel metal2 46322 8653 46322 8653 0 FrameData_O[30]
rlabel metal1 45908 7718 45908 7718 0 FrameData_O[31]
rlabel metal3 47938 2244 47938 2244 0 FrameData_O[3]
rlabel metal3 48444 2516 48444 2516 0 FrameData_O[4]
rlabel metal3 47938 2788 47938 2788 0 FrameData_O[5]
rlabel metal3 48122 3060 48122 3060 0 FrameData_O[6]
rlabel metal3 48030 3332 48030 3332 0 FrameData_O[7]
rlabel metal2 47334 3383 47334 3383 0 FrameData_O[8]
rlabel metal3 47938 3876 47938 3876 0 FrameData_O[9]
rlabel metal1 39514 7174 39514 7174 0 FrameStrobe[0]
rlabel metal2 43930 718 43930 718 0 FrameStrobe[10]
rlabel metal2 44298 259 44298 259 0 FrameStrobe[11]
rlabel metal1 43102 6766 43102 6766 0 FrameStrobe[12]
rlabel metal2 45034 718 45034 718 0 FrameStrobe[13]
rlabel metal1 44482 6290 44482 6290 0 FrameStrobe[14]
rlabel metal1 39790 7344 39790 7344 0 FrameStrobe[15]
rlabel metal2 46138 1401 46138 1401 0 FrameStrobe[16]
rlabel metal2 46506 1401 46506 1401 0 FrameStrobe[17]
rlabel metal2 46874 1401 46874 1401 0 FrameStrobe[18]
rlabel metal2 47380 5100 47380 5100 0 FrameStrobe[19]
rlabel metal1 39744 7242 39744 7242 0 FrameStrobe[1]
rlabel metal1 9982 7718 9982 7718 0 FrameStrobe[2]
rlabel metal1 10718 7310 10718 7310 0 FrameStrobe[3]
rlabel metal1 12052 7378 12052 7378 0 FrameStrobe[4]
rlabel metal1 14858 7344 14858 7344 0 FrameStrobe[5]
rlabel metal2 18078 6868 18078 6868 0 FrameStrobe[6]
rlabel metal2 20838 7650 20838 7650 0 FrameStrobe[7]
rlabel metal1 23690 7820 23690 7820 0 FrameStrobe[8]
rlabel metal2 36570 1768 36570 1768 0 FrameStrobe[9]
rlabel metal1 3818 8602 3818 8602 0 FrameStrobe_O[0]
rlabel metal1 26910 8602 26910 8602 0 FrameStrobe_O[10]
rlabel metal1 29118 8602 29118 8602 0 FrameStrobe_O[11]
rlabel metal1 31418 8602 31418 8602 0 FrameStrobe_O[12]
rlabel metal1 33718 8602 33718 8602 0 FrameStrobe_O[13]
rlabel metal1 36018 8602 36018 8602 0 FrameStrobe_O[14]
rlabel metal1 38318 8602 38318 8602 0 FrameStrobe_O[15]
rlabel metal1 40618 8602 40618 8602 0 FrameStrobe_O[16]
rlabel metal1 42918 8602 42918 8602 0 FrameStrobe_O[17]
rlabel metal1 45356 8602 45356 8602 0 FrameStrobe_O[18]
rlabel metal1 47196 8602 47196 8602 0 FrameStrobe_O[19]
rlabel metal1 6256 8602 6256 8602 0 FrameStrobe_O[1]
rlabel metal1 8464 8602 8464 8602 0 FrameStrobe_O[2]
rlabel metal1 10764 8602 10764 8602 0 FrameStrobe_O[3]
rlabel metal1 13064 8602 13064 8602 0 FrameStrobe_O[4]
rlabel metal1 15456 8602 15456 8602 0 FrameStrobe_O[5]
rlabel metal1 17618 8602 17618 8602 0 FrameStrobe_O[6]
rlabel metal1 19918 8602 19918 8602 0 FrameStrobe_O[7]
rlabel metal1 22218 8602 22218 8602 0 FrameStrobe_O[8]
rlabel metal1 24518 8602 24518 8602 0 FrameStrobe_O[9]
rlabel metal2 1610 3744 1610 3744 0 N1END[0]
rlabel metal2 1978 1279 1978 1279 0 N1END[1]
rlabel metal2 2346 2282 2346 2282 0 N1END[2]
rlabel metal2 2714 55 2714 55 0 N1END[3]
rlabel metal2 6026 1602 6026 1602 0 N2END[0]
rlabel metal2 6394 1738 6394 1738 0 N2END[1]
rlabel metal2 6762 2350 6762 2350 0 N2END[2]
rlabel metal2 7130 276 7130 276 0 N2END[3]
rlabel metal2 7498 2316 7498 2316 0 N2END[4]
rlabel metal2 7866 2078 7866 2078 0 N2END[5]
rlabel metal2 8234 1279 8234 1279 0 N2END[6]
rlabel metal2 8602 2078 8602 2078 0 N2END[7]
rlabel metal2 3082 55 3082 55 0 N2MID[0]
rlabel metal2 3450 242 3450 242 0 N2MID[1]
rlabel metal2 3818 3914 3818 3914 0 N2MID[2]
rlabel metal2 4186 3778 4186 3778 0 N2MID[3]
rlabel metal2 4554 2350 4554 2350 0 N2MID[4]
rlabel metal2 4922 2282 4922 2282 0 N2MID[5]
rlabel metal2 5290 2316 5290 2316 0 N2MID[6]
rlabel metal2 5658 2282 5658 2282 0 N2MID[7]
rlabel metal2 8970 106 8970 106 0 N4END[0]
rlabel metal1 10580 5678 10580 5678 0 N4END[10]
rlabel metal2 13018 55 13018 55 0 N4END[11]
rlabel metal2 13386 344 13386 344 0 N4END[12]
rlabel metal2 10442 4998 10442 4998 0 N4END[13]
rlabel metal2 14122 55 14122 55 0 N4END[14]
rlabel metal2 14490 55 14490 55 0 N4END[15]
rlabel metal2 9338 123 9338 123 0 N4END[1]
rlabel metal2 9706 106 9706 106 0 N4END[2]
rlabel metal2 10074 140 10074 140 0 N4END[3]
rlabel metal2 10442 174 10442 174 0 N4END[4]
rlabel metal2 10810 208 10810 208 0 N4END[5]
rlabel metal2 11178 259 11178 259 0 N4END[6]
rlabel metal2 11546 939 11546 939 0 N4END[7]
rlabel metal2 11914 2554 11914 2554 0 N4END[8]
rlabel metal2 12282 2112 12282 2112 0 N4END[9]
rlabel metal2 12374 4964 12374 4964 0 NN4END[0]
rlabel metal2 18538 191 18538 191 0 NN4END[10]
rlabel metal2 18906 1401 18906 1401 0 NN4END[11]
rlabel metal2 19274 2316 19274 2316 0 NN4END[12]
rlabel metal2 19642 3183 19642 3183 0 NN4END[13]
rlabel metal2 20010 55 20010 55 0 NN4END[14]
rlabel metal2 20378 310 20378 310 0 NN4END[15]
rlabel metal2 15226 55 15226 55 0 NN4END[1]
rlabel metal1 15410 5134 15410 5134 0 NN4END[2]
rlabel metal1 15272 5678 15272 5678 0 NN4END[3]
rlabel metal2 16330 1401 16330 1401 0 NN4END[4]
rlabel metal1 16514 5202 16514 5202 0 NN4END[5]
rlabel metal2 17066 2622 17066 2622 0 NN4END[6]
rlabel metal1 17480 5202 17480 5202 0 NN4END[7]
rlabel via2 17802 55 17802 55 0 NN4END[8]
rlabel metal2 18170 55 18170 55 0 NN4END[9]
rlabel metal2 20746 1160 20746 1160 0 S1BEG[0]
rlabel metal2 21114 55 21114 55 0 S1BEG[1]
rlabel metal2 21482 1160 21482 1160 0 S1BEG[2]
rlabel metal2 21850 1432 21850 1432 0 S1BEG[3]
rlabel metal2 22218 1160 22218 1160 0 S2BEG[0]
rlabel metal2 22586 1160 22586 1160 0 S2BEG[1]
rlabel metal2 22954 1160 22954 1160 0 S2BEG[2]
rlabel metal2 23322 1160 23322 1160 0 S2BEG[3]
rlabel metal2 23690 1160 23690 1160 0 S2BEG[4]
rlabel metal2 24058 1160 24058 1160 0 S2BEG[5]
rlabel metal2 24426 1160 24426 1160 0 S2BEG[6]
rlabel metal2 24794 1143 24794 1143 0 S2BEG[7]
rlabel metal2 25162 1160 25162 1160 0 S2BEGb[0]
rlabel metal2 25530 1160 25530 1160 0 S2BEGb[1]
rlabel metal2 25898 1160 25898 1160 0 S2BEGb[2]
rlabel metal2 26266 1160 26266 1160 0 S2BEGb[3]
rlabel metal2 26634 1160 26634 1160 0 S2BEGb[4]
rlabel metal2 27002 55 27002 55 0 S2BEGb[5]
rlabel metal2 27370 123 27370 123 0 S2BEGb[6]
rlabel metal2 27738 1160 27738 1160 0 S2BEGb[7]
rlabel metal2 28106 55 28106 55 0 S4BEG[0]
rlabel metal2 31786 718 31786 718 0 S4BEG[10]
rlabel metal2 32154 55 32154 55 0 S4BEG[11]
rlabel metal2 32522 599 32522 599 0 S4BEG[12]
rlabel metal2 32890 1330 32890 1330 0 S4BEG[13]
rlabel metal2 33258 55 33258 55 0 S4BEG[14]
rlabel metal1 33764 2822 33764 2822 0 S4BEG[15]
rlabel metal2 28474 55 28474 55 0 S4BEG[1]
rlabel metal2 28842 1296 28842 1296 0 S4BEG[2]
rlabel metal1 29670 2822 29670 2822 0 S4BEG[3]
rlabel metal2 29578 1194 29578 1194 0 S4BEG[4]
rlabel metal2 29946 55 29946 55 0 S4BEG[5]
rlabel metal2 30314 1330 30314 1330 0 S4BEG[6]
rlabel metal2 30682 1296 30682 1296 0 S4BEG[7]
rlabel metal1 31188 2822 31188 2822 0 S4BEG[8]
rlabel metal1 32338 2312 32338 2312 0 S4BEG[9]
rlabel metal2 33994 55 33994 55 0 SS4BEG[0]
rlabel metal2 37674 1330 37674 1330 0 SS4BEG[10]
rlabel metal2 38042 599 38042 599 0 SS4BEG[11]
rlabel metal2 38410 1296 38410 1296 0 SS4BEG[12]
rlabel metal1 38916 2822 38916 2822 0 SS4BEG[13]
rlabel metal2 39146 55 39146 55 0 SS4BEG[14]
rlabel metal2 39514 1296 39514 1296 0 SS4BEG[15]
rlabel metal2 34362 1296 34362 1296 0 SS4BEG[1]
rlabel metal2 34730 55 34730 55 0 SS4BEG[2]
rlabel metal2 35098 599 35098 599 0 SS4BEG[3]
rlabel metal2 35466 599 35466 599 0 SS4BEG[4]
rlabel metal2 35834 1296 35834 1296 0 SS4BEG[5]
rlabel metal2 36202 735 36202 735 0 SS4BEG[6]
rlabel metal2 36570 55 36570 55 0 SS4BEG[7]
rlabel metal2 36938 1296 36938 1296 0 SS4BEG[8]
rlabel metal2 37306 718 37306 718 0 SS4BEG[9]
rlabel metal1 38962 7786 38962 7786 0 UserCLK
rlabel metal1 1472 8602 1472 8602 0 UserCLKo
rlabel via2 2438 4029 2438 4029 0 net1
rlabel metal1 19826 4114 19826 4114 0 net10
rlabel metal1 38134 7718 38134 7718 0 net100
rlabel metal1 36570 3060 36570 3060 0 net101
rlabel metal1 39146 2482 39146 2482 0 net102
rlabel metal1 37444 2482 37444 2482 0 net103
rlabel metal2 38042 1938 38042 1938 0 net104
rlabel metal1 1702 8432 1702 8432 0 net105
rlabel metal2 42734 5882 42734 5882 0 net11
rlabel metal1 31878 4760 31878 4760 0 net12
rlabel metal1 31740 5576 31740 5576 0 net13
rlabel metal2 36570 7616 36570 7616 0 net14
rlabel metal1 27094 6868 27094 6868 0 net15
rlabel metal2 36570 6528 36570 6528 0 net16
rlabel metal2 26542 8432 26542 8432 0 net17
rlabel metal2 23966 8466 23966 8466 0 net18
rlabel metal2 19550 8602 19550 8602 0 net19
rlabel metal1 47150 4046 47150 4046 0 net2
rlabel metal1 22172 8058 22172 8058 0 net20
rlabel metal2 11822 7684 11822 7684 0 net21
rlabel metal1 21827 7922 21827 7922 0 net22
rlabel metal1 38870 2006 38870 2006 0 net23
rlabel metal2 18998 6188 18998 6188 0 net24
rlabel metal1 46138 6970 46138 6970 0 net25
rlabel metal1 46506 2482 46506 2482 0 net26
rlabel metal2 41630 3842 41630 3842 0 net27
rlabel metal1 46736 3026 46736 3026 0 net28
rlabel metal1 47104 2414 47104 2414 0 net29
rlabel metal2 37398 5882 37398 5882 0 net3
rlabel metal1 46966 3536 46966 3536 0 net30
rlabel metal1 47012 3026 47012 3026 0 net31
rlabel metal2 36478 7208 36478 7208 0 net32
rlabel metal1 4094 8908 4094 8908 0 net33
rlabel metal1 40020 6630 40020 6630 0 net34
rlabel metal1 29624 8058 29624 8058 0 net35
rlabel metal1 41354 6664 41354 6664 0 net36
rlabel metal2 40434 7752 40434 7752 0 net37
rlabel metal2 37214 7310 37214 7310 0 net38
rlabel metal2 39606 7990 39606 7990 0 net39
rlabel metal2 40066 5576 40066 5576 0 net4
rlabel metal1 40848 7514 40848 7514 0 net40
rlabel metal1 43884 6630 43884 6630 0 net41
rlabel metal1 46000 6630 46000 6630 0 net42
rlabel metal1 46736 7514 46736 7514 0 net43
rlabel metal2 6670 8704 6670 8704 0 net44
rlabel metal1 8372 8058 8372 8058 0 net45
rlabel metal1 10488 8058 10488 8058 0 net46
rlabel metal2 13018 7990 13018 7990 0 net47
rlabel metal1 15226 7514 15226 7514 0 net48
rlabel metal2 17894 7990 17894 7990 0 net49
rlabel metal2 23322 7072 23322 7072 0 net5
rlabel metal2 20654 8262 20654 8262 0 net50
rlabel metal2 23506 8262 23506 8262 0 net51
rlabel metal1 25990 8058 25990 8058 0 net52
rlabel metal2 2806 4352 2806 4352 0 net53
rlabel metal1 20884 2414 20884 2414 0 net54
rlabel metal1 18998 2448 18998 2448 0 net55
rlabel metal1 21390 3026 21390 3026 0 net56
rlabel metal2 5566 2856 5566 2856 0 net57
rlabel metal1 5750 4488 5750 4488 0 net58
rlabel metal2 5750 2754 5750 2754 0 net59
rlabel metal2 14582 3417 14582 3417 0 net6
rlabel metal2 7774 3264 7774 3264 0 net60
rlabel metal2 20562 7786 20562 7786 0 net61
rlabel metal1 21114 7752 21114 7752 0 net62
rlabel metal1 21712 4454 21712 4454 0 net63
rlabel metal1 24840 2414 24840 2414 0 net64
rlabel metal1 8878 3978 8878 3978 0 net65
rlabel metal1 20746 2584 20746 2584 0 net66
rlabel metal2 7590 3400 7590 3400 0 net67
rlabel metal2 9614 3128 9614 3128 0 net68
rlabel metal1 26818 2414 26818 2414 0 net69
rlabel metal1 26174 3094 26174 3094 0 net7
rlabel metal1 27002 2482 27002 2482 0 net70
rlabel metal1 25070 2380 25070 2380 0 net71
rlabel metal1 28106 2448 28106 2448 0 net72
rlabel metal1 28520 2414 28520 2414 0 net73
rlabel metal1 32614 2414 32614 2414 0 net74
rlabel metal2 32798 2244 32798 2244 0 net75
rlabel metal1 33258 2448 33258 2448 0 net76
rlabel metal1 33580 2414 33580 2414 0 net77
rlabel metal2 33994 2992 33994 2992 0 net78
rlabel metal1 32890 3026 32890 3026 0 net79
rlabel metal1 26174 2924 26174 2924 0 net8
rlabel metal2 11362 3332 11362 3332 0 net80
rlabel metal2 10626 3672 10626 3672 0 net81
rlabel metal1 28290 3060 28290 3060 0 net82
rlabel metal2 10534 3502 10534 3502 0 net83
rlabel metal2 8694 6154 8694 6154 0 net84
rlabel metal2 8510 4318 8510 4318 0 net85
rlabel metal2 11454 3638 11454 3638 0 net86
rlabel metal2 29762 2975 29762 2975 0 net87
rlabel metal2 32154 2210 32154 2210 0 net88
rlabel metal1 33718 3434 33718 3434 0 net89
rlabel metal2 46598 5814 46598 5814 0 net9
rlabel metal1 17572 5066 17572 5066 0 net90
rlabel metal2 38502 1989 38502 1989 0 net91
rlabel metal2 38870 2057 38870 2057 0 net92
rlabel metal2 15410 4352 15410 4352 0 net93
rlabel via2 39238 2397 39238 2397 0 net94
rlabel metal2 40066 2465 40066 2465 0 net95
rlabel metal1 34224 3366 34224 3366 0 net96
rlabel metal1 34730 6086 34730 6086 0 net97
rlabel metal2 35650 1972 35650 1972 0 net98
rlabel metal1 35880 7718 35880 7718 0 net99
<< properties >>
string FIXED_BBOX 0 0 49000 11250
<< end >>
