module DSP (Tile_X0Y0_UserCLKo,
    Tile_X0Y1_UserCLK,
    Tile_X0Y0_E1BEG,
    Tile_X0Y0_E1END,
    Tile_X0Y0_E2BEG,
    Tile_X0Y0_E2BEGb,
    Tile_X0Y0_E2END,
    Tile_X0Y0_E2MID,
    Tile_X0Y0_E6BEG,
    Tile_X0Y0_E6END,
    Tile_X0Y0_EE4BEG,
    Tile_X0Y0_EE4END,
    Tile_X0Y0_FrameData,
    Tile_X0Y0_FrameData_O,
    Tile_X0Y0_FrameStrobe_O,
    Tile_X0Y0_N1BEG,
    Tile_X0Y0_N2BEG,
    Tile_X0Y0_N2BEGb,
    Tile_X0Y0_N4BEG,
    Tile_X0Y0_NN4BEG,
    Tile_X0Y0_S1END,
    Tile_X0Y0_S2END,
    Tile_X0Y0_S2MID,
    Tile_X0Y0_S4END,
    Tile_X0Y0_SS4END,
    Tile_X0Y0_W1BEG,
    Tile_X0Y0_W1END,
    Tile_X0Y0_W2BEG,
    Tile_X0Y0_W2BEGb,
    Tile_X0Y0_W2END,
    Tile_X0Y0_W2MID,
    Tile_X0Y0_W6BEG,
    Tile_X0Y0_W6END,
    Tile_X0Y0_WW4BEG,
    Tile_X0Y0_WW4END,
    Tile_X0Y1_E1BEG,
    Tile_X0Y1_E1END,
    Tile_X0Y1_E2BEG,
    Tile_X0Y1_E2BEGb,
    Tile_X0Y1_E2END,
    Tile_X0Y1_E2MID,
    Tile_X0Y1_E6BEG,
    Tile_X0Y1_E6END,
    Tile_X0Y1_EE4BEG,
    Tile_X0Y1_EE4END,
    Tile_X0Y1_FrameData,
    Tile_X0Y1_FrameData_O,
    Tile_X0Y1_FrameStrobe,
    Tile_X0Y1_N1END,
    Tile_X0Y1_N2END,
    Tile_X0Y1_N2MID,
    Tile_X0Y1_N4END,
    Tile_X0Y1_NN4END,
    Tile_X0Y1_S1BEG,
    Tile_X0Y1_S2BEG,
    Tile_X0Y1_S2BEGb,
    Tile_X0Y1_S4BEG,
    Tile_X0Y1_SS4BEG,
    Tile_X0Y1_W1BEG,
    Tile_X0Y1_W1END,
    Tile_X0Y1_W2BEG,
    Tile_X0Y1_W2BEGb,
    Tile_X0Y1_W2END,
    Tile_X0Y1_W2MID,
    Tile_X0Y1_W6BEG,
    Tile_X0Y1_W6END,
    Tile_X0Y1_WW4BEG,
    Tile_X0Y1_WW4END);
 output Tile_X0Y0_UserCLKo;
 input Tile_X0Y1_UserCLK;
 output [3:0] Tile_X0Y0_E1BEG;
 input [3:0] Tile_X0Y0_E1END;
 output [7:0] Tile_X0Y0_E2BEG;
 output [7:0] Tile_X0Y0_E2BEGb;
 input [7:0] Tile_X0Y0_E2END;
 input [7:0] Tile_X0Y0_E2MID;
 output [11:0] Tile_X0Y0_E6BEG;
 input [11:0] Tile_X0Y0_E6END;
 output [15:0] Tile_X0Y0_EE4BEG;
 input [15:0] Tile_X0Y0_EE4END;
 input [31:0] Tile_X0Y0_FrameData;
 output [31:0] Tile_X0Y0_FrameData_O;
 output [19:0] Tile_X0Y0_FrameStrobe_O;
 output [3:0] Tile_X0Y0_N1BEG;
 output [7:0] Tile_X0Y0_N2BEG;
 output [7:0] Tile_X0Y0_N2BEGb;
 output [15:0] Tile_X0Y0_N4BEG;
 output [15:0] Tile_X0Y0_NN4BEG;
 input [3:0] Tile_X0Y0_S1END;
 input [7:0] Tile_X0Y0_S2END;
 input [7:0] Tile_X0Y0_S2MID;
 input [15:0] Tile_X0Y0_S4END;
 input [15:0] Tile_X0Y0_SS4END;
 output [3:0] Tile_X0Y0_W1BEG;
 input [3:0] Tile_X0Y0_W1END;
 output [7:0] Tile_X0Y0_W2BEG;
 output [7:0] Tile_X0Y0_W2BEGb;
 input [7:0] Tile_X0Y0_W2END;
 input [7:0] Tile_X0Y0_W2MID;
 output [11:0] Tile_X0Y0_W6BEG;
 input [11:0] Tile_X0Y0_W6END;
 output [15:0] Tile_X0Y0_WW4BEG;
 input [15:0] Tile_X0Y0_WW4END;
 output [3:0] Tile_X0Y1_E1BEG;
 input [3:0] Tile_X0Y1_E1END;
 output [7:0] Tile_X0Y1_E2BEG;
 output [7:0] Tile_X0Y1_E2BEGb;
 input [7:0] Tile_X0Y1_E2END;
 input [7:0] Tile_X0Y1_E2MID;
 output [11:0] Tile_X0Y1_E6BEG;
 input [11:0] Tile_X0Y1_E6END;
 output [15:0] Tile_X0Y1_EE4BEG;
 input [15:0] Tile_X0Y1_EE4END;
 input [31:0] Tile_X0Y1_FrameData;
 output [31:0] Tile_X0Y1_FrameData_O;
 input [19:0] Tile_X0Y1_FrameStrobe;
 input [3:0] Tile_X0Y1_N1END;
 input [7:0] Tile_X0Y1_N2END;
 input [7:0] Tile_X0Y1_N2MID;
 input [15:0] Tile_X0Y1_N4END;
 input [15:0] Tile_X0Y1_NN4END;
 output [3:0] Tile_X0Y1_S1BEG;
 output [7:0] Tile_X0Y1_S2BEG;
 output [7:0] Tile_X0Y1_S2BEGb;
 output [15:0] Tile_X0Y1_S4BEG;
 output [15:0] Tile_X0Y1_SS4BEG;
 output [3:0] Tile_X0Y1_W1BEG;
 input [3:0] Tile_X0Y1_W1END;
 output [7:0] Tile_X0Y1_W2BEG;
 output [7:0] Tile_X0Y1_W2BEGb;
 input [7:0] Tile_X0Y1_W2END;
 input [7:0] Tile_X0Y1_W2MID;
 output [11:0] Tile_X0Y1_W6BEG;
 input [11:0] Tile_X0Y1_W6END;
 output [15:0] Tile_X0Y1_WW4BEG;
 input [15:0] Tile_X0Y1_WW4END;

 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X ;
 wire \Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A ;
 wire \Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A ;
 wire \Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A ;
 wire \Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A ;
 wire \Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A ;
 wire \Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A ;
 wire \Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A ;
 wire \Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A ;
 wire net236;
 wire net237;
 wire net914;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net919;
 wire net874;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net928;
 wire net377;
 wire net866;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net946;
 wire net426;
 wire net827;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire \Tile_X0Y1_DSP_bot.A0 ;
 wire \Tile_X0Y1_DSP_bot.A1 ;
 wire \Tile_X0Y1_DSP_bot.A2 ;
 wire \Tile_X0Y1_DSP_bot.A3 ;
 wire \Tile_X0Y1_DSP_bot.B0 ;
 wire \Tile_X0Y1_DSP_bot.B1 ;
 wire \Tile_X0Y1_DSP_bot.B2 ;
 wire \Tile_X0Y1_DSP_bot.B3 ;
 wire \Tile_X0Y1_DSP_bot.C0 ;
 wire \Tile_X0Y1_DSP_bot.C1 ;
 wire \Tile_X0Y1_DSP_bot.C2 ;
 wire \Tile_X0Y1_DSP_bot.C3 ;
 wire \Tile_X0Y1_DSP_bot.C4 ;
 wire \Tile_X0Y1_DSP_bot.C5 ;
 wire \Tile_X0Y1_DSP_bot.C6 ;
 wire \Tile_X0Y1_DSP_bot.C7 ;
 wire \Tile_X0Y1_DSP_bot.C8 ;
 wire \Tile_X0Y1_DSP_bot.C9 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[0] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[10] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[11] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[12] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[13] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[14] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[15] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[16] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[17] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[18] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[19] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[1] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[2] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[3] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[4] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[5] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[6] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[7] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[8] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[9] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[0] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[1] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[2] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[3] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[4] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[5] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[6] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[7] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[0] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[1] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[2] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[3] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[4] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[5] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[6] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[7] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[0] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[10] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[11] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[12] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[13] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[14] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[15] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[16] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[17] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[18] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[19] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[1] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[2] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[3] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[4] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[5] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[6] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[7] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[8] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[9] ;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net875;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net660;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net651;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net911;
 wire net605;
 wire net606;
 wire net653;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net617;
 wire Tile_X0Y1_UserCLK_regs;
 wire clknet_0_Tile_X0Y1_UserCLK;
 wire clknet_1_0__leaf_Tile_X0Y1_UserCLK;
 wire clknet_0_Tile_X0Y1_UserCLK_regs;
 wire clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs;
 wire clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs;
 wire clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs;
 wire clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net652;
 wire net654;
 wire net655;
 wire net656;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net676;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net867;
 wire net868;
 wire net869;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net912;
 wire net913;
 wire net915;
 wire net918;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;

 sky130_fd_sc_hd__a21o_1 _2036_ (.A1(_0908_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q ),
    .B1(_0911_),
    .X(_0912_));
 sky130_fd_sc_hd__mux4_1 _2037_ (.A0(net1020),
    .A1(net1036),
    .A2(net1032),
    .A3(net983),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_0913_));
 sky130_fd_sc_hd__and2_1 _2038_ (.A(_0118_),
    .B(_0913_),
    .X(_0914_));
 sky130_fd_sc_hd__mux4_1 _2039_ (.A0(net1044),
    .A1(net1029),
    .A2(net1054),
    .A3(net1056),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_0915_));
 sky130_fd_sc_hd__a21bo_1 _2040_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ),
    .A2(_0915_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q ),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_4 _2041_ (.A0(_0414_),
    .A1(net193),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_0917_));
 sky130_fd_sc_hd__mux2_1 _2042_ (.A0(net1263),
    .A1(net12),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_0918_));
 sky130_fd_sc_hd__or2_1 _2043_ (.A(_0117_),
    .B(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__o211a_1 _2044_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .A2(_0917_),
    .B1(_0919_),
    .C1(_0118_),
    .X(_0920_));
 sky130_fd_sc_hd__mux2_1 _2045_ (.A0(net60),
    .A1(net68),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_0921_));
 sky130_fd_sc_hd__or2_1 _2046_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .B(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__mux2_1 _2047_ (.A0(net94),
    .A1(net1225),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_0923_));
 sky130_fd_sc_hd__o211a_1 _2048_ (.A1(_0117_),
    .A2(_0923_),
    .B1(_0922_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_0924_));
 sky130_fd_sc_hd__o32a_4 _2049_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q ),
    .A2(_0924_),
    .A3(_0920_),
    .B1(_0914_),
    .B2(_0916_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ));
 sky130_fd_sc_hd__mux4_2 _2050_ (.A0(net192),
    .A1(net228),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q ),
    .X(_0925_));
 sky130_fd_sc_hd__o21a_1 _2051_ (.A1(_0925_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ),
    .B1(_0912_),
    .X(_0926_));
 sky130_fd_sc_hd__mux2_4 _2052_ (.A0(_0926_),
    .A1(_0907_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q ),
    .X(\Tile_X0Y1_DSP_bot.A0 ));
 sky130_fd_sc_hd__nand2b_1 _2053_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[0] ),
    .B(net1059),
    .Y(_0927_));
 sky130_fd_sc_hd__o21ai_4 _2054_ (.A1(\Tile_X0Y1_DSP_bot.A0 ),
    .A2(net1059),
    .B1(_0927_),
    .Y(_0928_));
 sky130_fd_sc_hd__nor2_1 _2055_ (.A(net620),
    .B(_0667_),
    .Y(_0929_));
 sky130_fd_sc_hd__nand4b_1 _2056_ (.A_N(net620),
    .B(_0709_),
    .C(_0708_),
    .D(_0849_),
    .Y(_0930_));
 sky130_fd_sc_hd__nor2_1 _2057_ (.A(_0726_),
    .B(_0762_),
    .Y(_0931_));
 sky130_fd_sc_hd__a31o_1 _2058_ (.A1(_0708_),
    .A2(_0709_),
    .A3(_0847_),
    .B1(_0929_),
    .X(_0932_));
 sky130_fd_sc_hd__nand3_2 _2059_ (.A(_0930_),
    .B(_0931_),
    .C(_0932_),
    .Y(_0933_));
 sky130_fd_sc_hd__nand2_2 _2060_ (.A(_0930_),
    .B(_0933_),
    .Y(_0934_));
 sky130_fd_sc_hd__xnor2_1 _2061_ (.A(_0850_),
    .B(_0851_),
    .Y(_0935_));
 sky130_fd_sc_hd__and2b_1 _2062_ (.A_N(_0935_),
    .B(_0934_),
    .X(_0936_));
 sky130_fd_sc_hd__xor2_1 _2063_ (.A(_0934_),
    .B(_0935_),
    .X(_0937_));
 sky130_fd_sc_hd__or2_1 _2064_ (.A(net618),
    .B(_0878_),
    .X(_0938_));
 sky130_fd_sc_hd__nor2_4 _2065_ (.A(_0784_),
    .B(_0478_),
    .Y(_0939_));
 sky130_fd_sc_hd__and4_1 _2066_ (.A(_0611_),
    .B(_0612_),
    .C(_0782_),
    .D(_0783_),
    .X(_0940_));
 sky130_fd_sc_hd__xnor2_4 _2067_ (.A(_0939_),
    .B(_0881_),
    .Y(_0941_));
 sky130_fd_sc_hd__xnor2_4 _2068_ (.A(_0941_),
    .B(_0938_),
    .Y(_0942_));
 sky130_fd_sc_hd__nor2_4 _2069_ (.A(_0937_),
    .B(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__xor2_1 _2070_ (.A(_0855_),
    .B(_0883_),
    .X(_0944_));
 sky130_fd_sc_hd__o21ai_4 _2071_ (.A1(_0936_),
    .A2(_0943_),
    .B1(_0944_),
    .Y(_0945_));
 sky130_fd_sc_hd__o2bb2ai_1 _2072_ (.A1_N(_0881_),
    .A2_N(_0939_),
    .B1(_0941_),
    .B2(_0938_),
    .Y(_0946_));
 sky130_fd_sc_hd__or3_1 _2073_ (.A(_0936_),
    .B(_0943_),
    .C(_0944_),
    .X(_0947_));
 sky130_fd_sc_hd__nand2_2 _2074_ (.A(_0945_),
    .B(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__nand2b_2 _2075_ (.A_N(_0948_),
    .B(_0946_),
    .Y(_0949_));
 sky130_fd_sc_hd__xnor2_1 _2076_ (.A(_0887_),
    .B(_0888_),
    .Y(_0950_));
 sky130_fd_sc_hd__a21oi_4 _2077_ (.A1(_0949_),
    .A2(_0945_),
    .B1(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__xor2_1 _2078_ (.A(_0822_),
    .B(_0889_),
    .X(_0952_));
 sky130_fd_sc_hd__xnor2_2 _2079_ (.A(_0952_),
    .B(_0951_),
    .Y(_0953_));
 sky130_fd_sc_hd__inv_2 _2080_ (.A(_0953_),
    .Y(_0954_));
 sky130_fd_sc_hd__and3_1 _2081_ (.A(_0611_),
    .B(_0612_),
    .C(_0641_),
    .X(_0955_));
 sky130_fd_sc_hd__nor2_1 _2082_ (.A(_0478_),
    .B(_0640_),
    .Y(_0956_));
 sky130_fd_sc_hd__nor2_1 _2083_ (.A(_0799_),
    .B(_0878_),
    .Y(_0957_));
 sky130_fd_sc_hd__xor2_2 _2084_ (.A(_0940_),
    .B(_0956_),
    .X(_0958_));
 sky130_fd_sc_hd__a22o_1 _2085_ (.A1(_0940_),
    .A2(_0956_),
    .B1(_0957_),
    .B2(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__mux4_2 _2086_ (.A0(net180),
    .A1(net125),
    .A2(net71),
    .A3(net234),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q ),
    .X(_0960_));
 sky130_fd_sc_hd__mux2_1 _2087_ (.A0(_0960_),
    .A1(_0228_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ),
    .X(_0961_));
 sky130_fd_sc_hd__a211o_1 _2088_ (.A1(_0360_),
    .A2(_0361_),
    .B1(_0142_),
    .C1(_0386_),
    .X(_0962_));
 sky130_fd_sc_hd__a211o_1 _2089_ (.A1(_0561_),
    .A2(_0562_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .C1(_0556_),
    .X(_0963_));
 sky130_fd_sc_hd__mux2_1 _2090_ (.A0(net74),
    .A1(net211),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0964_));
 sky130_fd_sc_hd__a21o_1 _2091_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .A2(_0964_),
    .B1(_0144_),
    .X(_0965_));
 sky130_fd_sc_hd__a31o_1 _2092_ (.A1(_0143_),
    .A2(_0962_),
    .A3(_0963_),
    .B1(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__mux4_1 _2093_ (.A0(net175),
    .A1(net183),
    .A2(net120),
    .A3(net128),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0967_));
 sky130_fd_sc_hd__o21ba_1 _2094_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .A2(_0967_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_0968_));
 sky130_fd_sc_hd__mux4_2 _2095_ (.A0(net995),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .A2(net1005),
    .A3(net653),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0969_));
 sky130_fd_sc_hd__mux4_1 _2096_ (.A0(net655),
    .A1(net971),
    .A2(net981),
    .A3(net1000),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0970_));
 sky130_fd_sc_hd__or2_1 _2097_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .B(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__o211a_1 _2098_ (.A1(_0969_),
    .A2(_0144_),
    .B1(_0971_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_0972_));
 sky130_fd_sc_hd__a21o_1 _2099_ (.A1(_0968_),
    .A2(_0966_),
    .B1(_0972_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ));
 sky130_fd_sc_hd__a211o_1 _2100_ (.A1(_0966_),
    .A2(_0968_),
    .B1(_0141_),
    .C1(_0972_),
    .X(_0973_));
 sky130_fd_sc_hd__o21a_1 _2101_ (.A1(net224),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q ),
    .X(_0974_));
 sky130_fd_sc_hd__mux2_1 _2102_ (.A0(net188),
    .A1(net133),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .X(_0975_));
 sky130_fd_sc_hd__a221o_1 _2103_ (.A1(_0974_),
    .A2(_0973_),
    .B1(_0975_),
    .B2(_0145_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ),
    .X(_0976_));
 sky130_fd_sc_hd__mux4_2 _2104_ (.A0(net189),
    .A1(net134),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .A3(net225),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q ),
    .X(_0977_));
 sky130_fd_sc_hd__inv_2 _2105_ (.A(_0977_),
    .Y(_0978_));
 sky130_fd_sc_hd__a21oi_2 _2106_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ),
    .A2(_0978_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q ),
    .Y(_0979_));
 sky130_fd_sc_hd__a22o_4 _2107_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q ),
    .A2(_0961_),
    .B1(_0979_),
    .B2(_0976_),
    .X(\Tile_X0Y1_DSP_bot.B1 ));
 sky130_fd_sc_hd__nand2b_1 _2108_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[1] ),
    .B(net1061),
    .Y(_0980_));
 sky130_fd_sc_hd__o21ai_4 _2109_ (.A1(\Tile_X0Y1_DSP_bot.B1 ),
    .A2(net1061),
    .B1(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__nor2_2 _2110_ (.A(_0521_),
    .B(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__nand2_4 _2111_ (.A(_0959_),
    .B(_0982_),
    .Y(_0983_));
 sky130_fd_sc_hd__or2_1 _2112_ (.A(net622),
    .B(net620),
    .X(_0984_));
 sky130_fd_sc_hd__nor3_1 _2113_ (.A(_0710_),
    .B(_0848_),
    .C(_0984_),
    .Y(_0985_));
 sky130_fd_sc_hd__a21o_1 _2114_ (.A1(_0930_),
    .A2(_0932_),
    .B1(_0931_),
    .X(_0986_));
 sky130_fd_sc_hd__nand3_2 _2115_ (.A(_0933_),
    .B(_0985_),
    .C(_0986_),
    .Y(_0987_));
 sky130_fd_sc_hd__a21o_1 _2116_ (.A1(_0933_),
    .A2(_0986_),
    .B1(_0985_),
    .X(_0988_));
 sky130_fd_sc_hd__xor2_1 _2117_ (.A(_0957_),
    .B(_0958_),
    .X(_0989_));
 sky130_fd_sc_hd__nand3_2 _2118_ (.A(_0987_),
    .B(_0988_),
    .C(_0989_),
    .Y(_0990_));
 sky130_fd_sc_hd__nand2_1 _2119_ (.A(_0987_),
    .B(_0990_),
    .Y(_0991_));
 sky130_fd_sc_hd__xor2_2 _2120_ (.A(_0937_),
    .B(_0942_),
    .X(_0992_));
 sky130_fd_sc_hd__nand2_1 _2121_ (.A(_0991_),
    .B(_0992_),
    .Y(_0993_));
 sky130_fd_sc_hd__xnor2_1 _2122_ (.A(_0991_),
    .B(_0992_),
    .Y(_0994_));
 sky130_fd_sc_hd__xnor2_1 _2123_ (.A(_0959_),
    .B(_0982_),
    .Y(_0995_));
 sky130_fd_sc_hd__o21ai_2 _2124_ (.A1(_0994_),
    .A2(_0995_),
    .B1(_0993_),
    .Y(_0996_));
 sky130_fd_sc_hd__xnor2_1 _2125_ (.A(_0946_),
    .B(_0948_),
    .Y(_0997_));
 sky130_fd_sc_hd__and2_1 _2126_ (.A(_0996_),
    .B(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__xnor2_2 _2127_ (.A(_0996_),
    .B(_0997_),
    .Y(_0999_));
 sky130_fd_sc_hd__nor2_1 _2128_ (.A(_0983_),
    .B(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__xor2_4 _2129_ (.A(_0999_),
    .B(_0983_),
    .X(_1001_));
 sky130_fd_sc_hd__o22a_1 _2130_ (.A1(net622),
    .A2(_0848_),
    .B1(net620),
    .B2(_0710_),
    .X(_1002_));
 sky130_fd_sc_hd__or2_1 _2131_ (.A(_0985_),
    .B(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__nor2_1 _2132_ (.A(_0784_),
    .B(_0878_),
    .Y(_1004_));
 sky130_fd_sc_hd__nor2_4 _2133_ (.A(_0726_),
    .B(_0478_),
    .Y(_1005_));
 sky130_fd_sc_hd__xor2_2 _2134_ (.A(_0955_),
    .B(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__xnor2_2 _2135_ (.A(_1006_),
    .B(_1004_),
    .Y(_1007_));
 sky130_fd_sc_hd__nor2_1 _2136_ (.A(_1003_),
    .B(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__a21o_1 _2137_ (.A1(_0987_),
    .A2(_0988_),
    .B1(_0989_),
    .X(_1009_));
 sky130_fd_sc_hd__nand3_2 _2138_ (.A(_0990_),
    .B(_1008_),
    .C(_1009_),
    .Y(_1010_));
 sky130_fd_sc_hd__a21o_1 _2139_ (.A1(_0990_),
    .A2(_1009_),
    .B1(_1008_),
    .X(_1011_));
 sky130_fd_sc_hd__or2_1 _2140_ (.A(net618),
    .B(_0981_),
    .X(_1012_));
 sky130_fd_sc_hd__a22o_1 _2141_ (.A1(_0955_),
    .A2(_1005_),
    .B1(_1006_),
    .B2(_1004_),
    .X(_1013_));
 sky130_fd_sc_hd__mux2_1 _2142_ (.A0(net234),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q ),
    .X(_1014_));
 sky130_fd_sc_hd__mux2_1 _2143_ (.A0(net126),
    .A1(net92),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q ),
    .X(_1015_));
 sky130_fd_sc_hd__inv_1 _2144_ (.A(_1015_),
    .Y(_1016_));
 sky130_fd_sc_hd__o21ai_1 _2145_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q ),
    .A2(_1016_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .Y(_1017_));
 sky130_fd_sc_hd__a21o_1 _2146_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q ),
    .A2(_1014_),
    .B1(_1017_),
    .X(_1018_));
 sky130_fd_sc_hd__mux4_2 _2147_ (.A0(net205),
    .A1(net129),
    .A2(net75),
    .A3(net220),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q ),
    .X(_1019_));
 sky130_fd_sc_hd__or2_1 _2148_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .B(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__a211o_1 _2149_ (.A1(_0569_),
    .A2(_0567_),
    .B1(_0146_),
    .C1(_0541_),
    .X(_1021_));
 sky130_fd_sc_hd__o21a_1 _2150_ (.A1(net228),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .X(_1022_));
 sky130_fd_sc_hd__mux2_1 _2151_ (.A0(net137),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .X(_1023_));
 sky130_fd_sc_hd__a221o_1 _2152_ (.A1(_1022_),
    .A2(_1021_),
    .B1(_1023_),
    .B2(_0147_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .X(_1024_));
 sky130_fd_sc_hd__mux4_2 _2153_ (.A0(net193),
    .A1(net138),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ),
    .A3(net229),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q ),
    .X(_1025_));
 sky130_fd_sc_hd__inv_2 _2154_ (.A(_1025_),
    .Y(_1026_));
 sky130_fd_sc_hd__a21oi_2 _2155_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_1026_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q ),
    .Y(_1027_));
 sky130_fd_sc_hd__a32o_2 _2156_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q ),
    .A2(_1018_),
    .A3(_1020_),
    .B1(_1024_),
    .B2(_1027_),
    .X(\Tile_X0Y1_DSP_bot.B0 ));
 sky130_fd_sc_hd__nand2b_1 _2157_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[0] ),
    .B(net1061),
    .Y(_1028_));
 sky130_fd_sc_hd__o21ai_4 _2158_ (.A1(\Tile_X0Y1_DSP_bot.B0 ),
    .A2(net1061),
    .B1(_1028_),
    .Y(_1029_));
 sky130_fd_sc_hd__nor2_2 _2159_ (.A(_0521_),
    .B(net832),
    .Y(_1030_));
 sky130_fd_sc_hd__xnor2_1 _2160_ (.A(_1013_),
    .B(_1030_),
    .Y(_1031_));
 sky130_fd_sc_hd__xor2_1 _2161_ (.A(_1012_),
    .B(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__and3_4 _2162_ (.A(_1032_),
    .B(_1011_),
    .C(_1010_),
    .X(_1033_));
 sky130_fd_sc_hd__a31o_1 _2163_ (.A1(_0990_),
    .A2(_1008_),
    .A3(_1009_),
    .B1(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__xor2_1 _2164_ (.A(_0994_),
    .B(_0995_),
    .X(_1035_));
 sky130_fd_sc_hd__and2_1 _2165_ (.A(_1034_),
    .B(_1035_),
    .X(_1036_));
 sky130_fd_sc_hd__a2bb2o_1 _2166_ (.A1_N(_1012_),
    .A2_N(_1031_),
    .B1(_1030_),
    .B2(_1013_),
    .X(_1037_));
 sky130_fd_sc_hd__xor2_1 _2167_ (.A(_1034_),
    .B(_1035_),
    .X(_1038_));
 sky130_fd_sc_hd__a21oi_4 _2168_ (.A1(_1037_),
    .A2(_1038_),
    .B1(_1036_),
    .Y(_1039_));
 sky130_fd_sc_hd__and2b_1 _2169_ (.A_N(_1039_),
    .B(_1001_),
    .X(_1040_));
 sky130_fd_sc_hd__xnor2_4 _2170_ (.A(_1001_),
    .B(_1039_),
    .Y(_1041_));
 sky130_fd_sc_hd__xor2_1 _2171_ (.A(_1037_),
    .B(_1038_),
    .X(_1042_));
 sky130_fd_sc_hd__xor2_2 _2172_ (.A(_1007_),
    .B(_1003_),
    .X(_1043_));
 sky130_fd_sc_hd__nor2_8 _2173_ (.A(_0878_),
    .B(_0640_),
    .Y(_1044_));
 sky130_fd_sc_hd__nor2_1 _2174_ (.A(_0478_),
    .B(_0848_),
    .Y(_1045_));
 sky130_fd_sc_hd__a31o_1 _2175_ (.A1(_0725_),
    .A2(_0612_),
    .A3(_0611_),
    .B1(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__and3_4 _2176_ (.A(_0611_),
    .B(_0847_),
    .C(_0612_),
    .X(_1047_));
 sky130_fd_sc_hd__a21bo_4 _2177_ (.A1(_1047_),
    .A2(_1005_),
    .B1_N(_1046_),
    .X(_1048_));
 sky130_fd_sc_hd__xor2_4 _2178_ (.A(_1044_),
    .B(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__nor2_4 _2179_ (.A(_0984_),
    .B(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__nand2_4 _2180_ (.A(_1043_),
    .B(_1050_),
    .Y(_1051_));
 sky130_fd_sc_hd__xnor2_2 _2181_ (.A(_1043_),
    .B(_1050_),
    .Y(_1052_));
 sky130_fd_sc_hd__or2_4 _2182_ (.A(_0799_),
    .B(_0981_),
    .X(_1053_));
 sky130_fd_sc_hd__a22o_4 _2183_ (.A1(_1044_),
    .A2(_1046_),
    .B1(_1005_),
    .B2(_1047_),
    .X(_1054_));
 sky130_fd_sc_hd__nor2_1 _2184_ (.A(net618),
    .B(net832),
    .Y(_1055_));
 sky130_fd_sc_hd__nand2_1 _2185_ (.A(_1054_),
    .B(_1055_),
    .Y(_1056_));
 sky130_fd_sc_hd__xnor2_4 _2186_ (.A(_1055_),
    .B(_1054_),
    .Y(_1057_));
 sky130_fd_sc_hd__or2_4 _2187_ (.A(_1053_),
    .B(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__xnor2_2 _2188_ (.A(_1057_),
    .B(_1053_),
    .Y(_1059_));
 sky130_fd_sc_hd__or2_1 _2189_ (.A(_1052_),
    .B(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__a21oi_2 _2190_ (.A1(_1010_),
    .A2(_1011_),
    .B1(_1032_),
    .Y(_1061_));
 sky130_fd_sc_hd__a211oi_4 _2191_ (.A1(_1051_),
    .A2(_1060_),
    .B1(_1033_),
    .C1(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__o211a_1 _2192_ (.A1(_1033_),
    .A2(_1061_),
    .B1(_1060_),
    .C1(_1051_),
    .X(_1063_));
 sky130_fd_sc_hd__a211o_4 _2193_ (.A1(_1056_),
    .A2(_1058_),
    .B1(_1063_),
    .C1(_1062_),
    .X(_1064_));
 sky130_fd_sc_hd__and2b_1 _2194_ (.A_N(_1062_),
    .B(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__and2b_1 _2195_ (.A_N(_1065_),
    .B(_1042_),
    .X(_1066_));
 sky130_fd_sc_hd__xnor2_1 _2196_ (.A(_1042_),
    .B(_1065_),
    .Y(_1067_));
 sky130_fd_sc_hd__o211ai_2 _2197_ (.A1(_1063_),
    .A2(_1062_),
    .B1(_1056_),
    .C1(_1058_),
    .Y(_1068_));
 sky130_fd_sc_hd__xor2_2 _2198_ (.A(_1052_),
    .B(_1059_),
    .X(_1069_));
 sky130_fd_sc_hd__xnor2_2 _2199_ (.A(_0984_),
    .B(_1049_),
    .Y(_1070_));
 sky130_fd_sc_hd__nor2_8 _2200_ (.A(_0981_),
    .B(_0784_),
    .Y(_1071_));
 sky130_fd_sc_hd__and3b_1 _2201_ (.A_N(net620),
    .B(_0612_),
    .C(_0611_),
    .X(_1072_));
 sky130_fd_sc_hd__nor2_1 _2202_ (.A(_0478_),
    .B(_0928_),
    .Y(_1073_));
 sky130_fd_sc_hd__o211a_4 _2203_ (.A1(net1061),
    .A2(\Tile_X0Y1_DSP_bot.B2 ),
    .B1(_0877_),
    .C1(_0725_),
    .X(_1074_));
 sky130_fd_sc_hd__a31o_1 _2204_ (.A1(_0611_),
    .A2(_0612_),
    .A3(_0847_),
    .B1(_1073_),
    .X(_1075_));
 sky130_fd_sc_hd__a21boi_2 _2205_ (.A1(_1045_),
    .A2(_1072_),
    .B1_N(_1075_),
    .Y(_1076_));
 sky130_fd_sc_hd__a22o_1 _2206_ (.A1(_1045_),
    .A2(_1072_),
    .B1(_1074_),
    .B2(_1075_),
    .X(_1077_));
 sky130_fd_sc_hd__nor2_1 _2207_ (.A(_0799_),
    .B(net832),
    .Y(_1078_));
 sky130_fd_sc_hd__xor2_1 _2208_ (.A(_1077_),
    .B(_1078_),
    .X(_1079_));
 sky130_fd_sc_hd__xor2_2 _2209_ (.A(_1071_),
    .B(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__and2b_1 _2210_ (.A_N(_1070_),
    .B(_1080_),
    .X(_1081_));
 sky130_fd_sc_hd__and2_1 _2211_ (.A(_1069_),
    .B(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__a22oi_2 _2212_ (.A1(_1077_),
    .A2(_1078_),
    .B1(_1079_),
    .B2(_1071_),
    .Y(_1083_));
 sky130_fd_sc_hd__xnor2_2 _2213_ (.A(_1069_),
    .B(_1081_),
    .Y(_1084_));
 sky130_fd_sc_hd__nor2_1 _2214_ (.A(_1083_),
    .B(_1084_),
    .Y(_1085_));
 sky130_fd_sc_hd__a211oi_4 _2215_ (.A1(_1068_),
    .A2(_1064_),
    .B1(_1082_),
    .C1(_1085_),
    .Y(_1086_));
 sky130_fd_sc_hd__inv_2 _2216_ (.A(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__o211a_1 _2217_ (.A1(_1082_),
    .A2(_1085_),
    .B1(_1068_),
    .C1(_1064_),
    .X(_1088_));
 sky130_fd_sc_hd__xnor2_2 _2218_ (.A(_1083_),
    .B(_1084_),
    .Y(_1089_));
 sky130_fd_sc_hd__xnor2_2 _2219_ (.A(_1080_),
    .B(_1070_),
    .Y(_1090_));
 sky130_fd_sc_hd__xnor2_4 _2220_ (.A(_1074_),
    .B(_1076_),
    .Y(_1091_));
 sky130_fd_sc_hd__nor2_8 _2221_ (.A(_0640_),
    .B(_0981_),
    .Y(_1092_));
 sky130_fd_sc_hd__nor2_4 _2222_ (.A(_0878_),
    .B(_0928_),
    .Y(_1093_));
 sky130_fd_sc_hd__or3b_4 _2223_ (.A(_0878_),
    .B(_0928_),
    .C_N(_1047_),
    .X(_1094_));
 sky130_fd_sc_hd__nor2_8 _2224_ (.A(_0784_),
    .B(net832),
    .Y(_1095_));
 sky130_fd_sc_hd__xnor2_4 _2225_ (.A(_1095_),
    .B(_1094_),
    .Y(_1096_));
 sky130_fd_sc_hd__and2_1 _2226_ (.A(_1092_),
    .B(_1096_),
    .X(_1097_));
 sky130_fd_sc_hd__xnor2_4 _2227_ (.A(_1096_),
    .B(_1092_),
    .Y(_1098_));
 sky130_fd_sc_hd__nor2_4 _2228_ (.A(_1091_),
    .B(_1098_),
    .Y(_1099_));
 sky130_fd_sc_hd__a31o_1 _2229_ (.A1(_1047_),
    .A2(_1093_),
    .A3(_1095_),
    .B1(_1097_),
    .X(_1100_));
 sky130_fd_sc_hd__xnor2_2 _2230_ (.A(_1099_),
    .B(_1090_),
    .Y(_1101_));
 sky130_fd_sc_hd__nand2b_1 _2231_ (.A_N(_1101_),
    .B(_1100_),
    .Y(_1102_));
 sky130_fd_sc_hd__a21bo_1 _2232_ (.A1(_1090_),
    .A2(_1099_),
    .B1_N(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__and2b_1 _2233_ (.A_N(_1089_),
    .B(_1103_),
    .X(_1104_));
 sky130_fd_sc_hd__xnor2_2 _2234_ (.A(_1103_),
    .B(_1089_),
    .Y(_1105_));
 sky130_fd_sc_hd__xnor2_2 _2235_ (.A(_1101_),
    .B(_1100_),
    .Y(_1106_));
 sky130_fd_sc_hd__xor2_2 _2236_ (.A(_1091_),
    .B(_1098_),
    .X(_1107_));
 sky130_fd_sc_hd__o21bai_1 _2237_ (.A1(_0848_),
    .A2(_0878_),
    .B1_N(_1072_),
    .Y(_1108_));
 sky130_fd_sc_hd__nand2_1 _2238_ (.A(_1094_),
    .B(_1108_),
    .Y(_1109_));
 sky130_fd_sc_hd__nor2_4 _2239_ (.A(net832),
    .B(_0726_),
    .Y(_1110_));
 sky130_fd_sc_hd__and2_1 _2240_ (.A(_1092_),
    .B(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__o22a_1 _2241_ (.A1(_0726_),
    .A2(_0981_),
    .B1(net832),
    .B2(_0640_),
    .X(_1112_));
 sky130_fd_sc_hd__a21o_1 _2242_ (.A1(_1092_),
    .A2(_1110_),
    .B1(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__nor2_1 _2243_ (.A(_1109_),
    .B(_1113_),
    .Y(_1114_));
 sky130_fd_sc_hd__xor2_2 _2244_ (.A(_1107_),
    .B(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__o21ai_2 _2245_ (.A1(_1111_),
    .A2(_1114_),
    .B1(_1107_),
    .Y(_1116_));
 sky130_fd_sc_hd__and2b_1 _2246_ (.A_N(_1116_),
    .B(_1106_),
    .X(_1117_));
 sky130_fd_sc_hd__xnor2_4 _2247_ (.A(_1116_),
    .B(_1106_),
    .Y(_1118_));
 sky130_fd_sc_hd__xnor2_2 _2248_ (.A(_1115_),
    .B(_1111_),
    .Y(_1119_));
 sky130_fd_sc_hd__xor2_2 _2249_ (.A(_1113_),
    .B(_1109_),
    .X(_1120_));
 sky130_fd_sc_hd__nor2_2 _2250_ (.A(_0848_),
    .B(_0981_),
    .Y(_1121_));
 sky130_fd_sc_hd__xor2_1 _2251_ (.A(_1110_),
    .B(_1121_),
    .X(_1122_));
 sky130_fd_sc_hd__a22oi_2 _2252_ (.A1(_1110_),
    .A2(_1121_),
    .B1(_1122_),
    .B2(_1093_),
    .Y(_1123_));
 sky130_fd_sc_hd__and2b_1 _2253_ (.A_N(_1123_),
    .B(_1120_),
    .X(_1124_));
 sky130_fd_sc_hd__nor2_8 _2254_ (.A(_0928_),
    .B(net832),
    .Y(_1125_));
 sky130_fd_sc_hd__nand2_4 _2255_ (.A(_1121_),
    .B(net829),
    .Y(_1126_));
 sky130_fd_sc_hd__xor2_2 _2256_ (.A(_1093_),
    .B(_1122_),
    .X(_1127_));
 sky130_fd_sc_hd__and3_1 _2257_ (.A(_1121_),
    .B(_1125_),
    .C(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__xnor2_2 _2258_ (.A(_1120_),
    .B(_1123_),
    .Y(_1129_));
 sky130_fd_sc_hd__a21oi_1 _2259_ (.A1(_1128_),
    .A2(_1129_),
    .B1(_1124_),
    .Y(_1130_));
 sky130_fd_sc_hd__nor2_4 _2260_ (.A(_1119_),
    .B(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__a21o_1 _2261_ (.A1(_1131_),
    .A2(_1118_),
    .B1(_1117_),
    .X(_1132_));
 sky130_fd_sc_hd__a21o_1 _2262_ (.A1(_1105_),
    .A2(_1132_),
    .B1(_1104_),
    .X(_1133_));
 sky130_fd_sc_hd__a211o_1 _2263_ (.A1(_1105_),
    .A2(_1132_),
    .B1(_1104_),
    .C1(_1088_),
    .X(_1134_));
 sky130_fd_sc_hd__nor2_4 _2264_ (.A(_1088_),
    .B(_1086_),
    .Y(_1135_));
 sky130_fd_sc_hd__and3_1 _2265_ (.A(_1067_),
    .B(_1087_),
    .C(_1134_),
    .X(_1136_));
 sky130_fd_sc_hd__a31o_4 _2266_ (.A1(_1067_),
    .A2(_1134_),
    .A3(_1087_),
    .B1(_1066_),
    .X(_1137_));
 sky130_fd_sc_hd__a21o_4 _2267_ (.A1(_1041_),
    .A2(_1137_),
    .B1(_1040_),
    .X(_1138_));
 sky130_fd_sc_hd__and3_1 _2268_ (.A(_0945_),
    .B(_0949_),
    .C(_0950_),
    .X(_1139_));
 sky130_fd_sc_hd__nor2_2 _2269_ (.A(_0951_),
    .B(_1139_),
    .Y(_1140_));
 sky130_fd_sc_hd__o21a_1 _2270_ (.A1(_0998_),
    .A2(_1000_),
    .B1(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__nor3_1 _2271_ (.A(_0998_),
    .B(_1000_),
    .C(_1140_),
    .Y(_1142_));
 sky130_fd_sc_hd__nor2_4 _2272_ (.A(_1142_),
    .B(_1141_),
    .Y(_1143_));
 sky130_fd_sc_hd__and2_4 _2273_ (.A(_1143_),
    .B(_1138_),
    .X(_1144_));
 sky130_fd_sc_hd__o21a_1 _2274_ (.A1(_0951_),
    .A2(_1141_),
    .B1(_0952_),
    .X(_1145_));
 sky130_fd_sc_hd__a31oi_4 _2275_ (.A1(_0954_),
    .A2(_1138_),
    .A3(_1143_),
    .B1(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__nand2_2 _2276_ (.A(_0890_),
    .B(_0904_),
    .Y(_1147_));
 sky130_fd_sc_hd__and2b_1 _2277_ (.A_N(_0905_),
    .B(_1147_),
    .X(_1148_));
 sky130_fd_sc_hd__and2b_1 _2278_ (.A_N(_1146_),
    .B(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__or2_4 _2279_ (.A(_0667_),
    .B(_0521_),
    .X(_1150_));
 sky130_fd_sc_hd__o22ai_2 _2280_ (.A1(_0667_),
    .A2(net618),
    .B1(_0710_),
    .B2(_0521_),
    .Y(_1151_));
 sky130_fd_sc_hd__o21ai_4 _2281_ (.A1(_1150_),
    .A2(_0893_),
    .B1(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__o2bb2ai_1 _2282_ (.A1_N(_0810_),
    .A2_N(_0892_),
    .B1(_0894_),
    .B2(_0891_),
    .Y(_1153_));
 sky130_fd_sc_hd__nand2b_4 _2283_ (.A_N(_1152_),
    .B(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__xnor2_2 _2284_ (.A(_1152_),
    .B(_1153_),
    .Y(_1155_));
 sky130_fd_sc_hd__nand2_2 _2285_ (.A(_0896_),
    .B(_1155_),
    .Y(_1156_));
 sky130_fd_sc_hd__or2_1 _2286_ (.A(_0896_),
    .B(_1155_),
    .X(_1157_));
 sky130_fd_sc_hd__and2_4 _2287_ (.A(_1157_),
    .B(_1156_),
    .X(_1158_));
 sky130_fd_sc_hd__nor2_8 _2288_ (.A(_0903_),
    .B(_0900_),
    .Y(_1159_));
 sky130_fd_sc_hd__xnor2_4 _2289_ (.A(_1159_),
    .B(_1158_),
    .Y(_1160_));
 sky130_fd_sc_hd__o21a_1 _2290_ (.A1(_0905_),
    .A2(_1149_),
    .B1(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__and2_1 _2291_ (.A(_0903_),
    .B(_1158_),
    .X(_1162_));
 sky130_fd_sc_hd__nor2_1 _2292_ (.A(_0892_),
    .B(_1150_),
    .Y(_1163_));
 sky130_fd_sc_hd__xnor2_4 _2293_ (.A(_1163_),
    .B(_1154_),
    .Y(_1164_));
 sky130_fd_sc_hd__a21oi_4 _2294_ (.A1(_0900_),
    .A2(_1158_),
    .B1(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__and3_1 _2295_ (.A(_0896_),
    .B(_1155_),
    .C(_1164_),
    .X(_1166_));
 sky130_fd_sc_hd__a31o_1 _2296_ (.A1(_0900_),
    .A2(_1158_),
    .A3(_1164_),
    .B1(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__a21oi_4 _2297_ (.A1(_1165_),
    .A2(_1156_),
    .B1(_1167_),
    .Y(_1168_));
 sky130_fd_sc_hd__or3_4 _2298_ (.A(_1161_),
    .B(_1168_),
    .C(_1162_),
    .X(_1169_));
 sky130_fd_sc_hd__o21ai_4 _2299_ (.A1(_1162_),
    .A2(_1161_),
    .B1(_1168_),
    .Y(_1170_));
 sky130_fd_sc_hd__nand2_4 _2300_ (.A(_1169_),
    .B(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__and2b_1 _2301_ (.A_N(_1171_),
    .B(_0459_),
    .X(_1172_));
 sky130_fd_sc_hd__xnor2_4 _2302_ (.A(_0459_),
    .B(_1171_),
    .Y(_1173_));
 sky130_fd_sc_hd__mux4_1 _2303_ (.A0(net1019),
    .A1(net1039),
    .A2(net1035),
    .A3(net984),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_1174_));
 sky130_fd_sc_hd__nand2b_1 _2304_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ),
    .B(_1174_),
    .Y(_1175_));
 sky130_fd_sc_hd__mux4_1 _2305_ (.A0(net1044),
    .A1(net1030),
    .A2(net1048),
    .A3(net1058),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ),
    .X(_1176_));
 sky130_fd_sc_hd__nand2_1 _2306_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ),
    .B(_1176_),
    .Y(_1177_));
 sky130_fd_sc_hd__mux4_2 _2307_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .A1(net1264),
    .A2(net192),
    .A3(net11),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ),
    .X(_1178_));
 sky130_fd_sc_hd__mux4_1 _2308_ (.A0(net57),
    .A1(net59),
    .A2(net67),
    .A3(net1226),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_1179_));
 sky130_fd_sc_hd__mux2_2 _2309_ (.A0(_1178_),
    .A1(_1179_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ),
    .X(_1180_));
 sky130_fd_sc_hd__nor2_1 _2310_ (.A(_1180_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q ),
    .Y(_1181_));
 sky130_fd_sc_hd__a31o_1 _2311_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q ),
    .A2(_1175_),
    .A3(_1177_),
    .B1(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__inv_2 _2312_ (.A(_1182_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 ));
 sky130_fd_sc_hd__mux4_2 _2313_ (.A0(net13),
    .A1(net105),
    .A2(net69),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q ),
    .X(_1183_));
 sky130_fd_sc_hd__mux2_2 _2314_ (.A0(net868),
    .A1(net14),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q ),
    .X(_1184_));
 sky130_fd_sc_hd__nand2b_1 _2315_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q ),
    .B(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__mux2_1 _2316_ (.A0(net70),
    .A1(net106),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q ),
    .X(_1186_));
 sky130_fd_sc_hd__nand2_1 _2317_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q ),
    .B(_1186_),
    .Y(_1187_));
 sky130_fd_sc_hd__a31o_1 _2318_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q ),
    .A2(_1185_),
    .A3(_1187_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q ),
    .X(_1188_));
 sky130_fd_sc_hd__o21ba_1 _2319_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q ),
    .A2(_1183_),
    .B1_N(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__nand2_4 _2320_ (.A(_0494_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q ),
    .Y(_1190_));
 sky130_fd_sc_hd__o211a_1 _2321_ (.A1(net116),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q ),
    .C1(_1190_),
    .X(_1191_));
 sky130_fd_sc_hd__mux2_1 _2322_ (.A0(net26),
    .A1(net77),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q ),
    .X(_1192_));
 sky130_fd_sc_hd__inv_2 _2323_ (.A(_1192_),
    .Y(_1193_));
 sky130_fd_sc_hd__o21ai_1 _2324_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q ),
    .A2(_1193_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q ),
    .Y(_1194_));
 sky130_fd_sc_hd__mux4_2 _2325_ (.A0(net208),
    .A1(net6),
    .A2(net62),
    .A3(net98),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q ),
    .X(_1195_));
 sky130_fd_sc_hd__o221a_1 _2326_ (.A1(_1194_),
    .A2(_1191_),
    .B1(_1195_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q ),
    .X(_1196_));
 sky130_fd_sc_hd__or2_4 _2327_ (.A(_1196_),
    .B(_1189_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X ));
 sky130_fd_sc_hd__nor2_4 _2328_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X ),
    .B(net1064),
    .Y(_1197_));
 sky130_fd_sc_hd__a21o_1 _2329_ (.A1(net1064),
    .A2(_0171_),
    .B1(net1068),
    .X(_1198_));
 sky130_fd_sc_hd__o2bb2a_4 _2330_ (.A1_N(net1068),
    .A2_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[13] ),
    .B1(_1198_),
    .B2(_1197_),
    .X(_1199_));
 sky130_fd_sc_hd__nor3_2 _2331_ (.A(_0905_),
    .B(_1160_),
    .C(_1149_),
    .Y(_1200_));
 sky130_fd_sc_hd__or2_4 _2332_ (.A(_1200_),
    .B(_1161_),
    .X(_1201_));
 sky130_fd_sc_hd__nor2_1 _2333_ (.A(_1199_),
    .B(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__xor2_2 _2334_ (.A(_1201_),
    .B(_1199_),
    .X(_1203_));
 sky130_fd_sc_hd__mux4_2 _2335_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .A1(net16),
    .A2(net72),
    .A3(net108),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q ),
    .X(_1204_));
 sky130_fd_sc_hd__mux2_4 _2336_ (.A0(net79),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_1205_));
 sky130_fd_sc_hd__mux2_1 _2337_ (.A0(net208),
    .A1(net7),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_1206_));
 sky130_fd_sc_hd__inv_2 _2338_ (.A(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__mux4_1 _2339_ (.A0(net1019),
    .A1(net1038),
    .A2(net1034),
    .A3(net984),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1208_));
 sky130_fd_sc_hd__nand2b_1 _2340_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ),
    .B(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__mux4_1 _2341_ (.A0(net1043),
    .A1(net1030),
    .A2(net1047),
    .A3(net1057),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ),
    .X(_1210_));
 sky130_fd_sc_hd__nand2_1 _2342_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ),
    .B(_1210_),
    .Y(_1211_));
 sky130_fd_sc_hd__mux4_1 _2343_ (.A0(net57),
    .A1(net59),
    .A2(net67),
    .A3(net1226),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1212_));
 sky130_fd_sc_hd__mux4_1 _2344_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .A1(net1264),
    .A2(net192),
    .A3(net11),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ),
    .X(_1213_));
 sky130_fd_sc_hd__mux2_1 _2345_ (.A0(_1213_),
    .A1(_1212_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ),
    .X(_1214_));
 sky130_fd_sc_hd__nor2_1 _2346_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q ),
    .B(_1214_),
    .Y(_1215_));
 sky130_fd_sc_hd__a31o_2 _2347_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q ),
    .A2(_1209_),
    .A3(_1211_),
    .B1(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__inv_1 _2348_ (.A(_1216_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ));
 sky130_fd_sc_hd__mux4_2 _2349_ (.A0(net189),
    .A1(net8),
    .A2(net64),
    .A3(net116),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q ),
    .X(_1217_));
 sky130_fd_sc_hd__nand2b_1 _2350_ (.A_N(_1204_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q ),
    .Y(_1218_));
 sky130_fd_sc_hd__mux2_1 _2351_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .A1(net15),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q ),
    .X(_1219_));
 sky130_fd_sc_hd__nand2_1 _2352_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q ),
    .B(_1216_),
    .Y(_1220_));
 sky130_fd_sc_hd__o21a_1 _2353_ (.A1(net71),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q ),
    .X(_1221_));
 sky130_fd_sc_hd__a221o_1 _2354_ (.A1(_0110_),
    .A2(_1219_),
    .B1(_1220_),
    .B2(_1221_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q ),
    .X(_1222_));
 sky130_fd_sc_hd__o21ai_1 _2355_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q ),
    .A2(_1207_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q ),
    .Y(_1223_));
 sky130_fd_sc_hd__a21o_1 _2356_ (.A1(_1205_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q ),
    .B1(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__o211a_1 _2357_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q ),
    .A2(_1217_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q ),
    .C1(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__a31o_1 _2358_ (.A1(_0111_),
    .A2(_1218_),
    .A3(_1222_),
    .B1(_1225_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X ));
 sky130_fd_sc_hd__mux2_4 _2359_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[11] ),
    .S(net1064),
    .X(_1226_));
 sky130_fd_sc_hd__mux2_4 _2360_ (.A0(_1226_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[11] ),
    .S(net1069),
    .X(_1227_));
 sky130_fd_sc_hd__nor2_1 _2361_ (.A(_1141_),
    .B(_1144_),
    .Y(_1228_));
 sky130_fd_sc_hd__xnor2_1 _2362_ (.A(_0953_),
    .B(_1228_),
    .Y(_1229_));
 sky130_fd_sc_hd__and2b_1 _2363_ (.A_N(_1229_),
    .B(_1227_),
    .X(_1230_));
 sky130_fd_sc_hd__nand2b_1 _2364_ (.A_N(_1227_),
    .B(_1229_),
    .Y(_1231_));
 sky130_fd_sc_hd__nand2b_4 _2365_ (.A_N(_1230_),
    .B(_1231_),
    .Y(_1232_));
 sky130_fd_sc_hd__mux2_1 _2366_ (.A0(net100),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q ),
    .X(_1233_));
 sky130_fd_sc_hd__mux2_1 _2367_ (.A0(net201),
    .A1(net8),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q ),
    .X(_1234_));
 sky130_fd_sc_hd__inv_2 _2368_ (.A(_1234_),
    .Y(_1235_));
 sky130_fd_sc_hd__o21ai_1 _2369_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q ),
    .A2(_1235_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ),
    .Y(_1236_));
 sky130_fd_sc_hd__a21o_1 _2370_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q ),
    .A2(_1233_),
    .B1(_1236_),
    .X(_1237_));
 sky130_fd_sc_hd__mux4_1 _2371_ (.A0(net193),
    .A1(net25),
    .A2(net68),
    .A3(net104),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q ),
    .X(_1238_));
 sky130_fd_sc_hd__o21a_1 _2372_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ),
    .A2(_1238_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q ),
    .X(_1239_));
 sky130_fd_sc_hd__mux2_4 _2373_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .A1(net19),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ),
    .X(_1240_));
 sky130_fd_sc_hd__mux4_1 _2374_ (.A0(net1020),
    .A1(net1038),
    .A2(net1035),
    .A3(net985),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_1241_));
 sky130_fd_sc_hd__mux4_1 _2375_ (.A0(net1043),
    .A1(net1030),
    .A2(net1047),
    .A3(net1015),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_1242_));
 sky130_fd_sc_hd__mux2_1 _2376_ (.A0(_1241_),
    .A1(_1242_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ),
    .X(_1243_));
 sky130_fd_sc_hd__mux4_1 _2377_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .A1(net1264),
    .A2(net192),
    .A3(net11),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_1244_));
 sky130_fd_sc_hd__and2b_1 _2378_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ),
    .B(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__mux4_1 _2379_ (.A0(net59),
    .A1(net67),
    .A2(net93),
    .A3(net1226),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_1246_));
 sky130_fd_sc_hd__a211o_1 _2380_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ),
    .A2(_1246_),
    .B1(_1245_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q ),
    .X(_1247_));
 sky130_fd_sc_hd__o21ai_2 _2381_ (.A1(_0108_),
    .A2(_1243_),
    .B1(_1247_),
    .Y(_1248_));
 sky130_fd_sc_hd__inv_1 _2382_ (.A(_1248_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 ));
 sky130_fd_sc_hd__nand2_1 _2383_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ),
    .B(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hd__o211a_1 _2384_ (.A1(net111),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q ),
    .C1(_1249_),
    .X(_1250_));
 sky130_fd_sc_hd__a211o_1 _2385_ (.A1(_0109_),
    .A2(_1240_),
    .B1(_1250_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ),
    .X(_1251_));
 sky130_fd_sc_hd__a21oi_1 _2386_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ),
    .A2(_0560_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q ),
    .Y(_1252_));
 sky130_fd_sc_hd__a22o_1 _2387_ (.A1(_1237_),
    .A2(_1239_),
    .B1(_1252_),
    .B2(_1251_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X ));
 sky130_fd_sc_hd__mux2_4 _2388_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[10] ),
    .S(net1065),
    .X(_1253_));
 sky130_fd_sc_hd__mux2_4 _2389_ (.A0(_1253_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[10] ),
    .S(net1069),
    .X(_1254_));
 sky130_fd_sc_hd__nor2_4 _2390_ (.A(_1138_),
    .B(_1143_),
    .Y(_1255_));
 sky130_fd_sc_hd__nor2_8 _2391_ (.A(_1255_),
    .B(_1144_),
    .Y(_1256_));
 sky130_fd_sc_hd__nand2_1 _2392_ (.A(_1254_),
    .B(_1256_),
    .Y(_1257_));
 sky130_fd_sc_hd__xnor2_4 _2393_ (.A(_1256_),
    .B(_1254_),
    .Y(_1258_));
 sky130_fd_sc_hd__mux4_1 _2394_ (.A0(net922),
    .A1(net971),
    .A2(net981),
    .A3(net1000),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1259_));
 sky130_fd_sc_hd__and2b_1 _2395_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ),
    .B(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__mux4_1 _2396_ (.A0(net991),
    .A1(net1025),
    .A2(net1006),
    .A3(net1012),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1261_));
 sky130_fd_sc_hd__a21bo_1 _2397_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ),
    .A2(_1261_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q ),
    .X(_1262_));
 sky130_fd_sc_hd__mux4_2 _2398_ (.A0(_0442_),
    .A1(_0344_),
    .A2(net75),
    .A3(net1073),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1263_));
 sky130_fd_sc_hd__mux4_1 _2399_ (.A0(net176),
    .A1(net1224),
    .A2(net184),
    .A3(net129),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .X(_1264_));
 sky130_fd_sc_hd__mux2_4 _2400_ (.A0(_1264_),
    .A1(_1263_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ),
    .X(_1265_));
 sky130_fd_sc_hd__o22a_1 _2401_ (.A1(_1260_),
    .A2(_1262_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q ),
    .B2(_1265_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ));
 sky130_fd_sc_hd__nor2_1 _2402_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .B(_0442_),
    .Y(_1266_));
 sky130_fd_sc_hd__a211o_1 _2403_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(net630),
    .B1(_1266_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_1267_));
 sky130_fd_sc_hd__mux2_1 _2404_ (.A0(net89),
    .A1(net232),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1268_));
 sky130_fd_sc_hd__nand2_1 _2405_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .B(_1268_),
    .Y(_1269_));
 sky130_fd_sc_hd__and3_1 _2406_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .B(_1267_),
    .C(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__mux4_1 _2407_ (.A0(net174),
    .A1(net178),
    .A2(net119),
    .A3(net123),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_1271_));
 sky130_fd_sc_hd__nor2_1 _2408_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .B(_1271_),
    .Y(_1272_));
 sky130_fd_sc_hd__mux4_2 _2409_ (.A0(net991),
    .A1(net1023),
    .A2(net996),
    .A3(net812),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1273_));
 sky130_fd_sc_hd__nor2_1 _2410_ (.A(_1273_),
    .B(_0149_),
    .Y(_1274_));
 sky130_fd_sc_hd__mux4_1 _2411_ (.A0(net975),
    .A1(net972),
    .A2(net979),
    .A3(net831),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_1275_));
 sky130_fd_sc_hd__o21ai_1 _2412_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_1275_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q ),
    .Y(_1276_));
 sky130_fd_sc_hd__o32a_1 _2413_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q ),
    .A2(_1270_),
    .A3(_1272_),
    .B1(_1276_),
    .B2(_1274_),
    .X(_1277_));
 sky130_fd_sc_hd__inv_1 _2414_ (.A(_1277_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 ));
 sky130_fd_sc_hd__a21oi_2 _2415_ (.A1(_1277_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ),
    .Y(_1278_));
 sky130_fd_sc_hd__o21a_1 _2416_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .A2(net809),
    .B1(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__nand2_1 _2417_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .B(net629),
    .Y(_1280_));
 sky130_fd_sc_hd__o21ba_4 _2418_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .A2(_0442_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_1281_));
 sky130_fd_sc_hd__mux2_1 _2419_ (.A0(net75),
    .A1(net1073),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .X(_1282_));
 sky130_fd_sc_hd__a221o_1 _2420_ (.A1(_1281_),
    .A2(_1280_),
    .B1(_1282_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .C1(_0154_),
    .X(_1283_));
 sky130_fd_sc_hd__mux4_1 _2421_ (.A0(net176),
    .A1(net1224),
    .A2(net184),
    .A3(net129),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .X(_1284_));
 sky130_fd_sc_hd__o21ba_1 _2422_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .A2(_1284_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q ),
    .X(_1285_));
 sky130_fd_sc_hd__mux4_2 _2423_ (.A0(net990),
    .A1(net1023),
    .A2(net1004),
    .A3(net1011),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_1286_));
 sky130_fd_sc_hd__mux4_1 _2424_ (.A0(net974),
    .A1(net969),
    .A2(net978),
    .A3(net998),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_1287_));
 sky130_fd_sc_hd__or2_1 _2425_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .B(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__o21a_1 _2426_ (.A1(_0154_),
    .A2(_1286_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q ),
    .X(_1289_));
 sky130_fd_sc_hd__a22o_4 _2427_ (.A1(_1285_),
    .A2(_1283_),
    .B1(_1288_),
    .B2(_1289_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ));
 sky130_fd_sc_hd__mux4_1 _2428_ (.A0(_0442_),
    .A1(_0344_),
    .A2(net69),
    .A3(net210),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_1290_));
 sky130_fd_sc_hd__or2_1 _2429_ (.A(_0155_),
    .B(_1290_),
    .X(_1291_));
 sky130_fd_sc_hd__mux4_1 _2430_ (.A0(net174),
    .A1(net178),
    .A2(net119),
    .A3(net123),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_1292_));
 sky130_fd_sc_hd__o21ba_1 _2431_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q ),
    .A2(_1292_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q ),
    .X(_1293_));
 sky130_fd_sc_hd__mux4_1 _2432_ (.A0(net974),
    .A1(net972),
    .A2(net978),
    .A3(net831),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_1294_));
 sky130_fd_sc_hd__mux4_1 _2433_ (.A0(net990),
    .A1(net1024),
    .A2(net996),
    .A3(net1010),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .X(_1295_));
 sky130_fd_sc_hd__mux2_1 _2434_ (.A0(_1294_),
    .A1(_1295_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q ),
    .X(_1296_));
 sky130_fd_sc_hd__a221o_1 _2435_ (.A1(_1291_),
    .A2(_1293_),
    .B1(_1296_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q ),
    .C1(_0148_),
    .X(_1297_));
 sky130_fd_sc_hd__o211a_1 _2436_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ),
    .B1(_1297_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ),
    .X(_1298_));
 sky130_fd_sc_hd__or2_1 _2437_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .X(_1299_));
 sky130_fd_sc_hd__a21oi_1 _2438_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .A2(_0453_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ),
    .Y(_1300_));
 sky130_fd_sc_hd__mux4_1 _2439_ (.A0(net974),
    .A1(net972),
    .A2(net978),
    .A3(net831),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_1301_));
 sky130_fd_sc_hd__mux4_1 _2440_ (.A0(net989),
    .A1(net1023),
    .A2(net864),
    .A3(net1008),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_1302_));
 sky130_fd_sc_hd__or2_1 _2441_ (.A(_0152_),
    .B(_1302_),
    .X(_1303_));
 sky130_fd_sc_hd__o211a_1 _2442_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .A2(_1301_),
    .B1(_1303_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q ),
    .X(_1304_));
 sky130_fd_sc_hd__or2_1 _2443_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .B(_0442_),
    .X(_1305_));
 sky130_fd_sc_hd__a21oi_1 _2444_ (.A1(_0050_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .Y(_1306_));
 sky130_fd_sc_hd__mux2_1 _2445_ (.A0(net210),
    .A1(net1073),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_1307_));
 sky130_fd_sc_hd__a221o_1 _2446_ (.A1(_1305_),
    .A2(_1306_),
    .B1(_1307_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .C1(_0152_),
    .X(_1308_));
 sky130_fd_sc_hd__mux4_1 _2447_ (.A0(net174),
    .A1(net178),
    .A2(net119),
    .A3(net123),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_1309_));
 sky130_fd_sc_hd__or2_1 _2448_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .B(_1309_),
    .X(_1310_));
 sky130_fd_sc_hd__a31o_1 _2449_ (.A1(_0153_),
    .A2(_1308_),
    .A3(_1310_),
    .B1(_1304_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 ));
 sky130_fd_sc_hd__mux4_2 _2450_ (.A0(net974),
    .A1(net969),
    .A2(net979),
    .A3(net831),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_1311_));
 sky130_fd_sc_hd__mux4_1 _2451_ (.A0(net989),
    .A1(net1023),
    .A2(net1004),
    .A3(net1008),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_1312_));
 sky130_fd_sc_hd__o21a_1 _2452_ (.A1(_0151_),
    .A2(_1312_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_1313_));
 sky130_fd_sc_hd__o21ai_4 _2453_ (.A1(_1311_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .B1(_1313_),
    .Y(_1314_));
 sky130_fd_sc_hd__mux2_4 _2454_ (.A0(_0343_),
    .A1(_0068_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_1315_));
 sky130_fd_sc_hd__mux2_1 _2455_ (.A0(net210),
    .A1(net1073),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_1316_));
 sky130_fd_sc_hd__nand2_1 _2456_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .B(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__o211a_1 _2457_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .A2(_1315_),
    .B1(_1317_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .X(_1318_));
 sky130_fd_sc_hd__mux4_1 _2458_ (.A0(net176),
    .A1(net1224),
    .A2(net184),
    .A3(net129),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_1319_));
 sky130_fd_sc_hd__nor2_1 _2459_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .B(_1319_),
    .Y(_1320_));
 sky130_fd_sc_hd__o31ai_4 _2460_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q ),
    .A2(_1320_),
    .A3(_1318_),
    .B1(_1314_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ));
 sky130_fd_sc_hd__mux2_1 _2461_ (.A0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ),
    .S(_0148_),
    .X(_1321_));
 sky130_fd_sc_hd__a221o_1 _2462_ (.A1(_1299_),
    .A2(_1300_),
    .B1(_1321_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q ),
    .X(_1322_));
 sky130_fd_sc_hd__o31a_1 _2463_ (.A1(_0150_),
    .A2(_1279_),
    .A3(_1298_),
    .B1(_1322_),
    .X(\Tile_X0Y1_DSP_bot.C9 ));
 sky130_fd_sc_hd__mux2_4 _2464_ (.A0(\Tile_X0Y1_DSP_bot.C9 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[9] ),
    .S(net1063),
    .X(_1323_));
 sky130_fd_sc_hd__mux2_4 _2465_ (.A0(_1323_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[9] ),
    .S(net1067),
    .X(_1324_));
 sky130_fd_sc_hd__xor2_4 _2466_ (.A(_1137_),
    .B(_1041_),
    .X(_1325_));
 sky130_fd_sc_hd__nand2_4 _2467_ (.A(_1325_),
    .B(_1324_),
    .Y(_1326_));
 sky130_fd_sc_hd__nor2_1 _2468_ (.A(_1324_),
    .B(_1325_),
    .Y(_1327_));
 sky130_fd_sc_hd__or2_1 _2469_ (.A(_1324_),
    .B(_1325_),
    .X(_1328_));
 sky130_fd_sc_hd__and2_4 _2470_ (.A(_1326_),
    .B(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__nand2_2 _2471_ (.A(_0588_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .Y(_1330_));
 sky130_fd_sc_hd__o211a_1 _2472_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ),
    .B1(_0156_),
    .C1(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__mux4_2 _2473_ (.A0(net655),
    .A1(net971),
    .A2(net980),
    .A3(net1000),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_1332_));
 sky130_fd_sc_hd__or2_4 _2474_ (.A(_1332_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .X(_1333_));
 sky130_fd_sc_hd__mux4_2 _2475_ (.A0(net656),
    .A1(net1005),
    .A2(net995),
    .A3(net653),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_1334_));
 sky130_fd_sc_hd__or2_4 _2476_ (.A(_1334_),
    .B(_0157_),
    .X(_1335_));
 sky130_fd_sc_hd__mux2_1 _2477_ (.A0(_0563_),
    .A1(_0387_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_1336_));
 sky130_fd_sc_hd__and2b_1 _2478_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .B(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__mux2_1 _2479_ (.A0(net76),
    .A1(net1072),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_1338_));
 sky130_fd_sc_hd__a21o_1 _2480_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .A2(_1338_),
    .B1(_0157_),
    .X(_1339_));
 sky130_fd_sc_hd__mux4_1 _2481_ (.A0(net177),
    .A1(net185),
    .A2(net1223),
    .A3(net130),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_1340_));
 sky130_fd_sc_hd__o221a_1 _2482_ (.A1(_1337_),
    .A2(_1339_),
    .B1(_1340_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .C1(_0158_),
    .X(_1341_));
 sky130_fd_sc_hd__a31o_4 _2483_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q ),
    .A2(_1333_),
    .A3(_1335_),
    .B1(_1341_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ));
 sky130_fd_sc_hd__mux4_1 _2484_ (.A0(net974),
    .A1(net969),
    .A2(net978),
    .A3(net998),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_1342_));
 sky130_fd_sc_hd__mux4_1 _2485_ (.A0(net989),
    .A1(net1004),
    .A2(net864),
    .A3(net1008),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_1343_));
 sky130_fd_sc_hd__nor2_1 _2486_ (.A(_0162_),
    .B(_1343_),
    .Y(_1344_));
 sky130_fd_sc_hd__o21ai_1 _2487_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .A2(_1342_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q ),
    .Y(_1345_));
 sky130_fd_sc_hd__mux2_4 _2488_ (.A0(_0563_),
    .A1(_0387_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_1346_));
 sky130_fd_sc_hd__inv_2 _2489_ (.A(_1346_),
    .Y(_1347_));
 sky130_fd_sc_hd__mux2_1 _2490_ (.A0(net76),
    .A1(net1072),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_1348_));
 sky130_fd_sc_hd__nand2_1 _2491_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .B(_1348_),
    .Y(_1349_));
 sky130_fd_sc_hd__o211a_1 _2492_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .A2(_1347_),
    .B1(_1349_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .X(_1350_));
 sky130_fd_sc_hd__mux4_1 _2493_ (.A0(net177),
    .A1(net185),
    .A2(net1223),
    .A3(net130),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_1351_));
 sky130_fd_sc_hd__nor2_1 _2494_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .B(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__o32a_4 _2495_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q ),
    .A2(_1352_),
    .A3(_1350_),
    .B1(_1344_),
    .B2(_1345_),
    .X(_1353_));
 sky130_fd_sc_hd__inv_2 _2496_ (.A(_1353_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 ));
 sky130_fd_sc_hd__nand2_1 _2497_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .B(_1353_),
    .Y(_1354_));
 sky130_fd_sc_hd__o211a_1 _2498_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ),
    .B1(_1354_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ),
    .X(_1355_));
 sky130_fd_sc_hd__mux2_1 _2499_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .X(_1356_));
 sky130_fd_sc_hd__and2_1 _2500_ (.A(_0156_),
    .B(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__mux4_2 _2501_ (.A0(net974),
    .A1(net969),
    .A2(net978),
    .A3(net998),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_1358_));
 sky130_fd_sc_hd__mux4_1 _2502_ (.A0(net989),
    .A1(net1004),
    .A2(net994),
    .A3(net1011),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_1359_));
 sky130_fd_sc_hd__or2_1 _2503_ (.A(_0160_),
    .B(_1359_),
    .X(_1360_));
 sky130_fd_sc_hd__o211a_1 _2504_ (.A1(_1358_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .B1(_1360_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q ),
    .X(_1361_));
 sky130_fd_sc_hd__or2_1 _2505_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .B(_0387_),
    .X(_1362_));
 sky130_fd_sc_hd__a21oi_1 _2506_ (.A1(_0053_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .Y(_1363_));
 sky130_fd_sc_hd__mux2_1 _2507_ (.A0(net211),
    .A1(net1072),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_1364_));
 sky130_fd_sc_hd__a221o_1 _2508_ (.A1(_1362_),
    .A2(_1363_),
    .B1(_1364_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .C1(_0160_),
    .X(_1365_));
 sky130_fd_sc_hd__mux4_1 _2509_ (.A0(net177),
    .A1(net185),
    .A2(net1223),
    .A3(net130),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_1366_));
 sky130_fd_sc_hd__or2_1 _2510_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .B(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__a31o_4 _2511_ (.A1(_1365_),
    .A2(_0161_),
    .A3(_1367_),
    .B1(_1361_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ));
 sky130_fd_sc_hd__mux2_1 _2512_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .X(_1368_));
 sky130_fd_sc_hd__a21o_1 _2513_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ),
    .A2(_1368_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q ),
    .X(_1369_));
 sky130_fd_sc_hd__o32a_4 _2514_ (.A1(_0159_),
    .A2(_1331_),
    .A3(_1355_),
    .B1(_1357_),
    .B2(_1369_),
    .X(\Tile_X0Y1_DSP_bot.C8 ));
 sky130_fd_sc_hd__mux2_4 _2515_ (.A0(\Tile_X0Y1_DSP_bot.C8 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[8] ),
    .S(net1065),
    .X(_1370_));
 sky130_fd_sc_hd__mux2_4 _2516_ (.A0(_1370_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[8] ),
    .S(net1066),
    .X(_1371_));
 sky130_fd_sc_hd__a21oi_1 _2517_ (.A1(_1087_),
    .A2(_1134_),
    .B1(_1067_),
    .Y(_1372_));
 sky130_fd_sc_hd__nor2_1 _2518_ (.A(_1136_),
    .B(_1372_),
    .Y(_1373_));
 sky130_fd_sc_hd__and2_4 _2519_ (.A(_1371_),
    .B(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__xor2_4 _2520_ (.A(_1371_),
    .B(_1373_),
    .X(_1375_));
 sky130_fd_sc_hd__nand2_1 _2521_ (.A(net1066),
    .B(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[7] ),
    .Y(_1376_));
 sky130_fd_sc_hd__mux4_2 _2522_ (.A0(_0135_),
    .A1(_0134_),
    .A2(_0020_),
    .A3(_0588_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_1377_));
 sky130_fd_sc_hd__inv_4 _2523_ (.A(_1377_),
    .Y(_1378_));
 sky130_fd_sc_hd__nand2_1 _2524_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .B(_1377_),
    .Y(_1379_));
 sky130_fd_sc_hd__mux4_2 _2525_ (.A0(net179),
    .A1(net144),
    .A2(net70),
    .A3(net215),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q ),
    .X(_1380_));
 sky130_fd_sc_hd__o211a_1 _2526_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(_1380_),
    .B1(_1379_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q ),
    .X(_1381_));
 sky130_fd_sc_hd__nand2_2 _2527_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .B(_1353_),
    .Y(_1382_));
 sky130_fd_sc_hd__o21a_1 _2528_ (.A1(net222),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q ),
    .X(_1383_));
 sky130_fd_sc_hd__mux2_1 _2529_ (.A0(net186),
    .A1(net131),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .X(_1384_));
 sky130_fd_sc_hd__a221o_1 _2530_ (.A1(_1383_),
    .A2(_1382_),
    .B1(_1384_),
    .B2(_0163_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .X(_1385_));
 sky130_fd_sc_hd__mux2_1 _2531_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .A1(net223),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q ),
    .X(_1386_));
 sky130_fd_sc_hd__mux2_1 _2532_ (.A0(net187),
    .A1(net132),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q ),
    .X(_1387_));
 sky130_fd_sc_hd__inv_1 _2533_ (.A(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__o21ai_1 _2534_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q ),
    .A2(_1388_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .Y(_1389_));
 sky130_fd_sc_hd__a21o_1 _2535_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q ),
    .A2(_1386_),
    .B1(_1389_),
    .X(_1390_));
 sky130_fd_sc_hd__a31o_1 _2536_ (.A1(_1385_),
    .A2(_0164_),
    .A3(_1390_),
    .B1(_1381_),
    .X(\Tile_X0Y1_DSP_bot.C7 ));
 sky130_fd_sc_hd__mux2_4 _2537_ (.A0(\Tile_X0Y1_DSP_bot.C7 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[7] ),
    .S(net1063),
    .X(_1391_));
 sky130_fd_sc_hd__nand2b_4 _2538_ (.A_N(net1066),
    .B(_1391_),
    .Y(_1392_));
 sky130_fd_sc_hd__nand2_2 _2539_ (.A(_1376_),
    .B(_1392_),
    .Y(_1393_));
 sky130_fd_sc_hd__xnor2_4 _2540_ (.A(_1135_),
    .B(_1133_),
    .Y(_1394_));
 sky130_fd_sc_hd__a21oi_1 _2541_ (.A1(_1376_),
    .A2(_1392_),
    .B1(_1394_),
    .Y(_1395_));
 sky130_fd_sc_hd__xor2_2 _2542_ (.A(_1394_),
    .B(_1393_),
    .X(_1396_));
 sky130_fd_sc_hd__mux4_1 _2543_ (.A0(net1221),
    .A1(net82),
    .A2(net235),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_1397_));
 sky130_fd_sc_hd__mux4_2 _2544_ (.A0(net203),
    .A1(net128),
    .A2(net74),
    .A3(net219),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q ),
    .X(_1398_));
 sky130_fd_sc_hd__mux2_1 _2545_ (.A0(_1398_),
    .A1(_1397_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ),
    .X(_1399_));
 sky130_fd_sc_hd__mux4_2 _2546_ (.A0(net135),
    .A1(net226),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q ),
    .X(_1400_));
 sky130_fd_sc_hd__or2_1 _2547_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ),
    .B(_1400_),
    .X(_1401_));
 sky130_fd_sc_hd__mux4_1 _2548_ (.A0(net191),
    .A1(net136),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .A3(net227),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q ),
    .X(_1402_));
 sky130_fd_sc_hd__inv_1 _2549_ (.A(_1402_),
    .Y(_1403_));
 sky130_fd_sc_hd__a21oi_1 _2550_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(_1403_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q ),
    .Y(_1404_));
 sky130_fd_sc_hd__a22o_1 _2551_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q ),
    .A2(_1399_),
    .B1(_1401_),
    .B2(_1404_),
    .X(\Tile_X0Y1_DSP_bot.C6 ));
 sky130_fd_sc_hd__mux2_1 _2552_ (.A0(\Tile_X0Y1_DSP_bot.C6 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[6] ),
    .S(net1063),
    .X(_1405_));
 sky130_fd_sc_hd__mux2_1 _2553_ (.A0(_1405_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[6] ),
    .S(net1066),
    .X(_1406_));
 sky130_fd_sc_hd__xor2_2 _2554_ (.A(_1132_),
    .B(_1105_),
    .X(_1407_));
 sky130_fd_sc_hd__nand2_2 _2555_ (.A(_1407_),
    .B(_1406_),
    .Y(_1408_));
 sky130_fd_sc_hd__or2_1 _2556_ (.A(_1406_),
    .B(_1407_),
    .X(_1409_));
 sky130_fd_sc_hd__nand2_4 _2557_ (.A(_1408_),
    .B(_1409_),
    .Y(_1410_));
 sky130_fd_sc_hd__mux2_4 _2558_ (.A0(net216),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_1411_));
 sky130_fd_sc_hd__mux2_1 _2559_ (.A0(net196),
    .A1(net91),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_1412_));
 sky130_fd_sc_hd__inv_2 _2560_ (.A(_1412_),
    .Y(_1413_));
 sky130_fd_sc_hd__o21ai_1 _2561_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_1413_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ),
    .Y(_1414_));
 sky130_fd_sc_hd__a21o_1 _2562_ (.A1(_1411_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .B1(_1414_),
    .X(_1415_));
 sky130_fd_sc_hd__mux4_1 _2563_ (.A0(net181),
    .A1(net126),
    .A2(net89),
    .A3(net217),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q ),
    .X(_1416_));
 sky130_fd_sc_hd__o211a_1 _2564_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ),
    .A2(_1416_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q ),
    .C1(_1415_),
    .X(_1417_));
 sky130_fd_sc_hd__mux2_2 _2565_ (.A0(net224),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q ),
    .X(_1418_));
 sky130_fd_sc_hd__nand2_1 _2566_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q ),
    .B(_0677_),
    .Y(_1419_));
 sky130_fd_sc_hd__o21ba_1 _2567_ (.A1(net188),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q ),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q ),
    .X(_1420_));
 sky130_fd_sc_hd__a221o_1 _2568_ (.A1(_1418_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q ),
    .B1(_1419_),
    .B2(_1420_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ),
    .X(_1421_));
 sky130_fd_sc_hd__mux4_2 _2569_ (.A0(net189),
    .A1(net134),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .A3(net225),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q ),
    .X(_1422_));
 sky130_fd_sc_hd__nand2b_1 _2570_ (.A_N(_1422_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ),
    .Y(_1423_));
 sky130_fd_sc_hd__a31o_1 _2571_ (.A1(_1421_),
    .A2(_0165_),
    .A3(_1423_),
    .B1(_1417_),
    .X(\Tile_X0Y1_DSP_bot.C5 ));
 sky130_fd_sc_hd__nor2_2 _2572_ (.A(\Tile_X0Y1_DSP_bot.C5 ),
    .B(net1063),
    .Y(_1424_));
 sky130_fd_sc_hd__a21o_1 _2573_ (.A1(net1063),
    .A2(_0166_),
    .B1(net1066),
    .X(_1425_));
 sky130_fd_sc_hd__a2bb2o_4 _2574_ (.A1_N(_1425_),
    .A2_N(_1424_),
    .B1(net1066),
    .B2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[5] ),
    .X(_1426_));
 sky130_fd_sc_hd__xor2_4 _2575_ (.A(_1118_),
    .B(_1131_),
    .X(_1427_));
 sky130_fd_sc_hd__nand2_1 _2576_ (.A(_1426_),
    .B(_1427_),
    .Y(_1428_));
 sky130_fd_sc_hd__nor2_4 _2577_ (.A(_1427_),
    .B(_1426_),
    .Y(_1429_));
 sky130_fd_sc_hd__xor2_2 _2578_ (.A(_1426_),
    .B(_1427_),
    .X(_1430_));
 sky130_fd_sc_hd__mux2_1 _2579_ (.A0(net84),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_1431_));
 sky130_fd_sc_hd__mux2_1 _2580_ (.A0(net197),
    .A1(net141),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_1432_));
 sky130_fd_sc_hd__inv_1 _2581_ (.A(_1432_),
    .Y(_1433_));
 sky130_fd_sc_hd__o21ai_1 _2582_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(_1433_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ),
    .Y(_1434_));
 sky130_fd_sc_hd__a21o_1 _2583_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(_1431_),
    .B1(_1434_),
    .X(_1435_));
 sky130_fd_sc_hd__mux4_2 _2584_ (.A0(net185),
    .A1(net130),
    .A2(net76),
    .A3(net232),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q ),
    .X(_1436_));
 sky130_fd_sc_hd__or2_1 _2585_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ),
    .B(_1436_),
    .X(_1437_));
 sky130_fd_sc_hd__mux4_2 _2586_ (.A0(net192),
    .A1(net137),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q ),
    .X(_1438_));
 sky130_fd_sc_hd__mux4_1 _2587_ (.A0(net193),
    .A1(net138),
    .A2(net874),
    .A3(net229),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q ),
    .X(_1439_));
 sky130_fd_sc_hd__inv_2 _2588_ (.A(_1439_),
    .Y(_1440_));
 sky130_fd_sc_hd__a21oi_1 _2589_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ),
    .A2(_1440_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q ),
    .Y(_1441_));
 sky130_fd_sc_hd__o21a_1 _2590_ (.A1(_1438_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ),
    .B1(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__a31o_1 _2591_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q ),
    .A2(_1435_),
    .A3(_1437_),
    .B1(_1442_),
    .X(\Tile_X0Y1_DSP_bot.C4 ));
 sky130_fd_sc_hd__or2_4 _2592_ (.A(net1065),
    .B(\Tile_X0Y1_DSP_bot.C4 ),
    .X(_1443_));
 sky130_fd_sc_hd__a21oi_1 _2593_ (.A1(net1063),
    .A2(_0167_),
    .B1(net1066),
    .Y(_1444_));
 sky130_fd_sc_hd__a22o_4 _2594_ (.A1(net1067),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[4] ),
    .B1(_1444_),
    .B2(_1443_),
    .X(_1445_));
 sky130_fd_sc_hd__xor2_2 _2595_ (.A(_1119_),
    .B(_1130_),
    .X(_1446_));
 sky130_fd_sc_hd__nand2_1 _2596_ (.A(_1445_),
    .B(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__xnor2_4 _2597_ (.A(_1446_),
    .B(_1445_),
    .Y(_1448_));
 sky130_fd_sc_hd__mux2_1 _2598_ (.A0(net233),
    .A1(_0237_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q ),
    .X(_1449_));
 sky130_fd_sc_hd__mux2_1 _2599_ (.A0(net144),
    .A1(net81),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q ),
    .X(_1450_));
 sky130_fd_sc_hd__inv_2 _2600_ (.A(_1450_),
    .Y(_1451_));
 sky130_fd_sc_hd__o21ai_1 _2601_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q ),
    .A2(_1451_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .Y(_1452_));
 sky130_fd_sc_hd__a21o_1 _2602_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q ),
    .A2(_1449_),
    .B1(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__mux4_2 _2603_ (.A0(net204),
    .A1(net124),
    .A2(net70),
    .A3(net215),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q ),
    .X(_1454_));
 sky130_fd_sc_hd__or2_1 _2604_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .B(_1454_),
    .X(_1455_));
 sky130_fd_sc_hd__mux4_2 _2605_ (.A0(net131),
    .A1(net222),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q ),
    .X(_1456_));
 sky130_fd_sc_hd__mux4_2 _2606_ (.A0(net187),
    .A1(net132),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .A3(net223),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q ),
    .X(_1457_));
 sky130_fd_sc_hd__inv_2 _2607_ (.A(_1457_),
    .Y(_1458_));
 sky130_fd_sc_hd__a21oi_1 _2608_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .A2(_1458_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q ),
    .Y(_1459_));
 sky130_fd_sc_hd__o21a_1 _2609_ (.A1(_1456_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .B1(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__a31o_4 _2610_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q ),
    .A2(_1453_),
    .A3(_1455_),
    .B1(_1460_),
    .X(\Tile_X0Y1_DSP_bot.C3 ));
 sky130_fd_sc_hd__or2_4 _2611_ (.A(\Tile_X0Y1_DSP_bot.C3 ),
    .B(net1063),
    .X(_1461_));
 sky130_fd_sc_hd__a21oi_1 _2612_ (.A1(net1063),
    .A2(_0168_),
    .B1(net1066),
    .Y(_1462_));
 sky130_fd_sc_hd__a22oi_4 _2613_ (.A1(net1066),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[3] ),
    .B1(_1462_),
    .B2(_1461_),
    .Y(_1463_));
 sky130_fd_sc_hd__xnor2_2 _2614_ (.A(_1128_),
    .B(_1129_),
    .Y(_1464_));
 sky130_fd_sc_hd__xnor2_2 _2615_ (.A(_1464_),
    .B(_1463_),
    .Y(_1465_));
 sky130_fd_sc_hd__mux4_2 _2616_ (.A0(net183),
    .A1(net128),
    .A2(net90),
    .A3(net219),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q ),
    .X(_1466_));
 sky130_fd_sc_hd__o21ai_1 _2617_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ),
    .A2(_1466_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q ),
    .Y(_1467_));
 sky130_fd_sc_hd__a21o_1 _2618_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ),
    .A2(net660),
    .B1(_1467_),
    .X(_1468_));
 sky130_fd_sc_hd__mux2_4 _2619_ (.A0(net190),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_1469_));
 sky130_fd_sc_hd__and2b_1 _2620_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q ),
    .B(_1469_),
    .X(_1470_));
 sky130_fd_sc_hd__mux2_4 _2621_ (.A0(net226),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_1471_));
 sky130_fd_sc_hd__a21oi_4 _2622_ (.A1(_1471_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q ),
    .B1(_1470_),
    .Y(_1472_));
 sky130_fd_sc_hd__inv_2 _2623_ (.A(net632),
    .Y(_1473_));
 sky130_fd_sc_hd__mux2_1 _2624_ (.A0(net191),
    .A1(net136),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q ),
    .X(_1474_));
 sky130_fd_sc_hd__inv_1 _2625_ (.A(_1474_),
    .Y(_1475_));
 sky130_fd_sc_hd__mux2_2 _2626_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .A1(net227),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q ),
    .X(_1476_));
 sky130_fd_sc_hd__nand2_1 _2627_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q ),
    .B(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__o211a_1 _2628_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q ),
    .A2(_1475_),
    .B1(_1477_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ),
    .X(_1478_));
 sky130_fd_sc_hd__a211o_1 _2629_ (.A1(_1472_),
    .A2(_0169_),
    .B1(_1478_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q ),
    .X(_1479_));
 sky130_fd_sc_hd__nand2_2 _2630_ (.A(_1479_),
    .B(_1468_),
    .Y(\Tile_X0Y1_DSP_bot.C2 ));
 sky130_fd_sc_hd__mux2_4 _2631_ (.A0(\Tile_X0Y1_DSP_bot.C2 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[2] ),
    .S(net1063),
    .X(_1480_));
 sky130_fd_sc_hd__mux2_4 _2632_ (.A0(_1480_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[2] ),
    .S(net1066),
    .X(_1481_));
 sky130_fd_sc_hd__xnor2_4 _2633_ (.A(_1127_),
    .B(_1126_),
    .Y(_1482_));
 sky130_fd_sc_hd__nand2_2 _2634_ (.A(_1482_),
    .B(_1481_),
    .Y(_1483_));
 sky130_fd_sc_hd__xnor2_4 _2635_ (.A(_1482_),
    .B(_1481_),
    .Y(_1484_));
 sky130_fd_sc_hd__mux2_1 _2636_ (.A0(net83),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_1485_));
 sky130_fd_sc_hd__mux2_1 _2637_ (.A0(net204),
    .A1(net125),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_1486_));
 sky130_fd_sc_hd__o21a_1 _2638_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q ),
    .A2(_1486_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .X(_1487_));
 sky130_fd_sc_hd__o21ai_1 _2639_ (.A1(_0170_),
    .A2(_1485_),
    .B1(_1487_),
    .Y(_1488_));
 sky130_fd_sc_hd__mux4_1 _2640_ (.A0(net181),
    .A1(net126),
    .A2(net72),
    .A3(net233),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q ),
    .X(_1489_));
 sky130_fd_sc_hd__nand2b_1 _2641_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .B(_1489_),
    .Y(_1490_));
 sky130_fd_sc_hd__and3_1 _2642_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q ),
    .B(_1488_),
    .C(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__nand2_2 _2643_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q ),
    .Y(_1492_));
 sky130_fd_sc_hd__or2_1 _2644_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q ),
    .B(_0677_),
    .X(_1493_));
 sky130_fd_sc_hd__mux2_1 _2645_ (.A0(net188),
    .A1(net133),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q ),
    .X(_1494_));
 sky130_fd_sc_hd__nor2_1 _2646_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q ),
    .B(_1494_),
    .Y(_1495_));
 sky130_fd_sc_hd__a311o_1 _2647_ (.A1(_1492_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q ),
    .A3(_1493_),
    .B1(_1495_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .X(_1496_));
 sky130_fd_sc_hd__mux4_2 _2648_ (.A0(net189),
    .A1(net134),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .A3(net225),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q ),
    .X(_1497_));
 sky130_fd_sc_hd__a21oi_1 _2649_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_1497_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q ),
    .Y(_1498_));
 sky130_fd_sc_hd__a21oi_2 _2650_ (.A1(_1498_),
    .A2(_1496_),
    .B1(_1491_),
    .Y(\Tile_X0Y1_DSP_bot.C1 ));
 sky130_fd_sc_hd__mux2_4 _2651_ (.A0(\Tile_X0Y1_DSP_bot.C1 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[1] ),
    .S(net1063),
    .X(_1499_));
 sky130_fd_sc_hd__mux2_4 _2652_ (.A0(_1499_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[1] ),
    .S(net1067),
    .X(_1500_));
 sky130_fd_sc_hd__inv_6 _2653_ (.A(_1500_),
    .Y(_1501_));
 sky130_fd_sc_hd__o22a_1 _2654_ (.A1(_0928_),
    .A2(_0981_),
    .B1(net832),
    .B2(_0848_),
    .X(_1502_));
 sky130_fd_sc_hd__a21o_1 _2655_ (.A1(_1121_),
    .A2(_1125_),
    .B1(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__or2_1 _2656_ (.A(_1501_),
    .B(_1503_),
    .X(_1504_));
 sky130_fd_sc_hd__mux2_4 _2657_ (.A0(net217),
    .A1(net619),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q ),
    .X(_1505_));
 sky130_fd_sc_hd__mux2_1 _2658_ (.A0(net197),
    .A1(net126),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q ),
    .X(_1506_));
 sky130_fd_sc_hd__inv_1 _2659_ (.A(_1506_),
    .Y(_1507_));
 sky130_fd_sc_hd__o21ai_1 _2660_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q ),
    .A2(_1507_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .Y(_1508_));
 sky130_fd_sc_hd__a21o_1 _2661_ (.A1(_1505_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q ),
    .B1(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__mux4_1 _2662_ (.A0(net185),
    .A1(net143),
    .A2(net76),
    .A3(net221),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q ),
    .X(_1510_));
 sky130_fd_sc_hd__o211a_1 _2663_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .A2(_1510_),
    .B1(_1509_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q ),
    .X(_1511_));
 sky130_fd_sc_hd__mux2_4 _2664_ (.A0(net228),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .X(_1512_));
 sky130_fd_sc_hd__mux2_1 _2665_ (.A0(net192),
    .A1(net137),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .X(_1513_));
 sky130_fd_sc_hd__and2b_1 _2666_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q ),
    .B(_1513_),
    .X(_1514_));
 sky130_fd_sc_hd__a211o_1 _2667_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q ),
    .A2(_1512_),
    .B1(_1514_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .X(_1515_));
 sky130_fd_sc_hd__a21oi_2 _2668_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .A2(_0257_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q ),
    .Y(_1516_));
 sky130_fd_sc_hd__a21o_1 _2669_ (.A1(_1516_),
    .A2(_1515_),
    .B1(_1511_),
    .X(\Tile_X0Y1_DSP_bot.C0 ));
 sky130_fd_sc_hd__mux2_2 _2670_ (.A0(\Tile_X0Y1_DSP_bot.C0 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[0] ),
    .S(net1065),
    .X(_1517_));
 sky130_fd_sc_hd__mux2_4 _2671_ (.A0(_1517_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[0] ),
    .S(net1067),
    .X(_1518_));
 sky130_fd_sc_hd__and2_4 _2672_ (.A(net829),
    .B(_1518_),
    .X(_1519_));
 sky130_fd_sc_hd__inv_2 _2673_ (.A(_1519_),
    .Y(_1520_));
 sky130_fd_sc_hd__xnor2_4 _2674_ (.A(_1503_),
    .B(_1501_),
    .Y(_1521_));
 sky130_fd_sc_hd__o21a_1 _2675_ (.A1(_1520_),
    .A2(_1521_),
    .B1(_1504_),
    .X(_1522_));
 sky130_fd_sc_hd__or2_4 _2676_ (.A(_1522_),
    .B(_1484_),
    .X(_1523_));
 sky130_fd_sc_hd__a21oi_4 _2677_ (.A1(_1483_),
    .A2(_1523_),
    .B1(_1465_),
    .Y(_1524_));
 sky130_fd_sc_hd__o21ba_4 _2678_ (.A1(_1463_),
    .A2(_1464_),
    .B1_N(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__o21a_4 _2679_ (.A1(_1448_),
    .A2(_1525_),
    .B1(_1447_),
    .X(_1526_));
 sky130_fd_sc_hd__o21ai_4 _2680_ (.A1(_1526_),
    .A2(_1429_),
    .B1(_1428_),
    .Y(_1527_));
 sky130_fd_sc_hd__a21boi_4 _2681_ (.A1(_1527_),
    .A2(_1409_),
    .B1_N(_1408_),
    .Y(_1528_));
 sky130_fd_sc_hd__o21bai_4 _2682_ (.A1(_1528_),
    .A2(_1396_),
    .B1_N(_1395_),
    .Y(_1529_));
 sky130_fd_sc_hd__a21oi_4 _2683_ (.A1(_1375_),
    .A2(_1529_),
    .B1(_1374_),
    .Y(_1530_));
 sky130_fd_sc_hd__o21a_4 _2684_ (.A1(_1530_),
    .A2(_1327_),
    .B1(_1326_),
    .X(_1531_));
 sky130_fd_sc_hd__o21ai_4 _2685_ (.A1(_1531_),
    .A2(_1258_),
    .B1(_1257_),
    .Y(_1532_));
 sky130_fd_sc_hd__a21o_1 _2686_ (.A1(_1532_),
    .A2(_1231_),
    .B1(_1230_),
    .X(_1533_));
 sky130_fd_sc_hd__nand2_1 _2687_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q ),
    .B(_0554_),
    .Y(_1534_));
 sky130_fd_sc_hd__mux4_2 _2688_ (.A0(net191),
    .A1(net86),
    .A2(net10),
    .A3(net102),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q ),
    .X(_1535_));
 sky130_fd_sc_hd__or2_1 _2689_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q ),
    .B(_1535_),
    .X(_1536_));
 sky130_fd_sc_hd__mux4_2 _2690_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .A1(net109),
    .A2(net73),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_1537_));
 sky130_fd_sc_hd__nor2_1 _2691_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .Y(_1538_));
 sky130_fd_sc_hd__a211o_1 _2692_ (.A1(_0070_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q ),
    .C1(_1538_),
    .X(_1539_));
 sky130_fd_sc_hd__mux2_1 _2693_ (.A0(net74),
    .A1(net110),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q ),
    .X(_1540_));
 sky130_fd_sc_hd__nand2_1 _2694_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q ),
    .B(_1540_),
    .Y(_1541_));
 sky130_fd_sc_hd__a31o_1 _2695_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q ),
    .A2(_1539_),
    .A3(_1541_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q ),
    .X(_1542_));
 sky130_fd_sc_hd__o21ba_1 _2696_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q ),
    .A2(_1537_),
    .B1_N(_1542_),
    .X(_1543_));
 sky130_fd_sc_hd__a31o_1 _2697_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q ),
    .A2(_1534_),
    .A3(_1536_),
    .B1(_1543_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X ));
 sky130_fd_sc_hd__mux2_1 _2698_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[12] ),
    .S(net1064),
    .X(_1544_));
 sky130_fd_sc_hd__mux2_2 _2699_ (.A0(_1544_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[12] ),
    .S(net1068),
    .X(_1545_));
 sky130_fd_sc_hd__and2b_1 _2700_ (.A_N(_1148_),
    .B(_1146_),
    .X(_1546_));
 sky130_fd_sc_hd__nor2_2 _2701_ (.A(_1546_),
    .B(_1149_),
    .Y(_1547_));
 sky130_fd_sc_hd__nand2_2 _2702_ (.A(_1547_),
    .B(_1545_),
    .Y(_1548_));
 sky130_fd_sc_hd__or2_1 _2703_ (.A(_1545_),
    .B(_1547_),
    .X(_1549_));
 sky130_fd_sc_hd__and2_4 _2704_ (.A(_1548_),
    .B(_1549_),
    .X(_1550_));
 sky130_fd_sc_hd__a21oi_1 _2705_ (.A1(_1199_),
    .A2(_1201_),
    .B1(_1548_),
    .Y(_1551_));
 sky130_fd_sc_hd__a311o_1 _2706_ (.A1(_1533_),
    .A2(_1203_),
    .A3(_1550_),
    .B1(_1551_),
    .C1(_1202_),
    .X(_1552_));
 sky130_fd_sc_hd__xor2_1 _2707_ (.A(_1173_),
    .B(_1552_),
    .X(_1553_));
 sky130_fd_sc_hd__mux2_4 _2708_ (.A0(_1553_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[14] ),
    .S(net1071),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ));
 sky130_fd_sc_hd__nand2_2 _2709_ (.A(_1484_),
    .B(_1522_),
    .Y(_1554_));
 sky130_fd_sc_hd__and2_4 _2710_ (.A(_1554_),
    .B(_1523_),
    .X(_1555_));
 sky130_fd_sc_hd__mux2_4 _2711_ (.A0(_1555_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[2] ),
    .S(net1070),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ));
 sky130_fd_sc_hd__nor2_4 _2712_ (.A(_1518_),
    .B(net829),
    .Y(_1556_));
 sky130_fd_sc_hd__nor2_4 _2713_ (.A(_1556_),
    .B(_1519_),
    .Y(_1557_));
 sky130_fd_sc_hd__mux2_4 _2714_ (.A0(_1557_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[0] ),
    .S(net1070),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ));
 sky130_fd_sc_hd__xor2_1 _2715_ (.A(_1448_),
    .B(_1525_),
    .X(_1558_));
 sky130_fd_sc_hd__mux2_4 _2716_ (.A0(_1558_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[4] ),
    .S(net1070),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ));
 sky130_fd_sc_hd__and3_1 _2717_ (.A(_1465_),
    .B(_1483_),
    .C(_1523_),
    .X(_1559_));
 sky130_fd_sc_hd__nor2_2 _2718_ (.A(_1559_),
    .B(_1524_),
    .Y(_1560_));
 sky130_fd_sc_hd__mux2_4 _2719_ (.A0(_1560_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[3] ),
    .S(net1070),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ));
 sky130_fd_sc_hd__xnor2_2 _2720_ (.A(_1526_),
    .B(_1430_),
    .Y(_1561_));
 sky130_fd_sc_hd__mux2_4 _2721_ (.A0(_1561_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[5] ),
    .S(net1070),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ));
 sky130_fd_sc_hd__xnor2_2 _2722_ (.A(_1410_),
    .B(_1527_),
    .Y(_1562_));
 sky130_fd_sc_hd__mux2_4 _2723_ (.A0(_1562_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[6] ),
    .S(net1070),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ));
 sky130_fd_sc_hd__xor2_1 _2724_ (.A(_1396_),
    .B(_1528_),
    .X(_1563_));
 sky130_fd_sc_hd__mux2_4 _2725_ (.A0(_1563_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[7] ),
    .S(net1070),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ));
 sky130_fd_sc_hd__xnor2_2 _2726_ (.A(_1329_),
    .B(_1530_),
    .Y(_1564_));
 sky130_fd_sc_hd__mux2_4 _2727_ (.A0(_1564_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[9] ),
    .S(net1070),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ));
 sky130_fd_sc_hd__mux2_4 _2728_ (.A0(net987),
    .A1(net1013),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q ),
    .X(_1565_));
 sky130_fd_sc_hd__mux2_4 _2729_ (.A0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ),
    .A1(_1378_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q ),
    .X(_1566_));
 sky130_fd_sc_hd__mux2_8 _2730_ (.A0(_1565_),
    .A1(_1566_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ));
 sky130_fd_sc_hd__xor2_1 _2731_ (.A(_1531_),
    .B(_1258_),
    .X(_1567_));
 sky130_fd_sc_hd__mux2_4 _2732_ (.A0(_1567_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[10] ),
    .S(net1071),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ));
 sky130_fd_sc_hd__xnor2_2 _2733_ (.A(_1232_),
    .B(_1532_),
    .Y(_1568_));
 sky130_fd_sc_hd__mux2_4 _2734_ (.A0(_1568_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[11] ),
    .S(net1071),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ));
 sky130_fd_sc_hd__xor2_2 _2735_ (.A(_1533_),
    .B(_1550_),
    .X(_1569_));
 sky130_fd_sc_hd__mux2_4 _2736_ (.A0(_1569_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[12] ),
    .S(net1071),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ));
 sky130_fd_sc_hd__a21oi_2 _2737_ (.A1(_1173_),
    .A2(_1552_),
    .B1(_1172_),
    .Y(_1570_));
 sky130_fd_sc_hd__a21oi_1 _2738_ (.A1(_0893_),
    .A2(_1154_),
    .B1(_1150_),
    .Y(_1571_));
 sky130_fd_sc_hd__or3b_4 _2739_ (.A(_1167_),
    .B(_1571_),
    .C_N(_1170_),
    .X(_1572_));
 sky130_fd_sc_hd__mux4_1 _2740_ (.A0(net815),
    .A1(net1036),
    .A2(net1032),
    .A3(net985),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_1573_));
 sky130_fd_sc_hd__and2_1 _2741_ (.A(_0115_),
    .B(_1573_),
    .X(_1574_));
 sky130_fd_sc_hd__mux4_2 _2742_ (.A0(net1042),
    .A1(net1029),
    .A2(net1054),
    .A3(net669),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_1575_));
 sky130_fd_sc_hd__a21bo_1 _2743_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ),
    .A2(_1575_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q ),
    .X(_1576_));
 sky130_fd_sc_hd__mux2_4 _2744_ (.A0(net920),
    .A1(net193),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_1577_));
 sky130_fd_sc_hd__mux2_1 _2745_ (.A0(net1263),
    .A1(net12),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_1578_));
 sky130_fd_sc_hd__or2_1 _2746_ (.A(_0114_),
    .B(_1578_),
    .X(_1579_));
 sky130_fd_sc_hd__o211a_1 _2747_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .A2(_1577_),
    .B1(_1579_),
    .C1(_0115_),
    .X(_1580_));
 sky130_fd_sc_hd__mux2_1 _2748_ (.A0(net58),
    .A1(net60),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_1581_));
 sky130_fd_sc_hd__or2_1 _2749_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .B(_1581_),
    .X(_1582_));
 sky130_fd_sc_hd__mux2_1 _2750_ (.A0(net68),
    .A1(net1225),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_1583_));
 sky130_fd_sc_hd__o211a_1 _2751_ (.A1(_0114_),
    .A2(_1583_),
    .B1(_1582_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ),
    .X(_1584_));
 sky130_fd_sc_hd__o32a_4 _2752_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q ),
    .A2(_1580_),
    .A3(_1584_),
    .B1(_1574_),
    .B2(_1576_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ));
 sky130_fd_sc_hd__mux2_4 _2753_ (.A0(net107),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q ),
    .X(_1585_));
 sky130_fd_sc_hd__mux2_1 _2754_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .A1(net71),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q ),
    .X(_1586_));
 sky130_fd_sc_hd__and2b_1 _2755_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q ),
    .B(_1586_),
    .X(_1587_));
 sky130_fd_sc_hd__a211o_1 _2756_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q ),
    .A2(_1585_),
    .B1(_1587_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ),
    .X(_1588_));
 sky130_fd_sc_hd__nand2b_1 _2757_ (.A_N(net641),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ),
    .Y(_1589_));
 sky130_fd_sc_hd__nand2_2 _2758_ (.A(_0744_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q ),
    .Y(_1590_));
 sky130_fd_sc_hd__o211a_1 _2759_ (.A1(net99),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q ),
    .C1(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__mux2_1 _2760_ (.A0(net200),
    .A1(net87),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_1592_));
 sky130_fd_sc_hd__inv_2 _2761_ (.A(_1592_),
    .Y(_1593_));
 sky130_fd_sc_hd__o21ai_1 _2762_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_1593_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ),
    .Y(_1594_));
 sky130_fd_sc_hd__mux4_2 _2763_ (.A0(net189),
    .A1(net8),
    .A2(net85),
    .A3(net100),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q ),
    .X(_1595_));
 sky130_fd_sc_hd__o221a_1 _2764_ (.A1(_1591_),
    .A2(_1594_),
    .B1(_1595_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q ),
    .X(_1596_));
 sky130_fd_sc_hd__a31o_1 _2765_ (.A1(_0116_),
    .A2(_1588_),
    .A3(_1589_),
    .B1(_1596_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X ));
 sky130_fd_sc_hd__or2_4 _2766_ (.A(net1064),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X ),
    .X(_1597_));
 sky130_fd_sc_hd__a21oi_1 _2767_ (.A1(net1064),
    .A2(_0172_),
    .B1(net1068),
    .Y(_1598_));
 sky130_fd_sc_hd__a22o_1 _2768_ (.A1(net1068),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[15] ),
    .B1(_1597_),
    .B2(_1598_),
    .X(_1599_));
 sky130_fd_sc_hd__nand2_1 _2769_ (.A(_1572_),
    .B(_1599_),
    .Y(_1600_));
 sky130_fd_sc_hd__or2_4 _2770_ (.A(_1599_),
    .B(_1572_),
    .X(_1601_));
 sky130_fd_sc_hd__and2_1 _2771_ (.A(_1600_),
    .B(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__xnor2_2 _2772_ (.A(_1602_),
    .B(_1570_),
    .Y(_1603_));
 sky130_fd_sc_hd__mux2_4 _2773_ (.A0(_1603_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[15] ),
    .S(net1071),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ));
 sky130_fd_sc_hd__nand2_2 _2774_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q ),
    .B(_1572_),
    .Y(_1604_));
 sky130_fd_sc_hd__mux2_1 _2775_ (.A0(net118),
    .A1(net654),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q ),
    .X(_1605_));
 sky130_fd_sc_hd__nand2_1 _2776_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q ),
    .B(_1605_),
    .Y(_1606_));
 sky130_fd_sc_hd__mux2_1 _2777_ (.A0(net22),
    .A1(net78),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q ),
    .X(_1607_));
 sky130_fd_sc_hd__inv_2 _2778_ (.A(_1607_),
    .Y(_1608_));
 sky130_fd_sc_hd__o211a_1 _2779_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_1608_),
    .B1(_1606_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ),
    .X(_1609_));
 sky130_fd_sc_hd__mux4_2 _2780_ (.A0(net207),
    .A1(net66),
    .A2(net10),
    .A3(net102),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q ),
    .X(_1610_));
 sky130_fd_sc_hd__o21ai_1 _2781_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ),
    .A2(_1610_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q ),
    .Y(_1611_));
 sky130_fd_sc_hd__nor2_1 _2782_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .Y(_1612_));
 sky130_fd_sc_hd__a211o_1 _2783_ (.A1(_0070_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q ),
    .C1(_1612_),
    .X(_1613_));
 sky130_fd_sc_hd__mux2_1 _2784_ (.A0(net74),
    .A1(net110),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q ),
    .X(_1614_));
 sky130_fd_sc_hd__nand2_1 _2785_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q ),
    .B(_1614_),
    .Y(_1615_));
 sky130_fd_sc_hd__mux4_2 _2786_ (.A0(net17),
    .A1(net109),
    .A2(net73),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q ),
    .X(_1616_));
 sky130_fd_sc_hd__nor2_1 _2787_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ),
    .B(_1616_),
    .Y(_1617_));
 sky130_fd_sc_hd__a311o_1 _2788_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ),
    .A2(_1613_),
    .A3(_1615_),
    .B1(_1617_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q ),
    .X(_1618_));
 sky130_fd_sc_hd__o21ai_1 _2789_ (.A1(_1609_),
    .A2(_1611_),
    .B1(_1618_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X ));
 sky130_fd_sc_hd__mux2_1 _2790_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[16] ),
    .S(net1065),
    .X(_1619_));
 sky130_fd_sc_hd__and2b_1 _2791_ (.A_N(net1068),
    .B(_1619_),
    .X(_1620_));
 sky130_fd_sc_hd__a21oi_1 _2792_ (.A1(net1069),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[16] ),
    .B1(_1620_),
    .Y(_1621_));
 sky130_fd_sc_hd__nor2_1 _2793_ (.A(_1604_),
    .B(_1621_),
    .Y(_1622_));
 sky130_fd_sc_hd__xor2_1 _2794_ (.A(_1604_),
    .B(_1621_),
    .X(_1623_));
 sky130_fd_sc_hd__a221o_1 _2795_ (.A1(_1173_),
    .A2(_1552_),
    .B1(_1572_),
    .B2(_1599_),
    .C1(_1172_),
    .X(_1624_));
 sky130_fd_sc_hd__nand2_4 _2796_ (.A(_1601_),
    .B(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hd__xnor2_2 _2797_ (.A(_1623_),
    .B(_1625_),
    .Y(_1626_));
 sky130_fd_sc_hd__mux2_4 _2798_ (.A0(_1626_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[16] ),
    .S(net1071),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ));
 sky130_fd_sc_hd__a31o_1 _2799_ (.A1(_1601_),
    .A2(_1623_),
    .A3(_1624_),
    .B1(_1622_),
    .X(_1627_));
 sky130_fd_sc_hd__mux4_1 _2800_ (.A0(net187),
    .A1(net62),
    .A2(net26),
    .A3(net98),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q ),
    .X(_1628_));
 sky130_fd_sc_hd__mux2_1 _2801_ (.A0(_0317_),
    .A1(_1628_),
    .S(_0121_),
    .X(_1629_));
 sky130_fd_sc_hd__inv_1 _2802_ (.A(_1629_),
    .Y(_1630_));
 sky130_fd_sc_hd__mux4_2 _2803_ (.A0(net815),
    .A1(net1036),
    .A2(net1032),
    .A3(net983),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_1631_));
 sky130_fd_sc_hd__and2_4 _2804_ (.A(_1631_),
    .B(_0120_),
    .X(_1632_));
 sky130_fd_sc_hd__mux4_2 _2805_ (.A0(net1044),
    .A1(net1028),
    .A2(net1054),
    .A3(net669),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_1633_));
 sky130_fd_sc_hd__a21bo_1 _2806_ (.A1(_1633_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q ),
    .X(_1634_));
 sky130_fd_sc_hd__mux2_1 _2807_ (.A0(_0414_),
    .A1(net193),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_1635_));
 sky130_fd_sc_hd__mux2_1 _2808_ (.A0(net1263),
    .A1(net12),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_1636_));
 sky130_fd_sc_hd__or2_1 _2809_ (.A(_0119_),
    .B(_1636_),
    .X(_1637_));
 sky130_fd_sc_hd__o211a_1 _2810_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .A2(_1635_),
    .B1(_1637_),
    .C1(_0120_),
    .X(_1638_));
 sky130_fd_sc_hd__mux2_1 _2811_ (.A0(net58),
    .A1(net60),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_1639_));
 sky130_fd_sc_hd__or2_1 _2812_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .B(_1639_),
    .X(_1640_));
 sky130_fd_sc_hd__mux2_1 _2813_ (.A0(net68),
    .A1(net1225),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_1641_));
 sky130_fd_sc_hd__o211a_1 _2814_ (.A1(_0119_),
    .A2(_1641_),
    .B1(_1640_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ),
    .X(_1642_));
 sky130_fd_sc_hd__o32a_4 _2815_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q ),
    .A2(_1638_),
    .A3(_1642_),
    .B1(_1634_),
    .B2(_1632_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ));
 sky130_fd_sc_hd__mux2_4 _2816_ (.A0(net105),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q ),
    .X(_1643_));
 sky130_fd_sc_hd__mux2_2 _2817_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .A1(net13),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q ),
    .X(_1644_));
 sky130_fd_sc_hd__and2b_1 _2818_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q ),
    .B(_1644_),
    .X(_1645_));
 sky130_fd_sc_hd__a211o_1 _2819_ (.A1(_1643_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q ),
    .B1(_1645_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ),
    .X(_1646_));
 sky130_fd_sc_hd__mux4_1 _2820_ (.A0(net868),
    .A1(net70),
    .A2(net14),
    .A3(net106),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q ),
    .X(_1647_));
 sky130_fd_sc_hd__o21ai_1 _2821_ (.A1(_0121_),
    .A2(_1647_),
    .B1(_1646_),
    .Y(_1648_));
 sky130_fd_sc_hd__mux2_4 _2822_ (.A0(_1648_),
    .A1(_1630_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q ),
    .X(_1649_));
 sky130_fd_sc_hd__inv_2 _2823_ (.A(_1649_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X ));
 sky130_fd_sc_hd__mux2_4 _2824_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[17] ),
    .S(net1064),
    .X(_1650_));
 sky130_fd_sc_hd__mux2_4 _2825_ (.A0(_1650_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[17] ),
    .S(net1068),
    .X(_1651_));
 sky130_fd_sc_hd__inv_4 _2826_ (.A(_1651_),
    .Y(_1652_));
 sky130_fd_sc_hd__nand2_4 _2827_ (.A(_1604_),
    .B(_1652_),
    .Y(_1653_));
 sky130_fd_sc_hd__nor2_1 _2828_ (.A(_1604_),
    .B(_1652_),
    .Y(_1654_));
 sky130_fd_sc_hd__inv_1 _2829_ (.A(_1654_),
    .Y(_1655_));
 sky130_fd_sc_hd__nand2_4 _2830_ (.A(_1653_),
    .B(_1655_),
    .Y(_1656_));
 sky130_fd_sc_hd__xnor2_2 _2831_ (.A(_1627_),
    .B(_1656_),
    .Y(_1657_));
 sky130_fd_sc_hd__mux2_4 _2832_ (.A0(_1657_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[17] ),
    .S(net1071),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ));
 sky130_fd_sc_hd__mux2_4 _2833_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .X(_1658_));
 sky130_fd_sc_hd__nor2_4 _2834_ (.A(_1658_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ),
    .Y(_1659_));
 sky130_fd_sc_hd__nand2_1 _2835_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ),
    .Y(_1660_));
 sky130_fd_sc_hd__o211a_1 _2836_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .A2(_0744_),
    .B1(_1660_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ),
    .X(_1661_));
 sky130_fd_sc_hd__nand2_4 _2837_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ),
    .Y(_1662_));
 sky130_fd_sc_hd__o211a_1 _2838_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .A2(_0314_),
    .B1(_1662_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ),
    .X(_1663_));
 sky130_fd_sc_hd__mux2_1 _2839_ (.A0(net654),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .X(_1664_));
 sky130_fd_sc_hd__o21ai_1 _2840_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ),
    .A2(_1664_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q ),
    .Y(_1665_));
 sky130_fd_sc_hd__o32a_4 _2841_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q ),
    .A2(_1661_),
    .A3(_1659_),
    .B1(_1663_),
    .B2(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__inv_2 _2842_ (.A(_1666_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X ));
 sky130_fd_sc_hd__mux2_4 _2843_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[18] ),
    .S(net1064),
    .X(_1667_));
 sky130_fd_sc_hd__mux2_4 _2844_ (.A0(_1667_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[18] ),
    .S(net1068),
    .X(_1668_));
 sky130_fd_sc_hd__and3_4 _2845_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q ),
    .B(_1668_),
    .C(_1572_),
    .X(_1669_));
 sky130_fd_sc_hd__a21oi_1 _2846_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q ),
    .A2(_1572_),
    .B1(_1668_),
    .Y(_1670_));
 sky130_fd_sc_hd__nor2_8 _2847_ (.A(_1670_),
    .B(_1669_),
    .Y(_1671_));
 sky130_fd_sc_hd__a311o_1 _2848_ (.A1(_1601_),
    .A2(_1623_),
    .A3(_1624_),
    .B1(_1654_),
    .C1(_1622_),
    .X(_1672_));
 sky130_fd_sc_hd__nand2_1 _2849_ (.A(_1653_),
    .B(_1672_),
    .Y(_1673_));
 sky130_fd_sc_hd__a31o_1 _2850_ (.A1(_1653_),
    .A2(_1671_),
    .A3(_1672_),
    .B1(_1669_),
    .X(_1674_));
 sky130_fd_sc_hd__mux2_1 _2851_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .A1(net876),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_1675_));
 sky130_fd_sc_hd__mux4_1 _2852_ (.A0(net626),
    .A1(net186),
    .A2(net1),
    .A3(net5),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_1676_));
 sky130_fd_sc_hd__mux4_2 _2853_ (.A0(net57),
    .A1(net61),
    .A2(net59),
    .A3(net93),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ),
    .X(_1677_));
 sky130_fd_sc_hd__a21o_1 _2854_ (.A1(_1677_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q ),
    .X(_1678_));
 sky130_fd_sc_hd__a21oi_1 _2855_ (.A1(_0178_),
    .A2(_1676_),
    .B1(_1678_),
    .Y(_1679_));
 sky130_fd_sc_hd__mux4_1 _2856_ (.A0(net1020),
    .A1(net1038),
    .A2(net1034),
    .A3(net984),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_1680_));
 sky130_fd_sc_hd__mux4_1 _2857_ (.A0(net1043),
    .A1(net1047),
    .A2(net1055),
    .A3(net1057),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ),
    .X(_1681_));
 sky130_fd_sc_hd__mux2_1 _2858_ (.A0(_1680_),
    .A1(_1681_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ),
    .X(_1682_));
 sky130_fd_sc_hd__o21ai_1 _2859_ (.A1(_0179_),
    .A2(_1682_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .Y(_1683_));
 sky130_fd_sc_hd__o221a_1 _2860_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(_1182_),
    .B1(_1679_),
    .B2(_1683_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ),
    .X(_1684_));
 sky130_fd_sc_hd__o21ai_1 _2861_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ),
    .A2(_1675_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q ),
    .Y(_1685_));
 sky130_fd_sc_hd__mux4_1 _2862_ (.A0(net1019),
    .A1(net1038),
    .A2(net1034),
    .A3(net984),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_1686_));
 sky130_fd_sc_hd__and2_1 _2863_ (.A(_0177_),
    .B(_1686_),
    .X(_1687_));
 sky130_fd_sc_hd__mux4_1 _2864_ (.A0(net1043),
    .A1(net1047),
    .A2(net1055),
    .A3(net1057),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1688_));
 sky130_fd_sc_hd__a21bo_1 _2865_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_1688_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q ),
    .X(_1689_));
 sky130_fd_sc_hd__mux2_1 _2866_ (.A0(_0239_),
    .A1(net186),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1690_));
 sky130_fd_sc_hd__mux2_1 _2867_ (.A0(net1),
    .A1(net5),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1691_));
 sky130_fd_sc_hd__or2_1 _2868_ (.A(_0176_),
    .B(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__o211a_1 _2869_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .A2(_1690_),
    .B1(_1692_),
    .C1(_0177_),
    .X(_1693_));
 sky130_fd_sc_hd__mux2_1 _2870_ (.A0(net57),
    .A1(net59),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1694_));
 sky130_fd_sc_hd__or2_1 _2871_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .B(_1694_),
    .X(_1695_));
 sky130_fd_sc_hd__mux2_1 _2872_ (.A0(net85),
    .A1(net115),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1696_));
 sky130_fd_sc_hd__o211a_1 _2873_ (.A1(_0176_),
    .A2(_1696_),
    .B1(_1695_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_1697_));
 sky130_fd_sc_hd__o32a_1 _2874_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q ),
    .A2(_1693_),
    .A3(_1697_),
    .B1(_1687_),
    .B2(_1689_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 ));
 sky130_fd_sc_hd__nand2_1 _2875_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 ),
    .Y(_1698_));
 sky130_fd_sc_hd__o211a_1 _2876_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(_1216_),
    .B1(_1698_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ),
    .X(_1699_));
 sky130_fd_sc_hd__mux4_1 _2877_ (.A0(net1019),
    .A1(net1038),
    .A2(net1034),
    .A3(net984),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .X(_1700_));
 sky130_fd_sc_hd__and2_1 _2878_ (.A(_0175_),
    .B(_1700_),
    .X(_1701_));
 sky130_fd_sc_hd__mux4_1 _2879_ (.A0(net1043),
    .A1(net1047),
    .A2(net1055),
    .A3(net669),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_1702_));
 sky130_fd_sc_hd__a21bo_1 _2880_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ),
    .A2(_1702_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q ),
    .X(_1703_));
 sky130_fd_sc_hd__mux2_1 _2881_ (.A0(_0239_),
    .A1(net186),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_1704_));
 sky130_fd_sc_hd__mux2_1 _2882_ (.A0(net1),
    .A1(net23),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_1705_));
 sky130_fd_sc_hd__or2_1 _2883_ (.A(_0174_),
    .B(_1705_),
    .X(_1706_));
 sky130_fd_sc_hd__o211a_1 _2884_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .A2(_1704_),
    .B1(_1706_),
    .C1(_0175_),
    .X(_1707_));
 sky130_fd_sc_hd__mux2_1 _2885_ (.A0(net57),
    .A1(net61),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_1708_));
 sky130_fd_sc_hd__or2_1 _2886_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .B(_1708_),
    .X(_1709_));
 sky130_fd_sc_hd__mux2_1 _2887_ (.A0(net93),
    .A1(net1226),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_1710_));
 sky130_fd_sc_hd__o211a_1 _2888_ (.A1(_0174_),
    .A2(_1710_),
    .B1(_1709_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ),
    .X(_1711_));
 sky130_fd_sc_hd__o32a_1 _2889_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q ),
    .A2(_1707_),
    .A3(_1711_),
    .B1(_1701_),
    .B2(_1703_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 ));
 sky130_fd_sc_hd__a21oi_1 _2890_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ),
    .Y(_1712_));
 sky130_fd_sc_hd__o21a_1 _2891_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(_1248_),
    .B1(_1712_),
    .X(_1713_));
 sky130_fd_sc_hd__or3_1 _2892_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q ),
    .B(_1699_),
    .C(_1713_),
    .X(_1714_));
 sky130_fd_sc_hd__o21ai_2 _2893_ (.A1(_1685_),
    .A2(_1684_),
    .B1(_1714_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X ));
 sky130_fd_sc_hd__mux2_4 _2894_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[19] ),
    .S(net1064),
    .X(_1715_));
 sky130_fd_sc_hd__mux2_4 _2895_ (.A0(_1715_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[19] ),
    .S(net1068),
    .X(_1716_));
 sky130_fd_sc_hd__xor2_1 _2896_ (.A(_1604_),
    .B(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__xnor2_1 _2897_ (.A(_1717_),
    .B(_1674_),
    .Y(_1718_));
 sky130_fd_sc_hd__mux2_4 _2898_ (.A0(_1718_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[19] ),
    .S(net1071),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ));
 sky130_fd_sc_hd__a21boi_1 _2899_ (.A1(_1533_),
    .A2(_1550_),
    .B1_N(_1548_),
    .Y(_1719_));
 sky130_fd_sc_hd__xnor2_2 _2900_ (.A(_1719_),
    .B(_1203_),
    .Y(_1720_));
 sky130_fd_sc_hd__mux2_4 _2901_ (.A0(_1720_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[13] ),
    .S(net1071),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ));
 sky130_fd_sc_hd__xnor2_2 _2902_ (.A(_1673_),
    .B(_1671_),
    .Y(_1721_));
 sky130_fd_sc_hd__mux2_4 _2903_ (.A0(_1721_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[18] ),
    .S(net1071),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ));
 sky130_fd_sc_hd__xnor2_2 _2904_ (.A(_1521_),
    .B(_1519_),
    .Y(_1722_));
 sky130_fd_sc_hd__mux2_4 _2905_ (.A0(_1722_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[1] ),
    .S(net1070),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ));
 sky130_fd_sc_hd__xor2_1 _2906_ (.A(_1375_),
    .B(_1529_),
    .X(_1723_));
 sky130_fd_sc_hd__mux2_4 _2907_ (.A0(_1723_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[8] ),
    .S(net1070),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ));
 sky130_fd_sc_hd__mux4_1 _2908_ (.A0(net1020),
    .A1(net1038),
    .A2(net1034),
    .A3(net984),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_1724_));
 sky130_fd_sc_hd__mux4_1 _2909_ (.A0(net1043),
    .A1(net1030),
    .A2(net1047),
    .A3(net1015),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_1725_));
 sky130_fd_sc_hd__mux2_1 _2910_ (.A0(_1724_),
    .A1(_1725_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ),
    .X(_1726_));
 sky130_fd_sc_hd__mux4_2 _2911_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .A1(net3),
    .A2(net192),
    .A3(net11),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_1727_));
 sky130_fd_sc_hd__and2b_1 _2912_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ),
    .B(_1727_),
    .X(_1728_));
 sky130_fd_sc_hd__mux4_1 _2913_ (.A0(net59),
    .A1(net67),
    .A2(net93),
    .A3(net1226),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_1729_));
 sky130_fd_sc_hd__a21o_1 _2914_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ),
    .A2(_1729_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_1730_));
 sky130_fd_sc_hd__o22a_4 _2915_ (.A1(_0055_),
    .A2(_1726_),
    .B1(_1728_),
    .B2(_1730_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ));
 sky130_fd_sc_hd__mux4_2 _2916_ (.A0(_0414_),
    .A1(net6),
    .A2(net187),
    .A3(net1261),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_1731_));
 sky130_fd_sc_hd__or2_4 _2917_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ),
    .B(_1731_),
    .X(_1732_));
 sky130_fd_sc_hd__mux4_1 _2918_ (.A0(net62),
    .A1(net78),
    .A2(net98),
    .A3(net114),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_1733_));
 sky130_fd_sc_hd__inv_2 _2919_ (.A(_1733_),
    .Y(_1734_));
 sky130_fd_sc_hd__a21oi_1 _2920_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ),
    .A2(_1734_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q ),
    .Y(_1735_));
 sky130_fd_sc_hd__mux4_1 _2921_ (.A0(net1036),
    .A1(net1032),
    .A2(net983),
    .A3(net1044),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_1736_));
 sky130_fd_sc_hd__mux4_1 _2922_ (.A0(net1054),
    .A1(net1048),
    .A2(net1029),
    .A3(net1014),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_1737_));
 sky130_fd_sc_hd__mux2_1 _2923_ (.A0(_1736_),
    .A1(_1737_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ),
    .X(_1738_));
 sky130_fd_sc_hd__a221o_1 _2924_ (.A1(_1735_),
    .A2(_1732_),
    .B1(_1738_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q ),
    .X(_1739_));
 sky130_fd_sc_hd__nand2_1 _2925_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q ),
    .B(_0554_),
    .Y(_1740_));
 sky130_fd_sc_hd__nor2_1 _2926_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q ),
    .B(net983),
    .Y(_1741_));
 sky130_fd_sc_hd__a211oi_1 _2927_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q ),
    .A2(_0560_),
    .B1(_1741_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q ),
    .Y(_1742_));
 sky130_fd_sc_hd__a31o_4 _2928_ (.A1(_1739_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q ),
    .A3(_1740_),
    .B1(_1742_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 ));
 sky130_fd_sc_hd__mux2_4 _2929_ (.A0(net1042),
    .A1(net638),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q ),
    .X(_1743_));
 sky130_fd_sc_hd__mux2_1 _2930_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ),
    .A1(_0317_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q ),
    .X(_1744_));
 sky130_fd_sc_hd__mux2_4 _2931_ (.A0(_1743_),
    .A1(_1744_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 ));
 sky130_fd_sc_hd__o21ai_1 _2932_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q ),
    .Y(_1745_));
 sky130_fd_sc_hd__a21o_1 _2933_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q ),
    .A2(_0384_),
    .B1(_1745_),
    .X(_1746_));
 sky130_fd_sc_hd__nor2_1 _2934_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q ),
    .B(net1050),
    .Y(_1747_));
 sky130_fd_sc_hd__a211o_1 _2935_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q ),
    .A2(_0359_),
    .B1(_1747_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q ),
    .X(_1748_));
 sky130_fd_sc_hd__nand2_1 _2936_ (.A(_1746_),
    .B(_1748_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _2937_ (.A0(net188),
    .A1(net199),
    .A2(net1261),
    .A3(net1042),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2938_ (.A0(net189),
    .A1(net200),
    .A2(net1262),
    .A3(net1053),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _2939_ (.A0(net186),
    .A1(net201),
    .A2(net114),
    .A3(net1048),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _2940_ (.A0(net187),
    .A1(net113),
    .A2(net198),
    .A3(net1028),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 ));
 sky130_fd_sc_hd__mux2_1 _2941_ (.A0(net865),
    .A1(net670),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q ),
    .X(_1749_));
 sky130_fd_sc_hd__mux2_1 _2942_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ),
    .A1(_0429_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q ),
    .X(_1750_));
 sky130_fd_sc_hd__mux2_1 _2943_ (.A0(_1749_),
    .A1(_1750_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2944_ (.A0(net1036),
    .A1(net1032),
    .A2(net985),
    .A3(net1042),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_1751_));
 sky130_fd_sc_hd__or2_1 _2945_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ),
    .B(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__mux4_1 _2946_ (.A0(net1054),
    .A1(net1048),
    .A2(net1029),
    .A3(net1058),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_1753_));
 sky130_fd_sc_hd__o21a_1 _2947_ (.A1(_0081_),
    .A2(_1753_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_1754_));
 sky130_fd_sc_hd__mux4_1 _2948_ (.A0(net1261),
    .A1(net98),
    .A2(net86),
    .A3(net114),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ),
    .X(_1755_));
 sky130_fd_sc_hd__mux4_1 _2949_ (.A0(net187),
    .A1(net199),
    .A2(net1263),
    .A3(net6),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_1756_));
 sky130_fd_sc_hd__mux2_1 _2950_ (.A0(_1755_),
    .A1(_1756_),
    .S(_0081_),
    .X(_1757_));
 sky130_fd_sc_hd__a22o_1 _2951_ (.A1(_1752_),
    .A2(_1754_),
    .B1(_1757_),
    .B2(_0082_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 ));
 sky130_fd_sc_hd__o21ai_1 _2952_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q ),
    .Y(_1758_));
 sky130_fd_sc_hd__a21o_1 _2953_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q ),
    .A2(_0554_),
    .B1(_1758_),
    .X(_1759_));
 sky130_fd_sc_hd__nor2_1 _2954_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q ),
    .B(net1042),
    .Y(_1760_));
 sky130_fd_sc_hd__a211o_1 _2955_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q ),
    .A2(_0560_),
    .B1(_1760_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q ),
    .X(_1761_));
 sky130_fd_sc_hd__nand2_1 _2956_ (.A(_1759_),
    .B(_1761_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 ));
 sky130_fd_sc_hd__mux4_2 _2957_ (.A0(net1053),
    .A1(net641),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ),
    .A3(_0317_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 ));
 sky130_fd_sc_hd__o21ai_1 _2958_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q ),
    .Y(_1762_));
 sky130_fd_sc_hd__a21o_1 _2959_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ),
    .A2(_0384_),
    .B1(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__nor2_1 _2960_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ),
    .B(net828),
    .Y(_1764_));
 sky130_fd_sc_hd__a211o_1 _2961_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ),
    .A2(net621),
    .B1(_1764_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q ),
    .X(_1765_));
 sky130_fd_sc_hd__nand2_1 _2962_ (.A(_1763_),
    .B(_1765_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _2963_ (.A0(net22),
    .A1(net78),
    .A2(net63),
    .A3(net1019),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2964_ (.A0(net21),
    .A1(net79),
    .A2(net64),
    .A3(net1038),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _2965_ (.A0(net61),
    .A1(net114),
    .A2(net80),
    .A3(net1035),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _2966_ (.A0(net62),
    .A1(net77),
    .A2(net113),
    .A3(net986),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _2967_ (.A0(net1050),
    .A1(net670),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .A3(_0429_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2968_ (.A0(_0198_),
    .A1(_0560_),
    .A2(_0599_),
    .A3(_0554_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q ),
    .X(_1766_));
 sky130_fd_sc_hd__inv_1 _2969_ (.A(_1766_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 ));
 sky130_fd_sc_hd__mux4_1 _2970_ (.A0(net824),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .A2(net641),
    .A3(_0317_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _2971_ (.A0(_0199_),
    .A1(net621),
    .A2(_0677_),
    .A3(_0384_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q ),
    .X(_1767_));
 sky130_fd_sc_hd__inv_1 _2972_ (.A(_1767_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _2973_ (.A0(net637),
    .A1(net1264),
    .A2(net1226),
    .A3(net1034),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q ),
    .X(_1768_));
 sky130_fd_sc_hd__mux2_4 _2974_ (.A0(net1047),
    .A1(_0788_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ),
    .X(_1769_));
 sky130_fd_sc_hd__mux2_4 _2975_ (.A0(_0756_),
    .A1(_1595_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ),
    .X(_1770_));
 sky130_fd_sc_hd__mux2_1 _2976_ (.A0(_1769_),
    .A1(_1770_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q ),
    .X(_1771_));
 sky130_fd_sc_hd__mux2_1 _2977_ (.A0(_1768_),
    .A1(_1771_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 ));
 sky130_fd_sc_hd__nor2_1 _2978_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ),
    .B(net1030),
    .Y(_1772_));
 sky130_fd_sc_hd__a211oi_1 _2979_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ),
    .A2(_0571_),
    .B1(_1772_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ),
    .Y(_1773_));
 sky130_fd_sc_hd__mux2_4 _2980_ (.A0(_0700_),
    .A1(_1217_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ),
    .X(_1774_));
 sky130_fd_sc_hd__a21bo_1 _2981_ (.A1(_1774_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q ),
    .X(_1775_));
 sky130_fd_sc_hd__mux4_1 _2982_ (.A0(net920),
    .A1(net1225),
    .A2(net1263),
    .A3(net984),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ),
    .X(_1776_));
 sky130_fd_sc_hd__o22a_1 _2983_ (.A1(_1773_),
    .A2(_1775_),
    .B1(_1776_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 ));
 sky130_fd_sc_hd__or2_1 _2984_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .B(net626),
    .X(_1777_));
 sky130_fd_sc_hd__a21oi_1 _2985_ (.A1(_0027_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ),
    .Y(_1778_));
 sky130_fd_sc_hd__mux2_1 _2986_ (.A0(net93),
    .A1(net1043),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .X(_1779_));
 sky130_fd_sc_hd__a221o_1 _2987_ (.A1(_1777_),
    .A2(_1778_),
    .B1(_1779_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q ),
    .X(_1780_));
 sky130_fd_sc_hd__mux4_1 _2988_ (.A0(net1015),
    .A1(net641),
    .A2(_1204_),
    .A3(_0759_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .X(_1781_));
 sky130_fd_sc_hd__o21a_1 _2989_ (.A1(_0173_),
    .A2(_1781_),
    .B1(_1780_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 ));
 sky130_fd_sc_hd__mux2_4 _2990_ (.A0(net1057),
    .A1(net648),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ),
    .X(_1782_));
 sky130_fd_sc_hd__and2b_1 _2991_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ),
    .B(_1782_),
    .X(_1783_));
 sky130_fd_sc_hd__mux2_1 _2992_ (.A0(_1616_),
    .A1(_0796_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ),
    .X(_1784_));
 sky130_fd_sc_hd__a21bo_1 _2993_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ),
    .A2(_1784_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q ),
    .X(_1785_));
 sky130_fd_sc_hd__mux4_1 _2994_ (.A0(_0279_),
    .A1(net94),
    .A2(net2),
    .A3(net1055),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ),
    .X(_1786_));
 sky130_fd_sc_hd__o22a_1 _2995_ (.A1(_1785_),
    .A2(_1783_),
    .B1(_1786_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _2996_ (.A0(net637),
    .A1(net59),
    .A2(net1264),
    .A3(net1034),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ),
    .X(_1787_));
 sky130_fd_sc_hd__mux4_1 _2997_ (.A0(net1047),
    .A1(_0756_),
    .A2(_0788_),
    .A3(_0293_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ),
    .X(_1788_));
 sky130_fd_sc_hd__mux2_1 _2998_ (.A0(_1787_),
    .A1(_1788_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 ));
 sky130_fd_sc_hd__nor2_1 _2999_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ),
    .B(net1030),
    .Y(_1789_));
 sky130_fd_sc_hd__a211oi_1 _3000_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ),
    .A2(_0571_),
    .B1(_1789_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ),
    .Y(_1790_));
 sky130_fd_sc_hd__mux2_4 _3001_ (.A0(_0700_),
    .A1(_1238_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ),
    .X(_1791_));
 sky130_fd_sc_hd__a21bo_1 _3002_ (.A1(_1791_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q ),
    .X(_1792_));
 sky130_fd_sc_hd__mux4_1 _3003_ (.A0(_0414_),
    .A1(net1263),
    .A2(net60),
    .A3(net984),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ),
    .X(_1793_));
 sky130_fd_sc_hd__o22a_1 _3004_ (.A1(_1790_),
    .A2(_1792_),
    .B1(_1793_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 ));
 sky130_fd_sc_hd__or2_1 _3005_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ),
    .B(net626),
    .X(_1794_));
 sky130_fd_sc_hd__a21oi_1 _3006_ (.A1(_0027_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ),
    .Y(_1795_));
 sky130_fd_sc_hd__mux2_1 _3007_ (.A0(net57),
    .A1(net1043),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_1796_));
 sky130_fd_sc_hd__a221o_1 _3008_ (.A1(_1794_),
    .A2(_1795_),
    .B1(_1796_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q ),
    .X(_1797_));
 sky130_fd_sc_hd__mux4_1 _3009_ (.A0(net1015),
    .A1(net968),
    .A2(_1204_),
    .A3(_0471_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_1798_));
 sky130_fd_sc_hd__o21a_1 _3010_ (.A1(_0180_),
    .A2(_1798_),
    .B1(_1797_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 ));
 sky130_fd_sc_hd__mux2_4 _3011_ (.A0(net1057),
    .A1(net648),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_1799_));
 sky130_fd_sc_hd__and2b_1 _3012_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ),
    .B(_1799_),
    .X(_1800_));
 sky130_fd_sc_hd__mux2_4 _3013_ (.A0(_1616_),
    .A1(_0764_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_1801_));
 sky130_fd_sc_hd__a21bo_1 _3014_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ),
    .A2(_1801_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q ),
    .X(_1802_));
 sky130_fd_sc_hd__mux4_1 _3015_ (.A0(_0279_),
    .A1(net58),
    .A2(net2),
    .A3(net1055),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_1803_));
 sky130_fd_sc_hd__o22a_1 _3016_ (.A1(_1802_),
    .A2(_1800_),
    .B1(_1803_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _3017_ (.A0(net1263),
    .A1(net96),
    .A2(net1019),
    .A3(net1038),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_1804_));
 sky130_fd_sc_hd__or2_1 _3018_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ),
    .B(_1804_),
    .X(_1805_));
 sky130_fd_sc_hd__mux4_1 _3019_ (.A0(net1034),
    .A1(net984),
    .A2(net1043),
    .A3(net1055),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_1806_));
 sky130_fd_sc_hd__inv_1 _3020_ (.A(_1806_),
    .Y(_1807_));
 sky130_fd_sc_hd__a21oi_1 _3021_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(_1807_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q ),
    .Y(_1808_));
 sky130_fd_sc_hd__mux2_1 _3022_ (.A0(_1204_),
    .A1(net968),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_1809_));
 sky130_fd_sc_hd__mux2_1 _3023_ (.A0(_0788_),
    .A1(_0756_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_1810_));
 sky130_fd_sc_hd__mux2_4 _3024_ (.A0(_1810_),
    .A1(_1809_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_1811_));
 sky130_fd_sc_hd__mux4_1 _3025_ (.A0(net1047),
    .A1(net1030),
    .A2(net1015),
    .A3(net1057),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_1812_));
 sky130_fd_sc_hd__mux2_2 _3026_ (.A0(_1812_),
    .A1(_1811_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ),
    .X(_1813_));
 sky130_fd_sc_hd__a22o_1 _3027_ (.A1(_1805_),
    .A2(_1808_),
    .B1(_1813_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 ));
 sky130_fd_sc_hd__mux4_1 _3028_ (.A0(net1264),
    .A1(net1019),
    .A2(net1226),
    .A3(net1038),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .X(_1814_));
 sky130_fd_sc_hd__mux4_1 _3029_ (.A0(net1034),
    .A1(net984),
    .A2(net1043),
    .A3(net1055),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_1815_));
 sky130_fd_sc_hd__mux2_1 _3030_ (.A0(_1814_),
    .A1(_1815_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ),
    .X(_1816_));
 sky130_fd_sc_hd__mux2_1 _3031_ (.A0(_0571_),
    .A1(_0701_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .X(_1817_));
 sky130_fd_sc_hd__mux2_1 _3032_ (.A0(net648),
    .A1(_1616_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .X(_1818_));
 sky130_fd_sc_hd__nand2_2 _3033_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .B(_1818_),
    .Y(_1819_));
 sky130_fd_sc_hd__o211a_1 _3034_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .A2(_1817_),
    .B1(_1819_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ),
    .X(_1820_));
 sky130_fd_sc_hd__mux4_1 _3035_ (.A0(net1047),
    .A1(net1030),
    .A2(net1014),
    .A3(net1057),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_1821_));
 sky130_fd_sc_hd__o21ba_1 _3036_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_1821_),
    .B1_N(_1820_),
    .X(_1822_));
 sky130_fd_sc_hd__mux2_2 _3037_ (.A0(_1816_),
    .A1(_1822_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 ));
 sky130_fd_sc_hd__mux4_1 _3038_ (.A0(net1049),
    .A1(_0756_),
    .A2(_0788_),
    .A3(_1628_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ),
    .X(_1823_));
 sky130_fd_sc_hd__mux4_1 _3039_ (.A0(net637),
    .A1(net1264),
    .A2(net95),
    .A3(net1035),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q ),
    .X(_1824_));
 sky130_fd_sc_hd__mux2_1 _3040_ (.A0(_1824_),
    .A1(_1823_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 ));
 sky130_fd_sc_hd__mux2_4 _3041_ (.A0(_0700_),
    .A1(_1195_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ),
    .X(_1825_));
 sky130_fd_sc_hd__nor2_1 _3042_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ),
    .B(net1027),
    .Y(_1826_));
 sky130_fd_sc_hd__a211oi_1 _3043_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ),
    .A2(_0571_),
    .B1(_1826_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ),
    .Y(_1827_));
 sky130_fd_sc_hd__a21bo_1 _3044_ (.A1(_1825_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q ),
    .X(_1828_));
 sky130_fd_sc_hd__mux4_1 _3045_ (.A0(net920),
    .A1(net1225),
    .A2(net4),
    .A3(net986),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ),
    .X(_1829_));
 sky130_fd_sc_hd__o22a_1 _3046_ (.A1(_1827_),
    .A2(_1828_),
    .B1(_1829_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 ));
 sky130_fd_sc_hd__or2_1 _3047_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .B(_0239_),
    .X(_1830_));
 sky130_fd_sc_hd__a21oi_1 _3048_ (.A1(_0027_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ),
    .Y(_1831_));
 sky130_fd_sc_hd__mux2_1 _3049_ (.A0(net93),
    .A1(net1044),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .X(_1832_));
 sky130_fd_sc_hd__a221o_1 _3050_ (.A1(_1830_),
    .A2(_1831_),
    .B1(_1832_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q ),
    .X(_1833_));
 sky130_fd_sc_hd__mux2_1 _3051_ (.A0(net669),
    .A1(_1204_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .X(_1834_));
 sky130_fd_sc_hd__mux2_1 _3052_ (.A0(net968),
    .A1(_0659_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .X(_1835_));
 sky130_fd_sc_hd__mux2_1 _3053_ (.A0(_1834_),
    .A1(_1835_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ),
    .X(_1836_));
 sky130_fd_sc_hd__o21a_1 _3054_ (.A1(_0181_),
    .A2(_1836_),
    .B1(_1833_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 ));
 sky130_fd_sc_hd__mux2_4 _3055_ (.A0(net1057),
    .A1(net649),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ),
    .X(_1837_));
 sky130_fd_sc_hd__and2b_1 _3056_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ),
    .B(_1837_),
    .X(_1838_));
 sky130_fd_sc_hd__mux2_1 _3057_ (.A0(_1616_),
    .A1(_0518_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ),
    .X(_1839_));
 sky130_fd_sc_hd__a21bo_1 _3058_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ),
    .A2(_1839_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q ),
    .X(_1840_));
 sky130_fd_sc_hd__mux4_1 _3059_ (.A0(_0279_),
    .A1(net94),
    .A2(net2),
    .A3(net1055),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ),
    .X(_1841_));
 sky130_fd_sc_hd__o22a_1 _3060_ (.A1(_1838_),
    .A2(_1840_),
    .B1(_1841_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _3061_ (.A0(net1049),
    .A1(_0756_),
    .A2(_0788_),
    .A3(_1610_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ),
    .X(_1842_));
 sky130_fd_sc_hd__mux4_1 _3062_ (.A0(net637),
    .A1(net59),
    .A2(net1226),
    .A3(net1034),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ),
    .X(_1843_));
 sky130_fd_sc_hd__mux2_1 _3063_ (.A0(_1843_),
    .A1(_1842_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 ));
 sky130_fd_sc_hd__nor2_1 _3064_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ),
    .B(net1028),
    .Y(_1844_));
 sky130_fd_sc_hd__a211oi_1 _3065_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ),
    .A2(_0571_),
    .B1(_1844_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ),
    .Y(_1845_));
 sky130_fd_sc_hd__mux2_4 _3066_ (.A0(_0700_),
    .A1(_1535_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ),
    .X(_1846_));
 sky130_fd_sc_hd__a21bo_1 _3067_ (.A1(_1846_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q ),
    .X(_1847_));
 sky130_fd_sc_hd__mux4_1 _3068_ (.A0(net920),
    .A1(net1225),
    .A2(net60),
    .A3(net983),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ),
    .X(_1848_));
 sky130_fd_sc_hd__o22a_4 _3069_ (.A1(_1845_),
    .A2(_1847_),
    .B1(_1848_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 ));
 sky130_fd_sc_hd__or2_1 _3070_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .B(net626),
    .X(_1849_));
 sky130_fd_sc_hd__a21oi_1 _3071_ (.A1(_0041_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ),
    .Y(_1850_));
 sky130_fd_sc_hd__mux2_1 _3072_ (.A0(net93),
    .A1(net1044),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_1851_));
 sky130_fd_sc_hd__a221o_1 _3073_ (.A1(_1849_),
    .A2(_1850_),
    .B1(_1851_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q ),
    .X(_1852_));
 sky130_fd_sc_hd__mux2_1 _3074_ (.A0(net669),
    .A1(_1204_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_1853_));
 sky130_fd_sc_hd__mux2_1 _3075_ (.A0(net641),
    .A1(_0683_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_1854_));
 sky130_fd_sc_hd__mux2_2 _3076_ (.A0(_1853_),
    .A1(_1854_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ),
    .X(_1855_));
 sky130_fd_sc_hd__o21a_1 _3077_ (.A1(_0182_),
    .A2(_1855_),
    .B1(_1852_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 ));
 sky130_fd_sc_hd__mux2_1 _3078_ (.A0(net822),
    .A1(net647),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ),
    .X(_1856_));
 sky130_fd_sc_hd__and2b_1 _3079_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ),
    .B(_1856_),
    .X(_1857_));
 sky130_fd_sc_hd__mux2_4 _3080_ (.A0(_1616_),
    .A1(_0528_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ),
    .X(_1858_));
 sky130_fd_sc_hd__a21bo_1 _3081_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ),
    .A2(_1858_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q ),
    .X(_1859_));
 sky130_fd_sc_hd__mux4_1 _3082_ (.A0(_0279_),
    .A1(net94),
    .A2(net58),
    .A3(net1051),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ),
    .X(_1860_));
 sky130_fd_sc_hd__o22a_1 _3083_ (.A1(_1859_),
    .A2(_1857_),
    .B1(_1860_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _3084_ (.A0(net1263),
    .A1(net1225),
    .A2(net815),
    .A3(net1039),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .X(_1861_));
 sky130_fd_sc_hd__or2_1 _3085_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ),
    .B(_1861_),
    .X(_1862_));
 sky130_fd_sc_hd__mux4_1 _3086_ (.A0(net1033),
    .A1(net983),
    .A2(net1042),
    .A3(net1053),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .X(_1863_));
 sky130_fd_sc_hd__inv_1 _3087_ (.A(_1863_),
    .Y(_1864_));
 sky130_fd_sc_hd__a21oi_1 _3088_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_1864_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q ),
    .Y(_1865_));
 sky130_fd_sc_hd__mux4_2 _3089_ (.A0(_0788_),
    .A1(_1204_),
    .A2(_0756_),
    .A3(net968),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_1866_));
 sky130_fd_sc_hd__mux4_1 _3090_ (.A0(net1048),
    .A1(net1028),
    .A2(net1014),
    .A3(net822),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .X(_1867_));
 sky130_fd_sc_hd__mux2_4 _3091_ (.A0(_1867_),
    .A1(_1866_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ),
    .X(_1868_));
 sky130_fd_sc_hd__a22o_1 _3092_ (.A1(_1862_),
    .A2(_1865_),
    .B1(_1868_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 ));
 sky130_fd_sc_hd__mux2_1 _3093_ (.A0(_0571_),
    .A1(_0701_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_1869_));
 sky130_fd_sc_hd__mux2_1 _3094_ (.A0(net648),
    .A1(_1616_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_1870_));
 sky130_fd_sc_hd__nand2_1 _3095_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .B(_1870_),
    .Y(_1871_));
 sky130_fd_sc_hd__o211a_1 _3096_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .A2(_1869_),
    .B1(_1871_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ),
    .X(_1872_));
 sky130_fd_sc_hd__mux4_1 _3097_ (.A0(net1048),
    .A1(net1028),
    .A2(net1014),
    .A3(net1058),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .X(_1873_));
 sky130_fd_sc_hd__o21ba_1 _3098_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_1873_),
    .B1_N(_1872_),
    .X(_1874_));
 sky130_fd_sc_hd__mux4_1 _3099_ (.A0(net1264),
    .A1(net1018),
    .A2(net1226),
    .A3(net1039),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_1875_));
 sky130_fd_sc_hd__mux4_1 _3100_ (.A0(net1032),
    .A1(net983),
    .A2(net1042),
    .A3(net1053),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .X(_1876_));
 sky130_fd_sc_hd__mux2_1 _3101_ (.A0(_1875_),
    .A1(_1876_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ),
    .X(_1877_));
 sky130_fd_sc_hd__mux2_2 _3102_ (.A0(_1877_),
    .A1(_1874_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 ));
 sky130_fd_sc_hd__mux2_1 _3103_ (.A0(_0494_),
    .A1(_0428_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q ),
    .X(_1878_));
 sky130_fd_sc_hd__inv_1 _3104_ (.A(_1878_),
    .Y(_1879_));
 sky130_fd_sc_hd__mux2_1 _3105_ (.A0(net866),
    .A1(net670),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q ),
    .X(_1880_));
 sky130_fd_sc_hd__mux2_1 _3106_ (.A0(_1880_),
    .A1(_1879_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _3107_ (.A0(net180),
    .A1(net1221),
    .A2(net195),
    .A3(net989),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q ),
    .X(\Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A ));
 sky130_fd_sc_hd__mux4_1 _3108_ (.A0(net181),
    .A1(net1222),
    .A2(net196),
    .A3(net993),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q ),
    .X(\Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A ));
 sky130_fd_sc_hd__mux4_1 _3109_ (.A0(net178),
    .A1(net197),
    .A2(net231),
    .A3(net1023),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q ),
    .X(\Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A ));
 sky130_fd_sc_hd__mux4_1 _3110_ (.A0(net179),
    .A1(net194),
    .A2(net230),
    .A3(net1004),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q ),
    .X(\Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A ));
 sky130_fd_sc_hd__mux4_1 _3111_ (.A0(net1000),
    .A1(_0214_),
    .A2(net619),
    .A3(_0228_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 ));
 sky130_fd_sc_hd__o21ai_1 _3112_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q ),
    .Y(_1881_));
 sky130_fd_sc_hd__a21o_1 _3113_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q ),
    .A2(net661),
    .B1(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__nor2_1 _3114_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q ),
    .B(net991),
    .Y(_1883_));
 sky130_fd_sc_hd__a211o_1 _3115_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q ),
    .A2(_0257_),
    .B1(_1883_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q ),
    .X(_1884_));
 sky130_fd_sc_hd__nand2_1 _3116_ (.A(_1882_),
    .B(_1884_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 ));
 sky130_fd_sc_hd__mux4_1 _3117_ (.A0(net995),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .A2(net666),
    .A3(_1378_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _3118_ (.A0(net1025),
    .A1(net918),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .A3(_0405_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _3119_ (.A0(net987),
    .A1(_0214_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .A3(_0228_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _3120_ (.A0(net869),
    .A1(net664),
    .A2(net830),
    .A3(net988),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_1885_));
 sky130_fd_sc_hd__or2_1 _3121_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ),
    .B(_1885_),
    .X(_1886_));
 sky130_fd_sc_hd__mux4_1 _3122_ (.A0(net993),
    .A1(net1022),
    .A2(net1003),
    .A3(net1007),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_1887_));
 sky130_fd_sc_hd__o21a_1 _3123_ (.A1(_0183_),
    .A2(_1887_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q ),
    .X(_1888_));
 sky130_fd_sc_hd__mux4_1 _3124_ (.A0(net1221),
    .A1(net215),
    .A2(net70),
    .A3(net231),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_1889_));
 sky130_fd_sc_hd__mux4_1 _3125_ (.A0(net177),
    .A1(net179),
    .A2(net195),
    .A3(net142),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_1890_));
 sky130_fd_sc_hd__mux2_1 _3126_ (.A0(_1889_),
    .A1(_1890_),
    .S(_0183_),
    .X(_1891_));
 sky130_fd_sc_hd__a22o_1 _3127_ (.A1(_1886_),
    .A2(_1888_),
    .B1(_1891_),
    .B2(_0184_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 ));
 sky130_fd_sc_hd__o21ai_1 _3128_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q ),
    .Y(_1892_));
 sky130_fd_sc_hd__a21o_1 _3129_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(net662),
    .B1(_1892_),
    .X(_1893_));
 sky130_fd_sc_hd__nor2_1 _3130_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q ),
    .B(net992),
    .Y(_1894_));
 sky130_fd_sc_hd__a211o_1 _3131_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(net833),
    .B1(_1894_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q ),
    .X(_1895_));
 sky130_fd_sc_hd__nand2_1 _3132_ (.A(_1893_),
    .B(_1895_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 ));
 sky130_fd_sc_hd__mux2_1 _3133_ (.A0(net1022),
    .A1(net666),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q ),
    .X(_1896_));
 sky130_fd_sc_hd__mux2_1 _3134_ (.A0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ),
    .A1(_1378_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q ),
    .X(_1897_));
 sky130_fd_sc_hd__mux2_1 _3135_ (.A0(_1896_),
    .A1(_1897_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _3136_ (.A0(net1003),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ),
    .A2(_0413_),
    .A3(_0405_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _3137_ (.A0(net1221),
    .A1(net82),
    .A2(net71),
    .A3(net921),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _3138_ (.A0(net139),
    .A1(net72),
    .A2(net83),
    .A3(net971),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _3139_ (.A0(net69),
    .A1(net84),
    .A2(net231),
    .A3(net980),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _3140_ (.A0(net70),
    .A1(net81),
    .A2(net230),
    .A3(net1000),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _3141_ (.A0(net993),
    .A1(_0214_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .A3(_0228_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _3142_ (.A0(net869),
    .A1(net664),
    .A2(net830),
    .A3(net987),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_1898_));
 sky130_fd_sc_hd__or2_1 _3143_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .B(_1898_),
    .X(_1899_));
 sky130_fd_sc_hd__mux4_1 _3144_ (.A0(net992),
    .A1(net1021),
    .A2(net1002),
    .A3(net1010),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_1900_));
 sky130_fd_sc_hd__o21a_1 _3145_ (.A1(_0185_),
    .A2(_1900_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q ),
    .X(_1901_));
 sky130_fd_sc_hd__mux4_1 _3146_ (.A0(net70),
    .A1(net82),
    .A2(net215),
    .A3(net231),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_1902_));
 sky130_fd_sc_hd__mux4_1 _3147_ (.A0(net203),
    .A1(net1223),
    .A2(net124),
    .A3(net1221),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_1903_));
 sky130_fd_sc_hd__mux2_1 _3148_ (.A0(_1902_),
    .A1(_1903_),
    .S(_0185_),
    .X(_1904_));
 sky130_fd_sc_hd__a22o_1 _3149_ (.A1(_1899_),
    .A2(_1901_),
    .B1(_1904_),
    .B2(_0186_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 ));
 sky130_fd_sc_hd__o21ai_1 _3150_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q ),
    .Y(_1905_));
 sky130_fd_sc_hd__a21o_1 _3151_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q ),
    .A2(net662),
    .B1(_1905_),
    .X(_1906_));
 sky130_fd_sc_hd__nor2_1 _3152_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q ),
    .B(net1021),
    .Y(_1907_));
 sky130_fd_sc_hd__a211o_1 _3153_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q ),
    .A2(net833),
    .B1(_1907_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q ),
    .X(_1908_));
 sky130_fd_sc_hd__nand2_1 _3154_ (.A(_1906_),
    .B(_1908_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 ));
 sky130_fd_sc_hd__mux2_1 _3155_ (.A0(net1002),
    .A1(net666),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q ),
    .X(_1909_));
 sky130_fd_sc_hd__mux2_1 _3156_ (.A0(net665),
    .A1(_1378_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q ),
    .X(_1910_));
 sky130_fd_sc_hd__mux2_1 _3157_ (.A0(_1909_),
    .A1(_1910_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _3158_ (.A0(net975),
    .A1(net816),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ),
    .A3(_0405_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _3159_ (.A0(net176),
    .A1(net1224),
    .A2(net1073),
    .A3(net980),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ),
    .X(_1911_));
 sky130_fd_sc_hd__mux4_1 _3160_ (.A0(net1025),
    .A1(_0823_),
    .A2(_0977_),
    .A3(_1416_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ),
    .X(_1912_));
 sky130_fd_sc_hd__mux2_1 _3161_ (.A0(_1911_),
    .A1(_1912_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q ),
    .X(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A ));
 sky130_fd_sc_hd__mux4_1 _3162_ (.A0(net177),
    .A1(net1223),
    .A2(net1072),
    .A3(net830),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q ),
    .X(_1913_));
 sky130_fd_sc_hd__mux2_1 _3163_ (.A0(_0875_),
    .A1(_1489_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ),
    .X(_1914_));
 sky130_fd_sc_hd__mux2_1 _3164_ (.A0(net1006),
    .A1(_0712_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ),
    .X(_1915_));
 sky130_fd_sc_hd__mux2_1 _3165_ (.A0(_1915_),
    .A1(_1914_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q ),
    .X(_1916_));
 sky130_fd_sc_hd__mux2_1 _3166_ (.A0(_1913_),
    .A1(_1916_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q ),
    .X(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A ));
 sky130_fd_sc_hd__mux4_1 _3167_ (.A0(net1011),
    .A1(net1013),
    .A2(_1497_),
    .A3(_0960_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ),
    .X(_1917_));
 sky130_fd_sc_hd__mux4_1 _3168_ (.A0(net174),
    .A1(net119),
    .A2(net210),
    .A3(net990),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q ),
    .X(_1918_));
 sky130_fd_sc_hd__mux2_1 _3169_ (.A0(_1918_),
    .A1(_1917_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q ),
    .X(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A ));
 sky130_fd_sc_hd__mux4_1 _3170_ (.A0(net175),
    .A1(net211),
    .A2(net120),
    .A3(net996),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q ),
    .X(_1919_));
 sky130_fd_sc_hd__mux4_2 _3171_ (.A0(net1007),
    .A1(_1400_),
    .A2(_1473_),
    .A3(_0841_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q ),
    .X(_1920_));
 sky130_fd_sc_hd__mux2_1 _3172_ (.A0(_1919_),
    .A1(_1920_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q ),
    .X(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A ));
 sky130_fd_sc_hd__nand2b_1 _3173_ (.A_N(net980),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .Y(_1921_));
 sky130_fd_sc_hd__o211a_1 _3174_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .A2(_0344_),
    .B1(_1921_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ),
    .X(_1922_));
 sky130_fd_sc_hd__mux2_1 _3175_ (.A0(net176),
    .A1(net121),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .X(_1923_));
 sky130_fd_sc_hd__a21o_1 _3176_ (.A1(_0187_),
    .A2(_1923_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q ),
    .X(_1924_));
 sky130_fd_sc_hd__mux2_1 _3177_ (.A0(_0977_),
    .A1(_1436_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .X(_1925_));
 sky130_fd_sc_hd__mux2_1 _3178_ (.A0(net1025),
    .A1(_0823_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .X(_1926_));
 sky130_fd_sc_hd__mux2_1 _3179_ (.A0(_1925_),
    .A1(_1926_),
    .S(_0187_),
    .X(_1927_));
 sky130_fd_sc_hd__o22a_1 _3180_ (.A1(_1922_),
    .A2(_1924_),
    .B1(_1927_),
    .B2(_0188_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _3181_ (.A0(net177),
    .A1(net1223),
    .A2(_0387_),
    .A3(net1000),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ),
    .X(_1928_));
 sky130_fd_sc_hd__mux2_1 _3182_ (.A0(_0875_),
    .A1(_1510_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ),
    .X(_1929_));
 sky130_fd_sc_hd__nand2_1 _3183_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ),
    .B(_0711_),
    .Y(_1930_));
 sky130_fd_sc_hd__o21ba_1 _3184_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ),
    .A2(net1005),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ),
    .X(_1931_));
 sky130_fd_sc_hd__a221o_1 _3185_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ),
    .A2(_1929_),
    .B1(_1930_),
    .B2(_1931_),
    .C1(_0189_),
    .X(_1932_));
 sky130_fd_sc_hd__o21a_1 _3186_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q ),
    .A2(_1928_),
    .B1(_1932_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 ));
 sky130_fd_sc_hd__mux2_1 _3187_ (.A0(_0442_),
    .A1(net991),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .X(_1933_));
 sky130_fd_sc_hd__mux2_1 _3188_ (.A0(net174),
    .A1(net119),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .X(_1934_));
 sky130_fd_sc_hd__and2b_1 _3189_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ),
    .B(_1934_),
    .X(_1935_));
 sky130_fd_sc_hd__a211o_1 _3190_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ),
    .A2(_1933_),
    .B1(_1935_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q ),
    .X(_1936_));
 sky130_fd_sc_hd__mux4_1 _3191_ (.A0(net812),
    .A1(net666),
    .A2(_1497_),
    .A3(_1019_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .X(_1937_));
 sky130_fd_sc_hd__o21a_1 _3192_ (.A1(_0190_),
    .A2(_1937_),
    .B1(_1936_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 ));
 sky130_fd_sc_hd__nand2b_1 _3193_ (.A_N(_0906_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ),
    .Y(_1938_));
 sky130_fd_sc_hd__o211a_1 _3194_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ),
    .A2(_1400_),
    .B1(_1938_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_1939_));
 sky130_fd_sc_hd__nor2_1 _3195_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ),
    .B(net653),
    .Y(_1940_));
 sky130_fd_sc_hd__a211o_1 _3196_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ),
    .A2(net634),
    .B1(_1940_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_1941_));
 sky130_fd_sc_hd__nand2_1 _3197_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q ),
    .B(_1941_),
    .Y(_1942_));
 sky130_fd_sc_hd__mux4_2 _3198_ (.A0(net175),
    .A1(net120),
    .A2(_0563_),
    .A3(net995),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_1943_));
 sky130_fd_sc_hd__o22a_4 _3199_ (.A1(_1939_),
    .A2(_1942_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q ),
    .B2(_1943_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _3200_ (.A0(_0823_),
    .A1(_0977_),
    .A2(_1497_),
    .A3(net1013),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_1944_));
 sky130_fd_sc_hd__mux4_1 _3201_ (.A0(net1025),
    .A1(net1005),
    .A2(net812),
    .A3(net1009),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_1945_));
 sky130_fd_sc_hd__mux2_1 _3202_ (.A0(_1945_),
    .A1(_1944_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ),
    .X(_1946_));
 sky130_fd_sc_hd__mux4_1 _3203_ (.A0(net1223),
    .A1(net1072),
    .A2(net655),
    .A3(net971),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_1947_));
 sky130_fd_sc_hd__or2_1 _3204_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ),
    .B(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__mux4_1 _3205_ (.A0(net980),
    .A1(net656),
    .A2(net1000),
    .A3(net995),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .X(_1949_));
 sky130_fd_sc_hd__inv_1 _3206_ (.A(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__a21oi_1 _3207_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ),
    .A2(_1950_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q ),
    .Y(_1951_));
 sky130_fd_sc_hd__a22o_1 _3208_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q ),
    .A2(_1946_),
    .B1(_1948_),
    .B2(_1951_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 ));
 sky130_fd_sc_hd__mux4_1 _3209_ (.A0(net1224),
    .A1(net212),
    .A2(net924),
    .A3(net971),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_1952_));
 sky130_fd_sc_hd__mux4_1 _3210_ (.A0(net980),
    .A1(net656),
    .A2(net1000),
    .A3(net995),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_1953_));
 sky130_fd_sc_hd__mux2_1 _3211_ (.A0(_1952_),
    .A1(_1953_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ),
    .X(_1954_));
 sky130_fd_sc_hd__mux2_1 _3212_ (.A0(_1473_),
    .A1(_1400_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_1955_));
 sky130_fd_sc_hd__mux2_2 _3213_ (.A0(_0712_),
    .A1(_0875_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_1956_));
 sky130_fd_sc_hd__and2b_1 _3214_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .B(_1956_),
    .X(_1957_));
 sky130_fd_sc_hd__a21bo_1 _3215_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .A2(_1955_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ),
    .X(_1958_));
 sky130_fd_sc_hd__mux4_1 _3216_ (.A0(net1025),
    .A1(net1005),
    .A2(net812),
    .A3(net1009),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_1959_));
 sky130_fd_sc_hd__o22a_1 _3217_ (.A1(_1957_),
    .A2(_1958_),
    .B1(_1959_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ),
    .X(_1960_));
 sky130_fd_sc_hd__mux2_1 _3218_ (.A0(_1954_),
    .A1(_1960_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 ));
 sky130_fd_sc_hd__mux4_1 _3219_ (.A0(net176),
    .A1(net1224),
    .A2(net1073),
    .A3(net980),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ),
    .X(_1961_));
 sky130_fd_sc_hd__mux2_1 _3220_ (.A0(_0977_),
    .A1(_1380_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ),
    .X(_1962_));
 sky130_fd_sc_hd__mux2_1 _3221_ (.A0(net1025),
    .A1(_0823_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ),
    .X(_1963_));
 sky130_fd_sc_hd__mux2_1 _3222_ (.A0(_1963_),
    .A1(_1962_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ),
    .X(_1964_));
 sky130_fd_sc_hd__mux2_1 _3223_ (.A0(_1961_),
    .A1(_1964_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 ));
 sky130_fd_sc_hd__mux2_1 _3224_ (.A0(net1005),
    .A1(_0712_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ),
    .X(_1965_));
 sky130_fd_sc_hd__mux2_1 _3225_ (.A0(_0875_),
    .A1(_1454_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ),
    .X(_1966_));
 sky130_fd_sc_hd__mux2_1 _3226_ (.A0(_1965_),
    .A1(_1966_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ),
    .X(_1967_));
 sky130_fd_sc_hd__mux2_1 _3227_ (.A0(net177),
    .A1(net1223),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ),
    .X(_1968_));
 sky130_fd_sc_hd__and2b_1 _3228_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ),
    .B(_1968_),
    .X(_1969_));
 sky130_fd_sc_hd__mux2_1 _3229_ (.A0(net213),
    .A1(net1000),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ),
    .X(_1970_));
 sky130_fd_sc_hd__a211o_1 _3230_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ),
    .A2(_1970_),
    .B1(_1969_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q ),
    .X(_1971_));
 sky130_fd_sc_hd__o21a_1 _3231_ (.A1(_0191_),
    .A2(_1967_),
    .B1(_1971_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _3232_ (.A0(net812),
    .A1(net1013),
    .A2(_1497_),
    .A3(_0609_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ),
    .X(_1972_));
 sky130_fd_sc_hd__mux4_1 _3233_ (.A0(net174),
    .A1(net119),
    .A2(net210),
    .A3(net656),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ),
    .X(_1973_));
 sky130_fd_sc_hd__mux2_1 _3234_ (.A0(_1973_),
    .A1(_1972_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _3235_ (.A0(net175),
    .A1(net211),
    .A2(net120),
    .A3(net995),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ),
    .X(_1974_));
 sky130_fd_sc_hd__mux2_2 _3236_ (.A0(_1400_),
    .A1(_0637_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ),
    .X(_1975_));
 sky130_fd_sc_hd__nor2_1 _3237_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ),
    .B(net653),
    .Y(_1976_));
 sky130_fd_sc_hd__a211o_1 _3238_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ),
    .A2(net633),
    .B1(_1976_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ),
    .X(_1977_));
 sky130_fd_sc_hd__a21bo_1 _3239_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ),
    .A2(_1975_),
    .B1_N(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__mux2_2 _3240_ (.A0(_1974_),
    .A1(_1978_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 ));
 sky130_fd_sc_hd__nor2_1 _3241_ (.A(net176),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ),
    .Y(_1979_));
 sky130_fd_sc_hd__a211o_1 _3242_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ),
    .A2(net631),
    .B1(_1979_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ),
    .X(_1980_));
 sky130_fd_sc_hd__mux2_2 _3243_ (.A0(net1073),
    .A1(net979),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ),
    .X(_1981_));
 sky130_fd_sc_hd__a21oi_2 _3244_ (.A1(_1981_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q ),
    .Y(_1982_));
 sky130_fd_sc_hd__mux2_1 _3245_ (.A0(net1024),
    .A1(_0823_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ),
    .X(_1983_));
 sky130_fd_sc_hd__mux2_1 _3246_ (.A0(_0977_),
    .A1(_1398_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ),
    .X(_1984_));
 sky130_fd_sc_hd__mux2_1 _3247_ (.A0(_1983_),
    .A1(_1984_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ),
    .X(_1985_));
 sky130_fd_sc_hd__o2bb2a_4 _3248_ (.A1_N(_1982_),
    .A2_N(_1980_),
    .B1(_1985_),
    .B2(_0192_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _3249_ (.A0(net177),
    .A1(net1072),
    .A2(_0387_),
    .A3(net830),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ),
    .X(_1986_));
 sky130_fd_sc_hd__mux2_1 _3250_ (.A0(_0875_),
    .A1(_1466_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ),
    .X(_1987_));
 sky130_fd_sc_hd__nand2_1 _3251_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ),
    .B(_0711_),
    .Y(_1988_));
 sky130_fd_sc_hd__o21ba_1 _3252_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ),
    .A2(net1003),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ),
    .X(_1989_));
 sky130_fd_sc_hd__a221o_1 _3253_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ),
    .A2(_1987_),
    .B1(_1988_),
    .B2(_1989_),
    .C1(_0193_),
    .X(_1990_));
 sky130_fd_sc_hd__o21a_1 _3254_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q ),
    .A2(_1986_),
    .B1(_1990_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 ));
 sky130_fd_sc_hd__mux2_1 _3255_ (.A0(net174),
    .A1(_0442_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ),
    .X(_1991_));
 sky130_fd_sc_hd__and2b_1 _3256_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ),
    .B(_1991_),
    .X(_1992_));
 sky130_fd_sc_hd__mux2_1 _3257_ (.A0(net210),
    .A1(net989),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ),
    .X(_1993_));
 sky130_fd_sc_hd__a21o_1 _3258_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ),
    .A2(_1993_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q ),
    .X(_1994_));
 sky130_fd_sc_hd__mux2_1 _3259_ (.A0(net1011),
    .A1(_1497_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ),
    .X(_1995_));
 sky130_fd_sc_hd__mux2_1 _3260_ (.A0(net666),
    .A1(_0864_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ),
    .X(_1996_));
 sky130_fd_sc_hd__mux2_1 _3261_ (.A0(_1995_),
    .A1(_1996_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ),
    .X(_1997_));
 sky130_fd_sc_hd__o22a_1 _3262_ (.A1(_1992_),
    .A2(_1994_),
    .B1(_1997_),
    .B2(_0194_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 ));
 sky130_fd_sc_hd__mux4_2 _3263_ (.A0(net175),
    .A1(net211),
    .A2(_0563_),
    .A3(net864),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ),
    .X(_1998_));
 sky130_fd_sc_hd__mux2_4 _3264_ (.A0(_1400_),
    .A1(_0721_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ),
    .X(_1999_));
 sky130_fd_sc_hd__nand2_2 _3265_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ),
    .B(_1472_),
    .Y(_2000_));
 sky130_fd_sc_hd__o21ba_1 _3266_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ),
    .A2(net1007),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_2001_));
 sky130_fd_sc_hd__a221o_1 _3267_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ),
    .A2(_1999_),
    .B1(_2000_),
    .B2(_2001_),
    .C1(_0195_),
    .X(_2002_));
 sky130_fd_sc_hd__o21a_1 _3268_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q ),
    .A2(_1998_),
    .B1(_2002_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _3269_ (.A0(_0823_),
    .A1(_0977_),
    .A2(_1497_),
    .A3(net1013),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .X(_2003_));
 sky130_fd_sc_hd__mux4_1 _3270_ (.A0(net1023),
    .A1(net1004),
    .A2(net1010),
    .A3(net1008),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .X(_2004_));
 sky130_fd_sc_hd__mux2_1 _3271_ (.A0(_2004_),
    .A1(_2003_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ),
    .X(_2005_));
 sky130_fd_sc_hd__mux4_1 _3272_ (.A0(net1223),
    .A1(net1072),
    .A2(net974),
    .A3(net969),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .X(_2006_));
 sky130_fd_sc_hd__or2_1 _3273_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ),
    .B(_2006_),
    .X(_2007_));
 sky130_fd_sc_hd__mux4_1 _3274_ (.A0(net978),
    .A1(net990),
    .A2(net998),
    .A3(net864),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .X(_2008_));
 sky130_fd_sc_hd__inv_1 _3275_ (.A(_2008_),
    .Y(_2009_));
 sky130_fd_sc_hd__a21oi_1 _3276_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ),
    .A2(_2009_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q ),
    .Y(_2010_));
 sky130_fd_sc_hd__a22o_1 _3277_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q ),
    .A2(_2005_),
    .B1(_2007_),
    .B2(_2010_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 ));
 sky130_fd_sc_hd__mux2_1 _3278_ (.A0(_1473_),
    .A1(_1400_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_2011_));
 sky130_fd_sc_hd__mux2_2 _3279_ (.A0(_0712_),
    .A1(_0875_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_2012_));
 sky130_fd_sc_hd__and2b_1 _3280_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .B(_2012_),
    .X(_2013_));
 sky130_fd_sc_hd__a21bo_1 _3281_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .A2(_2011_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .X(_2014_));
 sky130_fd_sc_hd__mux4_1 _3282_ (.A0(net1023),
    .A1(net1004),
    .A2(net1011),
    .A3(net1008),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .X(_2015_));
 sky130_fd_sc_hd__o22a_1 _3283_ (.A1(_2013_),
    .A2(_2014_),
    .B1(_2015_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .X(_2016_));
 sky130_fd_sc_hd__mux4_1 _3284_ (.A0(net1224),
    .A1(net1073),
    .A2(net974),
    .A3(net969),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .X(_2017_));
 sky130_fd_sc_hd__mux4_1 _3285_ (.A0(net978),
    .A1(net990),
    .A2(net998),
    .A3(net994),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_2018_));
 sky130_fd_sc_hd__mux2_1 _3286_ (.A0(_2017_),
    .A1(_2018_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .X(_2019_));
 sky130_fd_sc_hd__mux2_1 _3287_ (.A0(_2019_),
    .A1(_2016_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 ));
 sky130_fd_sc_hd__mux2_4 _3288_ (.A0(net619),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .X(_2020_));
 sky130_fd_sc_hd__nor2_1 _3289_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .Y(_2021_));
 sky130_fd_sc_hd__a21o_1 _3290_ (.A1(net222),
    .A2(_2021_),
    .B1(_0197_),
    .X(_2022_));
 sky130_fd_sc_hd__a31o_1 _3291_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .A2(_0196_),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .B1(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__a21o_1 _3292_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(_2020_),
    .B1(_2023_),
    .X(_2024_));
 sky130_fd_sc_hd__nand2_1 _3293_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .B(_0599_),
    .Y(_2025_));
 sky130_fd_sc_hd__o211a_1 _3294_ (.A1(net137),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .C1(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__a31o_1 _3295_ (.A1(net131),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .A3(_0196_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .X(_2027_));
 sky130_fd_sc_hd__a211o_1 _3296_ (.A1(net192),
    .A2(_2021_),
    .B1(_2026_),
    .C1(_2027_),
    .X(_2028_));
 sky130_fd_sc_hd__and3b_1 _3297_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q ),
    .B(_2028_),
    .C(_2024_),
    .X(_2029_));
 sky130_fd_sc_hd__or2_1 _3298_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ),
    .X(_2030_));
 sky130_fd_sc_hd__a221o_1 _3299_ (.A1(net819),
    .A2(_2021_),
    .B1(_2030_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .C1(_0197_),
    .X(_2031_));
 sky130_fd_sc_hd__mux2_1 _3300_ (.A0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .X(_2032_));
 sky130_fd_sc_hd__a31o_1 _3301_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .A2(_0196_),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .X(_2033_));
 sky130_fd_sc_hd__a21o_1 _3302_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .A2(_2021_),
    .B1(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__a21o_1 _3303_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(_2032_),
    .B1(_2034_),
    .X(_2035_));
 sky130_fd_sc_hd__a31o_4 _3304_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q ),
    .A2(_2031_),
    .A3(_2035_),
    .B1(_2029_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ));
 sky130_fd_sc_hd__and2b_1 _3305_ (.A_N(net928),
    .B(_1557_),
    .X(_0000_));
 sky130_fd_sc_hd__and2b_1 _3306_ (.A_N(net966),
    .B(_1722_),
    .X(_0001_));
 sky130_fd_sc_hd__and2b_1 _3307_ (.A_N(net928),
    .B(_1555_),
    .X(_0002_));
 sky130_fd_sc_hd__and2b_1 _3308_ (.A_N(net966),
    .B(_1560_),
    .X(_0003_));
 sky130_fd_sc_hd__and2b_1 _3309_ (.A_N(net966),
    .B(_1558_),
    .X(_0004_));
 sky130_fd_sc_hd__and2b_1 _3310_ (.A_N(net928),
    .B(_1561_),
    .X(_0005_));
 sky130_fd_sc_hd__and2b_1 _3311_ (.A_N(net928),
    .B(_1562_),
    .X(_0006_));
 sky130_fd_sc_hd__and2b_1 _3312_ (.A_N(net928),
    .B(_1563_),
    .X(_0007_));
 sky130_fd_sc_hd__and2b_1 _3313_ (.A_N(net966),
    .B(_1723_),
    .X(_0008_));
 sky130_fd_sc_hd__and2b_1 _3314_ (.A_N(net966),
    .B(_1564_),
    .X(_0009_));
 sky130_fd_sc_hd__and2b_1 _3315_ (.A_N(net967),
    .B(_1567_),
    .X(_0010_));
 sky130_fd_sc_hd__and2b_1 _3316_ (.A_N(net967),
    .B(_1568_),
    .X(_0011_));
 sky130_fd_sc_hd__and2b_1 _3317_ (.A_N(net967),
    .B(_1569_),
    .X(_0012_));
 sky130_fd_sc_hd__and2b_1 _3318_ (.A_N(net967),
    .B(_1720_),
    .X(_0013_));
 sky130_fd_sc_hd__and2b_1 _3319_ (.A_N(net967),
    .B(_1553_),
    .X(_0014_));
 sky130_fd_sc_hd__and2b_1 _3320_ (.A_N(net967),
    .B(_1603_),
    .X(_0015_));
 sky130_fd_sc_hd__and2b_1 _3321_ (.A_N(net967),
    .B(_1626_),
    .X(_0016_));
 sky130_fd_sc_hd__and2b_1 _3322_ (.A_N(net967),
    .B(_1657_),
    .X(_0017_));
 sky130_fd_sc_hd__and2b_1 _3323_ (.A_N(net967),
    .B(_1721_),
    .X(_0018_));
 sky130_fd_sc_hd__and2b_1 _3324_ (.A_N(net967),
    .B(_1718_),
    .X(_0019_));
 sky130_fd_sc_hd__inv_2 _3325_ (.A(net1222),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _3326_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_1 _3327_ (.A(net190),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_1 _3328_ (.A(net101),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_1 _3329_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q ),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _3330_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_1 _3331_ (.A(net187),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _3332_ (.A(net1),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_1 _3333_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _3334_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q ),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _3335_ (.A(net223),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _3336_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q ),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _3337_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_1 _3338_ (.A(net218),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_1 _3339_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_1 _3340_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q ),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_1 _3341_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q ),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_1 _3342_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _3343_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q ),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _3344_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q ),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_1 _3345_ (.A(net186),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_1 _3346_ (.A(net57),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_1 _3347_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _3348_ (.A(net229),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _3349_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q ),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _3350_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_1 _3351_ (.A(net195),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_1 _3352_ (.A(net90),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _3353_ (.A(net189),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_1 _3354_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _3355_ (.A(net69),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _3356_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _3357_ (.A(net20),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _3358_ (.A(net76),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_1 _3359_ (.A(net191),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _3360_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q ),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _3361_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_1 _3362_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q ),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_1 _3363_ (.A(net199),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_1 _3364_ (.A(net86),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _3365_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _3366_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q ),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_1 _3367_ (.A(net188),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _3368_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_1 _3369_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q ),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_1 _3370_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _3371_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _3372_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _3373_ (.A(net75),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _3374_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .Y(_0069_));
 sky130_fd_sc_hd__clkinv_2 _3375_ (.A(net18),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _3376_ (.A(net74),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _3377_ (.A(net80),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _3378_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_1 _3379_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q ),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_1 _3380_ (.A(net209),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _3381_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_1 _3382_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q ),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_1 _3383_ (.A(net115),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_1 _3384_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_1 _3385_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q ),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _3386_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_1 _3387_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q ),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_1 _3388_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_1 _3389_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q ),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _3390_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_1 _3391_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _3392_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _3393_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _3394_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_1 _3395_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q ),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _3396_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _3397_ (.A(net17),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_1 _3398_ (.A(net109),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_1 _3399_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q ),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _3400_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _3401_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _3402_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _3403_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _3404_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _3405_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q ),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_1 _3406_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_1 _3407_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q ),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_1 _3408_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q ),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _3409_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _3410_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_1 _3411_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q ),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_1 _3412_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q ),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _3413_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q ),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_1 _3414_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q ),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_1 _3415_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q ),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_1 _3416_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q ),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _3417_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _3418_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _3419_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _3420_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_1 _3421_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q ),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _3422_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _3423_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _3424_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _3425_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _3426_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _3427_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_1 _3428_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_1 _3429_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_1 _3430_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q ),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_1 _3431_ (.A(net135),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_1 _3432_ (.A(net226),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_1 _3433_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_1 _3434_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q ),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _3435_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_1 _3436_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_1 _3437_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _3438_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_1 _3439_ (.A(net214),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_1 _3440_ (.A(net202),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_1 _3441_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_1 _3442_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q ),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _3443_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _3444_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_1 _3445_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q ),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _3446_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_1 _3447_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_1 _3448_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _3449_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_1 _3450_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q ),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _3451_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_1 _3452_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _3453_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_1 _3454_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_1 _3455_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q ),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_1 _3456_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _3457_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_1 _3458_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q ),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _3459_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_1 _3460_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q ),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _3461_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_2 _3462_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_1 _3463_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q ),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_1 _3464_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q ),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_2 _3465_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_1 _3466_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q ),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_1 _3467_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_1 _3468_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q ),
    .Y(_0163_));
 sky130_fd_sc_hd__inv_1 _3469_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q ),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_1 _3470_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q ),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_1 _3471_ (.A(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[5] ),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_1 _3472_ (.A(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[4] ),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_1 _3473_ (.A(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[3] ),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_1 _3474_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_1 _3475_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q ),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_1 _3476_ (.A(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[13] ),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_1 _3477_ (.A(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[15] ),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_1 _3478_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q ),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _3479_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _3480_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _3481_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _3482_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_1 _3483_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_1 _3484_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q ),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_1 _3485_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q ),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_1 _3486_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q ),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_1 _3487_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q ),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _3488_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_1 _3489_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q ),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_2 _3490_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_1 _3491_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q ),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _3492_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_1 _3493_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q ),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_1 _3494_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q ),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_1 _3495_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q ),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_1 _3496_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q ),
    .Y(_0191_));
 sky130_fd_sc_hd__inv_1 _3497_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q ),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_1 _3498_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q ),
    .Y(_0193_));
 sky130_fd_sc_hd__inv_1 _3499_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q ),
    .Y(_0194_));
 sky130_fd_sc_hd__inv_1 _3500_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q ),
    .Y(_0195_));
 sky130_fd_sc_hd__inv_2 _3501_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .Y(_0196_));
 sky130_fd_sc_hd__inv_2 _3502_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .Y(_0197_));
 sky130_fd_sc_hd__inv_1 _3503_ (.A(net1045),
    .Y(_0198_));
 sky130_fd_sc_hd__inv_1 _3504_ (.A(net1019),
    .Y(_0199_));
 sky130_fd_sc_hd__mux4_1 _3505_ (.A0(net1020),
    .A1(net1036),
    .A2(net1032),
    .A3(net985),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0200_));
 sky130_fd_sc_hd__and2_1 _3506_ (.A(_0097_),
    .B(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__mux4_1 _3507_ (.A0(net1053),
    .A1(net1048),
    .A2(net1029),
    .A3(net822),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0202_));
 sky130_fd_sc_hd__a21bo_1 _3508_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ),
    .A2(_0202_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q ),
    .X(_0203_));
 sky130_fd_sc_hd__mux4_2 _3509_ (.A0(net1018),
    .A1(net1033),
    .A2(net982),
    .A3(net1040),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0204_));
 sky130_fd_sc_hd__or2_4 _3510_ (.A(_0204_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_0205_));
 sky130_fd_sc_hd__mux4_2 _3511_ (.A0(net1050),
    .A1(net1045),
    .A2(net1026),
    .A3(net1016),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0206_));
 sky130_fd_sc_hd__o21a_1 _3512_ (.A1(_0028_),
    .A2(_0206_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q ),
    .X(_0207_));
 sky130_fd_sc_hd__mux4_1 _3513_ (.A0(net208),
    .A1(net1),
    .A2(net25),
    .A3(net1262),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0208_));
 sky130_fd_sc_hd__mux4_1 _3514_ (.A0(net79),
    .A1(net87),
    .A2(net99),
    .A3(net113),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _3515_ (.A0(_0208_),
    .A1(_0209_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_0210_));
 sky130_fd_sc_hd__a22o_4 _3516_ (.A1(_0207_),
    .A2(_0205_),
    .B1(_0210_),
    .B2(_0029_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ));
 sky130_fd_sc_hd__a221o_2 _3517_ (.A1(_0205_),
    .A2(_0207_),
    .B1(_0210_),
    .B2(_0029_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q ),
    .X(_0211_));
 sky130_fd_sc_hd__a21oi_1 _3518_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q ),
    .A2(_0030_),
    .B1(_0031_),
    .Y(_0212_));
 sky130_fd_sc_hd__mux2_1 _3519_ (.A0(net187),
    .A1(net132),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q ),
    .X(_0213_));
 sky130_fd_sc_hd__a22o_2 _3520_ (.A1(net651),
    .A2(_0212_),
    .B1(_0213_),
    .B2(_0031_),
    .X(_0214_));
 sky130_fd_sc_hd__inv_2 _3521_ (.A(_0214_),
    .Y(_0215_));
 sky130_fd_sc_hd__a221o_4 _3522_ (.A1(_0211_),
    .A2(_0212_),
    .B1(_0213_),
    .B2(_0031_),
    .C1(_0032_),
    .X(_0216_));
 sky130_fd_sc_hd__o21ba_4 _3523_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ),
    .A2(net979),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0217_));
 sky130_fd_sc_hd__mux4_2 _3524_ (.A0(net925),
    .A1(net970),
    .A2(net999),
    .A3(net987),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0218_));
 sky130_fd_sc_hd__or2_4 _3525_ (.A(_0218_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .X(_0219_));
 sky130_fd_sc_hd__mux4_1 _3526_ (.A0(net993),
    .A1(net1021),
    .A2(net1003),
    .A3(net1007),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0220_));
 sky130_fd_sc_hd__o21a_1 _3527_ (.A1(_0037_),
    .A2(_0220_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q ),
    .X(_0221_));
 sky130_fd_sc_hd__mux4_1 _3528_ (.A0(net175),
    .A1(net181),
    .A2(net197),
    .A3(net126),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0222_));
 sky130_fd_sc_hd__mux4_1 _3529_ (.A0(net1221),
    .A1(net72),
    .A2(net217),
    .A3(net231),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _3530_ (.A0(_0222_),
    .A1(_0223_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .X(_0224_));
 sky130_fd_sc_hd__a22o_4 _3531_ (.A1(net827),
    .A2(_0221_),
    .B1(_0224_),
    .B2(_0038_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ));
 sky130_fd_sc_hd__a221o_1 _3532_ (.A1(_0219_),
    .A2(_0221_),
    .B1(_0224_),
    .B2(_0038_),
    .C1(_0036_),
    .X(_0225_));
 sky130_fd_sc_hd__o21a_1 _3533_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q ),
    .A2(net221),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q ),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _3534_ (.A0(net196),
    .A1(net125),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q ),
    .X(_0227_));
 sky130_fd_sc_hd__a22o_2 _3535_ (.A1(net668),
    .A2(_0226_),
    .B1(_0227_),
    .B2(_0039_),
    .X(_0228_));
 sky130_fd_sc_hd__a221o_2 _3536_ (.A1(_0225_),
    .A2(_0226_),
    .B1(_0227_),
    .B2(_0039_),
    .C1(_0032_),
    .X(_0229_));
 sky130_fd_sc_hd__mux4_2 _3537_ (.A0(net811),
    .A1(net970),
    .A2(net664),
    .A3(net656),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0230_));
 sky130_fd_sc_hd__or2_4 _3538_ (.A(_0230_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ),
    .X(_0231_));
 sky130_fd_sc_hd__mux4_1 _3539_ (.A0(net992),
    .A1(net1022),
    .A2(net1002),
    .A3(net1010),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0232_));
 sky130_fd_sc_hd__o21a_1 _3540_ (.A1(_0034_),
    .A2(_0232_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0233_));
 sky130_fd_sc_hd__mux4_1 _3541_ (.A0(net176),
    .A1(net182),
    .A2(net127),
    .A3(net1222),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0234_));
 sky130_fd_sc_hd__mux4_1 _3542_ (.A0(net73),
    .A1(net81),
    .A2(net218),
    .A3(net230),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _3543_ (.A0(_0234_),
    .A1(_0235_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ),
    .X(_0236_));
 sky130_fd_sc_hd__a22o_4 _3544_ (.A1(_0233_),
    .A2(_0231_),
    .B1(_0236_),
    .B2(_0035_),
    .X(_0237_));
 sky130_fd_sc_hd__o21a_4 _3545_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ),
    .A2(_0237_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0238_));
 sky130_fd_sc_hd__a22o_4 _3546_ (.A1(_0216_),
    .A2(_0217_),
    .B1(net667),
    .B2(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__a221o_1 _3547_ (.A1(_0217_),
    .A2(_0216_),
    .B1(_0229_),
    .B2(_0238_),
    .C1(net617),
    .X(_0240_));
 sky130_fd_sc_hd__a21oi_1 _3548_ (.A1(_0040_),
    .A2(net617),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .Y(_0241_));
 sky130_fd_sc_hd__mux2_1 _3549_ (.A0(net1),
    .A1(net5),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_0242_));
 sky130_fd_sc_hd__a221o_1 _3550_ (.A1(_0241_),
    .A2(_0240_),
    .B1(_0242_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _3551_ (.A0(net57),
    .A1(net61),
    .S(net617),
    .X(_0244_));
 sky130_fd_sc_hd__inv_2 _3552_ (.A(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__mux2_1 _3553_ (.A0(net93),
    .A1(net1226),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_0246_));
 sky130_fd_sc_hd__nand2_1 _3554_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .B(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__o211a_1 _3555_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_0245_),
    .B1(_0247_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0248_));
 sky130_fd_sc_hd__nor2_1 _3556_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q ),
    .B(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__mux4_1 _3557_ (.A0(net867),
    .A1(net1045),
    .A2(net1050),
    .A3(net1016),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .S1(net617),
    .X(_0250_));
 sky130_fd_sc_hd__mux4_2 _3558_ (.A0(net1017),
    .A1(net1037),
    .A2(net1031),
    .A3(net982),
    .S0(net617),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0251_));
 sky130_fd_sc_hd__or2_4 _3559_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ),
    .B(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__o211a_1 _3560_ (.A1(_0042_),
    .A2(_0250_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q ),
    .C1(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__a21o_4 _3561_ (.A1(net825),
    .A2(_0249_),
    .B1(_0253_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ));
 sky130_fd_sc_hd__a211o_1 _3562_ (.A1(_0243_),
    .A2(_0249_),
    .B1(_0253_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .X(_0254_));
 sky130_fd_sc_hd__a21oi_2 _3563_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .A2(_0043_),
    .B1(_0044_),
    .Y(_0255_));
 sky130_fd_sc_hd__mux2_1 _3564_ (.A0(net193),
    .A1(net138),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .X(_0256_));
 sky130_fd_sc_hd__a22oi_4 _3565_ (.A1(net639),
    .A2(_0255_),
    .B1(_0256_),
    .B2(_0044_),
    .Y(_0257_));
 sky130_fd_sc_hd__a221o_1 _3566_ (.A1(_0255_),
    .A2(net834),
    .B1(_0256_),
    .B2(_0044_),
    .C1(_0045_),
    .X(_0258_));
 sky130_fd_sc_hd__o21ba_1 _3567_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ),
    .A2(net998),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q ),
    .X(_0259_));
 sky130_fd_sc_hd__mux4_1 _3568_ (.A0(net909),
    .A1(net970),
    .A2(net977),
    .A3(net987),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0260_));
 sky130_fd_sc_hd__and2b_1 _3569_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .B(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__mux4_1 _3570_ (.A0(net992),
    .A1(net1021),
    .A2(net1002),
    .A3(net1007),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0262_));
 sky130_fd_sc_hd__a21bo_1 _3571_ (.A1(_0262_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q ),
    .X(_0263_));
 sky130_fd_sc_hd__mux4_1 _3572_ (.A0(net182),
    .A1(net127),
    .A2(net1224),
    .A3(net1222),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0264_));
 sky130_fd_sc_hd__mux4_1 _3573_ (.A0(net73),
    .A1(net81),
    .A2(net218),
    .A3(net234),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _3574_ (.A0(_0264_),
    .A1(_0265_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .X(_0266_));
 sky130_fd_sc_hd__o22a_4 _3575_ (.A1(_0261_),
    .A2(_0263_),
    .B1(_0266_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ));
 sky130_fd_sc_hd__inv_4 _3576_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .Y(_0267_));
 sky130_fd_sc_hd__mux4_2 _3577_ (.A0(_0046_),
    .A1(_0047_),
    .A2(_0033_),
    .A3(_0267_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_0268_));
 sky130_fd_sc_hd__nand2_2 _3578_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ),
    .B(_0268_),
    .Y(_0269_));
 sky130_fd_sc_hd__mux4_2 _3579_ (.A0(net994),
    .A1(net1023),
    .A2(net1004),
    .A3(net1007),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0270_));
 sky130_fd_sc_hd__mux4_1 _3580_ (.A0(net969),
    .A1(net978),
    .A2(net998),
    .A3(net989),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0271_));
 sky130_fd_sc_hd__and2b_1 _3581_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .B(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__a21bo_1 _3582_ (.A1(_0270_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q ),
    .X(_0273_));
 sky130_fd_sc_hd__mux4_1 _3583_ (.A0(net70),
    .A1(net82),
    .A2(net215),
    .A3(net231),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0274_));
 sky130_fd_sc_hd__mux4_1 _3584_ (.A0(net177),
    .A1(net179),
    .A2(net124),
    .A3(net140),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _3585_ (.A0(_0275_),
    .A1(_0274_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .X(_0276_));
 sky130_fd_sc_hd__o22a_1 _3586_ (.A1(_0273_),
    .A2(_0272_),
    .B1(_0276_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q ),
    .X(_0277_));
 sky130_fd_sc_hd__o211a_4 _3587_ (.A1(_0277_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ),
    .B1(_0269_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q ),
    .X(_0278_));
 sky130_fd_sc_hd__a21o_4 _3588_ (.A1(net635),
    .A2(_0259_),
    .B1(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_4 _3589_ (.A0(_0279_),
    .A1(net191),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _3590_ (.A0(net2),
    .A1(net10),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .X(_0281_));
 sky130_fd_sc_hd__or2_1 _3591_ (.A(_0096_),
    .B(_0281_),
    .X(_0282_));
 sky130_fd_sc_hd__o211a_1 _3592_ (.A1(_0280_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .B1(_0282_),
    .C1(_0097_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _3593_ (.A0(net58),
    .A1(net66),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .X(_0284_));
 sky130_fd_sc_hd__or2_1 _3594_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .B(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _3595_ (.A0(net94),
    .A1(net1225),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .X(_0286_));
 sky130_fd_sc_hd__o211a_1 _3596_ (.A1(_0096_),
    .A2(_0286_),
    .B1(_0285_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ),
    .X(_0287_));
 sky130_fd_sc_hd__o32a_4 _3597_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0287_),
    .A3(_0283_),
    .B1(_0201_),
    .B2(_0203_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ));
 sky130_fd_sc_hd__mux2_4 _3598_ (.A0(net80),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _3599_ (.A0(net201),
    .A1(net23),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_0289_));
 sky130_fd_sc_hd__inv_2 _3600_ (.A(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__o21ai_1 _3601_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(_0290_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ),
    .Y(_0291_));
 sky130_fd_sc_hd__a21o_1 _3602_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(_0288_),
    .B1(_0291_),
    .X(_0292_));
 sky130_fd_sc_hd__mux4_1 _3603_ (.A0(net193),
    .A1(net68),
    .A2(net12),
    .A3(net115),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q ),
    .X(_0293_));
 sky130_fd_sc_hd__or2_1 _3604_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ),
    .B(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__mux4_1 _3605_ (.A0(net974),
    .A1(net969),
    .A2(net978),
    .A3(net998),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0295_));
 sky130_fd_sc_hd__mux4_2 _3606_ (.A0(net989),
    .A1(net1006),
    .A2(net864),
    .A3(net1010),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0296_));
 sky130_fd_sc_hd__or2_4 _3607_ (.A(_0087_),
    .B(_0296_),
    .X(_0297_));
 sky130_fd_sc_hd__o211a_1 _3608_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .A2(_0295_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q ),
    .C1(_0297_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _3609_ (.A0(net206),
    .A1(net1262),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_0299_));
 sky130_fd_sc_hd__nand2b_2 _3610_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q ),
    .B(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__mux4_2 _3611_ (.A0(net1017),
    .A1(net1037),
    .A2(net866),
    .A3(net865),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0301_));
 sky130_fd_sc_hd__mux4_2 _3612_ (.A0(net1051),
    .A1(net828),
    .A2(net1026),
    .A3(net1016),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0302_));
 sky130_fd_sc_hd__o21a_1 _3613_ (.A1(_0301_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0303_));
 sky130_fd_sc_hd__o21ai_4 _3614_ (.A1(_0065_),
    .A2(_0302_),
    .B1(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__a211o_4 _3615_ (.A1(net652),
    .A2(_0259_),
    .B1(_0278_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0305_));
 sky130_fd_sc_hd__a21oi_1 _3616_ (.A1(_0054_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .Y(_0306_));
 sky130_fd_sc_hd__mux2_1 _3617_ (.A0(net2),
    .A1(net10),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0307_));
 sky130_fd_sc_hd__a221oi_4 _3618_ (.A1(_0306_),
    .A2(_0305_),
    .B1(_0307_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ),
    .Y(_0308_));
 sky130_fd_sc_hd__mux2_1 _3619_ (.A0(net58),
    .A1(net60),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0309_));
 sky130_fd_sc_hd__inv_2 _3620_ (.A(_0309_),
    .Y(_0310_));
 sky130_fd_sc_hd__mux2_1 _3621_ (.A0(net66),
    .A1(net94),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0311_));
 sky130_fd_sc_hd__nand2_1 _3622_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .B(_0311_),
    .Y(_0312_));
 sky130_fd_sc_hd__o211a_1 _3623_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .A2(_0310_),
    .B1(_0312_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ),
    .X(_0313_));
 sky130_fd_sc_hd__o31a_4 _3624_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ),
    .A2(_0308_),
    .A3(_0313_),
    .B1(_0304_),
    .X(_0314_));
 sky130_fd_sc_hd__o311a_4 _3625_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ),
    .A2(_0313_),
    .A3(_0308_),
    .B1(_0304_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_0315_));
 sky130_fd_sc_hd__o21ai_2 _3626_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ),
    .A2(net97),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_0316_));
 sky130_fd_sc_hd__o21ai_4 _3627_ (.A1(_0315_),
    .A2(_0316_),
    .B1(_0300_),
    .Y(_0317_));
 sky130_fd_sc_hd__o211ai_4 _3628_ (.A1(_0316_),
    .A2(_0315_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ),
    .C1(_0300_),
    .Y(_0318_));
 sky130_fd_sc_hd__mux4_1 _3629_ (.A0(net1019),
    .A1(net1035),
    .A2(net986),
    .A3(net1041),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0319_));
 sky130_fd_sc_hd__and2_1 _3630_ (.A(_0067_),
    .B(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__mux4_2 _3631_ (.A0(net1052),
    .A1(net828),
    .A2(net1027),
    .A3(net1057),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0321_));
 sky130_fd_sc_hd__a21bo_1 _3632_ (.A1(_0321_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q ),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _3633_ (.A0(_0239_),
    .A1(net188),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _3634_ (.A0(net200),
    .A1(net7),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .X(_0324_));
 sky130_fd_sc_hd__or2_1 _3635_ (.A(_0066_),
    .B(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__o211a_1 _3636_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .A2(_0323_),
    .B1(_0325_),
    .C1(_0067_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _3637_ (.A0(net21),
    .A1(net63),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .X(_0327_));
 sky130_fd_sc_hd__or2_1 _3638_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .B(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _3639_ (.A0(net99),
    .A1(net118),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .X(_0329_));
 sky130_fd_sc_hd__o211a_1 _3640_ (.A1(_0066_),
    .A2(_0329_),
    .B1(_0328_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_0330_));
 sky130_fd_sc_hd__o32a_4 _3641_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q ),
    .A2(_0330_),
    .A3(_0326_),
    .B1(_0320_),
    .B2(_0322_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ));
 sky130_fd_sc_hd__o21ai_2 _3642_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q ),
    .Y(_0331_));
 sky130_fd_sc_hd__inv_2 _3643_ (.A(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__mux4_2 _3644_ (.A0(net909),
    .A1(net970),
    .A2(net977),
    .A3(net987),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0333_));
 sky130_fd_sc_hd__and2b_1 _3645_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q ),
    .B(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__mux4_1 _3646_ (.A0(net992),
    .A1(net1022),
    .A2(net1002),
    .A3(net1007),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0335_));
 sky130_fd_sc_hd__a21bo_1 _3647_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q ),
    .A2(_0335_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q ),
    .X(_0336_));
 sky130_fd_sc_hd__mux4_1 _3648_ (.A0(net182),
    .A1(net1224),
    .A2(net194),
    .A3(net127),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .X(_0337_));
 sky130_fd_sc_hd__mux4_1 _3649_ (.A0(net1222),
    .A1(net73),
    .A2(net218),
    .A3(net230),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _3650_ (.A0(_0337_),
    .A1(_0338_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q ),
    .X(_0339_));
 sky130_fd_sc_hd__o22a_4 _3651_ (.A1(_0336_),
    .A2(_0334_),
    .B1(_0339_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ));
 sky130_fd_sc_hd__mux4_2 _3652_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .A1(net16),
    .A2(net72),
    .A3(net108),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q ),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _3653_ (.A0(net1046),
    .A1(net968),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ),
    .X(_0341_));
 sky130_fd_sc_hd__and2b_1 _3654_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q ),
    .B(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__a21oi_4 _3655_ (.A1(_0332_),
    .A2(_0318_),
    .B1(net640),
    .Y(_0343_));
 sky130_fd_sc_hd__inv_6 _3656_ (.A(net629),
    .Y(_0344_));
 sky130_fd_sc_hd__a211o_1 _3657_ (.A1(_0318_),
    .A2(_0332_),
    .B1(_0342_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_0345_));
 sky130_fd_sc_hd__a21oi_1 _3658_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .A2(_0068_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .Y(_0346_));
 sky130_fd_sc_hd__mux2_1 _3659_ (.A0(net210),
    .A1(net1073),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_0347_));
 sky130_fd_sc_hd__a221o_1 _3660_ (.A1(_0346_),
    .A2(_0345_),
    .B1(_0347_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .C1(_0069_),
    .X(_0348_));
 sky130_fd_sc_hd__mux4_1 _3661_ (.A0(net176),
    .A1(net1224),
    .A2(net184),
    .A3(net129),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_0349_));
 sky130_fd_sc_hd__o21ba_1 _3662_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .A2(_0349_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q ),
    .X(_0350_));
 sky130_fd_sc_hd__mux4_2 _3663_ (.A0(net991),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .A2(net1005),
    .A3(net1009),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_0351_));
 sky130_fd_sc_hd__mux4_1 _3664_ (.A0(net655),
    .A1(net971),
    .A2(net980),
    .A3(net1001),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_0352_));
 sky130_fd_sc_hd__o21a_1 _3665_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .A2(_0352_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q ),
    .X(_0353_));
 sky130_fd_sc_hd__o21ai_2 _3666_ (.A1(_0069_),
    .A2(_0351_),
    .B1(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__inv_2 _3667_ (.A(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__a21o_4 _3668_ (.A1(_0348_),
    .A2(_0350_),
    .B1(_0355_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ));
 sky130_fd_sc_hd__a211o_4 _3669_ (.A1(_0348_),
    .A2(_0350_),
    .B1(_0355_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ),
    .X(_0356_));
 sky130_fd_sc_hd__a21oi_2 _3670_ (.A1(_0070_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ),
    .Y(_0357_));
 sky130_fd_sc_hd__mux2_1 _3671_ (.A0(net74),
    .A1(net110),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ),
    .X(_0358_));
 sky130_fd_sc_hd__a22oi_4 _3672_ (.A1(_0357_),
    .A2(_0356_),
    .B1(_0358_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ),
    .Y(_0359_));
 sky130_fd_sc_hd__a221o_2 _3673_ (.A1(_0357_),
    .A2(_0356_),
    .B1(_0358_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ),
    .C1(_0086_),
    .X(_0360_));
 sky130_fd_sc_hd__o21ba_1 _3674_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ),
    .A2(net1027),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q ),
    .X(_0361_));
 sky130_fd_sc_hd__a211o_1 _3675_ (.A1(net635),
    .A2(_0259_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .C1(_0278_),
    .X(_0362_));
 sky130_fd_sc_hd__a21oi_1 _3676_ (.A1(_0048_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .Y(_0363_));
 sky130_fd_sc_hd__mux2_1 _3677_ (.A0(net201),
    .A1(net8),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .X(_0364_));
 sky130_fd_sc_hd__a221o_1 _3678_ (.A1(_0363_),
    .A2(_0362_),
    .B1(_0364_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _3679_ (.A0(net1261),
    .A1(net64),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .X(_0366_));
 sky130_fd_sc_hd__inv_1 _3680_ (.A(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__mux2_1 _3681_ (.A0(net100),
    .A1(net114),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .X(_0368_));
 sky130_fd_sc_hd__nand2_1 _3682_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .B(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__o211a_1 _3683_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .A2(_0367_),
    .B1(_0369_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ),
    .X(_0370_));
 sky130_fd_sc_hd__nor2_1 _3684_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q ),
    .B(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__mux4_2 _3685_ (.A0(net1050),
    .A1(net1045),
    .A2(net1026),
    .A3(net1016),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0372_));
 sky130_fd_sc_hd__or2_4 _3686_ (.A(_0049_),
    .B(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__mux4_2 _3687_ (.A0(net1017),
    .A1(net823),
    .A2(net982),
    .A3(net867),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0374_));
 sky130_fd_sc_hd__o211a_1 _3688_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ),
    .A2(_0374_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q ),
    .C1(_0373_),
    .X(_0375_));
 sky130_fd_sc_hd__a21o_1 _3689_ (.A1(_0365_),
    .A2(_0371_),
    .B1(_0375_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ));
 sky130_fd_sc_hd__mux4_2 _3690_ (.A0(net1017),
    .A1(net1031),
    .A2(net982),
    .A3(net1042),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0376_));
 sky130_fd_sc_hd__or2_4 _3691_ (.A(_0376_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ),
    .X(_0377_));
 sky130_fd_sc_hd__mux4_1 _3692_ (.A0(net1053),
    .A1(net828),
    .A2(net1028),
    .A3(net1016),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0378_));
 sky130_fd_sc_hd__o21a_1 _3693_ (.A1(_0076_),
    .A2(_0378_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q ),
    .X(_0379_));
 sky130_fd_sc_hd__mux4_1 _3694_ (.A0(net1262),
    .A1(net99),
    .A2(net63),
    .A3(net113),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ),
    .X(_0380_));
 sky130_fd_sc_hd__mux4_1 _3695_ (.A0(net188),
    .A1(net1),
    .A2(net200),
    .A3(net7),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _3696_ (.A0(_0380_),
    .A1(_0381_),
    .S(_0076_),
    .X(_0382_));
 sky130_fd_sc_hd__a22o_4 _3697_ (.A1(_0379_),
    .A2(_0377_),
    .B1(_0382_),
    .B2(_0077_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ));
 sky130_fd_sc_hd__inv_2 _3698_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ),
    .Y(_0383_));
 sky130_fd_sc_hd__mux4_2 _3699_ (.A0(_0075_),
    .A1(_0078_),
    .A2(_0072_),
    .A3(_0383_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q ),
    .X(_0384_));
 sky130_fd_sc_hd__nand2_1 _3700_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ),
    .B(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__o211a_4 _3701_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ),
    .B1(_0385_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q ),
    .X(_0386_));
 sky130_fd_sc_hd__a21o_4 _3702_ (.A1(_0360_),
    .A2(_0361_),
    .B1(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__a211o_1 _3703_ (.A1(_0360_),
    .A2(_0361_),
    .B1(_0386_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0388_));
 sky130_fd_sc_hd__a21oi_1 _3704_ (.A1(_0053_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .Y(_0389_));
 sky130_fd_sc_hd__mux2_1 _3705_ (.A0(net211),
    .A1(net1072),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0390_));
 sky130_fd_sc_hd__a221o_1 _3706_ (.A1(_0388_),
    .A2(_0389_),
    .B1(_0390_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .C1(_0087_),
    .X(_0391_));
 sky130_fd_sc_hd__mux4_1 _3707_ (.A0(net177),
    .A1(net185),
    .A2(net122),
    .A3(net130),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0392_));
 sky130_fd_sc_hd__o21ba_1 _3708_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .A2(_0392_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q ),
    .X(_0393_));
 sky130_fd_sc_hd__a21o_4 _3709_ (.A1(_0391_),
    .A2(_0393_),
    .B1(_0298_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ));
 sky130_fd_sc_hd__mux4_1 _3710_ (.A0(net815),
    .A1(net1036),
    .A2(net1032),
    .A3(net985),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0394_));
 sky130_fd_sc_hd__and2_1 _3711_ (.A(_0113_),
    .B(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__mux4_2 _3712_ (.A0(net1042),
    .A1(net1028),
    .A2(net1053),
    .A3(net822),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0396_));
 sky130_fd_sc_hd__a21bo_1 _3713_ (.A1(_0396_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q ),
    .X(_0397_));
 sky130_fd_sc_hd__mux4_2 _3714_ (.A0(net973),
    .A1(net977),
    .A2(net997),
    .A3(net987),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0398_));
 sky130_fd_sc_hd__and2b_1 _3715_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .B(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__mux4_1 _3716_ (.A0(net992),
    .A1(net1021),
    .A2(net1002),
    .A3(net1007),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0400_));
 sky130_fd_sc_hd__a21bo_1 _3717_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .A2(_0400_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q ),
    .X(_0401_));
 sky130_fd_sc_hd__mux4_1 _3718_ (.A0(net180),
    .A1(net196),
    .A2(net119),
    .A3(net125),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0402_));
 sky130_fd_sc_hd__mux4_1 _3719_ (.A0(net1222),
    .A1(net71),
    .A2(net216),
    .A3(net230),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _3720_ (.A0(_0402_),
    .A1(_0403_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .X(_0404_));
 sky130_fd_sc_hd__o22a_4 _3721_ (.A1(_0399_),
    .A2(_0401_),
    .B1(_0404_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ));
 sky130_fd_sc_hd__mux4_2 _3722_ (.A0(net205),
    .A1(net232),
    .A2(net84),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q ),
    .X(_0405_));
 sky130_fd_sc_hd__mux4_1 _3723_ (.A0(net993),
    .A1(net1023),
    .A2(net1004),
    .A3(net1007),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0406_));
 sky130_fd_sc_hd__mux4_1 _3724_ (.A0(net973),
    .A1(net970),
    .A2(net997),
    .A3(net990),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _3725_ (.A0(_0406_),
    .A1(_0407_),
    .S(_0056_),
    .X(_0408_));
 sky130_fd_sc_hd__mux4_1 _3726_ (.A0(net72),
    .A1(net217),
    .A2(net84),
    .A3(net231),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .X(_0409_));
 sky130_fd_sc_hd__and2_1 _3727_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ),
    .B(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__mux4_1 _3728_ (.A0(net175),
    .A1(net181),
    .A2(net126),
    .A3(net1221),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0411_));
 sky130_fd_sc_hd__a21o_1 _3729_ (.A1(_0056_),
    .A2(_0411_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0412_));
 sky130_fd_sc_hd__o22a_2 _3730_ (.A1(_0057_),
    .A2(_0408_),
    .B1(_0410_),
    .B2(_0412_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ));
 sky130_fd_sc_hd__mux4_2 _3731_ (.A0(net191),
    .A1(net136),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .A3(net227),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q ),
    .X(_0413_));
 sky130_fd_sc_hd__mux4_2 _3732_ (.A0(net993),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ),
    .A2(_0413_),
    .A3(_0405_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q ),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _3733_ (.A0(_0414_),
    .A1(net193),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _3734_ (.A0(net1263),
    .A1(net12),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0416_));
 sky130_fd_sc_hd__or2_1 _3735_ (.A(_0112_),
    .B(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__o211a_1 _3736_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .A2(_0415_),
    .B1(_0417_),
    .C1(_0113_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _3737_ (.A0(net60),
    .A1(net68),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0419_));
 sky130_fd_sc_hd__or2_1 _3738_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .B(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _3739_ (.A0(net94),
    .A1(net1225),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0421_));
 sky130_fd_sc_hd__o211a_1 _3740_ (.A1(_0112_),
    .A2(_0421_),
    .B1(_0420_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ),
    .X(_0422_));
 sky130_fd_sc_hd__o32a_4 _3741_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0418_),
    .A3(_0422_),
    .B1(_0397_),
    .B2(_0395_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ));
 sky130_fd_sc_hd__mux4_1 _3742_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .A1(net19),
    .A2(net75),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q ),
    .X(_0423_));
 sky130_fd_sc_hd__a211o_1 _3743_ (.A1(_0371_),
    .A2(_0365_),
    .B1(_0375_),
    .C1(_0025_),
    .X(_0424_));
 sky130_fd_sc_hd__or2_1 _3744_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ),
    .B(net104),
    .X(_0425_));
 sky130_fd_sc_hd__o21ba_1 _3745_ (.A1(net200),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ),
    .X(_0426_));
 sky130_fd_sc_hd__o21a_1 _3746_ (.A1(net7),
    .A2(_0025_),
    .B1(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__a31oi_4 _3747_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ),
    .A2(_0424_),
    .A3(_0425_),
    .B1(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__inv_2 _3748_ (.A(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__a311o_1 _3749_ (.A1(_0424_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ),
    .A3(_0425_),
    .B1(_0427_),
    .C1(_0021_),
    .X(_0430_));
 sky130_fd_sc_hd__mux4_2 _3750_ (.A0(net1017),
    .A1(net823),
    .A2(net866),
    .A3(net867),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_0431_));
 sky130_fd_sc_hd__mux4_2 _3751_ (.A0(net1050),
    .A1(net1045),
    .A2(net824),
    .A3(net1056),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_4 _3752_ (.A0(_0431_),
    .A1(_0432_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ),
    .X(_0433_));
 sky130_fd_sc_hd__mux4_2 _3753_ (.A0(net637),
    .A1(net198),
    .A2(net190),
    .A3(net9),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ),
    .X(_0434_));
 sky130_fd_sc_hd__and2b_1 _3754_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ),
    .B(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__mux4_1 _3755_ (.A0(net1262),
    .A1(net65),
    .A2(net101),
    .A3(net113),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_0436_));
 sky130_fd_sc_hd__a21o_1 _3756_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ),
    .A2(_0436_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_0437_));
 sky130_fd_sc_hd__o22a_4 _3757_ (.A1(_0433_),
    .A2(_0024_),
    .B1(_0435_),
    .B2(_0437_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ));
 sky130_fd_sc_hd__or2_1 _3758_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ),
    .X(_0438_));
 sky130_fd_sc_hd__mux4_2 _3759_ (.A0(net868),
    .A1(net70),
    .A2(net14),
    .A3(net106),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q ),
    .X(_0439_));
 sky130_fd_sc_hd__o21ba_1 _3760_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ),
    .A2(net867),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ),
    .X(_0440_));
 sky130_fd_sc_hd__o21a_1 _3761_ (.A1(_0439_),
    .A2(_0021_),
    .B1(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__a31o_4 _3762_ (.A1(_0430_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ),
    .A3(_0438_),
    .B1(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__a311o_1 _3763_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ),
    .A2(_0430_),
    .A3(_0438_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .C1(_0441_),
    .X(_0443_));
 sky130_fd_sc_hd__a21oi_1 _3764_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .A2(_0050_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .Y(_0444_));
 sky130_fd_sc_hd__mux2_1 _3765_ (.A0(net210),
    .A1(net1073),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_0445_));
 sky130_fd_sc_hd__a221o_1 _3766_ (.A1(_0444_),
    .A2(_0443_),
    .B1(_0445_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .C1(_0051_),
    .X(_0446_));
 sky130_fd_sc_hd__mux4_1 _3767_ (.A0(net174),
    .A1(net178),
    .A2(net119),
    .A3(net141),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .X(_0447_));
 sky130_fd_sc_hd__o21ba_1 _3768_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .A2(_0447_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q ),
    .X(_0448_));
 sky130_fd_sc_hd__mux4_1 _3769_ (.A0(net974),
    .A1(net969),
    .A2(net979),
    .A3(net998),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .X(_0449_));
 sky130_fd_sc_hd__mux4_1 _3770_ (.A0(net989),
    .A1(net1024),
    .A2(net994),
    .A3(net1008),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_0450_));
 sky130_fd_sc_hd__or2_1 _3771_ (.A(_0051_),
    .B(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__o211a_4 _3772_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .A2(_0449_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q ),
    .C1(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__a21oi_4 _3773_ (.A1(net663),
    .A2(_0448_),
    .B1(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__inv_2 _3774_ (.A(_0453_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ));
 sky130_fd_sc_hd__mux4_2 _3775_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ),
    .A1(net76),
    .A2(net20),
    .A3(net112),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q ),
    .X(_0454_));
 sky130_fd_sc_hd__inv_2 _3776_ (.A(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__a21oi_1 _3777_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(_0455_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q ),
    .Y(_0456_));
 sky130_fd_sc_hd__o21a_1 _3778_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(_0423_),
    .B1(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__a31o_1 _3779_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q ),
    .A2(_0292_),
    .A3(_0294_),
    .B1(_0457_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X ));
 sky130_fd_sc_hd__mux2_4 _3780_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[14] ),
    .S(net1064),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_4 _3781_ (.A0(_0458_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[14] ),
    .S(net1068),
    .X(_0459_));
 sky130_fd_sc_hd__mux4_1 _3782_ (.A0(net1018),
    .A1(net1036),
    .A2(net983),
    .A3(net1042),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0460_));
 sky130_fd_sc_hd__or2_1 _3783_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ),
    .B(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__mux4_1 _3784_ (.A0(net1053),
    .A1(net1048),
    .A2(net1028),
    .A3(net1056),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0462_));
 sky130_fd_sc_hd__o21a_1 _3785_ (.A1(_0083_),
    .A2(_0462_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q ),
    .X(_0463_));
 sky130_fd_sc_hd__mux4_1 _3786_ (.A0(net189),
    .A1(net201),
    .A2(net2),
    .A3(net8),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0464_));
 sky130_fd_sc_hd__mux4_1 _3787_ (.A0(net1261),
    .A1(net64),
    .A2(net100),
    .A3(net116),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _3788_ (.A0(_0464_),
    .A1(_0465_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ),
    .X(_0466_));
 sky130_fd_sc_hd__a22o_1 _3789_ (.A1(_0461_),
    .A2(_0463_),
    .B1(_0466_),
    .B2(_0084_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ));
 sky130_fd_sc_hd__mux2_1 _3790_ (.A0(net117),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q ),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _3791_ (.A0(net8),
    .A1(net88),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q ),
    .X(_0468_));
 sky130_fd_sc_hd__and2b_1 _3792_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q ),
    .B(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__a211o_1 _3793_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q ),
    .A2(_0467_),
    .B1(_0469_),
    .C1(_0098_),
    .X(_0470_));
 sky130_fd_sc_hd__mux4_2 _3794_ (.A0(net209),
    .A1(net67),
    .A2(net11),
    .A3(net103),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q ),
    .X(_0471_));
 sky130_fd_sc_hd__or2_1 _3795_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ),
    .B(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__mux4_2 _3796_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ),
    .A1(net76),
    .A2(net20),
    .A3(net112),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ),
    .X(_0473_));
 sky130_fd_sc_hd__mux4_2 _3797_ (.A0(net19),
    .A1(net111),
    .A2(net75),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q ),
    .X(_0474_));
 sky130_fd_sc_hd__o21ba_1 _3798_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ),
    .A2(_0474_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q ),
    .X(_0475_));
 sky130_fd_sc_hd__o21a_1 _3799_ (.A1(_0098_),
    .A2(_0473_),
    .B1(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__a31o_4 _3800_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q ),
    .A2(_0470_),
    .A3(_0472_),
    .B1(_0476_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X ));
 sky130_fd_sc_hd__nand2b_1 _3801_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[4] ),
    .B(net1062),
    .Y(_0477_));
 sky130_fd_sc_hd__o21ai_4 _3802_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X ),
    .A2(net1062),
    .B1(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__mux4_1 _3803_ (.A0(net969),
    .A1(net978),
    .A2(net998),
    .A3(net989),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_0479_));
 sky130_fd_sc_hd__mux4_2 _3804_ (.A0(net994),
    .A1(net1023),
    .A2(net1004),
    .A3(net1011),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_4 _3805_ (.A0(_0479_),
    .A1(_0480_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .X(_0481_));
 sky130_fd_sc_hd__mux4_1 _3806_ (.A0(net179),
    .A1(net195),
    .A2(net1223),
    .A3(net124),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_0482_));
 sky130_fd_sc_hd__and2b_1 _3807_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .B(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__mux4_1 _3808_ (.A0(net1221),
    .A1(net215),
    .A2(net90),
    .A3(net231),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .X(_0484_));
 sky130_fd_sc_hd__a21o_1 _3809_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .A2(_0484_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_0485_));
 sky130_fd_sc_hd__o22a_4 _3810_ (.A1(_0481_),
    .A2(_0094_),
    .B1(_0483_),
    .B2(_0485_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ));
 sky130_fd_sc_hd__mux4_2 _3811_ (.A0(net1017),
    .A1(net823),
    .A2(net866),
    .A3(net1040),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0486_));
 sky130_fd_sc_hd__nor2_2 _3812_ (.A(_0486_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ),
    .Y(_0487_));
 sky130_fd_sc_hd__mux4_2 _3813_ (.A0(net1050),
    .A1(net1045),
    .A2(net1026),
    .A3(net1056),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0488_));
 sky130_fd_sc_hd__o21ai_2 _3814_ (.A1(_0488_),
    .A2(_0095_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q ),
    .Y(_0489_));
 sky130_fd_sc_hd__mux4_1 _3815_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .A1(net9),
    .A2(net190),
    .A3(net1262),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ),
    .X(_0490_));
 sky130_fd_sc_hd__nor2_1 _3816_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ),
    .B(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__mux4_1 _3817_ (.A0(net65),
    .A1(net101),
    .A2(net77),
    .A3(net113),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ),
    .X(_0492_));
 sky130_fd_sc_hd__nor2_1 _3818_ (.A(_0095_),
    .B(_0492_),
    .Y(_0493_));
 sky130_fd_sc_hd__o32a_4 _3819_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q ),
    .A2(_0491_),
    .A3(_0493_),
    .B1(_0487_),
    .B2(_0489_),
    .X(_0494_));
 sky130_fd_sc_hd__inv_1 _3820_ (.A(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__mux4_1 _3821_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .A1(net13),
    .A2(net69),
    .A3(_0495_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q ),
    .X(_0496_));
 sky130_fd_sc_hd__or2_1 _3822_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ),
    .B(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__mux4_1 _3823_ (.A0(net868),
    .A1(net70),
    .A2(net14),
    .A3(net106),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q ),
    .X(_0498_));
 sky130_fd_sc_hd__inv_1 _3824_ (.A(_0498_),
    .Y(_0499_));
 sky130_fd_sc_hd__a21oi_1 _3825_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ),
    .A2(_0499_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q ),
    .Y(_0500_));
 sky130_fd_sc_hd__mux4_2 _3826_ (.A0(net1017),
    .A1(net866),
    .A2(net865),
    .A3(net1041),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0501_));
 sky130_fd_sc_hd__mux4_1 _3827_ (.A0(net1051),
    .A1(net1046),
    .A2(net1027),
    .A3(net1056),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0502_));
 sky130_fd_sc_hd__or2_4 _3828_ (.A(_0063_),
    .B(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__o211a_1 _3829_ (.A1(_0501_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ),
    .B1(_0503_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q ),
    .X(_0504_));
 sky130_fd_sc_hd__or2_1 _3830_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .B(_0239_),
    .X(_0505_));
 sky130_fd_sc_hd__a21oi_1 _3831_ (.A1(_0062_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_0506_));
 sky130_fd_sc_hd__mux2_1 _3832_ (.A0(net7),
    .A1(net1262),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0507_));
 sky130_fd_sc_hd__a221o_1 _3833_ (.A1(_0505_),
    .A2(_0506_),
    .B1(_0507_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _3834_ (.A0(net63),
    .A1(net79),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0509_));
 sky130_fd_sc_hd__and2b_1 _3835_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .B(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _3836_ (.A0(net99),
    .A1(net113),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0511_));
 sky130_fd_sc_hd__a211o_1 _3837_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .A2(_0511_),
    .B1(_0510_),
    .C1(_0063_),
    .X(_0512_));
 sky130_fd_sc_hd__a31o_4 _3838_ (.A1(_0064_),
    .A2(_0508_),
    .A3(_0512_),
    .B1(_0504_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ));
 sky130_fd_sc_hd__mux2_4 _3839_ (.A0(net77),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _3840_ (.A0(net198),
    .A1(net1262),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ),
    .X(_0514_));
 sky130_fd_sc_hd__inv_2 _3841_ (.A(_0514_),
    .Y(_0515_));
 sky130_fd_sc_hd__o21ai_1 _3842_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q ),
    .A2(_0515_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ),
    .Y(_0516_));
 sky130_fd_sc_hd__a21o_1 _3843_ (.A1(_0513_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q ),
    .B1(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__mux4_2 _3844_ (.A0(net186),
    .A1(net5),
    .A2(net61),
    .A3(net118),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q ),
    .X(_0518_));
 sky130_fd_sc_hd__or2_1 _3845_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ),
    .B(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__a32o_2 _3846_ (.A1(_0517_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q ),
    .A3(_0519_),
    .B1(_0497_),
    .B2(_0500_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X ));
 sky130_fd_sc_hd__nand2b_1 _3847_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[7] ),
    .B(net1060),
    .Y(_0520_));
 sky130_fd_sc_hd__o21ai_4 _3848_ (.A1(net1060),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X ),
    .B1(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__or2_4 _3849_ (.A(_0478_),
    .B(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _3850_ (.A0(net114),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ),
    .X(_0523_));
 sky130_fd_sc_hd__and2_1 _3851_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q ),
    .B(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _3852_ (.A0(net199),
    .A1(net1261),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ),
    .X(_0525_));
 sky130_fd_sc_hd__inv_2 _3853_ (.A(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__o21ai_1 _3854_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q ),
    .A2(_0526_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ),
    .Y(_0527_));
 sky130_fd_sc_hd__mux4_2 _3855_ (.A0(net190),
    .A1(net65),
    .A2(net23),
    .A3(net101),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q ),
    .X(_0528_));
 sky130_fd_sc_hd__o221a_4 _3856_ (.A1(_0527_),
    .A2(_0524_),
    .B1(_0528_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q ),
    .X(_0529_));
 sky130_fd_sc_hd__mux4_2 _3857_ (.A0(net1050),
    .A1(net1045),
    .A2(net1026),
    .A3(net1016),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0530_));
 sky130_fd_sc_hd__mux4_1 _3858_ (.A0(net1017),
    .A1(net823),
    .A2(net1031),
    .A3(net1040),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_4 _3859_ (.A0(_0530_),
    .A1(_0531_),
    .S(_0060_),
    .X(_0532_));
 sky130_fd_sc_hd__mux4_1 _3860_ (.A0(net65),
    .A1(net101),
    .A2(net77),
    .A3(net117),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0533_));
 sky130_fd_sc_hd__and2_1 _3861_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ),
    .B(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__mux4_1 _3862_ (.A0(net190),
    .A1(net9),
    .A2(net1264),
    .A3(net1262),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0535_));
 sky130_fd_sc_hd__a21o_1 _3863_ (.A1(_0060_),
    .A2(_0535_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q ),
    .X(_0536_));
 sky130_fd_sc_hd__o22a_4 _3864_ (.A1(_0532_),
    .A2(_0061_),
    .B1(_0534_),
    .B2(_0536_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ));
 sky130_fd_sc_hd__inv_2 _3865_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .Y(_0537_));
 sky130_fd_sc_hd__mux4_1 _3866_ (.A0(net922),
    .A1(net971),
    .A2(net980),
    .A3(net1001),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0538_));
 sky130_fd_sc_hd__mux4_1 _3867_ (.A0(net995),
    .A1(net1025),
    .A2(net1005),
    .A3(net1012),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0539_));
 sky130_fd_sc_hd__or2_1 _3868_ (.A(_0091_),
    .B(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__o211a_1 _3869_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .A2(_0538_),
    .B1(_0540_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q ),
    .X(_0541_));
 sky130_fd_sc_hd__mux4_2 _3870_ (.A0(net1037),
    .A1(net1033),
    .A2(net865),
    .A3(net1040),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_0542_));
 sky130_fd_sc_hd__mux4_1 _3871_ (.A0(net1050),
    .A1(net1045),
    .A2(net824),
    .A3(net1016),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_0543_));
 sky130_fd_sc_hd__or2_1 _3872_ (.A(_0089_),
    .B(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__o211a_1 _3873_ (.A1(_0542_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ),
    .B1(_0544_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q ),
    .X(_0545_));
 sky130_fd_sc_hd__or2_4 _3874_ (.A(net813),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0546_));
 sky130_fd_sc_hd__a21oi_1 _3875_ (.A1(_0026_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .Y(_0547_));
 sky130_fd_sc_hd__mux2_1 _3876_ (.A0(net199),
    .A1(net24),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0548_));
 sky130_fd_sc_hd__a221o_1 _3877_ (.A1(_0547_),
    .A2(_0546_),
    .B1(_0548_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ),
    .X(_0549_));
 sky130_fd_sc_hd__mux2_1 _3878_ (.A0(net1261),
    .A1(net62),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0550_));
 sky130_fd_sc_hd__and2b_1 _3879_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .B(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_1 _3880_ (.A0(net98),
    .A1(net114),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0552_));
 sky130_fd_sc_hd__a211o_1 _3881_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .A2(_0552_),
    .B1(_0551_),
    .C1(_0089_),
    .X(_0553_));
 sky130_fd_sc_hd__a31o_4 _3882_ (.A1(_0090_),
    .A2(_0549_),
    .A3(_0553_),
    .B1(_0545_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 ));
 sky130_fd_sc_hd__mux4_2 _3883_ (.A0(_0058_),
    .A1(_0059_),
    .A2(_0023_),
    .A3(_0537_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_0554_));
 sky130_fd_sc_hd__nand2_1 _3884_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ),
    .B(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__o211a_4 _3885_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ),
    .B1(_0555_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q ),
    .X(_0556_));
 sky130_fd_sc_hd__a211o_4 _3886_ (.A1(_0448_),
    .A2(_0446_),
    .B1(_0452_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ),
    .X(_0557_));
 sky130_fd_sc_hd__a21oi_2 _3887_ (.A1(_0052_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ),
    .Y(_0558_));
 sky130_fd_sc_hd__mux2_1 _3888_ (.A0(net76),
    .A1(net112),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ),
    .X(_0559_));
 sky130_fd_sc_hd__a22oi_4 _3889_ (.A1(_0557_),
    .A2(_0558_),
    .B1(_0559_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ),
    .Y(_0560_));
 sky130_fd_sc_hd__a221o_2 _3890_ (.A1(_0558_),
    .A2(_0557_),
    .B1(_0559_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ),
    .C1(_0088_),
    .X(_0561_));
 sky130_fd_sc_hd__o21ba_1 _3891_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ),
    .A2(net1052),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q ),
    .X(_0562_));
 sky130_fd_sc_hd__a21o_4 _3892_ (.A1(_0561_),
    .A2(_0562_),
    .B1(_0556_),
    .X(_0563_));
 sky130_fd_sc_hd__a211o_1 _3893_ (.A1(_0562_),
    .A2(_0561_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .C1(_0556_),
    .X(_0564_));
 sky130_fd_sc_hd__a21oi_1 _3894_ (.A1(_0071_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .Y(_0565_));
 sky130_fd_sc_hd__mux2_1 _3895_ (.A0(net211),
    .A1(net1072),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .X(_0566_));
 sky130_fd_sc_hd__a221o_1 _3896_ (.A1(_0565_),
    .A2(_0564_),
    .B1(_0566_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .C1(_0091_),
    .X(_0567_));
 sky130_fd_sc_hd__mux4_1 _3897_ (.A0(net175),
    .A1(net183),
    .A2(net120),
    .A3(net128),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0568_));
 sky130_fd_sc_hd__o21ba_1 _3898_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .A2(_0568_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q ),
    .X(_0569_));
 sky130_fd_sc_hd__a21o_4 _3899_ (.A1(_0569_),
    .A2(_0567_),
    .B1(_0541_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ));
 sky130_fd_sc_hd__inv_1 _3900_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .Y(_0570_));
 sky130_fd_sc_hd__mux4_2 _3901_ (.A0(_0570_),
    .A1(_0093_),
    .A2(_0092_),
    .A3(_0537_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q ),
    .X(_0571_));
 sky130_fd_sc_hd__mux4_1 _3902_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .A1(net109),
    .A2(net17),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q ),
    .X(_0572_));
 sky130_fd_sc_hd__a21oi_1 _3903_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_0359_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q ),
    .Y(_0573_));
 sky130_fd_sc_hd__o21a_2 _3904_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_0572_),
    .B1(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__or2_1 _3905_ (.A(_0529_),
    .B(_0574_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X ));
 sky130_fd_sc_hd__nand2b_1 _3906_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[6] ),
    .B(net1060),
    .Y(_0575_));
 sky130_fd_sc_hd__o31ai_4 _3907_ (.A1(net1060),
    .A2(_0574_),
    .A3(_0529_),
    .B1(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__a211o_1 _3908_ (.A1(_0561_),
    .A2(_0562_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .C1(_0556_),
    .X(_0577_));
 sky130_fd_sc_hd__a211o_1 _3909_ (.A1(_0360_),
    .A2(_0361_),
    .B1(_0386_),
    .C1(_0131_),
    .X(_0578_));
 sky130_fd_sc_hd__mux2_1 _3910_ (.A0(net74),
    .A1(net211),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0579_));
 sky130_fd_sc_hd__a21o_1 _3911_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .A2(_0579_),
    .B1(_0133_),
    .X(_0580_));
 sky130_fd_sc_hd__a31o_4 _3912_ (.A1(_0578_),
    .A2(_0577_),
    .A3(_0132_),
    .B1(_0580_),
    .X(_0581_));
 sky130_fd_sc_hd__mux4_1 _3913_ (.A0(net175),
    .A1(net183),
    .A2(net120),
    .A3(net128),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0582_));
 sky130_fd_sc_hd__o21ba_1 _3914_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .A2(_0582_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0583_));
 sky130_fd_sc_hd__mux4_2 _3915_ (.A0(net995),
    .A1(net1025),
    .A2(net1005),
    .A3(net653),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0584_));
 sky130_fd_sc_hd__mux4_1 _3916_ (.A0(net655),
    .A1(net971),
    .A2(net980),
    .A3(net1001),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0585_));
 sky130_fd_sc_hd__or2_1 _3917_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .B(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__o211a_4 _3918_ (.A1(_0584_),
    .A2(_0133_),
    .B1(_0586_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0587_));
 sky130_fd_sc_hd__a21oi_4 _3919_ (.A1(_0581_),
    .A2(_0583_),
    .B1(_0587_),
    .Y(_0588_));
 sky130_fd_sc_hd__a211o_1 _3920_ (.A1(_0583_),
    .A2(_0581_),
    .B1(_0587_),
    .C1(_0130_),
    .X(_0589_));
 sky130_fd_sc_hd__or2_1 _3921_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .B(net222),
    .X(_0590_));
 sky130_fd_sc_hd__mux4_2 _3922_ (.A0(net1037),
    .A1(net1031),
    .A2(net982),
    .A3(net1040),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_0591_));
 sky130_fd_sc_hd__nor2_2 _3923_ (.A(_0591_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ),
    .Y(_0592_));
 sky130_fd_sc_hd__mux4_1 _3924_ (.A0(net1051),
    .A1(net1046),
    .A2(net824),
    .A3(net822),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_0593_));
 sky130_fd_sc_hd__o21ai_1 _3925_ (.A1(_0085_),
    .A2(_0593_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q ),
    .Y(_0594_));
 sky130_fd_sc_hd__mux4_1 _3926_ (.A0(net62),
    .A1(net78),
    .A2(net98),
    .A3(net114),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_0595_));
 sky130_fd_sc_hd__nor2_1 _3927_ (.A(_0085_),
    .B(_0595_),
    .Y(_0596_));
 sky130_fd_sc_hd__mux4_1 _3928_ (.A0(net207),
    .A1(net1263),
    .A2(net6),
    .A3(net1261),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_0597_));
 sky130_fd_sc_hd__nor2_1 _3929_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ),
    .B(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__o32a_4 _3930_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q ),
    .A2(_0596_),
    .A3(_0598_),
    .B1(_0594_),
    .B2(_0592_),
    .X(_0599_));
 sky130_fd_sc_hd__inv_2 _3931_ (.A(_0599_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ));
 sky130_fd_sc_hd__nor2_1 _3932_ (.A(net186),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .Y(_0600_));
 sky130_fd_sc_hd__a211oi_1 _3933_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .A2(_0599_),
    .B1(_0600_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .Y(_0601_));
 sky130_fd_sc_hd__a311o_1 _3934_ (.A1(_0589_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .A3(_0590_),
    .B1(_0601_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ),
    .X(_0602_));
 sky130_fd_sc_hd__a21oi_1 _3935_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ),
    .A2(_0215_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q ),
    .Y(_0603_));
 sky130_fd_sc_hd__mux2_1 _3936_ (.A0(net230),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_1 _3937_ (.A0(net194),
    .A1(net89),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .X(_0605_));
 sky130_fd_sc_hd__inv_2 _3938_ (.A(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__o21ai_1 _3939_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q ),
    .A2(_0606_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ),
    .Y(_0607_));
 sky130_fd_sc_hd__a21o_1 _3940_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q ),
    .A2(_0604_),
    .B1(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__mux4_2 _3941_ (.A0(net178),
    .A1(net69),
    .A2(net142),
    .A3(net214),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q ),
    .X(_0609_));
 sky130_fd_sc_hd__o211a_1 _3942_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ),
    .A2(_0609_),
    .B1(_0608_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q ),
    .X(_0610_));
 sky130_fd_sc_hd__a21o_1 _3943_ (.A1(_0602_),
    .A2(_0603_),
    .B1(_0610_),
    .X(\Tile_X0Y1_DSP_bot.B3 ));
 sky130_fd_sc_hd__a211o_4 _3944_ (.A1(_0603_),
    .A2(_0602_),
    .B1(_0610_),
    .C1(net1061),
    .X(_0611_));
 sky130_fd_sc_hd__nand2b_2 _3945_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[3] ),
    .B(net1061),
    .Y(_0612_));
 sky130_fd_sc_hd__nand2_1 _3946_ (.A(_0611_),
    .B(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hd__nor2_4 _3947_ (.A(_0613_),
    .B(_0576_),
    .Y(_0614_));
 sky130_fd_sc_hd__nor2_1 _3948_ (.A(_0478_),
    .B(_0576_),
    .Y(_0615_));
 sky130_fd_sc_hd__nor2_4 _3949_ (.A(_0613_),
    .B(_0521_),
    .Y(_0616_));
 sky130_fd_sc_hd__nand2_4 _3950_ (.A(_0615_),
    .B(_0616_),
    .Y(_0617_));
 sky130_fd_sc_hd__mux2_2 _3951_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .A1(net819),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _3952_ (.A0(net186),
    .A1(net131),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .X(_0619_));
 sky130_fd_sc_hd__and2b_1 _3953_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q ),
    .B(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__a211o_1 _3954_ (.A1(_0618_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q ),
    .B1(_0620_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ),
    .X(_0621_));
 sky130_fd_sc_hd__mux2_1 _3955_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .A1(net223),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q ),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_1 _3956_ (.A0(net187),
    .A1(net132),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q ),
    .X(_0623_));
 sky130_fd_sc_hd__and2b_1 _3957_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q ),
    .B(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__a211o_1 _3958_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q ),
    .A2(_0622_),
    .B1(_0624_),
    .C1(_0122_),
    .X(_0625_));
 sky130_fd_sc_hd__mux4_2 _3959_ (.A0(net973),
    .A1(net977),
    .A2(net830),
    .A3(net987),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0626_));
 sky130_fd_sc_hd__or2_4 _3960_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .B(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__mux4_1 _3961_ (.A0(net992),
    .A1(net1021),
    .A2(net1002),
    .A3(net1010),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0628_));
 sky130_fd_sc_hd__o21a_1 _3962_ (.A1(_0123_),
    .A2(_0628_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .X(_0629_));
 sky130_fd_sc_hd__mux4_1 _3963_ (.A0(net174),
    .A1(net180),
    .A2(net125),
    .A3(net1222),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0630_));
 sky130_fd_sc_hd__mux4_1 _3964_ (.A0(net71),
    .A1(net216),
    .A2(net83),
    .A3(net230),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_1 _3965_ (.A0(_0630_),
    .A1(_0631_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .X(_0632_));
 sky130_fd_sc_hd__a22o_1 _3966_ (.A1(_0629_),
    .A2(_0627_),
    .B1(_0632_),
    .B2(_0124_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ));
 sky130_fd_sc_hd__mux2_1 _3967_ (.A0(net81),
    .A1(net818),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q ),
    .X(_0633_));
 sky130_fd_sc_hd__or2_1 _3968_ (.A(net194),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q ),
    .X(_0634_));
 sky130_fd_sc_hd__a21oi_1 _3969_ (.A1(_0020_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q ),
    .Y(_0635_));
 sky130_fd_sc_hd__a221o_1 _3970_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q ),
    .A2(_0633_),
    .B1(_0634_),
    .B2(_0635_),
    .C1(_0122_),
    .X(_0636_));
 sky130_fd_sc_hd__mux4_2 _3971_ (.A0(net178),
    .A1(net69),
    .A2(net123),
    .A3(net235),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q ),
    .X(_0637_));
 sky130_fd_sc_hd__o211a_1 _3972_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ),
    .A2(_0637_),
    .B1(_0636_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q ),
    .X(_0638_));
 sky130_fd_sc_hd__a31o_4 _3973_ (.A1(_0621_),
    .A2(_0125_),
    .A3(_0625_),
    .B1(_0638_),
    .X(\Tile_X0Y1_DSP_bot.A3 ));
 sky130_fd_sc_hd__nand2b_1 _3974_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[3] ),
    .B(net1059),
    .Y(_0639_));
 sky130_fd_sc_hd__o21ai_4 _3975_ (.A1(net1059),
    .A2(\Tile_X0Y1_DSP_bot.A3 ),
    .B1(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__inv_2 _3976_ (.A(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__mux4_2 _3977_ (.A0(net1017),
    .A1(net823),
    .A2(net865),
    .A3(net867),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0642_));
 sky130_fd_sc_hd__mux4_2 _3978_ (.A0(net1050),
    .A1(net1045),
    .A2(net824),
    .A3(net1016),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0643_));
 sky130_fd_sc_hd__or2_4 _3979_ (.A(_0643_),
    .B(_0073_),
    .X(_0644_));
 sky130_fd_sc_hd__o211a_1 _3980_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ),
    .A2(_0642_),
    .B1(_0644_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0645_));
 sky130_fd_sc_hd__or2_1 _3981_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .B(_0279_),
    .X(_0646_));
 sky130_fd_sc_hd__a21oi_1 _3982_ (.A1(_0048_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .Y(_0647_));
 sky130_fd_sc_hd__mux2_1 _3983_ (.A0(net8),
    .A1(net1261),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .X(_0648_));
 sky130_fd_sc_hd__a221o_1 _3984_ (.A1(_0646_),
    .A2(_0647_),
    .B1(_0648_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ),
    .X(_0649_));
 sky130_fd_sc_hd__nor2_1 _3985_ (.A(net64),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .Y(_0650_));
 sky130_fd_sc_hd__a211oi_1 _3986_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .A2(_0072_),
    .B1(_0650_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .Y(_0651_));
 sky130_fd_sc_hd__mux2_1 _3987_ (.A0(net100),
    .A1(net114),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .X(_0652_));
 sky130_fd_sc_hd__a211o_1 _3988_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .A2(_0652_),
    .B1(_0651_),
    .C1(_0073_),
    .X(_0653_));
 sky130_fd_sc_hd__a31o_1 _3989_ (.A1(_0074_),
    .A2(_0649_),
    .A3(_0653_),
    .B1(_0645_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ));
 sky130_fd_sc_hd__mux2_4 _3990_ (.A0(net113),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _3991_ (.A0(net198),
    .A1(net85),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ),
    .X(_0655_));
 sky130_fd_sc_hd__inv_1 _3992_ (.A(_0655_),
    .Y(_0656_));
 sky130_fd_sc_hd__o21ai_1 _3993_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q ),
    .A2(_0656_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ),
    .Y(_0657_));
 sky130_fd_sc_hd__a21o_1 _3994_ (.A1(_0654_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q ),
    .B1(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__mux4_2 _3995_ (.A0(net186),
    .A1(net61),
    .A2(net24),
    .A3(net97),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q ),
    .X(_0659_));
 sky130_fd_sc_hd__o211a_1 _3996_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_0659_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q ),
    .C1(_0658_),
    .X(_0660_));
 sky130_fd_sc_hd__nand2_1 _3997_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q ),
    .B(_0314_),
    .Y(_0661_));
 sky130_fd_sc_hd__o21a_1 _3998_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q ),
    .A2(net105),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q ),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_1 _3999_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .A1(net69),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q ),
    .X(_0663_));
 sky130_fd_sc_hd__a221o_1 _4000_ (.A1(_0662_),
    .A2(_0661_),
    .B1(_0663_),
    .B2(_0106_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ),
    .X(_0664_));
 sky130_fd_sc_hd__nand2b_1 _4001_ (.A_N(_0439_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ),
    .Y(_0665_));
 sky130_fd_sc_hd__a31o_4 _4002_ (.A1(_0664_),
    .A2(_0107_),
    .A3(_0665_),
    .B1(_0660_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X ));
 sky130_fd_sc_hd__nand2b_1 _4003_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[7] ),
    .B(net1062),
    .Y(_0666_));
 sky130_fd_sc_hd__o21ai_4 _4004_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X ),
    .A2(net1062),
    .B1(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__nor2_8 _4005_ (.A(_0667_),
    .B(_0640_),
    .Y(_0668_));
 sky130_fd_sc_hd__mux4_1 _4006_ (.A0(net1019),
    .A1(net1038),
    .A2(net986),
    .A3(net1041),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0669_));
 sky130_fd_sc_hd__nand2b_1 _4007_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ),
    .B(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__mux4_1 _4008_ (.A0(net1052),
    .A1(net1046),
    .A2(net1027),
    .A3(net1057),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0671_));
 sky130_fd_sc_hd__nand2_1 _4009_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ),
    .B(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__mux4_1 _4010_ (.A0(net209),
    .A1(net2),
    .A2(net8),
    .A3(net1261),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0673_));
 sky130_fd_sc_hd__mux4_1 _4011_ (.A0(net64),
    .A1(net100),
    .A2(net80),
    .A3(net114),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _4012_ (.A0(_0673_),
    .A1(_0674_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ),
    .X(_0675_));
 sky130_fd_sc_hd__nor2_1 _4013_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q ),
    .B(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__a31o_4 _4014_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q ),
    .A2(_0670_),
    .A3(_0672_),
    .B1(_0676_),
    .X(_0677_));
 sky130_fd_sc_hd__inv_2 _4015_ (.A(_0677_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ));
 sky130_fd_sc_hd__nand2_1 _4016_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ),
    .B(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__o211a_1 _4017_ (.A1(net78),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q ),
    .C1(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_1 _4018_ (.A0(net207),
    .A1(net24),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ),
    .X(_0680_));
 sky130_fd_sc_hd__inv_2 _4019_ (.A(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hd__o21ai_1 _4020_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q ),
    .A2(_0681_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q ),
    .Y(_0682_));
 sky130_fd_sc_hd__mux4_2 _4021_ (.A0(net190),
    .A1(net9),
    .A2(net87),
    .A3(net101),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q ),
    .X(_0683_));
 sky130_fd_sc_hd__o221a_1 _4022_ (.A1(_0679_),
    .A2(_0682_),
    .B1(_0683_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q ),
    .X(_0684_));
 sky130_fd_sc_hd__mux4_2 _4023_ (.A0(net1018),
    .A1(net1036),
    .A2(net1032),
    .A3(net983),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0685_));
 sky130_fd_sc_hd__and2_4 _4024_ (.A(_0105_),
    .B(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__mux4_1 _4025_ (.A0(net1053),
    .A1(net1048),
    .A2(net1028),
    .A3(net1058),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0687_));
 sky130_fd_sc_hd__a21bo_1 _4026_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(_0687_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q ),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_4 _4027_ (.A0(_0279_),
    .A1(net191),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_1 _4028_ (.A0(net2),
    .A1(net10),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .X(_0690_));
 sky130_fd_sc_hd__or2_1 _4029_ (.A(_0104_),
    .B(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__o211a_1 _4030_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .A2(_0689_),
    .B1(_0691_),
    .C1(_0105_),
    .X(_0692_));
 sky130_fd_sc_hd__mux2_1 _4031_ (.A0(net58),
    .A1(net66),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .X(_0693_));
 sky130_fd_sc_hd__or2_1 _4032_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .B(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__mux2_1 _4033_ (.A0(net94),
    .A1(net1225),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .X(_0695_));
 sky130_fd_sc_hd__o211a_1 _4034_ (.A1(_0104_),
    .A2(_0695_),
    .B1(_0694_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ),
    .X(_0696_));
 sky130_fd_sc_hd__o32a_4 _4035_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q ),
    .A2(_0692_),
    .A3(_0696_),
    .B1(_0686_),
    .B2(_0688_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ));
 sky130_fd_sc_hd__mux2_1 _4036_ (.A0(net73),
    .A1(net654),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ),
    .X(_0697_));
 sky130_fd_sc_hd__a211o_1 _4037_ (.A1(_0569_),
    .A2(_0567_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ),
    .C1(_0541_),
    .X(_0698_));
 sky130_fd_sc_hd__a21oi_1 _4038_ (.A1(_0092_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q ),
    .Y(_0699_));
 sky130_fd_sc_hd__a22o_4 _4039_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q ),
    .A2(_0697_),
    .B1(_0699_),
    .B2(_0698_),
    .X(_0700_));
 sky130_fd_sc_hd__inv_2 _4040_ (.A(_0700_),
    .Y(_0701_));
 sky130_fd_sc_hd__a221o_1 _4041_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q ),
    .A2(_0697_),
    .B1(_0698_),
    .B2(_0699_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q ),
    .X(_0702_));
 sky130_fd_sc_hd__nor2_1 _4042_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .Y(_0703_));
 sky130_fd_sc_hd__a211o_1 _4043_ (.A1(_0070_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q ),
    .C1(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_1 _4044_ (.A0(net74),
    .A1(net110),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q ),
    .X(_0705_));
 sky130_fd_sc_hd__nand2_1 _4045_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q ),
    .B(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__a31oi_1 _4046_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q ),
    .A2(_0704_),
    .A3(_0706_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q ),
    .Y(_0707_));
 sky130_fd_sc_hd__a21o_1 _4047_ (.A1(_0702_),
    .A2(_0707_),
    .B1(_0684_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X ));
 sky130_fd_sc_hd__a211o_1 _4048_ (.A1(_0702_),
    .A2(_0707_),
    .B1(net1062),
    .C1(_0684_),
    .X(_0708_));
 sky130_fd_sc_hd__nand2b_1 _4049_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[6] ),
    .B(net1062),
    .Y(_0709_));
 sky130_fd_sc_hd__nand2_2 _4050_ (.A(_0708_),
    .B(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__mux4_2 _4051_ (.A0(_0022_),
    .A1(_0126_),
    .A2(_0127_),
    .A3(_0267_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q ),
    .X(_0711_));
 sky130_fd_sc_hd__mux4_2 _4052_ (.A0(net190),
    .A1(net135),
    .A2(net226),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q ),
    .X(_0712_));
 sky130_fd_sc_hd__mux4_2 _4053_ (.A0(net811),
    .A1(net664),
    .A2(net997),
    .A3(net987),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0713_));
 sky130_fd_sc_hd__or2_4 _4054_ (.A(_0713_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_0714_));
 sky130_fd_sc_hd__mux4_1 _4055_ (.A0(net992),
    .A1(net1021),
    .A2(net1002),
    .A3(net1007),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0715_));
 sky130_fd_sc_hd__o21a_1 _4056_ (.A1(_0128_),
    .A2(_0715_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q ),
    .X(_0716_));
 sky130_fd_sc_hd__mux4_1 _4057_ (.A0(net204),
    .A1(net143),
    .A2(net119),
    .A3(net1222),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .X(_0717_));
 sky130_fd_sc_hd__mux4_1 _4058_ (.A0(net83),
    .A1(net91),
    .A2(net216),
    .A3(net230),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0718_));
 sky130_fd_sc_hd__mux2_1 _4059_ (.A0(_0717_),
    .A1(_0718_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_0719_));
 sky130_fd_sc_hd__a22o_1 _4060_ (.A1(_0716_),
    .A2(_0714_),
    .B1(_0719_),
    .B2(_0129_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ));
 sky130_fd_sc_hd__mux4_2 _4061_ (.A0(net195),
    .A1(net231),
    .A2(net1221),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q ),
    .X(_0720_));
 sky130_fd_sc_hd__mux4_2 _4062_ (.A0(net182),
    .A1(net73),
    .A2(net141),
    .A3(net218),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q ),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_4 _4063_ (.A0(_0721_),
    .A1(_0720_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ),
    .X(_0722_));
 sky130_fd_sc_hd__mux2_1 _4064_ (.A0(_0712_),
    .A1(net816),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ),
    .X(_0723_));
 sky130_fd_sc_hd__mux2_4 _4065_ (.A0(_0723_),
    .A1(_0722_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q ),
    .X(\Tile_X0Y1_DSP_bot.A2 ));
 sky130_fd_sc_hd__and2b_1 _4066_ (.A_N(net1059),
    .B(\Tile_X0Y1_DSP_bot.A2 ),
    .X(_0724_));
 sky130_fd_sc_hd__a21o_1 _4067_ (.A1(net1059),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[2] ),
    .B1(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__a21oi_4 _4068_ (.A1(net1059),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[2] ),
    .B1(_0724_),
    .Y(_0726_));
 sky130_fd_sc_hd__and3_1 _4069_ (.A(_0708_),
    .B(_0709_),
    .C(_0725_),
    .X(_0727_));
 sky130_fd_sc_hd__and3_4 _4070_ (.A(_0641_),
    .B(_0708_),
    .C(_0709_),
    .X(_0728_));
 sky130_fd_sc_hd__nor2_1 _4071_ (.A(_0667_),
    .B(_0726_),
    .Y(_0729_));
 sky130_fd_sc_hd__mux4_2 _4072_ (.A0(net815),
    .A1(net1036),
    .A2(net1032),
    .A3(net983),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0730_));
 sky130_fd_sc_hd__nand2b_4 _4073_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ),
    .B(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__mux4_1 _4074_ (.A0(net1053),
    .A1(net1048),
    .A2(net1028),
    .A3(net1014),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0732_));
 sky130_fd_sc_hd__nand2_1 _4075_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ),
    .B(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__mux2_1 _4076_ (.A0(_0279_),
    .A1(net191),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0734_));
 sky130_fd_sc_hd__nor2_1 _4077_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .B(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__mux2_1 _4078_ (.A0(net2),
    .A1(net10),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0736_));
 sky130_fd_sc_hd__inv_1 _4079_ (.A(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__a211o_1 _4080_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .A2(_0737_),
    .B1(_0735_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _4081_ (.A0(net58),
    .A1(net60),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0739_));
 sky130_fd_sc_hd__or2_1 _4082_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .B(_0739_),
    .X(_0740_));
 sky130_fd_sc_hd__mux2_1 _4083_ (.A0(net66),
    .A1(net94),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0741_));
 sky130_fd_sc_hd__o211a_1 _4084_ (.A1(_0101_),
    .A2(_0741_),
    .B1(_0740_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ),
    .X(_0742_));
 sky130_fd_sc_hd__nor2_1 _4085_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q ),
    .B(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__a32o_2 _4086_ (.A1(_0733_),
    .A2(_0731_),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q ),
    .B1(_0738_),
    .B2(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__inv_1 _4087_ (.A(_0744_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ));
 sky130_fd_sc_hd__nand2_2 _4088_ (.A(_0744_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q ),
    .Y(_0745_));
 sky130_fd_sc_hd__o21a_1 _4089_ (.A1(net107),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q ),
    .X(_0746_));
 sky130_fd_sc_hd__mux4_1 _4090_ (.A0(net993),
    .A1(net1022),
    .A2(net1003),
    .A3(net1010),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0747_));
 sky130_fd_sc_hd__or2_1 _4091_ (.A(_0099_),
    .B(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__mux4_1 _4092_ (.A0(net975),
    .A1(net869),
    .A2(net999),
    .A3(net988),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0749_));
 sky130_fd_sc_hd__o21a_1 _4093_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .A2(_0749_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q ),
    .X(_0750_));
 sky130_fd_sc_hd__mux4_1 _4094_ (.A0(net140),
    .A1(net72),
    .A2(net217),
    .A3(net233),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0751_));
 sky130_fd_sc_hd__mux4_1 _4095_ (.A0(net181),
    .A1(net197),
    .A2(net120),
    .A3(net126),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0752_));
 sky130_fd_sc_hd__mux2_1 _4096_ (.A0(_0751_),
    .A1(_0752_),
    .S(_0099_),
    .X(_0753_));
 sky130_fd_sc_hd__a22o_4 _4097_ (.A1(_0748_),
    .A2(_0750_),
    .B1(_0753_),
    .B2(_0100_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ));
 sky130_fd_sc_hd__mux2_1 _4098_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .A1(net15),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q ),
    .X(_0754_));
 sky130_fd_sc_hd__a221o_1 _4099_ (.A1(_0746_),
    .A2(_0745_),
    .B1(_0754_),
    .B2(_0102_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ),
    .X(_0755_));
 sky130_fd_sc_hd__mux4_2 _4100_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .A1(net16),
    .A2(net72),
    .A3(net108),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q ),
    .X(_0756_));
 sky130_fd_sc_hd__nand2b_1 _4101_ (.A_N(_0756_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ),
    .Y(_0757_));
 sky130_fd_sc_hd__nand2_1 _4102_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ),
    .B(_0428_),
    .Y(_0758_));
 sky130_fd_sc_hd__mux4_2 _4103_ (.A0(net188),
    .A1(net63),
    .A2(net7),
    .A3(net117),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q ),
    .X(_0759_));
 sky130_fd_sc_hd__o211a_1 _4104_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ),
    .A2(_0759_),
    .B1(_0758_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q ),
    .X(_0760_));
 sky130_fd_sc_hd__a31o_4 _4105_ (.A1(_0755_),
    .A2(_0103_),
    .A3(_0757_),
    .B1(_0760_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X ));
 sky130_fd_sc_hd__nand2b_1 _4106_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[5] ),
    .B(net1062),
    .Y(_0761_));
 sky130_fd_sc_hd__o21ai_4 _4107_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X ),
    .A2(net1061),
    .B1(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__nand2_2 _4108_ (.A(_0384_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ),
    .Y(_0763_));
 sky130_fd_sc_hd__mux4_2 _4109_ (.A0(net192),
    .A1(net11),
    .A2(net88),
    .A3(net103),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q ),
    .X(_0764_));
 sky130_fd_sc_hd__o211a_1 _4110_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ),
    .A2(_0764_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q ),
    .C1(_0763_),
    .X(_0765_));
 sky130_fd_sc_hd__a211o_1 _4111_ (.A1(_0391_),
    .A2(_0393_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ),
    .C1(_0298_),
    .X(_0766_));
 sky130_fd_sc_hd__a21oi_1 _4112_ (.A1(_0068_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q ),
    .Y(_0767_));
 sky130_fd_sc_hd__mux4_1 _4113_ (.A0(net1017),
    .A1(net1037),
    .A2(net1031),
    .A3(net1041),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0768_));
 sky130_fd_sc_hd__or2_1 _4114_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ),
    .B(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__mux4_1 _4115_ (.A0(net1051),
    .A1(net1045),
    .A2(net1027),
    .A3(net1016),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0770_));
 sky130_fd_sc_hd__o21a_1 _4116_ (.A1(_0079_),
    .A2(_0770_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q ),
    .X(_0771_));
 sky130_fd_sc_hd__mux4_1 _4117_ (.A0(net190),
    .A1(net198),
    .A2(net1264),
    .A3(net9),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0772_));
 sky130_fd_sc_hd__mux4_1 _4118_ (.A0(net1262),
    .A1(net65),
    .A2(net101),
    .A3(net113),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0773_));
 sky130_fd_sc_hd__mux2_1 _4119_ (.A0(_0772_),
    .A1(_0773_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ),
    .X(_0774_));
 sky130_fd_sc_hd__a22o_2 _4120_ (.A1(_0769_),
    .A2(_0771_),
    .B1(_0774_),
    .B2(_0080_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ));
 sky130_fd_sc_hd__mux2_1 _4121_ (.A0(net111),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ),
    .X(_0775_));
 sky130_fd_sc_hd__a221o_1 _4122_ (.A1(_0766_),
    .A2(_0767_),
    .B1(_0775_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ),
    .X(_0776_));
 sky130_fd_sc_hd__mux2_1 _4123_ (.A0(_0453_),
    .A1(_0052_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q ),
    .X(_0777_));
 sky130_fd_sc_hd__mux2_1 _4124_ (.A0(net76),
    .A1(net112),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q ),
    .X(_0778_));
 sky130_fd_sc_hd__nand2_1 _4125_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q ),
    .B(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hd__o211a_1 _4126_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q ),
    .A2(_0777_),
    .B1(_0779_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ),
    .X(_0780_));
 sky130_fd_sc_hd__nor2_1 _4127_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q ),
    .B(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hd__a21o_1 _4128_ (.A1(_0776_),
    .A2(_0781_),
    .B1(_0765_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X ));
 sky130_fd_sc_hd__a211o_4 _4129_ (.A1(_0776_),
    .A2(_0781_),
    .B1(net1060),
    .C1(_0765_),
    .X(_0782_));
 sky130_fd_sc_hd__nand2b_1 _4130_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[4] ),
    .B(net1060),
    .Y(_0783_));
 sky130_fd_sc_hd__nand2_8 _4131_ (.A(_0782_),
    .B(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__or2_1 _4132_ (.A(net622),
    .B(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__xnor2_4 _4133_ (.A(_0729_),
    .B(_0728_),
    .Y(_0786_));
 sky130_fd_sc_hd__o2bb2a_4 _4134_ (.A1_N(_0728_),
    .A2_N(_0729_),
    .B1(_0785_),
    .B2(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__mux4_2 _4135_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .A1(net16),
    .A2(net72),
    .A3(net108),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q ),
    .X(_0788_));
 sky130_fd_sc_hd__mux4_1 _4136_ (.A0(net15),
    .A1(net107),
    .A2(net71),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q ),
    .X(_0789_));
 sky130_fd_sc_hd__mux2_1 _4137_ (.A0(_0789_),
    .A1(_0788_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ),
    .X(_0790_));
 sky130_fd_sc_hd__mux2_1 _4138_ (.A0(net104),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q ),
    .X(_0791_));
 sky130_fd_sc_hd__mux2_1 _4139_ (.A0(net25),
    .A1(net79),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q ),
    .X(_0792_));
 sky130_fd_sc_hd__inv_1 _4140_ (.A(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hd__o21ai_1 _4141_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q ),
    .A2(_0793_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ),
    .Y(_0794_));
 sky130_fd_sc_hd__a21o_1 _4142_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q ),
    .A2(_0791_),
    .B1(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__mux4_2 _4143_ (.A0(net206),
    .A1(net63),
    .A2(net7),
    .A3(net99),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q ),
    .X(_0796_));
 sky130_fd_sc_hd__o21a_1 _4144_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ),
    .A2(_0796_),
    .B1(_0795_),
    .X(_0797_));
 sky130_fd_sc_hd__mux2_2 _4145_ (.A0(_0790_),
    .A1(_0797_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X ));
 sky130_fd_sc_hd__nand2b_1 _4146_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[5] ),
    .B(net1059),
    .Y(_0798_));
 sky130_fd_sc_hd__o21ai_4 _4147_ (.A1(net1059),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X ),
    .B1(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__or2_4 _4148_ (.A(_0799_),
    .B(net622),
    .X(_0800_));
 sky130_fd_sc_hd__nor2_1 _4149_ (.A(_0710_),
    .B(_0784_),
    .Y(_0801_));
 sky130_fd_sc_hd__xnor2_4 _4150_ (.A(_0801_),
    .B(_0668_),
    .Y(_0802_));
 sky130_fd_sc_hd__xnor2_2 _4151_ (.A(_0802_),
    .B(_0800_),
    .Y(_0803_));
 sky130_fd_sc_hd__nor2_1 _4152_ (.A(_0803_),
    .B(_0787_),
    .Y(_0804_));
 sky130_fd_sc_hd__xnor2_1 _4153_ (.A(_0787_),
    .B(_0803_),
    .Y(_0805_));
 sky130_fd_sc_hd__or2_1 _4154_ (.A(_0615_),
    .B(_0616_),
    .X(_0806_));
 sky130_fd_sc_hd__nand2_4 _4155_ (.A(_0617_),
    .B(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__o21bai_4 _4156_ (.A1(_0805_),
    .A2(_0807_),
    .B1_N(_0804_),
    .Y(_0808_));
 sky130_fd_sc_hd__o2bb2ai_4 _4157_ (.A1_N(_0668_),
    .A2_N(_0801_),
    .B1(_0800_),
    .B2(_0802_),
    .Y(_0809_));
 sky130_fd_sc_hd__nor2_1 _4158_ (.A(_0667_),
    .B(_0799_),
    .Y(_0810_));
 sky130_fd_sc_hd__nand2_1 _4159_ (.A(_0801_),
    .B(_0810_),
    .Y(_0811_));
 sky130_fd_sc_hd__o22a_1 _4160_ (.A1(_0667_),
    .A2(_0784_),
    .B1(_0799_),
    .B2(_0710_),
    .X(_0812_));
 sky130_fd_sc_hd__a21o_1 _4161_ (.A1(_0801_),
    .A2(_0810_),
    .B1(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__or3_1 _4162_ (.A(_0576_),
    .B(_0762_),
    .C(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__o21ai_1 _4163_ (.A1(_0576_),
    .A2(_0762_),
    .B1(_0813_),
    .Y(_0815_));
 sky130_fd_sc_hd__nand2_1 _4164_ (.A(_0814_),
    .B(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__and3_1 _4165_ (.A(_0814_),
    .B(_0809_),
    .C(_0815_),
    .X(_0817_));
 sky130_fd_sc_hd__xor2_1 _4166_ (.A(_0809_),
    .B(_0816_),
    .X(_0818_));
 sky130_fd_sc_hd__xnor2_1 _4167_ (.A(_0522_),
    .B(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hd__and2b_1 _4168_ (.A_N(_0819_),
    .B(_0808_),
    .X(_0820_));
 sky130_fd_sc_hd__xnor2_4 _4169_ (.A(_0819_),
    .B(_0808_),
    .Y(_0821_));
 sky130_fd_sc_hd__xnor2_4 _4170_ (.A(_0821_),
    .B(_0617_),
    .Y(_0822_));
 sky130_fd_sc_hd__mux4_2 _4171_ (.A0(net189),
    .A1(net134),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .A3(net225),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q ),
    .X(_0823_));
 sky130_fd_sc_hd__mux4_2 _4172_ (.A0(net811),
    .A1(net664),
    .A2(net997),
    .A3(net987),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0824_));
 sky130_fd_sc_hd__or2_4 _4173_ (.A(_0824_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_0825_));
 sky130_fd_sc_hd__mux4_1 _4174_ (.A0(net992),
    .A1(net1021),
    .A2(net1002),
    .A3(net1010),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0826_));
 sky130_fd_sc_hd__o21a_1 _4175_ (.A1(_0136_),
    .A2(_0826_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q ),
    .X(_0827_));
 sky130_fd_sc_hd__mux4_1 _4176_ (.A0(net174),
    .A1(net180),
    .A2(net196),
    .A3(net125),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0828_));
 sky130_fd_sc_hd__mux4_1 _4177_ (.A0(net1222),
    .A1(net71),
    .A2(net216),
    .A3(net235),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0829_));
 sky130_fd_sc_hd__mux2_1 _4178_ (.A0(_0828_),
    .A1(_0829_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_0830_));
 sky130_fd_sc_hd__a22o_4 _4179_ (.A1(_0827_),
    .A2(_0825_),
    .B1(_0830_),
    .B2(_0137_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ));
 sky130_fd_sc_hd__mux2_2 _4180_ (.A0(net221),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ),
    .X(_0831_));
 sky130_fd_sc_hd__mux2_1 _4181_ (.A0(net143),
    .A1(net83),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ),
    .X(_0832_));
 sky130_fd_sc_hd__inv_2 _4182_ (.A(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__mux4_1 _4183_ (.A0(net992),
    .A1(net1021),
    .A2(net1003),
    .A3(net1010),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_0834_));
 sky130_fd_sc_hd__mux4_1 _4184_ (.A0(net811),
    .A1(net869),
    .A2(net977),
    .A3(net988),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_0835_));
 sky130_fd_sc_hd__and2b_1 _4185_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .B(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__a21bo_1 _4186_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .A2(_0834_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_0837_));
 sky130_fd_sc_hd__mux4_1 _4187_ (.A0(net176),
    .A1(net182),
    .A2(net194),
    .A3(net127),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_0838_));
 sky130_fd_sc_hd__mux4_1 _4188_ (.A0(net1222),
    .A1(net73),
    .A2(net218),
    .A3(net230),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_1 _4189_ (.A0(_0838_),
    .A1(_0839_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .X(_0840_));
 sky130_fd_sc_hd__o22a_4 _4190_ (.A1(_0837_),
    .A2(_0836_),
    .B1(_0840_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ));
 sky130_fd_sc_hd__mux4_1 _4191_ (.A0(net202),
    .A1(net71),
    .A2(net125),
    .A3(net216),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q ),
    .X(_0841_));
 sky130_fd_sc_hd__mux4_1 _4192_ (.A0(net133),
    .A1(net224),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q ),
    .X(_0842_));
 sky130_fd_sc_hd__mux2_1 _4193_ (.A0(_0842_),
    .A1(_0823_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ),
    .X(_0843_));
 sky130_fd_sc_hd__o21ai_1 _4194_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q ),
    .A2(_0833_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ),
    .Y(_0844_));
 sky130_fd_sc_hd__a21o_1 _4195_ (.A1(_0831_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q ),
    .B1(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__o21a_1 _4196_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_0841_),
    .B1(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__mux2_4 _4197_ (.A0(_0843_),
    .A1(_0846_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q ),
    .X(\Tile_X0Y1_DSP_bot.A1 ));
 sky130_fd_sc_hd__mux2_4 _4198_ (.A0(\Tile_X0Y1_DSP_bot.A1 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[1] ),
    .S(net1059),
    .X(_0847_));
 sky130_fd_sc_hd__clkinv_2 _4199_ (.A(_0847_),
    .Y(_0848_));
 sky130_fd_sc_hd__nor2_1 _4200_ (.A(_0667_),
    .B(_0848_),
    .Y(_0849_));
 sky130_fd_sc_hd__or2_1 _4201_ (.A(_0640_),
    .B(_0762_),
    .X(_0850_));
 sky130_fd_sc_hd__xnor2_1 _4202_ (.A(_0727_),
    .B(_0849_),
    .Y(_0851_));
 sky130_fd_sc_hd__o2bb2a_1 _4203_ (.A1_N(_0727_),
    .A2_N(_0849_),
    .B1(_0850_),
    .B2(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__xnor2_1 _4204_ (.A(_0785_),
    .B(_0786_),
    .Y(_0853_));
 sky130_fd_sc_hd__or2_1 _4205_ (.A(_0852_),
    .B(_0853_),
    .X(_0854_));
 sky130_fd_sc_hd__xnor2_1 _4206_ (.A(_0852_),
    .B(_0853_),
    .Y(_0855_));
 sky130_fd_sc_hd__mux4_2 _4207_ (.A0(net811),
    .A1(net869),
    .A2(net997),
    .A3(net988),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0856_));
 sky130_fd_sc_hd__or2_4 _4208_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .B(_0856_),
    .X(_0857_));
 sky130_fd_sc_hd__mux4_1 _4209_ (.A0(net993),
    .A1(net1021),
    .A2(net1002),
    .A3(net1010),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0858_));
 sky130_fd_sc_hd__o21a_1 _4210_ (.A1(_0139_),
    .A2(_0858_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q ),
    .X(_0859_));
 sky130_fd_sc_hd__mux4_1 _4211_ (.A0(net72),
    .A1(net217),
    .A2(net84),
    .A3(net231),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_0860_));
 sky130_fd_sc_hd__mux4_1 _4212_ (.A0(net205),
    .A1(net120),
    .A2(net126),
    .A3(net1221),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0861_));
 sky130_fd_sc_hd__mux2_1 _4213_ (.A0(_0860_),
    .A1(_0861_),
    .S(_0139_),
    .X(_0862_));
 sky130_fd_sc_hd__a22o_4 _4214_ (.A1(_0857_),
    .A2(_0859_),
    .B1(_0862_),
    .B2(_0140_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ));
 sky130_fd_sc_hd__mux4_2 _4215_ (.A0(net203),
    .A1(net142),
    .A2(net82),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q ),
    .X(_0863_));
 sky130_fd_sc_hd__mux4_2 _4216_ (.A0(net182),
    .A1(net127),
    .A2(net91),
    .A3(net218),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q ),
    .X(_0864_));
 sky130_fd_sc_hd__mux4_1 _4217_ (.A0(net923),
    .A1(net971),
    .A2(net981),
    .A3(net1000),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0865_));
 sky130_fd_sc_hd__or2_1 _4218_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .B(_0865_),
    .X(_0866_));
 sky130_fd_sc_hd__mux4_1 _4219_ (.A0(net995),
    .A1(net1025),
    .A2(net1005),
    .A3(net1012),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0867_));
 sky130_fd_sc_hd__or2_1 _4220_ (.A(_0138_),
    .B(_0867_),
    .X(_0868_));
 sky130_fd_sc_hd__a211o_1 _4221_ (.A1(_0561_),
    .A2(_0562_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .C1(_0556_),
    .X(_0869_));
 sky130_fd_sc_hd__a21oi_1 _4222_ (.A1(_0071_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .Y(_0870_));
 sky130_fd_sc_hd__mux2_1 _4223_ (.A0(net211),
    .A1(net1072),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .X(_0871_));
 sky130_fd_sc_hd__a221o_1 _4224_ (.A1(_0869_),
    .A2(_0870_),
    .B1(_0871_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .C1(_0138_),
    .X(_0872_));
 sky130_fd_sc_hd__mux4_1 _4225_ (.A0(net175),
    .A1(net183),
    .A2(net120),
    .A3(net128),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0873_));
 sky130_fd_sc_hd__o21ba_1 _4226_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(_0873_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q ),
    .X(_0874_));
 sky130_fd_sc_hd__a32o_4 _4227_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q ),
    .A2(_0866_),
    .A3(_0868_),
    .B1(_0872_),
    .B2(_0874_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ));
 sky130_fd_sc_hd__mux4_2 _4228_ (.A0(net190),
    .A1(net135),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .X(_0875_));
 sky130_fd_sc_hd__mux4_1 _4229_ (.A0(net191),
    .A1(net136),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .A3(net227),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q ),
    .X(_0876_));
 sky130_fd_sc_hd__mux4_2 _4230_ (.A0(_0875_),
    .A1(_0876_),
    .A2(_0864_),
    .A3(_0863_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q ),
    .X(\Tile_X0Y1_DSP_bot.B2 ));
 sky130_fd_sc_hd__nand2b_1 _4231_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[2] ),
    .B(net1061),
    .Y(_0877_));
 sky130_fd_sc_hd__o21ai_4 _4232_ (.A1(net1061),
    .A2(\Tile_X0Y1_DSP_bot.B2 ),
    .B1(_0877_),
    .Y(_0878_));
 sky130_fd_sc_hd__or2_1 _4233_ (.A(_0521_),
    .B(_0878_),
    .X(_0879_));
 sky130_fd_sc_hd__nor2_1 _4234_ (.A(_0478_),
    .B(_0799_),
    .Y(_0880_));
 sky130_fd_sc_hd__nor2_1 _4235_ (.A(_0613_),
    .B(_0799_),
    .Y(_0881_));
 sky130_fd_sc_hd__xnor2_2 _4236_ (.A(_0880_),
    .B(_0614_),
    .Y(_0882_));
 sky130_fd_sc_hd__xnor2_1 _4237_ (.A(_0879_),
    .B(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__o21a_1 _4238_ (.A1(_0855_),
    .A2(_0883_),
    .B1(_0854_),
    .X(_0884_));
 sky130_fd_sc_hd__xor2_2 _4239_ (.A(_0805_),
    .B(_0807_),
    .X(_0885_));
 sky130_fd_sc_hd__nand2b_1 _4240_ (.A_N(_0884_),
    .B(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__o2bb2ai_1 _4241_ (.A1_N(_0614_),
    .A2_N(_0880_),
    .B1(_0882_),
    .B2(_0879_),
    .Y(_0887_));
 sky130_fd_sc_hd__xnor2_1 _4242_ (.A(_0884_),
    .B(_0885_),
    .Y(_0888_));
 sky130_fd_sc_hd__a21bo_1 _4243_ (.A1(_0887_),
    .A2(_0888_),
    .B1_N(_0886_),
    .X(_0889_));
 sky130_fd_sc_hd__nand2_2 _4244_ (.A(_0889_),
    .B(_0822_),
    .Y(_0890_));
 sky130_fd_sc_hd__or2_1 _4245_ (.A(_0521_),
    .B(_0762_),
    .X(_0891_));
 sky130_fd_sc_hd__nor2_1 _4246_ (.A(_0576_),
    .B(_0710_),
    .Y(_0892_));
 sky130_fd_sc_hd__inv_2 _4247_ (.A(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__xnor2_1 _4248_ (.A(_0810_),
    .B(_0892_),
    .Y(_0894_));
 sky130_fd_sc_hd__xnor2_1 _4249_ (.A(_0891_),
    .B(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__a21oi_1 _4250_ (.A1(_0811_),
    .A2(_0814_),
    .B1(_0895_),
    .Y(_0896_));
 sky130_fd_sc_hd__and3_1 _4251_ (.A(_0811_),
    .B(_0814_),
    .C(_0895_),
    .X(_0897_));
 sky130_fd_sc_hd__or2_1 _4252_ (.A(_0896_),
    .B(_0897_),
    .X(_0898_));
 sky130_fd_sc_hd__o21ba_4 _4253_ (.A1(_0522_),
    .A2(_0818_),
    .B1_N(_0817_),
    .X(_0899_));
 sky130_fd_sc_hd__nor2_8 _4254_ (.A(_0899_),
    .B(_0898_),
    .Y(_0900_));
 sky130_fd_sc_hd__xnor2_1 _4255_ (.A(_0898_),
    .B(_0899_),
    .Y(_0901_));
 sky130_fd_sc_hd__a31oi_4 _4256_ (.A1(_0615_),
    .A2(_0616_),
    .A3(_0821_),
    .B1(_0820_),
    .Y(_0902_));
 sky130_fd_sc_hd__nor2_2 _4257_ (.A(_0901_),
    .B(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__xnor2_2 _4258_ (.A(_0901_),
    .B(_0902_),
    .Y(_0904_));
 sky130_fd_sc_hd__nor2_1 _4259_ (.A(_0890_),
    .B(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hd__mux4_2 _4260_ (.A0(net184),
    .A1(net129),
    .A2(net92),
    .A3(net220),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q ),
    .X(_0906_));
 sky130_fd_sc_hd__mux2_1 _4261_ (.A0(_0906_),
    .A1(_0405_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_0907_));
 sky130_fd_sc_hd__mux2_4 _4262_ (.A0(net875),
    .A1(net229),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ),
    .X(_0908_));
 sky130_fd_sc_hd__mux2_1 _4263_ (.A0(net193),
    .A1(net138),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ),
    .X(_0909_));
 sky130_fd_sc_hd__inv_1 _4264_ (.A(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__o21ai_1 _4265_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q ),
    .A2(_0910_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ),
    .Y(_0911_));
 sky130_fd_sc_hd__dlxtp_1 _4266_ (.D(net1234),
    .GATE(net1183),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4267_ (.D(net1235),
    .GATE(net1183),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4268_ (.D(net1237),
    .GATE(net1183),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4269_ (.D(net1238),
    .GATE(net1183),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4270_ (.D(net44),
    .GATE(net1184),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4271_ (.D(net43),
    .GATE(net1184),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4272_ (.D(net1242),
    .GATE(net1184),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4273_ (.D(net1243),
    .GATE(net1184),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4274_ (.D(net42),
    .GATE(net1183),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4275_ (.D(net1246),
    .GATE(net1185),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4276_ (.D(net1247),
    .GATE(net1182),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4277_ (.D(net1248),
    .GATE(net1182),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4278_ (.D(net37),
    .GATE(net1184),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4279_ (.D(net36),
    .GATE(net1184),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4280_ (.D(net1252),
    .GATE(net1184),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4281_ (.D(net1253),
    .GATE(net1184),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4282_ (.D(net1254),
    .GATE(net1182),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4283_ (.D(net1255),
    .GATE(net1182),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4284_ (.D(net1256),
    .GATE(net1183),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4285_ (.D(net30),
    .GATE(net1185),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4286_ (.D(net1258),
    .GATE(net1182),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4287_ (.D(net1259),
    .GATE(net1182),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4288_ (.D(net1227),
    .GATE(net1184),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4289_ (.D(net1228),
    .GATE(net1184),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4290_ (.D(net1229),
    .GATE(net1183),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4291_ (.D(net53),
    .GATE(net1185),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4292_ (.D(net1231),
    .GATE(net1182),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4293_ (.D(net1232),
    .GATE(net1182),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4294_ (.D(net1233),
    .GATE(net1183),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4295_ (.D(net1236),
    .GATE(net1183),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4296_ (.D(net1249),
    .GATE(net1182),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4297_ (.D(net1260),
    .GATE(net1182),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4298_ (.D(net1234),
    .GATE(net1149),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4299_ (.D(net1235),
    .GATE(net1149),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4300_ (.D(net46),
    .GATE(net1149),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4301_ (.D(net45),
    .GATE(net1149),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4302_ (.D(net1239),
    .GATE(net1148),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4303_ (.D(net1240),
    .GATE(net1148),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4304_ (.D(net1241),
    .GATE(net1148),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4305_ (.D(net1243),
    .GATE(net1148),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4306_ (.D(net42),
    .GATE(net1148),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4307_ (.D(net41),
    .GATE(net1149),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4308_ (.D(net40),
    .GATE(net1148),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4309_ (.D(net39),
    .GATE(net1149),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4310_ (.D(net1250),
    .GATE(net1147),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4311_ (.D(net1251),
    .GATE(net1147),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4312_ (.D(net1252),
    .GATE(net1147),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4313_ (.D(net1253),
    .GATE(net1146),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4314_ (.D(net1254),
    .GATE(net1146),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4315_ (.D(net1255),
    .GATE(net1146),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4316_ (.D(net1256),
    .GATE(net1146),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4317_ (.D(net1257),
    .GATE(net1146),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4318_ (.D(net1258),
    .GATE(net1146),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4319_ (.D(net1259),
    .GATE(net1146),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4320_ (.D(net1227),
    .GATE(net1146),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4321_ (.D(net1228),
    .GATE(net1146),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4322_ (.D(net1229),
    .GATE(net1147),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4323_ (.D(net1230),
    .GATE(net1147),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4324_ (.D(net1231),
    .GATE(net1146),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4325_ (.D(net1232),
    .GATE(net1147),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4326_ (.D(net50),
    .GATE(net1148),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4327_ (.D(net47),
    .GATE(net1148),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4328_ (.D(net1249),
    .GATE(net1148),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4329_ (.D(net1260),
    .GATE(net1148),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4330_ (.D(net1234),
    .GATE(net1137),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4331_ (.D(net1235),
    .GATE(net1137),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4332_ (.D(net1237),
    .GATE(net1137),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4333_ (.D(net1238),
    .GATE(net1140),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4334_ (.D(net1239),
    .GATE(net1140),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4335_ (.D(net1240),
    .GATE(net1140),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4336_ (.D(net1241),
    .GATE(net1140),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4337_ (.D(net1243),
    .GATE(net1140),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4338_ (.D(net1245),
    .GATE(net1141),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4339_ (.D(net1246),
    .GATE(net1140),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4340_ (.D(net1247),
    .GATE(net1141),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4341_ (.D(net1248),
    .GATE(net1141),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4342_ (.D(net1250),
    .GATE(net1140),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4343_ (.D(net1251),
    .GATE(net1140),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4344_ (.D(net35),
    .GATE(net1140),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4345_ (.D(net1253),
    .GATE(net1140),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4346_ (.D(net1254),
    .GATE(net1137),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4347_ (.D(net1255),
    .GATE(net1137),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4348_ (.D(net1256),
    .GATE(net1137),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4349_ (.D(net1257),
    .GATE(net1137),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4350_ (.D(net29),
    .GATE(net1139),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4351_ (.D(net28),
    .GATE(net1139),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4352_ (.D(net1227),
    .GATE(net1139),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4353_ (.D(net1228),
    .GATE(net1139),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4354_ (.D(net1229),
    .GATE(net1137),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4355_ (.D(net1230),
    .GATE(net1137),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4356_ (.D(net1231),
    .GATE(net1138),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4357_ (.D(net1232),
    .GATE(net1137),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4358_ (.D(net1233),
    .GATE(net1138),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4359_ (.D(net1236),
    .GATE(net1138),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4360_ (.D(net1249),
    .GATE(net1138),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4361_ (.D(net1260),
    .GATE(net1138),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4362_ (.D(net1234),
    .GATE(net1131),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4363_ (.D(net1235),
    .GATE(net1131),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4364_ (.D(net1237),
    .GATE(net1131),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4365_ (.D(net1238),
    .GATE(net1131),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4366_ (.D(net1239),
    .GATE(net1130),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4367_ (.D(net1240),
    .GATE(net1130),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4368_ (.D(net1241),
    .GATE(net1130),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4369_ (.D(net1243),
    .GATE(net1130),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4370_ (.D(net1245),
    .GATE(net1131),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4371_ (.D(net1246),
    .GATE(net1131),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4372_ (.D(net1247),
    .GATE(net1130),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4373_ (.D(net1248),
    .GATE(net1130),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4374_ (.D(net1250),
    .GATE(net1130),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4375_ (.D(net1251),
    .GATE(net1130),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4376_ (.D(net35),
    .GATE(net1130),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4377_ (.D(net1253),
    .GATE(net1130),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4378_ (.D(net1254),
    .GATE(net1128),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4379_ (.D(net1255),
    .GATE(net1128),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4380_ (.D(net1256),
    .GATE(net1128),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4381_ (.D(net1257),
    .GATE(net1128),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4382_ (.D(net1258),
    .GATE(net1128),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4383_ (.D(net1259),
    .GATE(net1128),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4384_ (.D(net1227),
    .GATE(net1128),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4385_ (.D(net1228),
    .GATE(net1128),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4386_ (.D(net1229),
    .GATE(net1129),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4387_ (.D(net1230),
    .GATE(net1129),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4388_ (.D(net52),
    .GATE(net1129),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4389_ (.D(net1232),
    .GATE(net1129),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4390_ (.D(net1233),
    .GATE(net1129),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4391_ (.D(net1236),
    .GATE(net1128),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4392_ (.D(net1249),
    .GATE(net1128),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4393_ (.D(net1260),
    .GATE(net1129),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4394_ (.D(net49),
    .GATE(net1122),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4395_ (.D(net48),
    .GATE(net1122),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4396_ (.D(net1237),
    .GATE(net1122),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4397_ (.D(net1238),
    .GATE(net1122),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4398_ (.D(net1239),
    .GATE(net1121),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4399_ (.D(net1240),
    .GATE(net1121),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4400_ (.D(net1241),
    .GATE(net1121),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4401_ (.D(net1243),
    .GATE(net1121),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4402_ (.D(net42),
    .GATE(net1122),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4403_ (.D(net41),
    .GATE(net1122),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4404_ (.D(net40),
    .GATE(net1122),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4405_ (.D(net39),
    .GATE(net1122),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4406_ (.D(net1250),
    .GATE(net1121),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4407_ (.D(net1251),
    .GATE(net1120),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4408_ (.D(net35),
    .GATE(net1120),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4409_ (.D(net1253),
    .GATE(net1120),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4410_ (.D(net1254),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4411_ (.D(net1255),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4412_ (.D(net1256),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4413_ (.D(net1257),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4414_ (.D(net1258),
    .GATE(net1120),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4415_ (.D(net1259),
    .GATE(net1120),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4416_ (.D(net56),
    .GATE(net1120),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4417_ (.D(net55),
    .GATE(net1120),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4418_ (.D(net54),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4419_ (.D(net1230),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4420_ (.D(net1231),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4421_ (.D(net1232),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4422_ (.D(net1233),
    .GATE(net1120),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4423_ (.D(net47),
    .GATE(net1120),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4424_ (.D(net1249),
    .GATE(net1121),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4425_ (.D(net1260),
    .GATE(net1120),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4426_ (.D(net1234),
    .GATE(net1114),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4427_ (.D(net1235),
    .GATE(net1114),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4428_ (.D(net1237),
    .GATE(net1113),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4429_ (.D(net1238),
    .GATE(net1113),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4430_ (.D(net1239),
    .GATE(net1114),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4431_ (.D(net1240),
    .GATE(net1114),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4432_ (.D(net1241),
    .GATE(net1115),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4433_ (.D(net1243),
    .GATE(net1115),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4434_ (.D(net1245),
    .GATE(net1112),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4435_ (.D(net1246),
    .GATE(net1112),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4436_ (.D(net1247),
    .GATE(net1113),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4437_ (.D(net1248),
    .GATE(net1113),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4438_ (.D(net1250),
    .GATE(net1114),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4439_ (.D(net1251),
    .GATE(net1114),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4440_ (.D(net35),
    .GATE(net1115),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4441_ (.D(net1253),
    .GATE(net1115),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4442_ (.D(net1254),
    .GATE(net1113),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4443_ (.D(net1255),
    .GATE(net1113),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4444_ (.D(net1256),
    .GATE(net1112),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4445_ (.D(net1257),
    .GATE(net1112),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4446_ (.D(net29),
    .GATE(net1114),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4447_ (.D(net28),
    .GATE(net1114),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4448_ (.D(net1227),
    .GATE(net1114),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4449_ (.D(net1228),
    .GATE(net1114),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4450_ (.D(net1229),
    .GATE(net1112),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4451_ (.D(net1230),
    .GATE(net1112),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4452_ (.D(net1231),
    .GATE(net1112),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4453_ (.D(net1232),
    .GATE(net1112),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4454_ (.D(net1233),
    .GATE(net1112),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4455_ (.D(net1236),
    .GATE(net1112),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4456_ (.D(net1249),
    .GATE(net1115),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4457_ (.D(net27),
    .GATE(net1115),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4458_ (.D(net1234),
    .GATE(net1104),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4459_ (.D(net1235),
    .GATE(net1104),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4460_ (.D(net1237),
    .GATE(net1105),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4461_ (.D(net1238),
    .GATE(net1105),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4462_ (.D(net1239),
    .GATE(net1103),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4463_ (.D(net1240),
    .GATE(net1103),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4464_ (.D(net1241),
    .GATE(net1103),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4465_ (.D(net1243),
    .GATE(net1103),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4466_ (.D(net42),
    .GATE(net1105),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4467_ (.D(net41),
    .GATE(net1105),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4468_ (.D(net1247),
    .GATE(net1105),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4469_ (.D(net1248),
    .GATE(net1105),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4470_ (.D(net1250),
    .GATE(net1103),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4471_ (.D(net1251),
    .GATE(net1103),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4472_ (.D(net1252),
    .GATE(net1102),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4473_ (.D(net1253),
    .GATE(net1102),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4474_ (.D(net1254),
    .GATE(net1102),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4475_ (.D(net1255),
    .GATE(net1102),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4476_ (.D(net1256),
    .GATE(net1102),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4477_ (.D(net30),
    .GATE(net1102),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4478_ (.D(net1258),
    .GATE(net1103),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4479_ (.D(net1259),
    .GATE(net1103),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4480_ (.D(net1227),
    .GATE(net1104),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4481_ (.D(net1228),
    .GATE(net1104),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4482_ (.D(net1229),
    .GATE(net1106),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4483_ (.D(net53),
    .GATE(net1106),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4484_ (.D(net52),
    .GATE(net1102),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4485_ (.D(net51),
    .GATE(net1102),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4486_ (.D(net50),
    .GATE(net1103),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4487_ (.D(net1236),
    .GATE(net1103),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4488_ (.D(net1249),
    .GATE(net1102),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4489_ (.D(net1260),
    .GATE(net1102),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4490_ (.D(net1234),
    .GATE(net1094),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4491_ (.D(net1235),
    .GATE(net1094),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4492_ (.D(net1237),
    .GATE(net1097),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4493_ (.D(net1238),
    .GATE(net1095),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4494_ (.D(net44),
    .GATE(net1096),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4495_ (.D(net43),
    .GATE(net1096),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4496_ (.D(net1241),
    .GATE(net1096),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4497_ (.D(net1243),
    .GATE(net1096),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4498_ (.D(net1245),
    .GATE(net1097),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4499_ (.D(net41),
    .GATE(net1097),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4500_ (.D(net40),
    .GATE(net1095),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4501_ (.D(net39),
    .GATE(net1095),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4502_ (.D(net37),
    .GATE(net1096),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4503_ (.D(net36),
    .GATE(net1096),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4504_ (.D(net1252),
    .GATE(net1096),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4505_ (.D(net1253),
    .GATE(net1096),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4506_ (.D(net1254),
    .GATE(net1094),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4507_ (.D(net1255),
    .GATE(net1094),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4508_ (.D(net31),
    .GATE(net1095),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4509_ (.D(net1257),
    .GATE(net1095),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4510_ (.D(net1258),
    .GATE(net1095),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4511_ (.D(net1259),
    .GATE(net1095),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4512_ (.D(net56),
    .GATE(net1096),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4513_ (.D(net55),
    .GATE(net1096),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4514_ (.D(net1229),
    .GATE(net1095),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4515_ (.D(net53),
    .GATE(net1095),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4516_ (.D(net1231),
    .GATE(net1094),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4517_ (.D(net1232),
    .GATE(net1094),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4518_ (.D(net1233),
    .GATE(net1094),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4519_ (.D(net1236),
    .GATE(net1094),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4520_ (.D(net1249),
    .GATE(net1094),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4521_ (.D(net1260),
    .GATE(net1094),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4522_ (.D(net49),
    .GATE(net1088),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4523_ (.D(net1235),
    .GATE(net1088),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4524_ (.D(net46),
    .GATE(net1088),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4525_ (.D(net45),
    .GATE(net1088),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4526_ (.D(net1239),
    .GATE(net1087),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4527_ (.D(net1240),
    .GATE(net1087),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4528_ (.D(net1241),
    .GATE(net1087),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4529_ (.D(net1244),
    .GATE(net1087),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4530_ (.D(net1245),
    .GATE(net1089),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4531_ (.D(net1246),
    .GATE(net1086),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4532_ (.D(net1247),
    .GATE(net1088),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4533_ (.D(net1248),
    .GATE(net1088),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4534_ (.D(net1250),
    .GATE(net1087),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4535_ (.D(net1251),
    .GATE(net1087),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4536_ (.D(net1252),
    .GATE(net1086),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4537_ (.D(net34),
    .GATE(net1086),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4538_ (.D(net33),
    .GATE(net1089),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4539_ (.D(net32),
    .GATE(net1089),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4540_ (.D(net1256),
    .GATE(net1088),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4541_ (.D(net1257),
    .GATE(net1088),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4542_ (.D(net1258),
    .GATE(net1087),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4543_ (.D(net1259),
    .GATE(net1087),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4544_ (.D(net1227),
    .GATE(net1086),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4545_ (.D(net1228),
    .GATE(net1086),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4546_ (.D(net1229),
    .GATE(net1086),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4547_ (.D(net1230),
    .GATE(net1086),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4548_ (.D(net1231),
    .GATE(net1086),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4549_ (.D(net51),
    .GATE(net1086),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4550_ (.D(net1233),
    .GATE(net1087),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4551_ (.D(net1236),
    .GATE(net1087),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4552_ (.D(net38),
    .GATE(net1086),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4553_ (.D(net27),
    .GATE(net1089),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4554_ (.D(net1234),
    .GATE(net1079),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4555_ (.D(net1235),
    .GATE(net1078),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4556_ (.D(net1237),
    .GATE(net1079),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4557_ (.D(net1238),
    .GATE(net1079),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4558_ (.D(net44),
    .GATE(net1079),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4559_ (.D(net43),
    .GATE(net1079),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4560_ (.D(net1241),
    .GATE(net1081),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4561_ (.D(net1243),
    .GATE(net1081),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4562_ (.D(net1245),
    .GATE(net1081),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4563_ (.D(net1246),
    .GATE(net1080),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4564_ (.D(net1247),
    .GATE(net1080),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4565_ (.D(net1248),
    .GATE(net1080),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4566_ (.D(net1250),
    .GATE(net1081),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4567_ (.D(net1251),
    .GATE(net1080),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4568_ (.D(net1252),
    .GATE(net1078),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4569_ (.D(net1253),
    .GATE(net1078),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4570_ (.D(net1254),
    .GATE(net1078),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4571_ (.D(net1255),
    .GATE(net1080),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4572_ (.D(net1256),
    .GATE(net1080),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4573_ (.D(net1257),
    .GATE(net1080),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4574_ (.D(net1258),
    .GATE(net1080),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4575_ (.D(net1259),
    .GATE(net1080),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4576_ (.D(net1227),
    .GATE(net1080),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4577_ (.D(net1228),
    .GATE(net1081),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4578_ (.D(net54),
    .GATE(net1081),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4579_ (.D(net1230),
    .GATE(net1081),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4580_ (.D(net1231),
    .GATE(net1078),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4581_ (.D(net1232),
    .GATE(net1078),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4582_ (.D(net1233),
    .GATE(net1078),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4583_ (.D(net1236),
    .GATE(net1078),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4584_ (.D(net1249),
    .GATE(net1078),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4585_ (.D(net1260),
    .GATE(net1078),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4586_ (.D(net1234),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4587_ (.D(net1235),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4588_ (.D(net1237),
    .GATE(net1176),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4589_ (.D(net1238),
    .GATE(net1176),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4590_ (.D(net1239),
    .GATE(net1177),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4591_ (.D(net43),
    .GATE(net1177),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4592_ (.D(net1242),
    .GATE(net1176),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4593_ (.D(net1244),
    .GATE(net1176),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4594_ (.D(net1245),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4595_ (.D(net1246),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4596_ (.D(net1247),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4597_ (.D(net1248),
    .GATE(net1177),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4598_ (.D(net37),
    .GATE(net1176),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4599_ (.D(net36),
    .GATE(net1176),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4600_ (.D(net1252),
    .GATE(net1174),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4601_ (.D(net34),
    .GATE(net1174),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4602_ (.D(net33),
    .GATE(net1176),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4603_ (.D(net32),
    .GATE(net1174),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4604_ (.D(net31),
    .GATE(net1174),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4605_ (.D(net30),
    .GATE(net1174),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4606_ (.D(net29),
    .GATE(net1174),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4607_ (.D(net28),
    .GATE(net1174),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4608_ (.D(net1227),
    .GATE(net1174),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4609_ (.D(net1228),
    .GATE(net1174),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4610_ (.D(net1229),
    .GATE(net1174),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4611_ (.D(net1230),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4612_ (.D(net1231),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4613_ (.D(net1232),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4614_ (.D(net1233),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4615_ (.D(net1236),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4616_ (.D(net38),
    .GATE(net1177),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4617_ (.D(net27),
    .GATE(net1177),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4618_ (.D(net49),
    .GATE(net1167),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4619_ (.D(net48),
    .GATE(net1166),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4620_ (.D(net46),
    .GATE(net1166),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4621_ (.D(net45),
    .GATE(net1167),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4622_ (.D(net44),
    .GATE(net1166),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4623_ (.D(net1240),
    .GATE(net1166),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4624_ (.D(net1242),
    .GATE(net1167),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4625_ (.D(net1244),
    .GATE(net1166),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4626_ (.D(net1245),
    .GATE(net1166),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4627_ (.D(net1246),
    .GATE(net1166),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4628_ (.D(net1247),
    .GATE(net1166),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4629_ (.D(net39),
    .GATE(net1166),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4630_ (.D(net1250),
    .GATE(net1164),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4631_ (.D(net1251),
    .GATE(net1164),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4632_ (.D(net1252),
    .GATE(net1164),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4633_ (.D(net34),
    .GATE(net1165),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4634_ (.D(net33),
    .GATE(net1164),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4635_ (.D(net32),
    .GATE(net1164),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4636_ (.D(net31),
    .GATE(net1168),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4637_ (.D(net30),
    .GATE(net1168),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4638_ (.D(net1258),
    .GATE(net1168),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4639_ (.D(net1259),
    .GATE(net1168),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4640_ (.D(net56),
    .GATE(net1164),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4641_ (.D(net55),
    .GATE(net1164),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4642_ (.D(net1229),
    .GATE(net1168),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4643_ (.D(net1230),
    .GATE(net1168),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4644_ (.D(net1231),
    .GATE(net1164),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4645_ (.D(net1232),
    .GATE(net1164),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4646_ (.D(net1233),
    .GATE(net1164),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4647_ (.D(net1236),
    .GATE(net1165),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4648_ (.D(net1249),
    .GATE(net1165),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4649_ (.D(net1260),
    .GATE(net1165),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4650_ (.D(net1234),
    .GATE(net1157),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4651_ (.D(net48),
    .GATE(net1157),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4652_ (.D(net46),
    .GATE(net1156),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4653_ (.D(net45),
    .GATE(net1156),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4654_ (.D(net1239),
    .GATE(net1158),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4655_ (.D(net1240),
    .GATE(net1158),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4656_ (.D(net1241),
    .GATE(net1156),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4657_ (.D(net1243),
    .GATE(net1156),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4658_ (.D(net1245),
    .GATE(net1157),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4659_ (.D(net1246),
    .GATE(net1157),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4660_ (.D(net1247),
    .GATE(net1156),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4661_ (.D(net1248),
    .GATE(net1156),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4662_ (.D(net1250),
    .GATE(net1156),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4663_ (.D(net1251),
    .GATE(net1156),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4664_ (.D(net1252),
    .GATE(net1159),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4665_ (.D(net1253),
    .GATE(net1159),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4666_ (.D(net1254),
    .GATE(net1156),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4667_ (.D(net1255),
    .GATE(net1159),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4668_ (.D(net1256),
    .GATE(net1157),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4669_ (.D(net1257),
    .GATE(net1156),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4670_ (.D(net1258),
    .GATE(net1159),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4671_ (.D(net1259),
    .GATE(net1159),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4672_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0000_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4673_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0001_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4674_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0002_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4675_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0003_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4676_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0004_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4677_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0005_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4678_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0006_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4679_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0007_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4680_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0008_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4681_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0009_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4682_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0010_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4683_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0011_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4684_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0012_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4685_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0013_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4686_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0014_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4687_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0015_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4688_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0016_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[16] ));
 sky130_fd_sc_hd__dfxtp_1 _4689_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0017_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[17] ));
 sky130_fd_sc_hd__dfxtp_1 _4690_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0018_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[18] ));
 sky130_fd_sc_hd__dfxtp_1 _4691_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0019_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[19] ));
 sky130_fd_sc_hd__dfxtp_1 _4692_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.A0 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4693_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.A1 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4694_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.A2 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4695_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.A3 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4696_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4697_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4698_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4699_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4700_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.B0 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4701_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.B1 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4702_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.B2 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4703_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.B3 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4704_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4705_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4706_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4707_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4708_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C0 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4709_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(net676),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4710_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C2 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4711_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C3 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4712_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C4 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4713_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C5 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4714_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C6 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4715_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C7 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4716_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C8 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4717_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C9 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4718_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4719_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4720_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4721_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4722_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4723_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4724_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[16] ));
 sky130_fd_sc_hd__dfxtp_1 _4725_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[17] ));
 sky130_fd_sc_hd__dfxtp_1 _4726_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[18] ));
 sky130_fd_sc_hd__dfxtp_1 _4727_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[19] ));
 sky130_fd_sc_hd__dlxtp_1 _4728_ (.D(net1193),
    .GATE(net1179),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4729_ (.D(net1194),
    .GATE(net1179),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4730_ (.D(net1196),
    .GATE(net1179),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4731_ (.D(net1197),
    .GATE(net1179),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4732_ (.D(net161),
    .GATE(net1180),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4733_ (.D(net1199),
    .GATE(net1180),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4734_ (.D(net159),
    .GATE(net1181),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4735_ (.D(net1202),
    .GATE(net1181),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4736_ (.D(net1203),
    .GATE(net1179),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4737_ (.D(net1205),
    .GATE(net1179),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4738_ (.D(net1207),
    .GATE(net1178),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4739_ (.D(net1208),
    .GATE(net1178),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4740_ (.D(net1210),
    .GATE(net1178),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4741_ (.D(net1211),
    .GATE(net1180),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4742_ (.D(net1212),
    .GATE(net1181),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4743_ (.D(net152),
    .GATE(net1181),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4744_ (.D(net151),
    .GATE(net1180),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4745_ (.D(net1215),
    .GATE(net1180),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4746_ (.D(net149),
    .GATE(net1180),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4747_ (.D(net1217),
    .GATE(net1178),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4748_ (.D(net1218),
    .GATE(net1178),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4749_ (.D(net1219),
    .GATE(net1178),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4750_ (.D(net1186),
    .GATE(net1181),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4751_ (.D(net172),
    .GATE(net1181),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4752_ (.D(net1188),
    .GATE(net1178),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4753_ (.D(net1189),
    .GATE(net1178),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4754_ (.D(net1190),
    .GATE(net1178),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4755_ (.D(net1191),
    .GATE(net1178),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4756_ (.D(net167),
    .GATE(net1179),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4757_ (.D(net164),
    .GATE(net1179),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4758_ (.D(net1209),
    .GATE(net1179),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4759_ (.D(net1220),
    .GATE(net1179),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4760_ (.D(net1193),
    .GATE(net1145),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4761_ (.D(net1194),
    .GATE(net1145),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4762_ (.D(net1196),
    .GATE(net1144),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4763_ (.D(net1197),
    .GATE(net1144),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4764_ (.D(net1198),
    .GATE(net1143),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4765_ (.D(net1199),
    .GATE(net1143),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4766_ (.D(net1200),
    .GATE(net1143),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4767_ (.D(net1202),
    .GATE(net1143),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4768_ (.D(net1204),
    .GATE(net1143),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4769_ (.D(net1206),
    .GATE(net1144),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4770_ (.D(net1207),
    .GATE(net1143),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4771_ (.D(net1208),
    .GATE(net1144),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4772_ (.D(net155),
    .GATE(net1145),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4773_ (.D(net154),
    .GATE(net1145),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4774_ (.D(net153),
    .GATE(net1145),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4775_ (.D(net152),
    .GATE(net1145),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4776_ (.D(net1214),
    .GATE(net1142),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4777_ (.D(net1215),
    .GATE(net1142),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4778_ (.D(net1216),
    .GATE(net1142),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4779_ (.D(net1217),
    .GATE(net1142),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4780_ (.D(net1218),
    .GATE(net1142),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4781_ (.D(net1219),
    .GATE(net1142),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4782_ (.D(net1186),
    .GATE(net1150),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4783_ (.D(net1187),
    .GATE(net1150),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4784_ (.D(net1188),
    .GATE(net1142),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4785_ (.D(net1189),
    .GATE(net1142),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4786_ (.D(net1190),
    .GATE(net1142),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4787_ (.D(net1191),
    .GATE(net1142),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4788_ (.D(net1192),
    .GATE(net1143),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4789_ (.D(net1195),
    .GATE(net1143),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4790_ (.D(net1209),
    .GATE(net1143),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4791_ (.D(net1220),
    .GATE(net1143),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4792_ (.D(net1193),
    .GATE(net1135),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4793_ (.D(net1194),
    .GATE(net1135),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4794_ (.D(net1196),
    .GATE(net1135),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4795_ (.D(net1197),
    .GATE(net1135),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4796_ (.D(net1198),
    .GATE(net1135),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4797_ (.D(net1199),
    .GATE(net1135),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4798_ (.D(net1200),
    .GATE(net1135),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4799_ (.D(net1202),
    .GATE(net1135),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4800_ (.D(net1204),
    .GATE(net1136),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4801_ (.D(net1206),
    .GATE(net1136),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4802_ (.D(net1207),
    .GATE(net1135),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4803_ (.D(net1208),
    .GATE(net1135),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4804_ (.D(net1210),
    .GATE(net1136),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4805_ (.D(net1211),
    .GATE(net1136),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4806_ (.D(net1212),
    .GATE(net1136),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4807_ (.D(net1213),
    .GATE(net1136),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4808_ (.D(net1214),
    .GATE(net1134),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4809_ (.D(net1215),
    .GATE(net1134),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4810_ (.D(net1216),
    .GATE(net1133),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4811_ (.D(net1217),
    .GATE(net1133),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4812_ (.D(net1218),
    .GATE(net1134),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4813_ (.D(net1219),
    .GATE(net1134),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4814_ (.D(net1186),
    .GATE(net1134),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4815_ (.D(net1187),
    .GATE(net1134),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4816_ (.D(net1188),
    .GATE(net1133),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4817_ (.D(net1189),
    .GATE(net1133),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4818_ (.D(net1190),
    .GATE(net1133),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4819_ (.D(net1191),
    .GATE(net1133),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4820_ (.D(net1192),
    .GATE(net1133),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4821_ (.D(net1195),
    .GATE(net1133),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4822_ (.D(net1209),
    .GATE(net1133),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4823_ (.D(net1220),
    .GATE(net1133),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4824_ (.D(net1193),
    .GATE(net1127),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4825_ (.D(net1194),
    .GATE(net1132),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4826_ (.D(net1196),
    .GATE(net1127),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4827_ (.D(net1197),
    .GATE(net1127),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4828_ (.D(net1198),
    .GATE(net1126),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4829_ (.D(net160),
    .GATE(net1126),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4830_ (.D(net159),
    .GATE(net1126),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4831_ (.D(net1201),
    .GATE(net1126),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4832_ (.D(net1203),
    .GATE(net1127),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4833_ (.D(net1205),
    .GATE(net1127),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4834_ (.D(net1207),
    .GATE(net1132),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4835_ (.D(net1208),
    .GATE(net1127),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4836_ (.D(net1210),
    .GATE(net1127),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4837_ (.D(net154),
    .GATE(net1127),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4838_ (.D(net1212),
    .GATE(net1127),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4839_ (.D(net1213),
    .GATE(net1127),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4840_ (.D(net1214),
    .GATE(net1124),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4841_ (.D(net1215),
    .GATE(net1124),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4842_ (.D(net1216),
    .GATE(net1124),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4843_ (.D(net1217),
    .GATE(net1124),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4844_ (.D(net1218),
    .GATE(net1125),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4845_ (.D(net1219),
    .GATE(net1124),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4846_ (.D(net1186),
    .GATE(net1125),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4847_ (.D(net1187),
    .GATE(net1124),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4848_ (.D(net1188),
    .GATE(net1124),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4849_ (.D(net1189),
    .GATE(net1124),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4850_ (.D(net1190),
    .GATE(net1124),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4851_ (.D(net1191),
    .GATE(net1124),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4852_ (.D(net1192),
    .GATE(net1125),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4853_ (.D(net1195),
    .GATE(net1125),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4854_ (.D(net1209),
    .GATE(net1125),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4855_ (.D(net1220),
    .GATE(net1125),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4856_ (.D(net1193),
    .GATE(net1118),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4857_ (.D(net1194),
    .GATE(net1118),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4858_ (.D(net1196),
    .GATE(net1117),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4859_ (.D(net1197),
    .GATE(net1117),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4860_ (.D(net1198),
    .GATE(net1117),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4861_ (.D(net1199),
    .GATE(net1117),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4862_ (.D(net1200),
    .GATE(net1117),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4863_ (.D(net1202),
    .GATE(net1117),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4864_ (.D(net1204),
    .GATE(net1119),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4865_ (.D(net1206),
    .GATE(net1118),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4866_ (.D(net158),
    .GATE(net1118),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4867_ (.D(net1208),
    .GATE(net1118),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4868_ (.D(net1210),
    .GATE(net1118),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4869_ (.D(net154),
    .GATE(net1118),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4870_ (.D(net153),
    .GATE(net1118),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4871_ (.D(net152),
    .GATE(net1118),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4872_ (.D(net1214),
    .GATE(net1116),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4873_ (.D(net1215),
    .GATE(net1116),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4874_ (.D(net1216),
    .GATE(net1116),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4875_ (.D(net1217),
    .GATE(net1116),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4876_ (.D(net1218),
    .GATE(net1119),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4877_ (.D(net1219),
    .GATE(net1119),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4878_ (.D(net1186),
    .GATE(net1116),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4879_ (.D(net1187),
    .GATE(net1116),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4880_ (.D(net1188),
    .GATE(net1116),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4881_ (.D(net1189),
    .GATE(net1116),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4882_ (.D(net1190),
    .GATE(net1116),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4883_ (.D(net1191),
    .GATE(net1116),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4884_ (.D(net1192),
    .GATE(net1117),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4885_ (.D(net1195),
    .GATE(net1117),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4886_ (.D(net1209),
    .GATE(net1117),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4887_ (.D(net1220),
    .GATE(net1117),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4888_ (.D(net1193),
    .GATE(net1107),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4889_ (.D(net1194),
    .GATE(net1107),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4890_ (.D(net1196),
    .GATE(net1109),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4891_ (.D(net1197),
    .GATE(net1109),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4892_ (.D(net161),
    .GATE(net1109),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4893_ (.D(net160),
    .GATE(net1109),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4894_ (.D(net159),
    .GATE(net1109),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4895_ (.D(net1201),
    .GATE(net1109),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4896_ (.D(net1204),
    .GATE(net1107),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4897_ (.D(net1206),
    .GATE(net1107),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4898_ (.D(net1207),
    .GATE(net1109),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4899_ (.D(net1208),
    .GATE(net1109),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4900_ (.D(net1210),
    .GATE(net1110),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4901_ (.D(net1211),
    .GATE(net1110),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4902_ (.D(net153),
    .GATE(net1109),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4903_ (.D(net1213),
    .GATE(net1109),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4904_ (.D(net1214),
    .GATE(net1107),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4905_ (.D(net1215),
    .GATE(net1107),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4906_ (.D(net1216),
    .GATE(net1108),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4907_ (.D(net1217),
    .GATE(net1108),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4908_ (.D(net1218),
    .GATE(net1108),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4909_ (.D(net1219),
    .GATE(net1108),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4910_ (.D(net173),
    .GATE(net1111),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4911_ (.D(net1187),
    .GATE(net1111),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4912_ (.D(net1188),
    .GATE(net1107),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4913_ (.D(net1189),
    .GATE(net1107),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4914_ (.D(net1190),
    .GATE(net1108),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4915_ (.D(net1191),
    .GATE(net1108),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4916_ (.D(net1192),
    .GATE(net1107),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4917_ (.D(net1195),
    .GATE(net1107),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4918_ (.D(net156),
    .GATE(net1111),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4919_ (.D(net145),
    .GATE(net1111),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4920_ (.D(net166),
    .GATE(net1099),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4921_ (.D(net165),
    .GATE(net1099),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4922_ (.D(net163),
    .GATE(net1099),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4923_ (.D(net162),
    .GATE(net1099),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4924_ (.D(net1198),
    .GATE(net1098),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4925_ (.D(net1199),
    .GATE(net1100),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4926_ (.D(net1200),
    .GATE(net1101),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4927_ (.D(net1201),
    .GATE(net1101),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4928_ (.D(net1203),
    .GATE(net1099),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4929_ (.D(net1205),
    .GATE(net1099),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4930_ (.D(net158),
    .GATE(net1100),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4931_ (.D(net157),
    .GATE(net1099),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4932_ (.D(net1210),
    .GATE(net1098),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4933_ (.D(net1211),
    .GATE(net1098),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4934_ (.D(net1212),
    .GATE(net1101),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4935_ (.D(net1213),
    .GATE(net1101),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4936_ (.D(net1214),
    .GATE(net1098),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4937_ (.D(net1215),
    .GATE(net1101),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4938_ (.D(net1216),
    .GATE(net1099),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4939_ (.D(net148),
    .GATE(net1099),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4940_ (.D(net1218),
    .GATE(net1098),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4941_ (.D(net1219),
    .GATE(net1098),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4942_ (.D(net173),
    .GATE(net1101),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4943_ (.D(net1187),
    .GATE(net1101),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4944_ (.D(net1188),
    .GATE(net1098),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4945_ (.D(net1189),
    .GATE(net1098),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4946_ (.D(net169),
    .GATE(net1100),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4947_ (.D(net168),
    .GATE(net1099),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4948_ (.D(net1192),
    .GATE(net1098),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4949_ (.D(net1195),
    .GATE(net1098),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4950_ (.D(net156),
    .GATE(net1101),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4951_ (.D(net1220),
    .GATE(net1101),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4952_ (.D(net166),
    .GATE(net1091),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4953_ (.D(net165),
    .GATE(net1091),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4954_ (.D(net1196),
    .GATE(net1090),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4955_ (.D(net1197),
    .GATE(net1090),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4956_ (.D(net161),
    .GATE(net1091),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4957_ (.D(net1199),
    .GATE(net1091),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4958_ (.D(net159),
    .GATE(net1092),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4959_ (.D(net1201),
    .GATE(net1092),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4960_ (.D(net1203),
    .GATE(net1090),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4961_ (.D(net1205),
    .GATE(net1090),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4962_ (.D(net1207),
    .GATE(net1091),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4963_ (.D(net1208),
    .GATE(net1091),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4964_ (.D(net1210),
    .GATE(net1093),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4965_ (.D(net1211),
    .GATE(net1093),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4966_ (.D(net1212),
    .GATE(net1092),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4967_ (.D(net1213),
    .GATE(net1092),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4968_ (.D(net151),
    .GATE(net1092),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4969_ (.D(net150),
    .GATE(net1092),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4970_ (.D(net149),
    .GATE(net1090),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4971_ (.D(net1217),
    .GATE(net1090),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4972_ (.D(net147),
    .GATE(net1092),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4973_ (.D(net146),
    .GATE(net1092),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4974_ (.D(net173),
    .GATE(net1092),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4975_ (.D(net172),
    .GATE(net1092),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4976_ (.D(net1188),
    .GATE(net1090),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4977_ (.D(net1189),
    .GATE(net1090),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4978_ (.D(net1190),
    .GATE(net1090),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4979_ (.D(net1191),
    .GATE(net1090),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4980_ (.D(net1192),
    .GATE(net1091),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4981_ (.D(net1195),
    .GATE(net1091),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4982_ (.D(net1209),
    .GATE(net1093),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4983_ (.D(net1220),
    .GATE(net1093),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4984_ (.D(net166),
    .GATE(net1083),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4985_ (.D(net165),
    .GATE(net1083),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4986_ (.D(net163),
    .GATE(net1083),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4987_ (.D(net162),
    .GATE(net1083),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4988_ (.D(net1198),
    .GATE(net1084),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4989_ (.D(net1199),
    .GATE(net1084),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4990_ (.D(net1200),
    .GATE(net1084),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4991_ (.D(net1201),
    .GATE(net1084),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4992_ (.D(net1203),
    .GATE(net1084),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4993_ (.D(net1205),
    .GATE(net1085),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4994_ (.D(net158),
    .GATE(net1083),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4995_ (.D(net157),
    .GATE(net1083),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4996_ (.D(net155),
    .GATE(net1083),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4997_ (.D(net1211),
    .GATE(net1082),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4998_ (.D(net1212),
    .GATE(net1082),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4999_ (.D(net1213),
    .GATE(net1083),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5000_ (.D(net1214),
    .GATE(net1084),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5001_ (.D(net150),
    .GATE(net1085),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5002_ (.D(net1216),
    .GATE(net1082),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5003_ (.D(net148),
    .GATE(net1082),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5004_ (.D(net1218),
    .GATE(net1082),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5005_ (.D(net1219),
    .GATE(net1082),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5006_ (.D(net1186),
    .GATE(net1082),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5007_ (.D(net1187),
    .GATE(net1082),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5008_ (.D(net171),
    .GATE(net1084),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5009_ (.D(net170),
    .GATE(net1085),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5010_ (.D(net169),
    .GATE(net1084),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5011_ (.D(net168),
    .GATE(net1084),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5012_ (.D(net1192),
    .GATE(net1082),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5013_ (.D(net164),
    .GATE(net1082),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5014_ (.D(net156),
    .GATE(net1084),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5015_ (.D(net145),
    .GATE(net1085),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5016_ (.D(net166),
    .GATE(net1076),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5017_ (.D(net1194),
    .GATE(net1076),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5018_ (.D(net1196),
    .GATE(net1075),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5019_ (.D(net1197),
    .GATE(net1075),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5020_ (.D(net1198),
    .GATE(net1075),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5021_ (.D(net1199),
    .GATE(net1074),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5022_ (.D(net1200),
    .GATE(net1077),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5023_ (.D(net1201),
    .GATE(net1077),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5024_ (.D(net1203),
    .GATE(net1076),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5025_ (.D(net1205),
    .GATE(net1077),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5026_ (.D(net1207),
    .GATE(net1074),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5027_ (.D(net1208),
    .GATE(net1074),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5028_ (.D(net1210),
    .GATE(net1074),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5029_ (.D(net1211),
    .GATE(net1074),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5030_ (.D(net1212),
    .GATE(net1074),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5031_ (.D(net1213),
    .GATE(net1074),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5032_ (.D(net1214),
    .GATE(net1076),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5033_ (.D(net1215),
    .GATE(net1076),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5034_ (.D(net1216),
    .GATE(net1074),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5035_ (.D(net1217),
    .GATE(net1074),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5036_ (.D(net1218),
    .GATE(net1074),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5037_ (.D(net1219),
    .GATE(net1076),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5038_ (.D(net1186),
    .GATE(net1076),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5039_ (.D(net1187),
    .GATE(net1076),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5040_ (.D(net1188),
    .GATE(net1075),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5041_ (.D(net1189),
    .GATE(net1075),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5042_ (.D(net1190),
    .GATE(net1075),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5043_ (.D(net1191),
    .GATE(net1075),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5044_ (.D(net1192),
    .GATE(net1076),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5045_ (.D(net1195),
    .GATE(net1076),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5046_ (.D(net1209),
    .GATE(net1075),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5047_ (.D(net1220),
    .GATE(net1075),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5048_ (.D(net1193),
    .GATE(net1169),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5049_ (.D(net1194),
    .GATE(net1169),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5050_ (.D(net1196),
    .GATE(net1169),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5051_ (.D(net1197),
    .GATE(net1169),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5052_ (.D(net1198),
    .GATE(net1170),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5053_ (.D(net1199),
    .GATE(net1170),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5054_ (.D(net1200),
    .GATE(net1173),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5055_ (.D(net1201),
    .GATE(net1173),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5056_ (.D(net1203),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5057_ (.D(net1205),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5058_ (.D(net1207),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5059_ (.D(net1208),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5060_ (.D(net155),
    .GATE(net1172),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5061_ (.D(net1211),
    .GATE(net1172),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5062_ (.D(net1212),
    .GATE(net1172),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5063_ (.D(net1213),
    .GATE(net1172),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5064_ (.D(net151),
    .GATE(net1172),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5065_ (.D(net150),
    .GATE(net1172),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5066_ (.D(net1216),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5067_ (.D(net148),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5068_ (.D(net147),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5069_ (.D(net146),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5070_ (.D(net1186),
    .GATE(net1170),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5071_ (.D(net1187),
    .GATE(net1170),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5072_ (.D(net171),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5073_ (.D(net170),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5074_ (.D(net1190),
    .GATE(net1169),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5075_ (.D(net1191),
    .GATE(net1169),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5076_ (.D(net1192),
    .GATE(net1169),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5077_ (.D(net1195),
    .GATE(net1169),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5078_ (.D(net1209),
    .GATE(net1169),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5079_ (.D(net1220),
    .GATE(net1169),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5080_ (.D(net1193),
    .GATE(net1162),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5081_ (.D(net1194),
    .GATE(net1162),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5082_ (.D(net163),
    .GATE(net1160),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5083_ (.D(net162),
    .GATE(net1160),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5084_ (.D(net161),
    .GATE(net1160),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5085_ (.D(net160),
    .GATE(net1160),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5086_ (.D(net1200),
    .GATE(net1160),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5087_ (.D(net1201),
    .GATE(net1160),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5088_ (.D(net1203),
    .GATE(net1161),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5089_ (.D(net1205),
    .GATE(net1161),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5090_ (.D(net1207),
    .GATE(net1160),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5091_ (.D(net157),
    .GATE(net1160),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5092_ (.D(net155),
    .GATE(net1160),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5093_ (.D(net1211),
    .GATE(net1163),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5094_ (.D(net1212),
    .GATE(net1163),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5095_ (.D(net1213),
    .GATE(net1163),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5096_ (.D(net1214),
    .GATE(net1162),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5097_ (.D(net1215),
    .GATE(net1162),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5098_ (.D(net1216),
    .GATE(net1162),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5099_ (.D(net148),
    .GATE(net1160),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5100_ (.D(net147),
    .GATE(net1161),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5101_ (.D(net146),
    .GATE(net1161),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5102_ (.D(net173),
    .GATE(net1161),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5103_ (.D(net172),
    .GATE(net1162),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5104_ (.D(net171),
    .GATE(net1161),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5105_ (.D(net170),
    .GATE(net1161),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5106_ (.D(net169),
    .GATE(net1162),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5107_ (.D(net168),
    .GATE(net1162),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5108_ (.D(net167),
    .GATE(net1161),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5109_ (.D(net1195),
    .GATE(net1161),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5110_ (.D(net1209),
    .GATE(net1163),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5111_ (.D(net1220),
    .GATE(net1162),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5112_ (.D(net1193),
    .GATE(net1151),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5113_ (.D(net1194),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5114_ (.D(net1196),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5115_ (.D(net1197),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5116_ (.D(net1198),
    .GATE(net1151),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5117_ (.D(net1199),
    .GATE(net1151),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5118_ (.D(net1200),
    .GATE(net1152),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5119_ (.D(net1201),
    .GATE(net1153),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5120_ (.D(net1203),
    .GATE(net1153),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5121_ (.D(net1205),
    .GATE(net1153),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5122_ (.D(net1207),
    .GATE(net1151),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5123_ (.D(net1208),
    .GATE(net1151),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5124_ (.D(net1210),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5125_ (.D(net1211),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5126_ (.D(net1212),
    .GATE(net1151),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5127_ (.D(net1213),
    .GATE(net1151),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5128_ (.D(net1214),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5129_ (.D(net1215),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5130_ (.D(net149),
    .GATE(net1152),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5131_ (.D(net1217),
    .GATE(net1151),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5132_ (.D(net1218),
    .GATE(net1152),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5133_ (.D(net1219),
    .GATE(net1152),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5134_ (.D(net1186),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5135_ (.D(net1187),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5136_ (.D(net1188),
    .GATE(net1151),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5137_ (.D(net1189),
    .GATE(net1151),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5138_ (.D(net169),
    .GATE(net1155),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5139_ (.D(net168),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5140_ (.D(net167),
    .GATE(net1153),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5141_ (.D(net164),
    .GATE(net1153),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5142_ (.D(net156),
    .GATE(net1155),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _5143_ (.D(net145),
    .GATE(net1155),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ));
 sky130_fd_sc_hd__buf_2 _5144_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 ),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 _5145_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 ),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_1 rebuffer297 (.A(net915),
    .X(net914));
 sky130_fd_sc_hd__clkbuf_2 _5147_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 ),
    .X(net239));
 sky130_fd_sc_hd__buf_4 _5148_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 ),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 _5149_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ),
    .X(net241));
 sky130_fd_sc_hd__buf_2 _5150_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ),
    .X(net242));
 sky130_fd_sc_hd__buf_4 _5151_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_2 _5152_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ),
    .X(net244));
 sky130_fd_sc_hd__buf_1 _5153_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ),
    .X(net245));
 sky130_fd_sc_hd__buf_6 _5154_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ),
    .X(net246));
 sky130_fd_sc_hd__buf_1 _5155_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 ),
    .X(net247));
 sky130_fd_sc_hd__buf_1 _5156_ (.A(net13),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_2 _5157_ (.A(net14),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 _5158_ (.A(net15),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_2 _5159_ (.A(net16),
    .X(net251));
 sky130_fd_sc_hd__buf_1 _5160_ (.A(net17),
    .X(net252));
 sky130_fd_sc_hd__buf_1 _5161_ (.A(net18),
    .X(net253));
 sky130_fd_sc_hd__buf_1 _5162_ (.A(net19),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_2 _5163_ (.A(net20),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_1 _5164_ (.A(Tile_X0Y0_E6END[2]),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_1 _5165_ (.A(Tile_X0Y0_E6END[3]),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_1 _5166_ (.A(Tile_X0Y0_E6END[4]),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 _5167_ (.A(Tile_X0Y0_E6END[5]),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 _5168_ (.A(Tile_X0Y0_E6END[6]),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_1 _5169_ (.A(Tile_X0Y0_E6END[7]),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_1 _5170_ (.A(Tile_X0Y0_E6END[8]),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_1 _5171_ (.A(Tile_X0Y0_E6END[9]),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 _5172_ (.A(Tile_X0Y0_E6END[10]),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_1 _5173_ (.A(Tile_X0Y0_E6END[11]),
    .X(net267));
 sky130_fd_sc_hd__buf_6 _5174_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 ),
    .X(net257));
 sky130_fd_sc_hd__buf_6 _5175_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 ),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_1 _5176_ (.A(Tile_X0Y0_EE4END[4]),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 _5177_ (.A(Tile_X0Y0_EE4END[5]),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_1 _5178_ (.A(Tile_X0Y0_EE4END[6]),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_1 _5179_ (.A(Tile_X0Y0_EE4END[7]),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_1 _5180_ (.A(Tile_X0Y0_EE4END[8]),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_1 _5181_ (.A(Tile_X0Y0_EE4END[9]),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_1 _5182_ (.A(Tile_X0Y0_EE4END[10]),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_1 _5183_ (.A(Tile_X0Y0_EE4END[11]),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_1 _5184_ (.A(Tile_X0Y0_EE4END[12]),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_1 _5185_ (.A(Tile_X0Y0_EE4END[13]),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_1 _5186_ (.A(Tile_X0Y0_EE4END[14]),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_1 _5187_ (.A(Tile_X0Y0_EE4END[15]),
    .X(net270));
 sky130_fd_sc_hd__buf_1 _5188_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 ),
    .X(net271));
 sky130_fd_sc_hd__buf_6 _5189_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 ),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_1 _5190_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 ),
    .X(net273));
 sky130_fd_sc_hd__buf_6 _5191_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 ),
    .X(net274));
 sky130_fd_sc_hd__buf_4 _5192_ (.A(net1260),
    .X(net284));
 sky130_fd_sc_hd__buf_1 _5193_ (.A(net38),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_2 _5194_ (.A(net47),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_2 _5195_ (.A(net50),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_2 _5196_ (.A(net51),
    .X(net310));
 sky130_fd_sc_hd__buf_2 _5197_ (.A(net52),
    .X(net311));
 sky130_fd_sc_hd__buf_4 _5198_ (.A(net1230),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_2 _5199_ (.A(net54),
    .X(net313));
 sky130_fd_sc_hd__buf_4 _5200_ (.A(net1228),
    .X(net314));
 sky130_fd_sc_hd__buf_4 _5201_ (.A(net1227),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_2 _5202_ (.A(net28),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_2 _5203_ (.A(net29),
    .X(net286));
 sky130_fd_sc_hd__buf_4 _5204_ (.A(net1257),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_2 _5205_ (.A(net31),
    .X(net288));
 sky130_fd_sc_hd__buf_1 _5206_ (.A(net32),
    .X(net289));
 sky130_fd_sc_hd__buf_1 _5207_ (.A(net33),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_1 _5208_ (.A(net34),
    .X(net291));
 sky130_fd_sc_hd__buf_2 _5209_ (.A(net1252),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_2 _5210_ (.A(net36),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_2 _5211_ (.A(net37),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_2 _5212_ (.A(net1248),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_2 _5213_ (.A(net40),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_2 _5214_ (.A(net1246),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_2 _5215_ (.A(net1245),
    .X(net299));
 sky130_fd_sc_hd__buf_1 _5216_ (.A(net1244),
    .X(net300));
 sky130_fd_sc_hd__buf_1 _5217_ (.A(net1242),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_2 _5218_ (.A(net1240),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_2 _5219_ (.A(net1239),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_2 _5220_ (.A(net1238),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_2 _5221_ (.A(net1237),
    .X(net305));
 sky130_fd_sc_hd__buf_1 _5222_ (.A(net48),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_1 _5223_ (.A(net49),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_2 _5224_ (.A(net1185),
    .X(net316));
 sky130_fd_sc_hd__buf_1 _5225_ (.A(net1149),
    .X(net327));
 sky130_fd_sc_hd__buf_4 _5226_ (.A(net1141),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_1 _5227_ (.A(net1131),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_2 _5228_ (.A(net1122),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_2 _5229_ (.A(net1115),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_2 _5230_ (.A(net1105),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_2 _5231_ (.A(net1097),
    .X(net333));
 sky130_fd_sc_hd__buf_1 _5232_ (.A(net1088),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_2 _5233_ (.A(net1081),
    .X(net335));
 sky130_fd_sc_hd__buf_1 _5234_ (.A(net1176),
    .X(net317));
 sky130_fd_sc_hd__buf_1 _5235_ (.A(net1166),
    .X(net318));
 sky130_fd_sc_hd__buf_1 _5236_ (.A(net1158),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_1 _5237_ (.A(Tile_X0Y1_FrameStrobe[13]),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_1 _5238_ (.A(Tile_X0Y1_FrameStrobe[14]),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_1 _5239_ (.A(Tile_X0Y1_FrameStrobe[15]),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_1 _5240_ (.A(Tile_X0Y1_FrameStrobe[16]),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_1 _5241_ (.A(Tile_X0Y1_FrameStrobe[17]),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_1 _5242_ (.A(Tile_X0Y1_FrameStrobe[18]),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_1 _5243_ (.A(Tile_X0Y1_FrameStrobe[19]),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_2 _5244_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 ),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer302 (.A(_1566_),
    .X(net919));
 sky130_fd_sc_hd__buf_6 rebuffer257 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_2 _5247_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 ),
    .X(net339));
 sky130_fd_sc_hd__buf_1 _5248_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 ),
    .X(net340));
 sky130_fd_sc_hd__buf_1 _5249_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ),
    .X(net341));
 sky130_fd_sc_hd__buf_1 _5250_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 _5251_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_1 _5252_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_2 _5253_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 ),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_1 _5254_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_2 _5255_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 ),
    .X(net347));
 sky130_fd_sc_hd__buf_2 _5256_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .X(net348));
 sky130_fd_sc_hd__buf_6 _5257_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .X(net349));
 sky130_fd_sc_hd__buf_4 _5258_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .X(net350));
 sky130_fd_sc_hd__buf_4 _5259_ (.A(net619),
    .X(net351));
 sky130_fd_sc_hd__buf_6 _5260_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .X(net352));
 sky130_fd_sc_hd__buf_4 _5261_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_2 _5262_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .X(net354));
 sky130_fd_sc_hd__buf_2 _5263_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_1 _5264_ (.A(Tile_X0Y1_N4END[8]),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_1 _5265_ (.A(Tile_X0Y1_N4END[9]),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_1 _5266_ (.A(Tile_X0Y1_N4END[10]),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_1 _5267_ (.A(Tile_X0Y1_N4END[11]),
    .X(net365));
 sky130_fd_sc_hd__buf_1 _5268_ (.A(Tile_X0Y1_N4END[12]),
    .X(net366));
 sky130_fd_sc_hd__buf_1 _5269_ (.A(Tile_X0Y1_N4END[13]),
    .X(net367));
 sky130_fd_sc_hd__buf_1 _5270_ (.A(Tile_X0Y1_N4END[14]),
    .X(net368));
 sky130_fd_sc_hd__buf_1 _5271_ (.A(Tile_X0Y1_N4END[15]),
    .X(net369));
 sky130_fd_sc_hd__buf_4 _5272_ (.A(\Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A ),
    .X(net370));
 sky130_fd_sc_hd__buf_4 _5273_ (.A(\Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A ),
    .X(net371));
 sky130_fd_sc_hd__buf_4 _5274_ (.A(\Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A ),
    .X(net357));
 sky130_fd_sc_hd__buf_4 _5275_ (.A(\Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A ),
    .X(net358));
 sky130_fd_sc_hd__buf_1 _5276_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 ),
    .X(net359));
 sky130_fd_sc_hd__buf_1 _5277_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 ),
    .X(net360));
 sky130_fd_sc_hd__buf_1 _5278_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 ),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_2 _5279_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 ),
    .X(net362));
 sky130_fd_sc_hd__buf_1 _5280_ (.A(Tile_X0Y1_NN4END[8]),
    .X(net372));
 sky130_fd_sc_hd__buf_1 _5281_ (.A(Tile_X0Y1_NN4END[9]),
    .X(net379));
 sky130_fd_sc_hd__buf_1 _5282_ (.A(Tile_X0Y1_NN4END[10]),
    .X(net380));
 sky130_fd_sc_hd__buf_1 _5283_ (.A(Tile_X0Y1_NN4END[11]),
    .X(net381));
 sky130_fd_sc_hd__buf_1 _5284_ (.A(Tile_X0Y1_NN4END[12]),
    .X(net382));
 sky130_fd_sc_hd__buf_1 _5285_ (.A(Tile_X0Y1_NN4END[13]),
    .X(net383));
 sky130_fd_sc_hd__buf_1 _5286_ (.A(Tile_X0Y1_NN4END[14]),
    .X(net384));
 sky130_fd_sc_hd__buf_4 _5287_ (.A(Tile_X0Y1_NN4END[15]),
    .X(net385));
 sky130_fd_sc_hd__buf_6 _5288_ (.A(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A ),
    .X(net386));
 sky130_fd_sc_hd__buf_4 _5289_ (.A(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A ),
    .X(net387));
 sky130_fd_sc_hd__buf_4 _5290_ (.A(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A ),
    .X(net373));
 sky130_fd_sc_hd__buf_6 _5291_ (.A(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A ),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_2 _5292_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 ),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_1 clone311 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .X(net928));
 sky130_fd_sc_hd__buf_4 _5294_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 ),
    .X(net377));
 sky130_fd_sc_hd__buf_8 clone249 (.A(net1033),
    .X(net866));
 sky130_fd_sc_hd__buf_2 _5296_ (.A(clknet_1_0__leaf_Tile_X0Y1_UserCLK),
    .X(net388));
 sky130_fd_sc_hd__buf_1 _5297_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 ),
    .X(net389));
 sky130_fd_sc_hd__buf_1 _5298_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 ),
    .X(net390));
 sky130_fd_sc_hd__buf_6 _5299_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 ),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_2 _5300_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 ),
    .X(net392));
 sky130_fd_sc_hd__buf_1 _5301_ (.A(net97),
    .X(net393));
 sky130_fd_sc_hd__buf_1 _5302_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ),
    .X(net394));
 sky130_fd_sc_hd__buf_1 _5303_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_2 _5304_ (.A(net100),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_1 _5305_ (.A(net101),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_2 _5306_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 ),
    .X(net398));
 sky130_fd_sc_hd__buf_4 _5307_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_2 _5308_ (.A(net104),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_2 _5309_ (.A(net105),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_2 _5310_ (.A(net106),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_2 _5311_ (.A(net107),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_2 _5312_ (.A(net108),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_2 _5313_ (.A(net109),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_2 _5314_ (.A(net110),
    .X(net406));
 sky130_fd_sc_hd__buf_1 _5315_ (.A(net111),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_2 _5316_ (.A(net112),
    .X(net408));
 sky130_fd_sc_hd__buf_4 _5317_ (.A(Tile_X0Y0_W6END[2]),
    .X(net409));
 sky130_fd_sc_hd__buf_4 _5318_ (.A(Tile_X0Y0_W6END[3]),
    .X(net412));
 sky130_fd_sc_hd__buf_4 _5319_ (.A(Tile_X0Y0_W6END[4]),
    .X(net413));
 sky130_fd_sc_hd__buf_4 _5320_ (.A(Tile_X0Y0_W6END[5]),
    .X(net414));
 sky130_fd_sc_hd__buf_4 _5321_ (.A(Tile_X0Y0_W6END[6]),
    .X(net415));
 sky130_fd_sc_hd__buf_4 _5322_ (.A(Tile_X0Y0_W6END[7]),
    .X(net416));
 sky130_fd_sc_hd__buf_4 _5323_ (.A(Tile_X0Y0_W6END[8]),
    .X(net417));
 sky130_fd_sc_hd__buf_4 _5324_ (.A(Tile_X0Y0_W6END[9]),
    .X(net418));
 sky130_fd_sc_hd__buf_4 _5325_ (.A(Tile_X0Y0_W6END[10]),
    .X(net419));
 sky130_fd_sc_hd__buf_4 _5326_ (.A(Tile_X0Y0_W6END[11]),
    .X(net420));
 sky130_fd_sc_hd__buf_6 _5327_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 ),
    .X(net410));
 sky130_fd_sc_hd__buf_6 _5328_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 ),
    .X(net411));
 sky130_fd_sc_hd__buf_4 _5329_ (.A(Tile_X0Y0_WW4END[4]),
    .X(net421));
 sky130_fd_sc_hd__buf_4 _5330_ (.A(Tile_X0Y0_WW4END[5]),
    .X(net428));
 sky130_fd_sc_hd__buf_4 _5331_ (.A(Tile_X0Y0_WW4END[6]),
    .X(net429));
 sky130_fd_sc_hd__buf_4 _5332_ (.A(Tile_X0Y0_WW4END[7]),
    .X(net430));
 sky130_fd_sc_hd__buf_4 _5333_ (.A(Tile_X0Y0_WW4END[8]),
    .X(net431));
 sky130_fd_sc_hd__buf_4 _5334_ (.A(Tile_X0Y0_WW4END[9]),
    .X(net432));
 sky130_fd_sc_hd__buf_4 _5335_ (.A(Tile_X0Y0_WW4END[10]),
    .X(net433));
 sky130_fd_sc_hd__buf_4 _5336_ (.A(Tile_X0Y0_WW4END[11]),
    .X(net434));
 sky130_fd_sc_hd__buf_4 _5337_ (.A(Tile_X0Y0_WW4END[12]),
    .X(net435));
 sky130_fd_sc_hd__buf_4 _5338_ (.A(Tile_X0Y0_WW4END[13]),
    .X(net436));
 sky130_fd_sc_hd__buf_4 _5339_ (.A(Tile_X0Y0_WW4END[14]),
    .X(net422));
 sky130_fd_sc_hd__buf_4 _5340_ (.A(Tile_X0Y0_WW4END[15]),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_2 _5341_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 ),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_2 rebuffer329 (.A(net947),
    .X(net946));
 sky130_fd_sc_hd__buf_6 _5343_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer210 (.A(_0219_),
    .X(net827));
 sky130_fd_sc_hd__buf_1 _5345_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 ),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_2 _5346_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 ),
    .X(net438));
 sky130_fd_sc_hd__buf_1 _5347_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 ),
    .X(net439));
 sky130_fd_sc_hd__buf_1 _5348_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 ),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_2 _5349_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 ),
    .X(net441));
 sky130_fd_sc_hd__buf_1 _5350_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_2 _5351_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_2 _5352_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .X(net444));
 sky130_fd_sc_hd__buf_1 _5353_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_1 _5354_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_1 _5355_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_2 rebuffer258 (.A(net874),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_2 _5357_ (.A(net131),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_2 _5358_ (.A(net132),
    .X(net450));
 sky130_fd_sc_hd__buf_1 _5359_ (.A(net133),
    .X(net451));
 sky130_fd_sc_hd__buf_1 _5360_ (.A(net134),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_2 _5361_ (.A(net135),
    .X(net453));
 sky130_fd_sc_hd__buf_1 _5362_ (.A(net136),
    .X(net454));
 sky130_fd_sc_hd__buf_1 _5363_ (.A(net137),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_2 _5364_ (.A(net138),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_1 _5365_ (.A(Tile_X0Y1_E6END[2]),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_1 _5366_ (.A(Tile_X0Y1_E6END[3]),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_1 _5367_ (.A(Tile_X0Y1_E6END[4]),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_1 _5368_ (.A(Tile_X0Y1_E6END[5]),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_1 _5369_ (.A(Tile_X0Y1_E6END[6]),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_1 _5370_ (.A(Tile_X0Y1_E6END[7]),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_1 _5371_ (.A(Tile_X0Y1_E6END[8]),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_1 _5372_ (.A(Tile_X0Y1_E6END[9]),
    .X(net466));
 sky130_fd_sc_hd__clkbuf_1 _5373_ (.A(Tile_X0Y1_E6END[10]),
    .X(net467));
 sky130_fd_sc_hd__clkbuf_1 _5374_ (.A(Tile_X0Y1_E6END[11]),
    .X(net468));
 sky130_fd_sc_hd__clkbuf_1 _5375_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 ),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_2 _5376_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 ),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_1 _5377_ (.A(Tile_X0Y1_EE4END[4]),
    .X(net469));
 sky130_fd_sc_hd__clkbuf_1 _5378_ (.A(Tile_X0Y1_EE4END[5]),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_1 _5379_ (.A(Tile_X0Y1_EE4END[6]),
    .X(net477));
 sky130_fd_sc_hd__clkbuf_1 _5380_ (.A(Tile_X0Y1_EE4END[7]),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_1 _5381_ (.A(Tile_X0Y1_EE4END[8]),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_1 _5382_ (.A(Tile_X0Y1_EE4END[9]),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_1 _5383_ (.A(Tile_X0Y1_EE4END[10]),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_1 _5384_ (.A(Tile_X0Y1_EE4END[11]),
    .X(net482));
 sky130_fd_sc_hd__clkbuf_1 _5385_ (.A(Tile_X0Y1_EE4END[12]),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_1 _5386_ (.A(Tile_X0Y1_EE4END[13]),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_1 _5387_ (.A(Tile_X0Y1_EE4END[14]),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_1 _5388_ (.A(Tile_X0Y1_EE4END[15]),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_1 _5389_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 ),
    .X(net472));
 sky130_fd_sc_hd__clkbuf_2 _5390_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 ),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_2 _5391_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer43 (.A(_0268_),
    .X(net660));
 sky130_fd_sc_hd__buf_1 _5393_ (.A(net145),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_2 _5394_ (.A(net1209),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_1 _5395_ (.A(net164),
    .X(net507));
 sky130_fd_sc_hd__buf_1 _5396_ (.A(net167),
    .X(net510));
 sky130_fd_sc_hd__buf_4 _5397_ (.A(net1191),
    .X(net511));
 sky130_fd_sc_hd__buf_4 _5398_ (.A(net1190),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_2 _5399_ (.A(net170),
    .X(net513));
 sky130_fd_sc_hd__clkbuf_2 _5400_ (.A(net171),
    .X(net514));
 sky130_fd_sc_hd__buf_1 _5401_ (.A(net172),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_2 _5402_ (.A(net1186),
    .X(net516));
 sky130_fd_sc_hd__buf_1 _5403_ (.A(net146),
    .X(net486));
 sky130_fd_sc_hd__buf_1 _5404_ (.A(net147),
    .X(net487));
 sky130_fd_sc_hd__buf_2 _5405_ (.A(net1217),
    .X(net488));
 sky130_fd_sc_hd__buf_4 _5406_ (.A(net149),
    .X(net489));
 sky130_fd_sc_hd__buf_1 _5407_ (.A(net150),
    .X(net490));
 sky130_fd_sc_hd__buf_1 _5408_ (.A(net151),
    .X(net491));
 sky130_fd_sc_hd__buf_1 _5409_ (.A(net152),
    .X(net492));
 sky130_fd_sc_hd__buf_1 _5410_ (.A(net153),
    .X(net493));
 sky130_fd_sc_hd__buf_1 _5411_ (.A(net154),
    .X(net494));
 sky130_fd_sc_hd__buf_1 _5412_ (.A(net1210),
    .X(net495));
 sky130_fd_sc_hd__clkbuf_2 _5413_ (.A(net157),
    .X(net497));
 sky130_fd_sc_hd__clkbuf_2 _5414_ (.A(net158),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_2 _5415_ (.A(net1205),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_2 _5416_ (.A(net1203),
    .X(net500));
 sky130_fd_sc_hd__buf_1 _5417_ (.A(net1201),
    .X(net501));
 sky130_fd_sc_hd__buf_1 _5418_ (.A(net1200),
    .X(net502));
 sky130_fd_sc_hd__buf_1 _5419_ (.A(net160),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_2 _5420_ (.A(net1198),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_2 _5421_ (.A(net162),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_2 _5422_ (.A(net163),
    .X(net506));
 sky130_fd_sc_hd__clkbuf_2 _5423_ (.A(net165),
    .X(net508));
 sky130_fd_sc_hd__buf_4 _5424_ (.A(net1193),
    .X(net509));
 sky130_fd_sc_hd__clkbuf_1 _5425_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 ),
    .X(net517));
 sky130_fd_sc_hd__buf_4 _5426_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 ),
    .X(net518));
 sky130_fd_sc_hd__buf_1 _5427_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 ),
    .X(net519));
 sky130_fd_sc_hd__buf_1 _5428_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 ),
    .X(net520));
 sky130_fd_sc_hd__clkbuf_2 _5429_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 ),
    .X(net521));
 sky130_fd_sc_hd__buf_1 _5430_ (.A(net665),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_1 _5431_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ),
    .X(net523));
 sky130_fd_sc_hd__buf_1 _5432_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .X(net524));
 sky130_fd_sc_hd__buf_1 _5433_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ),
    .X(net525));
 sky130_fd_sc_hd__clkbuf_1 _5434_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ),
    .X(net526));
 sky130_fd_sc_hd__buf_1 _5435_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ),
    .X(net527));
 sky130_fd_sc_hd__buf_1 _5436_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 ),
    .X(net528));
 sky130_fd_sc_hd__clkbuf_1 _5437_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .X(net529));
 sky130_fd_sc_hd__clkbuf_1 _5438_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .X(net530));
 sky130_fd_sc_hd__buf_1 _5439_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ),
    .X(net531));
 sky130_fd_sc_hd__buf_2 _5440_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .X(net532));
 sky130_fd_sc_hd__buf_1 _5441_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .X(net533));
 sky130_fd_sc_hd__buf_4 _5442_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .X(net534));
 sky130_fd_sc_hd__buf_8 _5443_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .X(net535));
 sky130_fd_sc_hd__buf_6 _5444_ (.A(net876),
    .X(net536));
 sky130_fd_sc_hd__buf_1 _5445_ (.A(Tile_X0Y0_S4END[8]),
    .X(net537));
 sky130_fd_sc_hd__buf_1 _5446_ (.A(Tile_X0Y0_S4END[9]),
    .X(net544));
 sky130_fd_sc_hd__buf_1 _5447_ (.A(Tile_X0Y0_S4END[10]),
    .X(net545));
 sky130_fd_sc_hd__buf_1 _5448_ (.A(Tile_X0Y0_S4END[11]),
    .X(net546));
 sky130_fd_sc_hd__buf_1 _5449_ (.A(Tile_X0Y0_S4END[12]),
    .X(net547));
 sky130_fd_sc_hd__buf_1 _5450_ (.A(Tile_X0Y0_S4END[13]),
    .X(net548));
 sky130_fd_sc_hd__buf_1 _5451_ (.A(Tile_X0Y0_S4END[14]),
    .X(net549));
 sky130_fd_sc_hd__buf_4 _5452_ (.A(Tile_X0Y0_S4END[15]),
    .X(net550));
 sky130_fd_sc_hd__buf_4 _5453_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 ),
    .X(net551));
 sky130_fd_sc_hd__buf_4 _5454_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 ),
    .X(net552));
 sky130_fd_sc_hd__buf_4 _5455_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 ),
    .X(net538));
 sky130_fd_sc_hd__buf_4 _5456_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 ),
    .X(net539));
 sky130_fd_sc_hd__buf_1 _5457_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 ),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_2 _5458_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 ),
    .X(net541));
 sky130_fd_sc_hd__buf_1 _5459_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 ),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_1 _5460_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 ),
    .X(net543));
 sky130_fd_sc_hd__buf_4 _5461_ (.A(Tile_X0Y0_SS4END[8]),
    .X(net553));
 sky130_fd_sc_hd__buf_4 _5462_ (.A(Tile_X0Y0_SS4END[9]),
    .X(net560));
 sky130_fd_sc_hd__buf_4 _5463_ (.A(Tile_X0Y0_SS4END[10]),
    .X(net561));
 sky130_fd_sc_hd__buf_4 _5464_ (.A(Tile_X0Y0_SS4END[11]),
    .X(net562));
 sky130_fd_sc_hd__buf_4 _5465_ (.A(Tile_X0Y0_SS4END[12]),
    .X(net563));
 sky130_fd_sc_hd__buf_4 _5466_ (.A(Tile_X0Y0_SS4END[13]),
    .X(net564));
 sky130_fd_sc_hd__buf_4 _5467_ (.A(Tile_X0Y0_SS4END[14]),
    .X(net565));
 sky130_fd_sc_hd__buf_4 _5468_ (.A(Tile_X0Y0_SS4END[15]),
    .X(net566));
 sky130_fd_sc_hd__buf_4 _5469_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 ),
    .X(net567));
 sky130_fd_sc_hd__buf_6 _5470_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 ),
    .X(net568));
 sky130_fd_sc_hd__buf_4 _5471_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 ),
    .X(net554));
 sky130_fd_sc_hd__buf_8 _5472_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 ),
    .X(net555));
 sky130_fd_sc_hd__buf_1 _5473_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 ),
    .X(net556));
 sky130_fd_sc_hd__clkbuf_1 _5474_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 ),
    .X(net557));
 sky130_fd_sc_hd__buf_1 _5475_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(_0211_),
    .X(net651));
 sky130_fd_sc_hd__buf_1 _5477_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 ),
    .X(net569));
 sky130_fd_sc_hd__buf_4 _5478_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 ),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_1 _5479_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 ),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_2 _5480_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 ),
    .X(net572));
 sky130_fd_sc_hd__buf_1 _5481_ (.A(net214),
    .X(net573));
 sky130_fd_sc_hd__clkbuf_1 _5482_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ),
    .X(net574));
 sky130_fd_sc_hd__buf_1 _5483_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_2 _5484_ (.A(net217),
    .X(net576));
 sky130_fd_sc_hd__buf_1 _5485_ (.A(net218),
    .X(net577));
 sky130_fd_sc_hd__buf_6 _5486_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ),
    .X(net578));
 sky130_fd_sc_hd__buf_6 _5487_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 ),
    .X(net579));
 sky130_fd_sc_hd__buf_1 _5488_ (.A(net221),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_2 _5489_ (.A(net222),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_2 _5490_ (.A(net223),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_2 _5491_ (.A(net224),
    .X(net583));
 sky130_fd_sc_hd__buf_4 _5492_ (.A(net225),
    .X(net584));
 sky130_fd_sc_hd__buf_1 _5493_ (.A(net226),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_2 _5494_ (.A(net227),
    .X(net586));
 sky130_fd_sc_hd__buf_4 _5495_ (.A(net228),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_2 _5496_ (.A(net229),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_2 _5497_ (.A(Tile_X0Y1_W6END[2]),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_2 _5498_ (.A(Tile_X0Y1_W6END[3]),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_2 _5499_ (.A(Tile_X0Y1_W6END[4]),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_2 _5500_ (.A(Tile_X0Y1_W6END[5]),
    .X(net594));
 sky130_fd_sc_hd__clkbuf_2 _5501_ (.A(Tile_X0Y1_W6END[6]),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_2 _5502_ (.A(Tile_X0Y1_W6END[7]),
    .X(net596));
 sky130_fd_sc_hd__buf_2 _5503_ (.A(Tile_X0Y1_W6END[8]),
    .X(net597));
 sky130_fd_sc_hd__buf_4 _5504_ (.A(Tile_X0Y1_W6END[9]),
    .X(net598));
 sky130_fd_sc_hd__buf_4 _5505_ (.A(Tile_X0Y1_W6END[10]),
    .X(net599));
 sky130_fd_sc_hd__buf_4 _5506_ (.A(Tile_X0Y1_W6END[11]),
    .X(net600));
 sky130_fd_sc_hd__buf_1 _5507_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 ),
    .X(net590));
 sky130_fd_sc_hd__buf_1 _5508_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 ),
    .X(net591));
 sky130_fd_sc_hd__buf_4 _5509_ (.A(Tile_X0Y1_WW4END[4]),
    .X(net601));
 sky130_fd_sc_hd__buf_4 _5510_ (.A(Tile_X0Y1_WW4END[5]),
    .X(net608));
 sky130_fd_sc_hd__buf_4 _5511_ (.A(Tile_X0Y1_WW4END[6]),
    .X(net609));
 sky130_fd_sc_hd__buf_4 _5512_ (.A(Tile_X0Y1_WW4END[7]),
    .X(net610));
 sky130_fd_sc_hd__buf_4 _5513_ (.A(Tile_X0Y1_WW4END[8]),
    .X(net611));
 sky130_fd_sc_hd__buf_4 _5514_ (.A(Tile_X0Y1_WW4END[9]),
    .X(net612));
 sky130_fd_sc_hd__buf_4 _5515_ (.A(Tile_X0Y1_WW4END[10]),
    .X(net613));
 sky130_fd_sc_hd__buf_4 _5516_ (.A(Tile_X0Y1_WW4END[11]),
    .X(net614));
 sky130_fd_sc_hd__buf_2 _5517_ (.A(Tile_X0Y1_WW4END[12]),
    .X(net615));
 sky130_fd_sc_hd__buf_2 _5518_ (.A(Tile_X0Y1_WW4END[13]),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_2 _5519_ (.A(Tile_X0Y1_WW4END[14]),
    .X(net602));
 sky130_fd_sc_hd__clkbuf_2 _5520_ (.A(Tile_X0Y1_WW4END[15]),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_2 rebuffer294 (.A(net913),
    .X(net911));
 sky130_fd_sc_hd__buf_1 _5522_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 ),
    .X(net605));
 sky130_fd_sc_hd__buf_1 _5523_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 ),
    .X(net606));
 sky130_fd_sc_hd__buf_8 clone36 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .X(net653));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Left_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1585 ();
 sky130_fd_sc_hd__buf_8 fanout966 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .X(net966));
 sky130_fd_sc_hd__clkbuf_2 fanout967 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .X(net967));
 sky130_fd_sc_hd__buf_8 fanout968 (.A(_0340_),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_4 fanout969 (.A(net972),
    .X(net969));
 sky130_fd_sc_hd__buf_8 fanout970 (.A(net972),
    .X(net970));
 sky130_fd_sc_hd__clkbuf_4 fanout971 (.A(net972),
    .X(net971));
 sky130_fd_sc_hd__buf_8 fanout972 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .X(net972));
 sky130_fd_sc_hd__buf_8 fanout973 (.A(net975),
    .X(net973));
 sky130_fd_sc_hd__buf_2 fanout974 (.A(net975),
    .X(net974));
 sky130_fd_sc_hd__buf_8 fanout975 (.A(net976),
    .X(net975));
 sky130_fd_sc_hd__buf_8 fanout976 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .X(net976));
 sky130_fd_sc_hd__buf_8 fanout977 (.A(net979),
    .X(net977));
 sky130_fd_sc_hd__buf_6 fanout978 (.A(net979),
    .X(net978));
 sky130_fd_sc_hd__buf_12 fanout979 (.A(net981),
    .X(net979));
 sky130_fd_sc_hd__buf_2 fanout980 (.A(net981),
    .X(net980));
 sky130_fd_sc_hd__buf_8 fanout981 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .X(net981));
 sky130_fd_sc_hd__buf_8 fanout982 (.A(net986),
    .X(net982));
 sky130_fd_sc_hd__buf_2 fanout983 (.A(net985),
    .X(net983));
 sky130_fd_sc_hd__buf_2 fanout984 (.A(net985),
    .X(net984));
 sky130_fd_sc_hd__buf_2 fanout985 (.A(net986),
    .X(net985));
 sky130_fd_sc_hd__buf_8 fanout986 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .X(net986));
 sky130_fd_sc_hd__buf_6 fanout987 (.A(net988),
    .X(net987));
 sky130_fd_sc_hd__buf_8 fanout988 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .X(net988));
 sky130_fd_sc_hd__buf_2 fanout989 (.A(net990),
    .X(net989));
 sky130_fd_sc_hd__clkbuf_2 fanout990 (.A(net991),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_2 fanout991 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .X(net991));
 sky130_fd_sc_hd__buf_6 fanout992 (.A(net993),
    .X(net992));
 sky130_fd_sc_hd__buf_6 fanout993 (.A(net996),
    .X(net993));
 sky130_fd_sc_hd__buf_8 fanout994 (.A(net996),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_4 fanout995 (.A(net996),
    .X(net995));
 sky130_fd_sc_hd__buf_8 fanout996 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .X(net996));
 sky130_fd_sc_hd__buf_8 fanout997 (.A(net999),
    .X(net997));
 sky130_fd_sc_hd__buf_2 fanout998 (.A(net999),
    .X(net998));
 sky130_fd_sc_hd__buf_8 fanout999 (.A(net1001),
    .X(net999));
 sky130_fd_sc_hd__clkbuf_4 fanout1000 (.A(net1001),
    .X(net1000));
 sky130_fd_sc_hd__buf_8 fanout1001 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .X(net1001));
 sky130_fd_sc_hd__buf_6 fanout1002 (.A(net1003),
    .X(net1002));
 sky130_fd_sc_hd__buf_6 fanout1003 (.A(net1006),
    .X(net1003));
 sky130_fd_sc_hd__buf_2 fanout1004 (.A(net1006),
    .X(net1004));
 sky130_fd_sc_hd__clkbuf_4 fanout1005 (.A(net1006),
    .X(net1005));
 sky130_fd_sc_hd__buf_8 fanout1006 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .X(net1006));
 sky130_fd_sc_hd__clkbuf_4 fanout1007 (.A(net1009),
    .X(net1007));
 sky130_fd_sc_hd__buf_4 fanout1008 (.A(net1009),
    .X(net1008));
 sky130_fd_sc_hd__buf_8 fanout1009 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .X(net1009));
 sky130_fd_sc_hd__clkbuf_4 fanout1010 (.A(net1012),
    .X(net1010));
 sky130_fd_sc_hd__buf_6 fanout1011 (.A(net1012),
    .X(net1011));
 sky130_fd_sc_hd__buf_8 fanout1012 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .X(net1012));
 sky130_fd_sc_hd__buf_8 fanout1013 (.A(_1422_),
    .X(net1013));
 sky130_fd_sc_hd__buf_8 fanout1014 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .X(net1014));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1015 (.A(net1016),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_4 fanout1016 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .X(net1016));
 sky130_fd_sc_hd__buf_8 fanout1017 (.A(net1018),
    .X(net1017));
 sky130_fd_sc_hd__buf_8 fanout1018 (.A(net1020),
    .X(net1018));
 sky130_fd_sc_hd__clkbuf_4 fanout1019 (.A(net1020),
    .X(net1019));
 sky130_fd_sc_hd__buf_8 fanout1020 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .X(net1020));
 sky130_fd_sc_hd__buf_2 fanout1021 (.A(net1022),
    .X(net1021));
 sky130_fd_sc_hd__clkbuf_2 fanout1022 (.A(net1024),
    .X(net1022));
 sky130_fd_sc_hd__buf_2 fanout1023 (.A(net1024),
    .X(net1023));
 sky130_fd_sc_hd__buf_2 fanout1024 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .X(net1024));
 sky130_fd_sc_hd__buf_2 fanout1025 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .X(net1025));
 sky130_fd_sc_hd__buf_8 fanout1026 (.A(net1027),
    .X(net1026));
 sky130_fd_sc_hd__buf_12 fanout1027 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .X(net1027));
 sky130_fd_sc_hd__buf_2 fanout1028 (.A(net1030),
    .X(net1028));
 sky130_fd_sc_hd__buf_1 fanout1029 (.A(net1030),
    .X(net1029));
 sky130_fd_sc_hd__clkbuf_4 fanout1030 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .X(net1030));
 sky130_fd_sc_hd__buf_8 fanout1031 (.A(net1033),
    .X(net1031));
 sky130_fd_sc_hd__buf_4 fanout1032 (.A(net1033),
    .X(net1032));
 sky130_fd_sc_hd__buf_8 fanout1033 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .X(net1033));
 sky130_fd_sc_hd__buf_2 fanout1034 (.A(net1035),
    .X(net1034));
 sky130_fd_sc_hd__clkbuf_2 fanout1035 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .X(net1035));
 sky130_fd_sc_hd__buf_2 fanout1036 (.A(net1039),
    .X(net1036));
 sky130_fd_sc_hd__buf_8 fanout1037 (.A(net1039),
    .X(net1037));
 sky130_fd_sc_hd__clkbuf_4 fanout1038 (.A(net1039),
    .X(net1038));
 sky130_fd_sc_hd__buf_12 fanout1039 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .X(net1039));
 sky130_fd_sc_hd__buf_8 fanout1040 (.A(net1041),
    .X(net1040));
 sky130_fd_sc_hd__buf_8 fanout1041 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .X(net1041));
 sky130_fd_sc_hd__buf_2 fanout1042 (.A(net1044),
    .X(net1042));
 sky130_fd_sc_hd__buf_2 fanout1043 (.A(net1044),
    .X(net1043));
 sky130_fd_sc_hd__clkbuf_4 fanout1044 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .X(net1044));
 sky130_fd_sc_hd__buf_8 fanout1045 (.A(net1046),
    .X(net1045));
 sky130_fd_sc_hd__buf_8 fanout1046 (.A(net1049),
    .X(net1046));
 sky130_fd_sc_hd__buf_2 fanout1047 (.A(net1049),
    .X(net1047));
 sky130_fd_sc_hd__buf_2 fanout1048 (.A(net1049),
    .X(net1048));
 sky130_fd_sc_hd__buf_8 fanout1049 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .X(net1049));
 sky130_fd_sc_hd__buf_6 fanout1050 (.A(net1052),
    .X(net1050));
 sky130_fd_sc_hd__buf_6 fanout1051 (.A(net1052),
    .X(net1051));
 sky130_fd_sc_hd__buf_8 fanout1052 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .X(net1052));
 sky130_fd_sc_hd__buf_2 fanout1053 (.A(net1055),
    .X(net1053));
 sky130_fd_sc_hd__buf_1 fanout1054 (.A(net1055),
    .X(net1054));
 sky130_fd_sc_hd__buf_2 fanout1055 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .X(net1055));
 sky130_fd_sc_hd__buf_8 fanout1056 (.A(net1058),
    .X(net1056));
 sky130_fd_sc_hd__clkbuf_4 fanout1057 (.A(net1058),
    .X(net1057));
 sky130_fd_sc_hd__buf_8 fanout1058 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .X(net1058));
 sky130_fd_sc_hd__buf_4 fanout1059 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .X(net1059));
 sky130_fd_sc_hd__buf_2 fanout1060 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .X(net1060));
 sky130_fd_sc_hd__clkbuf_8 fanout1061 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ),
    .X(net1061));
 sky130_fd_sc_hd__clkbuf_4 fanout1062 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ),
    .X(net1062));
 sky130_fd_sc_hd__clkbuf_4 fanout1063 (.A(net1065),
    .X(net1063));
 sky130_fd_sc_hd__clkbuf_4 fanout1064 (.A(net1065),
    .X(net1064));
 sky130_fd_sc_hd__clkbuf_4 fanout1065 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .X(net1065));
 sky130_fd_sc_hd__buf_2 fanout1066 (.A(net1067),
    .X(net1066));
 sky130_fd_sc_hd__clkbuf_2 fanout1067 (.A(net1069),
    .X(net1067));
 sky130_fd_sc_hd__buf_2 fanout1068 (.A(net1069),
    .X(net1068));
 sky130_fd_sc_hd__clkbuf_4 fanout1069 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .X(net1069));
 sky130_fd_sc_hd__clkbuf_4 fanout1070 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .X(net1070));
 sky130_fd_sc_hd__clkbuf_4 fanout1071 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .X(net1071));
 sky130_fd_sc_hd__buf_4 fanout1072 (.A(net213),
    .X(net1072));
 sky130_fd_sc_hd__clkbuf_4 fanout1073 (.A(net212),
    .X(net1073));
 sky130_fd_sc_hd__clkbuf_2 fanout1074 (.A(net1075),
    .X(net1074));
 sky130_fd_sc_hd__buf_2 fanout1075 (.A(net1077),
    .X(net1075));
 sky130_fd_sc_hd__buf_2 fanout1076 (.A(net1077),
    .X(net1076));
 sky130_fd_sc_hd__clkbuf_2 fanout1077 (.A(Tile_X0Y1_FrameStrobe[9]),
    .X(net1077));
 sky130_fd_sc_hd__buf_2 fanout1078 (.A(Tile_X0Y1_FrameStrobe[9]),
    .X(net1078));
 sky130_fd_sc_hd__clkbuf_2 fanout1079 (.A(Tile_X0Y1_FrameStrobe[9]),
    .X(net1079));
 sky130_fd_sc_hd__clkbuf_4 fanout1080 (.A(net1081),
    .X(net1080));
 sky130_fd_sc_hd__buf_2 fanout1081 (.A(Tile_X0Y1_FrameStrobe[9]),
    .X(net1081));
 sky130_fd_sc_hd__buf_2 fanout1082 (.A(net1085),
    .X(net1082));
 sky130_fd_sc_hd__clkbuf_2 fanout1083 (.A(net1085),
    .X(net1083));
 sky130_fd_sc_hd__buf_2 fanout1084 (.A(net1085),
    .X(net1084));
 sky130_fd_sc_hd__buf_2 fanout1085 (.A(Tile_X0Y1_FrameStrobe[8]),
    .X(net1085));
 sky130_fd_sc_hd__buf_2 fanout1086 (.A(net1089),
    .X(net1086));
 sky130_fd_sc_hd__buf_2 fanout1087 (.A(net1088),
    .X(net1087));
 sky130_fd_sc_hd__buf_2 fanout1088 (.A(net1089),
    .X(net1088));
 sky130_fd_sc_hd__clkbuf_2 fanout1089 (.A(Tile_X0Y1_FrameStrobe[8]),
    .X(net1089));
 sky130_fd_sc_hd__clkbuf_2 fanout1090 (.A(net1091),
    .X(net1090));
 sky130_fd_sc_hd__clkbuf_4 fanout1091 (.A(Tile_X0Y1_FrameStrobe[7]),
    .X(net1091));
 sky130_fd_sc_hd__buf_2 fanout1092 (.A(net1093),
    .X(net1092));
 sky130_fd_sc_hd__clkbuf_2 fanout1093 (.A(Tile_X0Y1_FrameStrobe[7]),
    .X(net1093));
 sky130_fd_sc_hd__buf_2 fanout1094 (.A(net1095),
    .X(net1094));
 sky130_fd_sc_hd__buf_2 fanout1095 (.A(net1097),
    .X(net1095));
 sky130_fd_sc_hd__clkbuf_2 fanout1096 (.A(net1097),
    .X(net1096));
 sky130_fd_sc_hd__clkbuf_2 fanout1097 (.A(Tile_X0Y1_FrameStrobe[7]),
    .X(net1097));
 sky130_fd_sc_hd__clkbuf_4 fanout1098 (.A(net1100),
    .X(net1098));
 sky130_fd_sc_hd__clkbuf_2 fanout1099 (.A(net1100),
    .X(net1099));
 sky130_fd_sc_hd__clkbuf_2 fanout1100 (.A(net1101),
    .X(net1100));
 sky130_fd_sc_hd__clkbuf_4 fanout1101 (.A(net1106),
    .X(net1101));
 sky130_fd_sc_hd__clkbuf_2 fanout1102 (.A(net1106),
    .X(net1102));
 sky130_fd_sc_hd__buf_2 fanout1103 (.A(net1104),
    .X(net1103));
 sky130_fd_sc_hd__buf_1 fanout1104 (.A(net1105),
    .X(net1104));
 sky130_fd_sc_hd__clkbuf_2 fanout1105 (.A(net1106),
    .X(net1105));
 sky130_fd_sc_hd__buf_1 fanout1106 (.A(Tile_X0Y1_FrameStrobe[6]),
    .X(net1106));
 sky130_fd_sc_hd__clkbuf_2 fanout1107 (.A(net1110),
    .X(net1107));
 sky130_fd_sc_hd__buf_1 fanout1108 (.A(net1110),
    .X(net1108));
 sky130_fd_sc_hd__clkbuf_2 fanout1109 (.A(net1110),
    .X(net1109));
 sky130_fd_sc_hd__clkbuf_2 fanout1110 (.A(net1111),
    .X(net1110));
 sky130_fd_sc_hd__clkbuf_2 fanout1111 (.A(Tile_X0Y1_FrameStrobe[5]),
    .X(net1111));
 sky130_fd_sc_hd__buf_2 fanout1112 (.A(Tile_X0Y1_FrameStrobe[5]),
    .X(net1112));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1113 (.A(Tile_X0Y1_FrameStrobe[5]),
    .X(net1113));
 sky130_fd_sc_hd__buf_2 fanout1114 (.A(net1115),
    .X(net1114));
 sky130_fd_sc_hd__clkbuf_2 fanout1115 (.A(Tile_X0Y1_FrameStrobe[5]),
    .X(net1115));
 sky130_fd_sc_hd__clkbuf_2 fanout1116 (.A(net1119),
    .X(net1116));
 sky130_fd_sc_hd__clkbuf_2 fanout1117 (.A(net1118),
    .X(net1117));
 sky130_fd_sc_hd__buf_2 fanout1118 (.A(net1119),
    .X(net1118));
 sky130_fd_sc_hd__clkbuf_2 fanout1119 (.A(Tile_X0Y1_FrameStrobe[4]),
    .X(net1119));
 sky130_fd_sc_hd__clkbuf_2 fanout1120 (.A(net1121),
    .X(net1120));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1121 (.A(net1122),
    .X(net1121));
 sky130_fd_sc_hd__clkbuf_4 fanout1122 (.A(net1123),
    .X(net1122));
 sky130_fd_sc_hd__buf_2 fanout1123 (.A(Tile_X0Y1_FrameStrobe[4]),
    .X(net1123));
 sky130_fd_sc_hd__buf_2 fanout1124 (.A(net1126),
    .X(net1124));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1125 (.A(net1126),
    .X(net1125));
 sky130_fd_sc_hd__clkbuf_2 fanout1126 (.A(net1132),
    .X(net1126));
 sky130_fd_sc_hd__buf_2 fanout1127 (.A(net1132),
    .X(net1127));
 sky130_fd_sc_hd__clkbuf_2 fanout1128 (.A(net1129),
    .X(net1128));
 sky130_fd_sc_hd__clkbuf_2 fanout1129 (.A(net1132),
    .X(net1129));
 sky130_fd_sc_hd__clkbuf_4 fanout1130 (.A(net1132),
    .X(net1130));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1131 (.A(net1132),
    .X(net1131));
 sky130_fd_sc_hd__clkbuf_4 fanout1132 (.A(Tile_X0Y1_FrameStrobe[3]),
    .X(net1132));
 sky130_fd_sc_hd__buf_2 fanout1133 (.A(net1134),
    .X(net1133));
 sky130_fd_sc_hd__clkbuf_2 fanout1134 (.A(Tile_X0Y1_FrameStrobe[2]),
    .X(net1134));
 sky130_fd_sc_hd__clkbuf_2 fanout1135 (.A(net1136),
    .X(net1135));
 sky130_fd_sc_hd__clkbuf_2 fanout1136 (.A(Tile_X0Y1_FrameStrobe[2]),
    .X(net1136));
 sky130_fd_sc_hd__clkbuf_2 fanout1137 (.A(net1138),
    .X(net1137));
 sky130_fd_sc_hd__clkbuf_2 fanout1138 (.A(net1139),
    .X(net1138));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1139 (.A(net1141),
    .X(net1139));
 sky130_fd_sc_hd__clkbuf_4 fanout1140 (.A(net1141),
    .X(net1140));
 sky130_fd_sc_hd__buf_2 fanout1141 (.A(Tile_X0Y1_FrameStrobe[2]),
    .X(net1141));
 sky130_fd_sc_hd__buf_2 fanout1142 (.A(net1150),
    .X(net1142));
 sky130_fd_sc_hd__clkbuf_2 fanout1143 (.A(net1144),
    .X(net1143));
 sky130_fd_sc_hd__buf_1 fanout1144 (.A(net1145),
    .X(net1144));
 sky130_fd_sc_hd__buf_2 fanout1145 (.A(net1150),
    .X(net1145));
 sky130_fd_sc_hd__clkbuf_2 fanout1146 (.A(net1150),
    .X(net1146));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1147 (.A(net1150),
    .X(net1147));
 sky130_fd_sc_hd__buf_2 fanout1148 (.A(net1150),
    .X(net1148));
 sky130_fd_sc_hd__clkbuf_2 fanout1149 (.A(net1150),
    .X(net1149));
 sky130_fd_sc_hd__buf_4 fanout1150 (.A(Tile_X0Y1_FrameStrobe[1]),
    .X(net1150));
 sky130_fd_sc_hd__clkbuf_2 fanout1151 (.A(net1152),
    .X(net1151));
 sky130_fd_sc_hd__clkbuf_2 fanout1152 (.A(net1153),
    .X(net1152));
 sky130_fd_sc_hd__clkbuf_2 fanout1153 (.A(net1155),
    .X(net1153));
 sky130_fd_sc_hd__clkbuf_4 fanout1154 (.A(net1155),
    .X(net1154));
 sky130_fd_sc_hd__clkbuf_1 fanout1155 (.A(Tile_X0Y1_FrameStrobe[12]),
    .X(net1155));
 sky130_fd_sc_hd__buf_2 fanout1156 (.A(net1158),
    .X(net1156));
 sky130_fd_sc_hd__clkbuf_2 fanout1157 (.A(net1158),
    .X(net1157));
 sky130_fd_sc_hd__buf_1 fanout1158 (.A(net1159),
    .X(net1158));
 sky130_fd_sc_hd__buf_2 fanout1159 (.A(Tile_X0Y1_FrameStrobe[12]),
    .X(net1159));
 sky130_fd_sc_hd__buf_2 fanout1160 (.A(net1161),
    .X(net1160));
 sky130_fd_sc_hd__clkbuf_4 fanout1161 (.A(net1162),
    .X(net1161));
 sky130_fd_sc_hd__clkbuf_4 fanout1162 (.A(net1163),
    .X(net1162));
 sky130_fd_sc_hd__clkbuf_2 fanout1163 (.A(Tile_X0Y1_FrameStrobe[11]),
    .X(net1163));
 sky130_fd_sc_hd__buf_2 fanout1164 (.A(net1165),
    .X(net1164));
 sky130_fd_sc_hd__buf_1 fanout1165 (.A(net1167),
    .X(net1165));
 sky130_fd_sc_hd__clkbuf_2 fanout1166 (.A(net1167),
    .X(net1166));
 sky130_fd_sc_hd__clkbuf_2 fanout1167 (.A(net1168),
    .X(net1167));
 sky130_fd_sc_hd__buf_2 fanout1168 (.A(Tile_X0Y1_FrameStrobe[11]),
    .X(net1168));
 sky130_fd_sc_hd__buf_2 fanout1169 (.A(net1170),
    .X(net1169));
 sky130_fd_sc_hd__buf_1 fanout1170 (.A(net1173),
    .X(net1170));
 sky130_fd_sc_hd__buf_2 fanout1171 (.A(net1173),
    .X(net1171));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1172 (.A(net1173),
    .X(net1172));
 sky130_fd_sc_hd__clkbuf_4 fanout1173 (.A(Tile_X0Y1_FrameStrobe[10]),
    .X(net1173));
 sky130_fd_sc_hd__buf_2 fanout1174 (.A(net1176),
    .X(net1174));
 sky130_fd_sc_hd__clkbuf_4 fanout1175 (.A(net1176),
    .X(net1175));
 sky130_fd_sc_hd__buf_2 fanout1176 (.A(Tile_X0Y1_FrameStrobe[10]),
    .X(net1176));
 sky130_fd_sc_hd__clkbuf_2 fanout1177 (.A(Tile_X0Y1_FrameStrobe[10]),
    .X(net1177));
 sky130_fd_sc_hd__buf_2 fanout1178 (.A(net1180),
    .X(net1178));
 sky130_fd_sc_hd__buf_2 fanout1179 (.A(net1180),
    .X(net1179));
 sky130_fd_sc_hd__clkbuf_2 fanout1180 (.A(net1181),
    .X(net1180));
 sky130_fd_sc_hd__clkbuf_2 fanout1181 (.A(Tile_X0Y1_FrameStrobe[0]),
    .X(net1181));
 sky130_fd_sc_hd__buf_2 fanout1182 (.A(net1183),
    .X(net1182));
 sky130_fd_sc_hd__buf_2 fanout1183 (.A(net1185),
    .X(net1183));
 sky130_fd_sc_hd__buf_2 fanout1184 (.A(net1185),
    .X(net1184));
 sky130_fd_sc_hd__clkbuf_2 fanout1185 (.A(Tile_X0Y1_FrameStrobe[0]),
    .X(net1185));
 sky130_fd_sc_hd__clkbuf_4 fanout1186 (.A(net173),
    .X(net1186));
 sky130_fd_sc_hd__clkbuf_4 fanout1187 (.A(net172),
    .X(net1187));
 sky130_fd_sc_hd__clkbuf_4 fanout1188 (.A(net171),
    .X(net1188));
 sky130_fd_sc_hd__clkbuf_4 fanout1189 (.A(net170),
    .X(net1189));
 sky130_fd_sc_hd__buf_4 fanout1190 (.A(net169),
    .X(net1190));
 sky130_fd_sc_hd__clkbuf_4 fanout1191 (.A(net168),
    .X(net1191));
 sky130_fd_sc_hd__buf_4 fanout1192 (.A(net167),
    .X(net1192));
 sky130_fd_sc_hd__buf_4 fanout1193 (.A(net166),
    .X(net1193));
 sky130_fd_sc_hd__buf_4 fanout1194 (.A(net165),
    .X(net1194));
 sky130_fd_sc_hd__clkbuf_4 fanout1195 (.A(net164),
    .X(net1195));
 sky130_fd_sc_hd__buf_4 fanout1196 (.A(net163),
    .X(net1196));
 sky130_fd_sc_hd__clkbuf_4 fanout1197 (.A(net162),
    .X(net1197));
 sky130_fd_sc_hd__buf_4 fanout1198 (.A(net161),
    .X(net1198));
 sky130_fd_sc_hd__clkbuf_4 fanout1199 (.A(net160),
    .X(net1199));
 sky130_fd_sc_hd__buf_4 fanout1200 (.A(net159),
    .X(net1200));
 sky130_fd_sc_hd__clkbuf_4 fanout1201 (.A(net1202),
    .X(net1201));
 sky130_fd_sc_hd__clkbuf_2 fanout1202 (.A(Tile_X0Y1_FrameData[24]),
    .X(net1202));
 sky130_fd_sc_hd__clkbuf_4 fanout1203 (.A(net1204),
    .X(net1203));
 sky130_fd_sc_hd__clkbuf_2 fanout1204 (.A(Tile_X0Y1_FrameData[23]),
    .X(net1204));
 sky130_fd_sc_hd__buf_4 fanout1205 (.A(net1206),
    .X(net1205));
 sky130_fd_sc_hd__clkbuf_2 fanout1206 (.A(Tile_X0Y1_FrameData[22]),
    .X(net1206));
 sky130_fd_sc_hd__buf_4 fanout1207 (.A(net158),
    .X(net1207));
 sky130_fd_sc_hd__buf_4 fanout1208 (.A(net157),
    .X(net1208));
 sky130_fd_sc_hd__buf_4 fanout1209 (.A(net156),
    .X(net1209));
 sky130_fd_sc_hd__buf_4 fanout1210 (.A(net155),
    .X(net1210));
 sky130_fd_sc_hd__buf_4 fanout1211 (.A(net154),
    .X(net1211));
 sky130_fd_sc_hd__buf_4 fanout1212 (.A(net153),
    .X(net1212));
 sky130_fd_sc_hd__buf_4 fanout1213 (.A(net152),
    .X(net1213));
 sky130_fd_sc_hd__buf_4 fanout1214 (.A(net151),
    .X(net1214));
 sky130_fd_sc_hd__clkbuf_4 fanout1215 (.A(net150),
    .X(net1215));
 sky130_fd_sc_hd__clkbuf_4 fanout1216 (.A(net149),
    .X(net1216));
 sky130_fd_sc_hd__buf_4 fanout1217 (.A(net148),
    .X(net1217));
 sky130_fd_sc_hd__buf_4 fanout1218 (.A(net147),
    .X(net1218));
 sky130_fd_sc_hd__clkbuf_4 fanout1219 (.A(net146),
    .X(net1219));
 sky130_fd_sc_hd__buf_4 fanout1220 (.A(net145),
    .X(net1220));
 sky130_fd_sc_hd__buf_2 fanout1221 (.A(net140),
    .X(net1221));
 sky130_fd_sc_hd__clkbuf_4 fanout1222 (.A(net139),
    .X(net1222));
 sky130_fd_sc_hd__buf_4 fanout1223 (.A(net122),
    .X(net1223));
 sky130_fd_sc_hd__clkbuf_4 fanout1224 (.A(net121),
    .X(net1224));
 sky130_fd_sc_hd__clkbuf_4 fanout1225 (.A(net96),
    .X(net1225));
 sky130_fd_sc_hd__clkbuf_4 fanout1226 (.A(net95),
    .X(net1226));
 sky130_fd_sc_hd__clkbuf_4 fanout1227 (.A(net56),
    .X(net1227));
 sky130_fd_sc_hd__clkbuf_4 fanout1228 (.A(net55),
    .X(net1228));
 sky130_fd_sc_hd__clkbuf_4 fanout1229 (.A(net54),
    .X(net1229));
 sky130_fd_sc_hd__buf_4 fanout1230 (.A(net53),
    .X(net1230));
 sky130_fd_sc_hd__buf_4 fanout1231 (.A(net52),
    .X(net1231));
 sky130_fd_sc_hd__buf_4 fanout1232 (.A(net51),
    .X(net1232));
 sky130_fd_sc_hd__clkbuf_4 fanout1233 (.A(net50),
    .X(net1233));
 sky130_fd_sc_hd__buf_4 fanout1234 (.A(net49),
    .X(net1234));
 sky130_fd_sc_hd__clkbuf_4 fanout1235 (.A(net48),
    .X(net1235));
 sky130_fd_sc_hd__buf_4 fanout1236 (.A(net47),
    .X(net1236));
 sky130_fd_sc_hd__buf_4 fanout1237 (.A(net46),
    .X(net1237));
 sky130_fd_sc_hd__buf_4 fanout1238 (.A(net45),
    .X(net1238));
 sky130_fd_sc_hd__buf_4 fanout1239 (.A(net44),
    .X(net1239));
 sky130_fd_sc_hd__buf_2 fanout1240 (.A(net43),
    .X(net1240));
 sky130_fd_sc_hd__buf_4 fanout1241 (.A(net1242),
    .X(net1241));
 sky130_fd_sc_hd__clkbuf_2 fanout1242 (.A(Tile_X0Y0_FrameData[25]),
    .X(net1242));
 sky130_fd_sc_hd__buf_4 fanout1243 (.A(net1244),
    .X(net1243));
 sky130_fd_sc_hd__clkbuf_2 fanout1244 (.A(Tile_X0Y0_FrameData[24]),
    .X(net1244));
 sky130_fd_sc_hd__buf_4 fanout1245 (.A(net42),
    .X(net1245));
 sky130_fd_sc_hd__clkbuf_4 fanout1246 (.A(net41),
    .X(net1246));
 sky130_fd_sc_hd__clkbuf_4 fanout1247 (.A(net40),
    .X(net1247));
 sky130_fd_sc_hd__buf_4 fanout1248 (.A(net39),
    .X(net1248));
 sky130_fd_sc_hd__buf_4 fanout1249 (.A(net38),
    .X(net1249));
 sky130_fd_sc_hd__clkbuf_4 fanout1250 (.A(net37),
    .X(net1250));
 sky130_fd_sc_hd__clkbuf_4 fanout1251 (.A(net36),
    .X(net1251));
 sky130_fd_sc_hd__buf_4 fanout1252 (.A(net35),
    .X(net1252));
 sky130_fd_sc_hd__buf_4 fanout1253 (.A(net34),
    .X(net1253));
 sky130_fd_sc_hd__clkbuf_4 fanout1254 (.A(net33),
    .X(net1254));
 sky130_fd_sc_hd__clkbuf_4 fanout1255 (.A(net32),
    .X(net1255));
 sky130_fd_sc_hd__buf_4 fanout1256 (.A(net31),
    .X(net1256));
 sky130_fd_sc_hd__buf_4 fanout1257 (.A(net30),
    .X(net1257));
 sky130_fd_sc_hd__clkbuf_4 fanout1258 (.A(net29),
    .X(net1258));
 sky130_fd_sc_hd__clkbuf_4 fanout1259 (.A(net28),
    .X(net1259));
 sky130_fd_sc_hd__buf_4 fanout1260 (.A(net27),
    .X(net1260));
 sky130_fd_sc_hd__clkbuf_4 fanout1261 (.A(net22),
    .X(net1261));
 sky130_fd_sc_hd__clkbuf_4 fanout1262 (.A(net21),
    .X(net1262));
 sky130_fd_sc_hd__clkbuf_4 fanout1263 (.A(net4),
    .X(net1263));
 sky130_fd_sc_hd__buf_4 fanout1264 (.A(net3),
    .X(net1264));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(Tile_X0Y0_E1END[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(Tile_X0Y0_E1END[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(Tile_X0Y0_E1END[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(Tile_X0Y0_E1END[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(Tile_X0Y0_E2END[0]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(Tile_X0Y0_E2END[1]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(Tile_X0Y0_E2END[2]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(Tile_X0Y0_E2END[3]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(Tile_X0Y0_E2END[4]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(Tile_X0Y0_E2END[5]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(Tile_X0Y0_E2END[6]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(Tile_X0Y0_E2END[7]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(Tile_X0Y0_E2MID[0]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(Tile_X0Y0_E2MID[1]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(Tile_X0Y0_E2MID[2]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(Tile_X0Y0_E2MID[3]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(Tile_X0Y0_E2MID[4]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(Tile_X0Y0_E2MID[5]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(Tile_X0Y0_E2MID[6]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input20 (.A(Tile_X0Y0_E2MID[7]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(Tile_X0Y0_E6END[0]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(Tile_X0Y0_E6END[1]),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input23 (.A(Tile_X0Y0_EE4END[0]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(Tile_X0Y0_EE4END[1]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(Tile_X0Y0_EE4END[2]),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(Tile_X0Y0_EE4END[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_2 input27 (.A(Tile_X0Y0_FrameData[0]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(Tile_X0Y0_FrameData[10]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(Tile_X0Y0_FrameData[11]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input30 (.A(Tile_X0Y0_FrameData[12]),
    .X(net30));
 sky130_fd_sc_hd__buf_2 input31 (.A(Tile_X0Y0_FrameData[13]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input32 (.A(Tile_X0Y0_FrameData[14]),
    .X(net32));
 sky130_fd_sc_hd__buf_2 input33 (.A(Tile_X0Y0_FrameData[15]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(Tile_X0Y0_FrameData[16]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(Tile_X0Y0_FrameData[17]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(Tile_X0Y0_FrameData[18]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(Tile_X0Y0_FrameData[19]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 input38 (.A(Tile_X0Y0_FrameData[1]),
    .X(net38));
 sky130_fd_sc_hd__buf_2 input39 (.A(Tile_X0Y0_FrameData[20]),
    .X(net39));
 sky130_fd_sc_hd__buf_2 input40 (.A(Tile_X0Y0_FrameData[21]),
    .X(net40));
 sky130_fd_sc_hd__buf_2 input41 (.A(Tile_X0Y0_FrameData[22]),
    .X(net41));
 sky130_fd_sc_hd__buf_2 input42 (.A(Tile_X0Y0_FrameData[23]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(Tile_X0Y0_FrameData[26]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 input44 (.A(Tile_X0Y0_FrameData[27]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 input45 (.A(Tile_X0Y0_FrameData[28]),
    .X(net45));
 sky130_fd_sc_hd__buf_2 input46 (.A(Tile_X0Y0_FrameData[29]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(Tile_X0Y0_FrameData[2]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(Tile_X0Y0_FrameData[30]),
    .X(net48));
 sky130_fd_sc_hd__buf_2 input49 (.A(Tile_X0Y0_FrameData[31]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(Tile_X0Y0_FrameData[3]),
    .X(net50));
 sky130_fd_sc_hd__buf_2 input51 (.A(Tile_X0Y0_FrameData[4]),
    .X(net51));
 sky130_fd_sc_hd__buf_2 input52 (.A(Tile_X0Y0_FrameData[5]),
    .X(net52));
 sky130_fd_sc_hd__buf_2 input53 (.A(Tile_X0Y0_FrameData[6]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(Tile_X0Y0_FrameData[7]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(Tile_X0Y0_FrameData[8]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(Tile_X0Y0_FrameData[9]),
    .X(net56));
 sky130_fd_sc_hd__buf_6 input57 (.A(Tile_X0Y0_S1END[0]),
    .X(net57));
 sky130_fd_sc_hd__buf_2 input58 (.A(Tile_X0Y0_S1END[1]),
    .X(net58));
 sky130_fd_sc_hd__buf_6 input59 (.A(Tile_X0Y0_S1END[2]),
    .X(net59));
 sky130_fd_sc_hd__buf_2 input60 (.A(Tile_X0Y0_S1END[3]),
    .X(net60));
 sky130_fd_sc_hd__buf_6 input61 (.A(Tile_X0Y0_S2END[0]),
    .X(net61));
 sky130_fd_sc_hd__buf_2 input62 (.A(Tile_X0Y0_S2END[1]),
    .X(net62));
 sky130_fd_sc_hd__buf_2 input63 (.A(Tile_X0Y0_S2END[2]),
    .X(net63));
 sky130_fd_sc_hd__buf_2 input64 (.A(Tile_X0Y0_S2END[3]),
    .X(net64));
 sky130_fd_sc_hd__buf_2 input65 (.A(Tile_X0Y0_S2END[4]),
    .X(net65));
 sky130_fd_sc_hd__buf_2 input66 (.A(Tile_X0Y0_S2END[5]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 input67 (.A(Tile_X0Y0_S2END[6]),
    .X(net67));
 sky130_fd_sc_hd__buf_2 input68 (.A(Tile_X0Y0_S2END[7]),
    .X(net68));
 sky130_fd_sc_hd__buf_4 input69 (.A(Tile_X0Y0_S2MID[0]),
    .X(net69));
 sky130_fd_sc_hd__buf_4 input70 (.A(Tile_X0Y0_S2MID[1]),
    .X(net70));
 sky130_fd_sc_hd__buf_4 input71 (.A(Tile_X0Y0_S2MID[2]),
    .X(net71));
 sky130_fd_sc_hd__buf_4 input72 (.A(Tile_X0Y0_S2MID[3]),
    .X(net72));
 sky130_fd_sc_hd__buf_4 input73 (.A(Tile_X0Y0_S2MID[4]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_4 input74 (.A(Tile_X0Y0_S2MID[5]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_4 input75 (.A(Tile_X0Y0_S2MID[6]),
    .X(net75));
 sky130_fd_sc_hd__buf_4 input76 (.A(Tile_X0Y0_S2MID[7]),
    .X(net76));
 sky130_fd_sc_hd__buf_2 input77 (.A(Tile_X0Y0_S4END[0]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_4 input78 (.A(Tile_X0Y0_S4END[1]),
    .X(net78));
 sky130_fd_sc_hd__buf_2 input79 (.A(Tile_X0Y0_S4END[2]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(Tile_X0Y0_S4END[3]),
    .X(net80));
 sky130_fd_sc_hd__buf_4 input81 (.A(Tile_X0Y0_S4END[4]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 input82 (.A(Tile_X0Y0_S4END[5]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 input83 (.A(Tile_X0Y0_S4END[6]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 input84 (.A(Tile_X0Y0_S4END[7]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(Tile_X0Y0_SS4END[0]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(Tile_X0Y0_SS4END[1]),
    .X(net86));
 sky130_fd_sc_hd__buf_2 input87 (.A(Tile_X0Y0_SS4END[2]),
    .X(net87));
 sky130_fd_sc_hd__dlymetal6s2s_1 input88 (.A(Tile_X0Y0_SS4END[3]),
    .X(net88));
 sky130_fd_sc_hd__buf_2 input89 (.A(Tile_X0Y0_SS4END[4]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 input90 (.A(Tile_X0Y0_SS4END[5]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_4 input91 (.A(Tile_X0Y0_SS4END[6]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 input92 (.A(Tile_X0Y0_SS4END[7]),
    .X(net92));
 sky130_fd_sc_hd__buf_12 input93 (.A(Tile_X0Y0_W1END[0]),
    .X(net93));
 sky130_fd_sc_hd__buf_4 input94 (.A(Tile_X0Y0_W1END[1]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(Tile_X0Y0_W1END[2]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 input96 (.A(Tile_X0Y0_W1END[3]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(Tile_X0Y0_W2END[0]),
    .X(net97));
 sky130_fd_sc_hd__buf_2 input98 (.A(Tile_X0Y0_W2END[1]),
    .X(net98));
 sky130_fd_sc_hd__buf_2 input99 (.A(Tile_X0Y0_W2END[2]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_4 input100 (.A(Tile_X0Y0_W2END[3]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_4 input101 (.A(Tile_X0Y0_W2END[4]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 input102 (.A(Tile_X0Y0_W2END[5]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 input103 (.A(Tile_X0Y0_W2END[6]),
    .X(net103));
 sky130_fd_sc_hd__buf_2 input104 (.A(Tile_X0Y0_W2END[7]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 input105 (.A(Tile_X0Y0_W2MID[0]),
    .X(net105));
 sky130_fd_sc_hd__dlymetal6s2s_1 input106 (.A(Tile_X0Y0_W2MID[1]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 input107 (.A(Tile_X0Y0_W2MID[2]),
    .X(net107));
 sky130_fd_sc_hd__buf_2 input108 (.A(Tile_X0Y0_W2MID[3]),
    .X(net108));
 sky130_fd_sc_hd__dlymetal6s2s_1 input109 (.A(Tile_X0Y0_W2MID[4]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input110 (.A(Tile_X0Y0_W2MID[5]),
    .X(net110));
 sky130_fd_sc_hd__buf_2 input111 (.A(Tile_X0Y0_W2MID[6]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 input112 (.A(Tile_X0Y0_W2MID[7]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 input113 (.A(Tile_X0Y0_W6END[0]),
    .X(net113));
 sky130_fd_sc_hd__buf_4 input114 (.A(Tile_X0Y0_W6END[1]),
    .X(net114));
 sky130_fd_sc_hd__buf_2 input115 (.A(Tile_X0Y0_WW4END[0]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 input116 (.A(Tile_X0Y0_WW4END[1]),
    .X(net116));
 sky130_fd_sc_hd__buf_2 input117 (.A(Tile_X0Y0_WW4END[2]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 input118 (.A(Tile_X0Y0_WW4END[3]),
    .X(net118));
 sky130_fd_sc_hd__buf_2 input119 (.A(Tile_X0Y1_E1END[0]),
    .X(net119));
 sky130_fd_sc_hd__buf_4 input120 (.A(Tile_X0Y1_E1END[1]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 input121 (.A(Tile_X0Y1_E1END[2]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 input122 (.A(Tile_X0Y1_E1END[3]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 input123 (.A(Tile_X0Y1_E2END[0]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input124 (.A(Tile_X0Y1_E2END[1]),
    .X(net124));
 sky130_fd_sc_hd__buf_2 input125 (.A(Tile_X0Y1_E2END[2]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_4 input126 (.A(Tile_X0Y1_E2END[3]),
    .X(net126));
 sky130_fd_sc_hd__buf_1 input127 (.A(Tile_X0Y1_E2END[4]),
    .X(net127));
 sky130_fd_sc_hd__buf_2 input128 (.A(Tile_X0Y1_E2END[5]),
    .X(net128));
 sky130_fd_sc_hd__buf_2 input129 (.A(Tile_X0Y1_E2END[6]),
    .X(net129));
 sky130_fd_sc_hd__buf_2 input130 (.A(Tile_X0Y1_E2END[7]),
    .X(net130));
 sky130_fd_sc_hd__buf_2 input131 (.A(Tile_X0Y1_E2MID[0]),
    .X(net131));
 sky130_fd_sc_hd__buf_2 input132 (.A(Tile_X0Y1_E2MID[1]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 input133 (.A(Tile_X0Y1_E2MID[2]),
    .X(net133));
 sky130_fd_sc_hd__buf_2 input134 (.A(Tile_X0Y1_E2MID[3]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 input135 (.A(Tile_X0Y1_E2MID[4]),
    .X(net135));
 sky130_fd_sc_hd__buf_2 input136 (.A(Tile_X0Y1_E2MID[5]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_4 input137 (.A(Tile_X0Y1_E2MID[6]),
    .X(net137));
 sky130_fd_sc_hd__buf_2 input138 (.A(Tile_X0Y1_E2MID[7]),
    .X(net138));
 sky130_fd_sc_hd__buf_1 input139 (.A(Tile_X0Y1_E6END[0]),
    .X(net139));
 sky130_fd_sc_hd__buf_1 input140 (.A(Tile_X0Y1_E6END[1]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_2 input141 (.A(Tile_X0Y1_EE4END[0]),
    .X(net141));
 sky130_fd_sc_hd__dlymetal6s2s_1 input142 (.A(Tile_X0Y1_EE4END[1]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 input143 (.A(Tile_X0Y1_EE4END[2]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 input144 (.A(Tile_X0Y1_EE4END[3]),
    .X(net144));
 sky130_fd_sc_hd__buf_2 input145 (.A(Tile_X0Y1_FrameData[0]),
    .X(net145));
 sky130_fd_sc_hd__buf_2 input146 (.A(Tile_X0Y1_FrameData[10]),
    .X(net146));
 sky130_fd_sc_hd__buf_2 input147 (.A(Tile_X0Y1_FrameData[11]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 input148 (.A(Tile_X0Y1_FrameData[12]),
    .X(net148));
 sky130_fd_sc_hd__buf_2 input149 (.A(Tile_X0Y1_FrameData[13]),
    .X(net149));
 sky130_fd_sc_hd__buf_2 input150 (.A(Tile_X0Y1_FrameData[14]),
    .X(net150));
 sky130_fd_sc_hd__buf_2 input151 (.A(Tile_X0Y1_FrameData[15]),
    .X(net151));
 sky130_fd_sc_hd__buf_2 input152 (.A(Tile_X0Y1_FrameData[16]),
    .X(net152));
 sky130_fd_sc_hd__buf_2 input153 (.A(Tile_X0Y1_FrameData[17]),
    .X(net153));
 sky130_fd_sc_hd__buf_2 input154 (.A(Tile_X0Y1_FrameData[18]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_4 input155 (.A(Tile_X0Y1_FrameData[19]),
    .X(net155));
 sky130_fd_sc_hd__buf_2 input156 (.A(Tile_X0Y1_FrameData[1]),
    .X(net156));
 sky130_fd_sc_hd__buf_2 input157 (.A(Tile_X0Y1_FrameData[20]),
    .X(net157));
 sky130_fd_sc_hd__buf_2 input158 (.A(Tile_X0Y1_FrameData[21]),
    .X(net158));
 sky130_fd_sc_hd__buf_2 input159 (.A(Tile_X0Y1_FrameData[25]),
    .X(net159));
 sky130_fd_sc_hd__buf_2 input160 (.A(Tile_X0Y1_FrameData[26]),
    .X(net160));
 sky130_fd_sc_hd__buf_2 input161 (.A(Tile_X0Y1_FrameData[27]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 input162 (.A(Tile_X0Y1_FrameData[28]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_4 input163 (.A(Tile_X0Y1_FrameData[29]),
    .X(net163));
 sky130_fd_sc_hd__buf_2 input164 (.A(Tile_X0Y1_FrameData[2]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_4 input165 (.A(Tile_X0Y1_FrameData[30]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_4 input166 (.A(Tile_X0Y1_FrameData[31]),
    .X(net166));
 sky130_fd_sc_hd__buf_2 input167 (.A(Tile_X0Y1_FrameData[3]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_4 input168 (.A(Tile_X0Y1_FrameData[4]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_4 input169 (.A(Tile_X0Y1_FrameData[5]),
    .X(net169));
 sky130_fd_sc_hd__buf_2 input170 (.A(Tile_X0Y1_FrameData[6]),
    .X(net170));
 sky130_fd_sc_hd__buf_2 input171 (.A(Tile_X0Y1_FrameData[7]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 input172 (.A(Tile_X0Y1_FrameData[8]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_2 input173 (.A(Tile_X0Y1_FrameData[9]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_4 input174 (.A(Tile_X0Y1_N1END[0]),
    .X(net174));
 sky130_fd_sc_hd__buf_4 input175 (.A(Tile_X0Y1_N1END[1]),
    .X(net175));
 sky130_fd_sc_hd__buf_4 input176 (.A(Tile_X0Y1_N1END[2]),
    .X(net176));
 sky130_fd_sc_hd__buf_4 input177 (.A(Tile_X0Y1_N1END[3]),
    .X(net177));
 sky130_fd_sc_hd__buf_2 input178 (.A(Tile_X0Y1_N2END[0]),
    .X(net178));
 sky130_fd_sc_hd__buf_2 input179 (.A(Tile_X0Y1_N2END[1]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 input180 (.A(Tile_X0Y1_N2END[2]),
    .X(net180));
 sky130_fd_sc_hd__buf_2 input181 (.A(Tile_X0Y1_N2END[3]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_2 input182 (.A(Tile_X0Y1_N2END[4]),
    .X(net182));
 sky130_fd_sc_hd__buf_2 input183 (.A(Tile_X0Y1_N2END[5]),
    .X(net183));
 sky130_fd_sc_hd__buf_2 input184 (.A(Tile_X0Y1_N2END[6]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_4 input185 (.A(Tile_X0Y1_N2END[7]),
    .X(net185));
 sky130_fd_sc_hd__buf_6 input186 (.A(Tile_X0Y1_N2MID[0]),
    .X(net186));
 sky130_fd_sc_hd__buf_4 input187 (.A(Tile_X0Y1_N2MID[1]),
    .X(net187));
 sky130_fd_sc_hd__buf_4 input188 (.A(Tile_X0Y1_N2MID[2]),
    .X(net188));
 sky130_fd_sc_hd__buf_4 input189 (.A(Tile_X0Y1_N2MID[3]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_4 input190 (.A(Tile_X0Y1_N2MID[4]),
    .X(net190));
 sky130_fd_sc_hd__buf_4 input191 (.A(Tile_X0Y1_N2MID[5]),
    .X(net191));
 sky130_fd_sc_hd__buf_4 input192 (.A(Tile_X0Y1_N2MID[6]),
    .X(net192));
 sky130_fd_sc_hd__buf_4 input193 (.A(Tile_X0Y1_N2MID[7]),
    .X(net193));
 sky130_fd_sc_hd__buf_2 input194 (.A(Tile_X0Y1_N4END[0]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 input195 (.A(Tile_X0Y1_N4END[1]),
    .X(net195));
 sky130_fd_sc_hd__buf_2 input196 (.A(Tile_X0Y1_N4END[2]),
    .X(net196));
 sky130_fd_sc_hd__buf_2 input197 (.A(Tile_X0Y1_N4END[3]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_4 input198 (.A(Tile_X0Y1_N4END[4]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_4 input199 (.A(Tile_X0Y1_N4END[5]),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_4 input200 (.A(Tile_X0Y1_N4END[6]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_4 input201 (.A(Tile_X0Y1_N4END[7]),
    .X(net201));
 sky130_fd_sc_hd__buf_1 input202 (.A(Tile_X0Y1_NN4END[0]),
    .X(net202));
 sky130_fd_sc_hd__buf_2 input203 (.A(Tile_X0Y1_NN4END[1]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 input204 (.A(Tile_X0Y1_NN4END[2]),
    .X(net204));
 sky130_fd_sc_hd__buf_2 input205 (.A(Tile_X0Y1_NN4END[3]),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_2 input206 (.A(Tile_X0Y1_NN4END[4]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_4 input207 (.A(Tile_X0Y1_NN4END[5]),
    .X(net207));
 sky130_fd_sc_hd__buf_2 input208 (.A(Tile_X0Y1_NN4END[6]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_4 input209 (.A(Tile_X0Y1_NN4END[7]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_4 input210 (.A(Tile_X0Y1_W1END[0]),
    .X(net210));
 sky130_fd_sc_hd__buf_4 input211 (.A(Tile_X0Y1_W1END[1]),
    .X(net211));
 sky130_fd_sc_hd__buf_1 input212 (.A(Tile_X0Y1_W1END[2]),
    .X(net212));
 sky130_fd_sc_hd__buf_1 input213 (.A(Tile_X0Y1_W1END[3]),
    .X(net213));
 sky130_fd_sc_hd__dlymetal6s2s_1 input214 (.A(Tile_X0Y1_W2END[0]),
    .X(net214));
 sky130_fd_sc_hd__buf_2 input215 (.A(Tile_X0Y1_W2END[1]),
    .X(net215));
 sky130_fd_sc_hd__buf_2 input216 (.A(Tile_X0Y1_W2END[2]),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_4 input217 (.A(Tile_X0Y1_W2END[3]),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_4 input218 (.A(Tile_X0Y1_W2END[4]),
    .X(net218));
 sky130_fd_sc_hd__dlymetal6s2s_1 input219 (.A(Tile_X0Y1_W2END[5]),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 input220 (.A(Tile_X0Y1_W2END[6]),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_2 input221 (.A(Tile_X0Y1_W2END[7]),
    .X(net221));
 sky130_fd_sc_hd__buf_2 input222 (.A(Tile_X0Y1_W2MID[0]),
    .X(net222));
 sky130_fd_sc_hd__buf_2 input223 (.A(Tile_X0Y1_W2MID[1]),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_2 input224 (.A(Tile_X0Y1_W2MID[2]),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_2 input225 (.A(Tile_X0Y1_W2MID[3]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_2 input226 (.A(Tile_X0Y1_W2MID[4]),
    .X(net226));
 sky130_fd_sc_hd__dlymetal6s2s_1 input227 (.A(Tile_X0Y1_W2MID[5]),
    .X(net227));
 sky130_fd_sc_hd__buf_2 input228 (.A(Tile_X0Y1_W2MID[6]),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_4 input229 (.A(Tile_X0Y1_W2MID[7]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_4 input230 (.A(Tile_X0Y1_W6END[0]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_4 input231 (.A(Tile_X0Y1_W6END[1]),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 input232 (.A(Tile_X0Y1_WW4END[0]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_2 input233 (.A(Tile_X0Y1_WW4END[1]),
    .X(net233));
 sky130_fd_sc_hd__buf_2 input234 (.A(Tile_X0Y1_WW4END[2]),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_2 input235 (.A(Tile_X0Y1_WW4END[3]),
    .X(net235));
 sky130_fd_sc_hd__buf_2 output236 (.A(net236),
    .X(Tile_X0Y0_E1BEG[0]));
 sky130_fd_sc_hd__buf_2 output237 (.A(net237),
    .X(Tile_X0Y0_E1BEG[1]));
 sky130_fd_sc_hd__buf_8 output238 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 ),
    .X(Tile_X0Y0_E1BEG[2]));
 sky130_fd_sc_hd__buf_2 output239 (.A(net239),
    .X(Tile_X0Y0_E1BEG[3]));
 sky130_fd_sc_hd__buf_2 output240 (.A(net240),
    .X(Tile_X0Y0_E2BEG[0]));
 sky130_fd_sc_hd__buf_2 output241 (.A(net241),
    .X(Tile_X0Y0_E2BEG[1]));
 sky130_fd_sc_hd__buf_4 output242 (.A(net242),
    .X(Tile_X0Y0_E2BEG[2]));
 sky130_fd_sc_hd__buf_2 output243 (.A(net243),
    .X(Tile_X0Y0_E2BEG[3]));
 sky130_fd_sc_hd__buf_2 output244 (.A(net244),
    .X(Tile_X0Y0_E2BEG[4]));
 sky130_fd_sc_hd__buf_2 output245 (.A(net245),
    .X(Tile_X0Y0_E2BEG[5]));
 sky130_fd_sc_hd__buf_8 output246 (.A(net246),
    .X(Tile_X0Y0_E2BEG[6]));
 sky130_fd_sc_hd__buf_2 output247 (.A(net247),
    .X(Tile_X0Y0_E2BEG[7]));
 sky130_fd_sc_hd__buf_2 output248 (.A(net248),
    .X(Tile_X0Y0_E2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output249 (.A(net249),
    .X(Tile_X0Y0_E2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output250 (.A(net250),
    .X(Tile_X0Y0_E2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output251 (.A(net251),
    .X(Tile_X0Y0_E2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output252 (.A(net252),
    .X(Tile_X0Y0_E2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output253 (.A(net253),
    .X(Tile_X0Y0_E2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output254 (.A(net254),
    .X(Tile_X0Y0_E2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output255 (.A(net255),
    .X(Tile_X0Y0_E2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output256 (.A(net256),
    .X(Tile_X0Y0_E6BEG[0]));
 sky130_fd_sc_hd__buf_8 output257 (.A(net257),
    .X(Tile_X0Y0_E6BEG[10]));
 sky130_fd_sc_hd__buf_6 output258 (.A(net258),
    .X(Tile_X0Y0_E6BEG[11]));
 sky130_fd_sc_hd__buf_2 output259 (.A(net259),
    .X(Tile_X0Y0_E6BEG[1]));
 sky130_fd_sc_hd__buf_2 output260 (.A(net260),
    .X(Tile_X0Y0_E6BEG[2]));
 sky130_fd_sc_hd__buf_2 output261 (.A(net261),
    .X(Tile_X0Y0_E6BEG[3]));
 sky130_fd_sc_hd__buf_2 output262 (.A(net262),
    .X(Tile_X0Y0_E6BEG[4]));
 sky130_fd_sc_hd__buf_2 output263 (.A(net263),
    .X(Tile_X0Y0_E6BEG[5]));
 sky130_fd_sc_hd__buf_2 output264 (.A(net264),
    .X(Tile_X0Y0_E6BEG[6]));
 sky130_fd_sc_hd__buf_2 output265 (.A(net265),
    .X(Tile_X0Y0_E6BEG[7]));
 sky130_fd_sc_hd__buf_2 output266 (.A(net266),
    .X(Tile_X0Y0_E6BEG[8]));
 sky130_fd_sc_hd__buf_2 output267 (.A(net267),
    .X(Tile_X0Y0_E6BEG[9]));
 sky130_fd_sc_hd__buf_2 output268 (.A(net268),
    .X(Tile_X0Y0_EE4BEG[0]));
 sky130_fd_sc_hd__buf_2 output269 (.A(net269),
    .X(Tile_X0Y0_EE4BEG[10]));
 sky130_fd_sc_hd__buf_2 output270 (.A(net270),
    .X(Tile_X0Y0_EE4BEG[11]));
 sky130_fd_sc_hd__buf_2 output271 (.A(net271),
    .X(Tile_X0Y0_EE4BEG[12]));
 sky130_fd_sc_hd__buf_8 output272 (.A(net272),
    .X(Tile_X0Y0_EE4BEG[13]));
 sky130_fd_sc_hd__buf_2 output273 (.A(net273),
    .X(Tile_X0Y0_EE4BEG[14]));
 sky130_fd_sc_hd__buf_8 output274 (.A(net274),
    .X(Tile_X0Y0_EE4BEG[15]));
 sky130_fd_sc_hd__buf_2 output275 (.A(net275),
    .X(Tile_X0Y0_EE4BEG[1]));
 sky130_fd_sc_hd__buf_2 output276 (.A(net276),
    .X(Tile_X0Y0_EE4BEG[2]));
 sky130_fd_sc_hd__buf_2 output277 (.A(net277),
    .X(Tile_X0Y0_EE4BEG[3]));
 sky130_fd_sc_hd__buf_2 output278 (.A(net278),
    .X(Tile_X0Y0_EE4BEG[4]));
 sky130_fd_sc_hd__buf_2 output279 (.A(net279),
    .X(Tile_X0Y0_EE4BEG[5]));
 sky130_fd_sc_hd__buf_2 output280 (.A(net280),
    .X(Tile_X0Y0_EE4BEG[6]));
 sky130_fd_sc_hd__buf_2 output281 (.A(net281),
    .X(Tile_X0Y0_EE4BEG[7]));
 sky130_fd_sc_hd__buf_2 output282 (.A(net282),
    .X(Tile_X0Y0_EE4BEG[8]));
 sky130_fd_sc_hd__buf_2 output283 (.A(net283),
    .X(Tile_X0Y0_EE4BEG[9]));
 sky130_fd_sc_hd__buf_2 output284 (.A(net284),
    .X(Tile_X0Y0_FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output285 (.A(net285),
    .X(Tile_X0Y0_FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output286 (.A(net286),
    .X(Tile_X0Y0_FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output287 (.A(net287),
    .X(Tile_X0Y0_FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output288 (.A(net288),
    .X(Tile_X0Y0_FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .X(Tile_X0Y0_FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output290 (.A(net290),
    .X(Tile_X0Y0_FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output291 (.A(net291),
    .X(Tile_X0Y0_FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output292 (.A(net292),
    .X(Tile_X0Y0_FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output293 (.A(net293),
    .X(Tile_X0Y0_FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output294 (.A(net294),
    .X(Tile_X0Y0_FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output295 (.A(net295),
    .X(Tile_X0Y0_FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output296 (.A(net296),
    .X(Tile_X0Y0_FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output297 (.A(net297),
    .X(Tile_X0Y0_FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output298 (.A(net298),
    .X(Tile_X0Y0_FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output299 (.A(net299),
    .X(Tile_X0Y0_FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output300 (.A(net300),
    .X(Tile_X0Y0_FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output301 (.A(net301),
    .X(Tile_X0Y0_FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output302 (.A(net302),
    .X(Tile_X0Y0_FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output303 (.A(net303),
    .X(Tile_X0Y0_FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output304 (.A(net304),
    .X(Tile_X0Y0_FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output305 (.A(net305),
    .X(Tile_X0Y0_FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output306 (.A(net306),
    .X(Tile_X0Y0_FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output307 (.A(net307),
    .X(Tile_X0Y0_FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output308 (.A(net308),
    .X(Tile_X0Y0_FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output309 (.A(net309),
    .X(Tile_X0Y0_FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output310 (.A(net310),
    .X(Tile_X0Y0_FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output311 (.A(net311),
    .X(Tile_X0Y0_FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output312 (.A(net312),
    .X(Tile_X0Y0_FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output313 (.A(net313),
    .X(Tile_X0Y0_FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output314 (.A(net314),
    .X(Tile_X0Y0_FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output315 (.A(net315),
    .X(Tile_X0Y0_FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output316 (.A(net316),
    .X(Tile_X0Y0_FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output317 (.A(net317),
    .X(Tile_X0Y0_FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output318 (.A(net318),
    .X(Tile_X0Y0_FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output319 (.A(net319),
    .X(Tile_X0Y0_FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output320 (.A(net320),
    .X(Tile_X0Y0_FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output321 (.A(net321),
    .X(Tile_X0Y0_FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output322 (.A(net322),
    .X(Tile_X0Y0_FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output323 (.A(net323),
    .X(Tile_X0Y0_FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output324 (.A(net324),
    .X(Tile_X0Y0_FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output325 (.A(net325),
    .X(Tile_X0Y0_FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output326 (.A(net326),
    .X(Tile_X0Y0_FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output327 (.A(net327),
    .X(Tile_X0Y0_FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output328 (.A(net328),
    .X(Tile_X0Y0_FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output329 (.A(net329),
    .X(Tile_X0Y0_FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output330 (.A(net330),
    .X(Tile_X0Y0_FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output331 (.A(net331),
    .X(Tile_X0Y0_FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output332 (.A(net332),
    .X(Tile_X0Y0_FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output333 (.A(net333),
    .X(Tile_X0Y0_FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output334 (.A(net334),
    .X(Tile_X0Y0_FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output335 (.A(net335),
    .X(Tile_X0Y0_FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_2 output336 (.A(net336),
    .X(Tile_X0Y0_N1BEG[0]));
 sky130_fd_sc_hd__buf_8 output337 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 ),
    .X(Tile_X0Y0_N1BEG[1]));
 sky130_fd_sc_hd__buf_8 output338 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 ),
    .X(Tile_X0Y0_N1BEG[2]));
 sky130_fd_sc_hd__buf_2 output339 (.A(net339),
    .X(Tile_X0Y0_N1BEG[3]));
 sky130_fd_sc_hd__buf_2 output340 (.A(net340),
    .X(Tile_X0Y0_N2BEG[0]));
 sky130_fd_sc_hd__buf_2 output341 (.A(net341),
    .X(Tile_X0Y0_N2BEG[1]));
 sky130_fd_sc_hd__buf_2 output342 (.A(net342),
    .X(Tile_X0Y0_N2BEG[2]));
 sky130_fd_sc_hd__buf_2 output343 (.A(net343),
    .X(Tile_X0Y0_N2BEG[3]));
 sky130_fd_sc_hd__buf_2 output344 (.A(net344),
    .X(Tile_X0Y0_N2BEG[4]));
 sky130_fd_sc_hd__buf_2 output345 (.A(net345),
    .X(Tile_X0Y0_N2BEG[5]));
 sky130_fd_sc_hd__buf_2 output346 (.A(net346),
    .X(Tile_X0Y0_N2BEG[6]));
 sky130_fd_sc_hd__buf_2 output347 (.A(net347),
    .X(Tile_X0Y0_N2BEG[7]));
 sky130_fd_sc_hd__buf_2 output348 (.A(net348),
    .X(Tile_X0Y0_N2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output349 (.A(net349),
    .X(Tile_X0Y0_N2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output350 (.A(net350),
    .X(Tile_X0Y0_N2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output351 (.A(net351),
    .X(Tile_X0Y0_N2BEGb[3]));
 sky130_fd_sc_hd__buf_6 output352 (.A(net352),
    .X(Tile_X0Y0_N2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output353 (.A(net353),
    .X(Tile_X0Y0_N2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output354 (.A(net354),
    .X(Tile_X0Y0_N2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output355 (.A(net355),
    .X(Tile_X0Y0_N2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output356 (.A(net356),
    .X(Tile_X0Y0_N4BEG[0]));
 sky130_fd_sc_hd__buf_2 output357 (.A(net357),
    .X(Tile_X0Y0_N4BEG[10]));
 sky130_fd_sc_hd__buf_2 output358 (.A(net358),
    .X(Tile_X0Y0_N4BEG[11]));
 sky130_fd_sc_hd__buf_2 output359 (.A(net359),
    .X(Tile_X0Y0_N4BEG[12]));
 sky130_fd_sc_hd__buf_2 output360 (.A(net360),
    .X(Tile_X0Y0_N4BEG[13]));
 sky130_fd_sc_hd__buf_2 output361 (.A(net361),
    .X(Tile_X0Y0_N4BEG[14]));
 sky130_fd_sc_hd__buf_2 output362 (.A(net362),
    .X(Tile_X0Y0_N4BEG[15]));
 sky130_fd_sc_hd__buf_2 output363 (.A(net363),
    .X(Tile_X0Y0_N4BEG[1]));
 sky130_fd_sc_hd__buf_2 output364 (.A(net364),
    .X(Tile_X0Y0_N4BEG[2]));
 sky130_fd_sc_hd__buf_2 output365 (.A(net365),
    .X(Tile_X0Y0_N4BEG[3]));
 sky130_fd_sc_hd__buf_2 output366 (.A(net366),
    .X(Tile_X0Y0_N4BEG[4]));
 sky130_fd_sc_hd__buf_2 output367 (.A(net367),
    .X(Tile_X0Y0_N4BEG[5]));
 sky130_fd_sc_hd__buf_2 output368 (.A(net368),
    .X(Tile_X0Y0_N4BEG[6]));
 sky130_fd_sc_hd__buf_2 output369 (.A(net369),
    .X(Tile_X0Y0_N4BEG[7]));
 sky130_fd_sc_hd__buf_2 output370 (.A(net370),
    .X(Tile_X0Y0_N4BEG[8]));
 sky130_fd_sc_hd__buf_2 output371 (.A(net371),
    .X(Tile_X0Y0_N4BEG[9]));
 sky130_fd_sc_hd__buf_2 output372 (.A(net372),
    .X(Tile_X0Y0_NN4BEG[0]));
 sky130_fd_sc_hd__buf_2 output373 (.A(net373),
    .X(Tile_X0Y0_NN4BEG[10]));
 sky130_fd_sc_hd__buf_8 output374 (.A(net374),
    .X(Tile_X0Y0_NN4BEG[11]));
 sky130_fd_sc_hd__buf_6 output375 (.A(net375),
    .X(Tile_X0Y0_NN4BEG[12]));
 sky130_fd_sc_hd__buf_6 output376 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 ),
    .X(Tile_X0Y0_NN4BEG[13]));
 sky130_fd_sc_hd__buf_8 output377 (.A(net377),
    .X(Tile_X0Y0_NN4BEG[14]));
 sky130_fd_sc_hd__buf_6 output378 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 ),
    .X(Tile_X0Y0_NN4BEG[15]));
 sky130_fd_sc_hd__buf_2 output379 (.A(net379),
    .X(Tile_X0Y0_NN4BEG[1]));
 sky130_fd_sc_hd__buf_2 output380 (.A(net380),
    .X(Tile_X0Y0_NN4BEG[2]));
 sky130_fd_sc_hd__buf_2 output381 (.A(net381),
    .X(Tile_X0Y0_NN4BEG[3]));
 sky130_fd_sc_hd__buf_2 output382 (.A(net382),
    .X(Tile_X0Y0_NN4BEG[4]));
 sky130_fd_sc_hd__buf_2 output383 (.A(net383),
    .X(Tile_X0Y0_NN4BEG[5]));
 sky130_fd_sc_hd__buf_2 output384 (.A(net384),
    .X(Tile_X0Y0_NN4BEG[6]));
 sky130_fd_sc_hd__buf_2 output385 (.A(net385),
    .X(Tile_X0Y0_NN4BEG[7]));
 sky130_fd_sc_hd__buf_2 output386 (.A(net386),
    .X(Tile_X0Y0_NN4BEG[8]));
 sky130_fd_sc_hd__buf_4 output387 (.A(net387),
    .X(Tile_X0Y0_NN4BEG[9]));
 sky130_fd_sc_hd__buf_1 output388 (.A(net388),
    .X(Tile_X0Y0_UserCLKo));
 sky130_fd_sc_hd__buf_2 output389 (.A(net389),
    .X(Tile_X0Y0_W1BEG[0]));
 sky130_fd_sc_hd__buf_2 output390 (.A(net390),
    .X(Tile_X0Y0_W1BEG[1]));
 sky130_fd_sc_hd__buf_6 output391 (.A(net391),
    .X(Tile_X0Y0_W1BEG[2]));
 sky130_fd_sc_hd__buf_2 output392 (.A(net392),
    .X(Tile_X0Y0_W1BEG[3]));
 sky130_fd_sc_hd__buf_2 output393 (.A(net393),
    .X(Tile_X0Y0_W2BEG[0]));
 sky130_fd_sc_hd__buf_2 output394 (.A(net394),
    .X(Tile_X0Y0_W2BEG[1]));
 sky130_fd_sc_hd__buf_2 output395 (.A(net395),
    .X(Tile_X0Y0_W2BEG[2]));
 sky130_fd_sc_hd__buf_2 output396 (.A(net396),
    .X(Tile_X0Y0_W2BEG[3]));
 sky130_fd_sc_hd__buf_2 output397 (.A(net397),
    .X(Tile_X0Y0_W2BEG[4]));
 sky130_fd_sc_hd__buf_2 output398 (.A(net398),
    .X(Tile_X0Y0_W2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output399 (.A(net399),
    .X(Tile_X0Y0_W2BEG[6]));
 sky130_fd_sc_hd__buf_2 output400 (.A(net400),
    .X(Tile_X0Y0_W2BEG[7]));
 sky130_fd_sc_hd__buf_2 output401 (.A(net401),
    .X(Tile_X0Y0_W2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output402 (.A(net402),
    .X(Tile_X0Y0_W2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output403 (.A(net403),
    .X(Tile_X0Y0_W2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output404 (.A(net404),
    .X(Tile_X0Y0_W2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output405 (.A(net405),
    .X(Tile_X0Y0_W2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output406 (.A(net406),
    .X(Tile_X0Y0_W2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output407 (.A(net407),
    .X(Tile_X0Y0_W2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output408 (.A(net408),
    .X(Tile_X0Y0_W2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output409 (.A(net409),
    .X(Tile_X0Y0_W6BEG[0]));
 sky130_fd_sc_hd__buf_8 output410 (.A(net410),
    .X(Tile_X0Y0_W6BEG[10]));
 sky130_fd_sc_hd__buf_6 output411 (.A(net411),
    .X(Tile_X0Y0_W6BEG[11]));
 sky130_fd_sc_hd__buf_2 output412 (.A(net412),
    .X(Tile_X0Y0_W6BEG[1]));
 sky130_fd_sc_hd__buf_2 output413 (.A(net413),
    .X(Tile_X0Y0_W6BEG[2]));
 sky130_fd_sc_hd__buf_2 output414 (.A(net414),
    .X(Tile_X0Y0_W6BEG[3]));
 sky130_fd_sc_hd__buf_2 output415 (.A(net415),
    .X(Tile_X0Y0_W6BEG[4]));
 sky130_fd_sc_hd__buf_2 output416 (.A(net416),
    .X(Tile_X0Y0_W6BEG[5]));
 sky130_fd_sc_hd__buf_2 output417 (.A(net417),
    .X(Tile_X0Y0_W6BEG[6]));
 sky130_fd_sc_hd__buf_2 output418 (.A(net418),
    .X(Tile_X0Y0_W6BEG[7]));
 sky130_fd_sc_hd__buf_2 output419 (.A(net419),
    .X(Tile_X0Y0_W6BEG[8]));
 sky130_fd_sc_hd__buf_2 output420 (.A(net420),
    .X(Tile_X0Y0_W6BEG[9]));
 sky130_fd_sc_hd__buf_2 output421 (.A(net421),
    .X(Tile_X0Y0_WW4BEG[0]));
 sky130_fd_sc_hd__buf_2 output422 (.A(net422),
    .X(Tile_X0Y0_WW4BEG[10]));
 sky130_fd_sc_hd__buf_2 output423 (.A(net423),
    .X(Tile_X0Y0_WW4BEG[11]));
 sky130_fd_sc_hd__buf_2 output424 (.A(net424),
    .X(Tile_X0Y0_WW4BEG[12]));
 sky130_fd_sc_hd__buf_8 output425 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 ),
    .X(Tile_X0Y0_WW4BEG[13]));
 sky130_fd_sc_hd__buf_8 output426 (.A(net426),
    .X(Tile_X0Y0_WW4BEG[14]));
 sky130_fd_sc_hd__buf_6 output427 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 ),
    .X(Tile_X0Y0_WW4BEG[15]));
 sky130_fd_sc_hd__buf_2 output428 (.A(net428),
    .X(Tile_X0Y0_WW4BEG[1]));
 sky130_fd_sc_hd__buf_2 output429 (.A(net429),
    .X(Tile_X0Y0_WW4BEG[2]));
 sky130_fd_sc_hd__buf_2 output430 (.A(net430),
    .X(Tile_X0Y0_WW4BEG[3]));
 sky130_fd_sc_hd__buf_2 output431 (.A(net431),
    .X(Tile_X0Y0_WW4BEG[4]));
 sky130_fd_sc_hd__buf_2 output432 (.A(net432),
    .X(Tile_X0Y0_WW4BEG[5]));
 sky130_fd_sc_hd__buf_2 output433 (.A(net433),
    .X(Tile_X0Y0_WW4BEG[6]));
 sky130_fd_sc_hd__buf_2 output434 (.A(net434),
    .X(Tile_X0Y0_WW4BEG[7]));
 sky130_fd_sc_hd__buf_2 output435 (.A(net435),
    .X(Tile_X0Y0_WW4BEG[8]));
 sky130_fd_sc_hd__buf_2 output436 (.A(net436),
    .X(Tile_X0Y0_WW4BEG[9]));
 sky130_fd_sc_hd__buf_2 output437 (.A(net437),
    .X(Tile_X0Y1_E1BEG[0]));
 sky130_fd_sc_hd__buf_6 output438 (.A(net438),
    .X(Tile_X0Y1_E1BEG[1]));
 sky130_fd_sc_hd__buf_2 output439 (.A(net439),
    .X(Tile_X0Y1_E1BEG[2]));
 sky130_fd_sc_hd__buf_2 output440 (.A(net440),
    .X(Tile_X0Y1_E1BEG[3]));
 sky130_fd_sc_hd__buf_2 output441 (.A(net441),
    .X(Tile_X0Y1_E2BEG[0]));
 sky130_fd_sc_hd__buf_2 output442 (.A(net442),
    .X(Tile_X0Y1_E2BEG[1]));
 sky130_fd_sc_hd__buf_2 output443 (.A(net443),
    .X(Tile_X0Y1_E2BEG[2]));
 sky130_fd_sc_hd__buf_2 output444 (.A(net444),
    .X(Tile_X0Y1_E2BEG[3]));
 sky130_fd_sc_hd__buf_2 output445 (.A(net445),
    .X(Tile_X0Y1_E2BEG[4]));
 sky130_fd_sc_hd__buf_2 output446 (.A(net446),
    .X(Tile_X0Y1_E2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output447 (.A(net447),
    .X(Tile_X0Y1_E2BEG[6]));
 sky130_fd_sc_hd__buf_6 output448 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 ),
    .X(Tile_X0Y1_E2BEG[7]));
 sky130_fd_sc_hd__buf_2 output449 (.A(net449),
    .X(Tile_X0Y1_E2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output450 (.A(net450),
    .X(Tile_X0Y1_E2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output451 (.A(net451),
    .X(Tile_X0Y1_E2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output452 (.A(net452),
    .X(Tile_X0Y1_E2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output453 (.A(net453),
    .X(Tile_X0Y1_E2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output454 (.A(net454),
    .X(Tile_X0Y1_E2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output455 (.A(net455),
    .X(Tile_X0Y1_E2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output456 (.A(net456),
    .X(Tile_X0Y1_E2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output457 (.A(net457),
    .X(Tile_X0Y1_E6BEG[0]));
 sky130_fd_sc_hd__buf_2 output458 (.A(net458),
    .X(Tile_X0Y1_E6BEG[10]));
 sky130_fd_sc_hd__buf_6 output459 (.A(net459),
    .X(Tile_X0Y1_E6BEG[11]));
 sky130_fd_sc_hd__buf_2 output460 (.A(net460),
    .X(Tile_X0Y1_E6BEG[1]));
 sky130_fd_sc_hd__buf_2 output461 (.A(net461),
    .X(Tile_X0Y1_E6BEG[2]));
 sky130_fd_sc_hd__buf_2 output462 (.A(net462),
    .X(Tile_X0Y1_E6BEG[3]));
 sky130_fd_sc_hd__buf_2 output463 (.A(net463),
    .X(Tile_X0Y1_E6BEG[4]));
 sky130_fd_sc_hd__buf_2 output464 (.A(net464),
    .X(Tile_X0Y1_E6BEG[5]));
 sky130_fd_sc_hd__buf_2 output465 (.A(net465),
    .X(Tile_X0Y1_E6BEG[6]));
 sky130_fd_sc_hd__buf_2 output466 (.A(net466),
    .X(Tile_X0Y1_E6BEG[7]));
 sky130_fd_sc_hd__buf_2 output467 (.A(net467),
    .X(Tile_X0Y1_E6BEG[8]));
 sky130_fd_sc_hd__buf_2 output468 (.A(net468),
    .X(Tile_X0Y1_E6BEG[9]));
 sky130_fd_sc_hd__buf_2 output469 (.A(net469),
    .X(Tile_X0Y1_EE4BEG[0]));
 sky130_fd_sc_hd__buf_2 output470 (.A(net470),
    .X(Tile_X0Y1_EE4BEG[10]));
 sky130_fd_sc_hd__buf_2 output471 (.A(net471),
    .X(Tile_X0Y1_EE4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output472 (.A(net472),
    .X(Tile_X0Y1_EE4BEG[12]));
 sky130_fd_sc_hd__buf_4 output473 (.A(net473),
    .X(Tile_X0Y1_EE4BEG[13]));
 sky130_fd_sc_hd__buf_2 output474 (.A(net474),
    .X(Tile_X0Y1_EE4BEG[14]));
 sky130_fd_sc_hd__buf_8 output475 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 ),
    .X(Tile_X0Y1_EE4BEG[15]));
 sky130_fd_sc_hd__buf_2 output476 (.A(net476),
    .X(Tile_X0Y1_EE4BEG[1]));
 sky130_fd_sc_hd__buf_2 output477 (.A(net477),
    .X(Tile_X0Y1_EE4BEG[2]));
 sky130_fd_sc_hd__buf_2 output478 (.A(net478),
    .X(Tile_X0Y1_EE4BEG[3]));
 sky130_fd_sc_hd__buf_2 output479 (.A(net479),
    .X(Tile_X0Y1_EE4BEG[4]));
 sky130_fd_sc_hd__buf_2 output480 (.A(net480),
    .X(Tile_X0Y1_EE4BEG[5]));
 sky130_fd_sc_hd__buf_2 output481 (.A(net481),
    .X(Tile_X0Y1_EE4BEG[6]));
 sky130_fd_sc_hd__buf_2 output482 (.A(net482),
    .X(Tile_X0Y1_EE4BEG[7]));
 sky130_fd_sc_hd__buf_2 output483 (.A(net483),
    .X(Tile_X0Y1_EE4BEG[8]));
 sky130_fd_sc_hd__buf_2 output484 (.A(net484),
    .X(Tile_X0Y1_EE4BEG[9]));
 sky130_fd_sc_hd__buf_2 output485 (.A(net485),
    .X(Tile_X0Y1_FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output486 (.A(net486),
    .X(Tile_X0Y1_FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output487 (.A(net487),
    .X(Tile_X0Y1_FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output488 (.A(net488),
    .X(Tile_X0Y1_FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output489 (.A(net489),
    .X(Tile_X0Y1_FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output490 (.A(net490),
    .X(Tile_X0Y1_FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output491 (.A(net491),
    .X(Tile_X0Y1_FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output492 (.A(net492),
    .X(Tile_X0Y1_FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output493 (.A(net493),
    .X(Tile_X0Y1_FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output494 (.A(net494),
    .X(Tile_X0Y1_FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output495 (.A(net495),
    .X(Tile_X0Y1_FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output496 (.A(net496),
    .X(Tile_X0Y1_FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output497 (.A(net497),
    .X(Tile_X0Y1_FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output498 (.A(net498),
    .X(Tile_X0Y1_FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output499 (.A(net499),
    .X(Tile_X0Y1_FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output500 (.A(net500),
    .X(Tile_X0Y1_FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output501 (.A(net501),
    .X(Tile_X0Y1_FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output502 (.A(net502),
    .X(Tile_X0Y1_FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output503 (.A(net503),
    .X(Tile_X0Y1_FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output504 (.A(net504),
    .X(Tile_X0Y1_FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output505 (.A(net505),
    .X(Tile_X0Y1_FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output506 (.A(net506),
    .X(Tile_X0Y1_FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output507 (.A(net507),
    .X(Tile_X0Y1_FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output508 (.A(net508),
    .X(Tile_X0Y1_FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output509 (.A(net509),
    .X(Tile_X0Y1_FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output510 (.A(net510),
    .X(Tile_X0Y1_FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output511 (.A(net511),
    .X(Tile_X0Y1_FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output512 (.A(net512),
    .X(Tile_X0Y1_FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output513 (.A(net513),
    .X(Tile_X0Y1_FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output514 (.A(net514),
    .X(Tile_X0Y1_FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output515 (.A(net515),
    .X(Tile_X0Y1_FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output516 (.A(net516),
    .X(Tile_X0Y1_FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output517 (.A(net517),
    .X(Tile_X0Y1_S1BEG[0]));
 sky130_fd_sc_hd__buf_8 output518 (.A(net518),
    .X(Tile_X0Y1_S1BEG[1]));
 sky130_fd_sc_hd__buf_2 output519 (.A(net519),
    .X(Tile_X0Y1_S1BEG[2]));
 sky130_fd_sc_hd__buf_2 output520 (.A(net520),
    .X(Tile_X0Y1_S1BEG[3]));
 sky130_fd_sc_hd__buf_2 output521 (.A(net521),
    .X(Tile_X0Y1_S2BEG[0]));
 sky130_fd_sc_hd__buf_2 output522 (.A(net522),
    .X(Tile_X0Y1_S2BEG[1]));
 sky130_fd_sc_hd__buf_2 output523 (.A(net523),
    .X(Tile_X0Y1_S2BEG[2]));
 sky130_fd_sc_hd__buf_2 output524 (.A(net524),
    .X(Tile_X0Y1_S2BEG[3]));
 sky130_fd_sc_hd__buf_4 output525 (.A(net525),
    .X(Tile_X0Y1_S2BEG[4]));
 sky130_fd_sc_hd__buf_6 output526 (.A(net526),
    .X(Tile_X0Y1_S2BEG[5]));
 sky130_fd_sc_hd__buf_2 output527 (.A(net527),
    .X(Tile_X0Y1_S2BEG[6]));
 sky130_fd_sc_hd__buf_2 output528 (.A(net528),
    .X(Tile_X0Y1_S2BEG[7]));
 sky130_fd_sc_hd__buf_2 output529 (.A(net529),
    .X(Tile_X0Y1_S2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output530 (.A(net530),
    .X(Tile_X0Y1_S2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output531 (.A(net531),
    .X(Tile_X0Y1_S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output532 (.A(net532),
    .X(Tile_X0Y1_S2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output533 (.A(net533),
    .X(Tile_X0Y1_S2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output534 (.A(net534),
    .X(Tile_X0Y1_S2BEGb[5]));
 sky130_fd_sc_hd__buf_8 output535 (.A(net535),
    .X(Tile_X0Y1_S2BEGb[6]));
 sky130_fd_sc_hd__buf_8 output536 (.A(net536),
    .X(Tile_X0Y1_S2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output537 (.A(net537),
    .X(Tile_X0Y1_S4BEG[0]));
 sky130_fd_sc_hd__buf_2 output538 (.A(net538),
    .X(Tile_X0Y1_S4BEG[10]));
 sky130_fd_sc_hd__buf_2 output539 (.A(net539),
    .X(Tile_X0Y1_S4BEG[11]));
 sky130_fd_sc_hd__buf_2 output540 (.A(net540),
    .X(Tile_X0Y1_S4BEG[12]));
 sky130_fd_sc_hd__buf_2 output541 (.A(net541),
    .X(Tile_X0Y1_S4BEG[13]));
 sky130_fd_sc_hd__buf_2 output542 (.A(net542),
    .X(Tile_X0Y1_S4BEG[14]));
 sky130_fd_sc_hd__buf_2 output543 (.A(net543),
    .X(Tile_X0Y1_S4BEG[15]));
 sky130_fd_sc_hd__buf_2 output544 (.A(net544),
    .X(Tile_X0Y1_S4BEG[1]));
 sky130_fd_sc_hd__buf_2 output545 (.A(net545),
    .X(Tile_X0Y1_S4BEG[2]));
 sky130_fd_sc_hd__buf_2 output546 (.A(net546),
    .X(Tile_X0Y1_S4BEG[3]));
 sky130_fd_sc_hd__buf_2 output547 (.A(net547),
    .X(Tile_X0Y1_S4BEG[4]));
 sky130_fd_sc_hd__buf_2 output548 (.A(net548),
    .X(Tile_X0Y1_S4BEG[5]));
 sky130_fd_sc_hd__buf_2 output549 (.A(net549),
    .X(Tile_X0Y1_S4BEG[6]));
 sky130_fd_sc_hd__buf_2 output550 (.A(net550),
    .X(Tile_X0Y1_S4BEG[7]));
 sky130_fd_sc_hd__buf_2 output551 (.A(net551),
    .X(Tile_X0Y1_S4BEG[8]));
 sky130_fd_sc_hd__buf_2 output552 (.A(net552),
    .X(Tile_X0Y1_S4BEG[9]));
 sky130_fd_sc_hd__buf_2 output553 (.A(net553),
    .X(Tile_X0Y1_SS4BEG[0]));
 sky130_fd_sc_hd__buf_2 output554 (.A(net554),
    .X(Tile_X0Y1_SS4BEG[10]));
 sky130_fd_sc_hd__buf_8 output555 (.A(net555),
    .X(Tile_X0Y1_SS4BEG[11]));
 sky130_fd_sc_hd__buf_2 output556 (.A(net556),
    .X(Tile_X0Y1_SS4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output557 (.A(net557),
    .X(Tile_X0Y1_SS4BEG[13]));
 sky130_fd_sc_hd__buf_2 output558 (.A(net558),
    .X(Tile_X0Y1_SS4BEG[14]));
 sky130_fd_sc_hd__buf_6 output559 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 ),
    .X(Tile_X0Y1_SS4BEG[15]));
 sky130_fd_sc_hd__buf_2 output560 (.A(net560),
    .X(Tile_X0Y1_SS4BEG[1]));
 sky130_fd_sc_hd__buf_2 output561 (.A(net561),
    .X(Tile_X0Y1_SS4BEG[2]));
 sky130_fd_sc_hd__buf_2 output562 (.A(net562),
    .X(Tile_X0Y1_SS4BEG[3]));
 sky130_fd_sc_hd__buf_2 output563 (.A(net563),
    .X(Tile_X0Y1_SS4BEG[4]));
 sky130_fd_sc_hd__buf_2 output564 (.A(net564),
    .X(Tile_X0Y1_SS4BEG[5]));
 sky130_fd_sc_hd__buf_2 output565 (.A(net565),
    .X(Tile_X0Y1_SS4BEG[6]));
 sky130_fd_sc_hd__buf_2 output566 (.A(net566),
    .X(Tile_X0Y1_SS4BEG[7]));
 sky130_fd_sc_hd__buf_2 output567 (.A(net567),
    .X(Tile_X0Y1_SS4BEG[8]));
 sky130_fd_sc_hd__buf_8 output568 (.A(net568),
    .X(Tile_X0Y1_SS4BEG[9]));
 sky130_fd_sc_hd__buf_2 output569 (.A(net569),
    .X(Tile_X0Y1_W1BEG[0]));
 sky130_fd_sc_hd__buf_8 output570 (.A(net570),
    .X(Tile_X0Y1_W1BEG[1]));
 sky130_fd_sc_hd__buf_2 output571 (.A(net571),
    .X(Tile_X0Y1_W1BEG[2]));
 sky130_fd_sc_hd__buf_2 output572 (.A(net572),
    .X(Tile_X0Y1_W1BEG[3]));
 sky130_fd_sc_hd__buf_2 output573 (.A(net573),
    .X(Tile_X0Y1_W2BEG[0]));
 sky130_fd_sc_hd__buf_2 output574 (.A(net574),
    .X(Tile_X0Y1_W2BEG[1]));
 sky130_fd_sc_hd__buf_2 output575 (.A(net575),
    .X(Tile_X0Y1_W2BEG[2]));
 sky130_fd_sc_hd__buf_2 output576 (.A(net576),
    .X(Tile_X0Y1_W2BEG[3]));
 sky130_fd_sc_hd__buf_2 output577 (.A(net577),
    .X(Tile_X0Y1_W2BEG[4]));
 sky130_fd_sc_hd__buf_8 output578 (.A(net578),
    .X(Tile_X0Y1_W2BEG[5]));
 sky130_fd_sc_hd__buf_8 output579 (.A(net579),
    .X(Tile_X0Y1_W2BEG[6]));
 sky130_fd_sc_hd__buf_2 output580 (.A(net580),
    .X(Tile_X0Y1_W2BEG[7]));
 sky130_fd_sc_hd__buf_2 output581 (.A(net581),
    .X(Tile_X0Y1_W2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output582 (.A(net582),
    .X(Tile_X0Y1_W2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output583 (.A(net583),
    .X(Tile_X0Y1_W2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output584 (.A(net584),
    .X(Tile_X0Y1_W2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output585 (.A(net585),
    .X(Tile_X0Y1_W2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output586 (.A(net586),
    .X(Tile_X0Y1_W2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output587 (.A(net587),
    .X(Tile_X0Y1_W2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output588 (.A(net588),
    .X(Tile_X0Y1_W2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output589 (.A(net589),
    .X(Tile_X0Y1_W6BEG[0]));
 sky130_fd_sc_hd__buf_2 output590 (.A(net590),
    .X(Tile_X0Y1_W6BEG[10]));
 sky130_fd_sc_hd__buf_4 output591 (.A(net591),
    .X(Tile_X0Y1_W6BEG[11]));
 sky130_fd_sc_hd__buf_2 output592 (.A(net592),
    .X(Tile_X0Y1_W6BEG[1]));
 sky130_fd_sc_hd__buf_2 output593 (.A(net593),
    .X(Tile_X0Y1_W6BEG[2]));
 sky130_fd_sc_hd__buf_2 output594 (.A(net594),
    .X(Tile_X0Y1_W6BEG[3]));
 sky130_fd_sc_hd__buf_2 output595 (.A(net595),
    .X(Tile_X0Y1_W6BEG[4]));
 sky130_fd_sc_hd__buf_2 output596 (.A(net596),
    .X(Tile_X0Y1_W6BEG[5]));
 sky130_fd_sc_hd__buf_2 output597 (.A(net597),
    .X(Tile_X0Y1_W6BEG[6]));
 sky130_fd_sc_hd__buf_2 output598 (.A(net598),
    .X(Tile_X0Y1_W6BEG[7]));
 sky130_fd_sc_hd__buf_2 output599 (.A(net599),
    .X(Tile_X0Y1_W6BEG[8]));
 sky130_fd_sc_hd__buf_2 output600 (.A(net600),
    .X(Tile_X0Y1_W6BEG[9]));
 sky130_fd_sc_hd__buf_2 output601 (.A(net601),
    .X(Tile_X0Y1_WW4BEG[0]));
 sky130_fd_sc_hd__buf_2 output602 (.A(net602),
    .X(Tile_X0Y1_WW4BEG[10]));
 sky130_fd_sc_hd__buf_2 output603 (.A(net603),
    .X(Tile_X0Y1_WW4BEG[11]));
 sky130_fd_sc_hd__buf_6 output604 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 ),
    .X(Tile_X0Y1_WW4BEG[12]));
 sky130_fd_sc_hd__buf_4 output605 (.A(net605),
    .X(Tile_X0Y1_WW4BEG[13]));
 sky130_fd_sc_hd__buf_2 output606 (.A(net606),
    .X(Tile_X0Y1_WW4BEG[14]));
 sky130_fd_sc_hd__buf_6 output607 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 ),
    .X(Tile_X0Y1_WW4BEG[15]));
 sky130_fd_sc_hd__buf_2 output608 (.A(net608),
    .X(Tile_X0Y1_WW4BEG[1]));
 sky130_fd_sc_hd__buf_2 output609 (.A(net609),
    .X(Tile_X0Y1_WW4BEG[2]));
 sky130_fd_sc_hd__buf_2 output610 (.A(net610),
    .X(Tile_X0Y1_WW4BEG[3]));
 sky130_fd_sc_hd__buf_2 output611 (.A(net611),
    .X(Tile_X0Y1_WW4BEG[4]));
 sky130_fd_sc_hd__buf_2 output612 (.A(net612),
    .X(Tile_X0Y1_WW4BEG[5]));
 sky130_fd_sc_hd__buf_2 output613 (.A(net613),
    .X(Tile_X0Y1_WW4BEG[6]));
 sky130_fd_sc_hd__buf_2 output614 (.A(net614),
    .X(Tile_X0Y1_WW4BEG[7]));
 sky130_fd_sc_hd__buf_2 output615 (.A(net615),
    .X(Tile_X0Y1_WW4BEG[8]));
 sky130_fd_sc_hd__buf_2 output616 (.A(net616),
    .X(Tile_X0Y1_WW4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 max_cap617 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_regs_0_Tile_X0Y1_UserCLK (.A(Tile_X0Y1_UserCLK),
    .X(Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_Tile_X0Y1_UserCLK (.A(Tile_X0Y1_UserCLK),
    .X(clknet_0_Tile_X0Y1_UserCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_Tile_X0Y1_UserCLK (.A(clknet_0_Tile_X0Y1_UserCLK),
    .X(clknet_1_0__leaf_Tile_X0Y1_UserCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_Tile_X0Y1_UserCLK_regs (.A(Tile_X0Y1_UserCLK_regs),
    .X(clknet_0_Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_Tile_X0Y1_UserCLK_regs (.A(clknet_0_Tile_X0Y1_UserCLK_regs),
    .X(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_Tile_X0Y1_UserCLK_regs (.A(clknet_0_Tile_X0Y1_UserCLK_regs),
    .X(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_Tile_X0Y1_UserCLK_regs (.A(clknet_0_Tile_X0Y1_UserCLK_regs),
    .X(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_Tile_X0Y1_UserCLK_regs (.A(clknet_0_Tile_X0Y1_UserCLK_regs),
    .X(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__inv_8 clkload0 (.A(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__clkinv_4 clkload1 (.A(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload2 (.A(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__o31ai_4 clone1 (.A1(net1060),
    .A2(_0529_),
    .A3(_0574_),
    .B1(_0575_),
    .Y(net618));
 sky130_fd_sc_hd__o22a_4 clone2 (.A1(net636),
    .A2(_0336_),
    .B1(_0339_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q ),
    .X(net619));
 sky130_fd_sc_hd__o21ai_4 clone3 (.A1(\Tile_X0Y1_DSP_bot.A0 ),
    .A2(net1059),
    .B1(_0927_),
    .Y(net620));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(_0359_),
    .X(net621));
 sky130_fd_sc_hd__o21ai_4 clone5 (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X ),
    .A2(net1061),
    .B1(_0761_),
    .Y(net622));
 sky130_fd_sc_hd__a22o_1 clone9 (.A1(net628),
    .A2(net821),
    .B1(net627),
    .B2(net650),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net667),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(_0216_),
    .X(net628));
 sky130_fd_sc_hd__buf_6 rebuffer12 (.A(_0343_),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net629),
    .X(net630));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer14 (.A(net630),
    .X(net631));
 sky130_fd_sc_hd__buf_6 rebuffer15 (.A(_1472_),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net632),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net633),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_2 rebuffer18 (.A(_0258_),
    .X(net635));
 sky130_fd_sc_hd__buf_6 rebuffer19 (.A(_0334_),
    .X(net636));
 sky130_fd_sc_hd__mux2_4 clone20 (.A0(_1565_),
    .A1(net817),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q ),
    .X(net637));
 sky130_fd_sc_hd__buf_6 rebuffer21 (.A(net912),
    .X(net638));
 sky130_fd_sc_hd__buf_6 rebuffer22 (.A(net820),
    .X(net639));
 sky130_fd_sc_hd__buf_6 rebuffer23 (.A(_0342_),
    .X(net640));
 sky130_fd_sc_hd__buf_8 clone24 (.A(net642),
    .X(net641));
 sky130_fd_sc_hd__buf_6 rebuffer25 (.A(net911),
    .X(net642));
 sky130_fd_sc_hd__buf_6 rebuffer30 (.A(_1537_),
    .X(net647));
 sky130_fd_sc_hd__buf_6 rebuffer31 (.A(_1537_),
    .X(net648));
 sky130_fd_sc_hd__clkbuf_2 rebuffer32 (.A(net648),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(_0238_),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(_0258_),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .X(net654));
 sky130_fd_sc_hd__buf_6 clone38 (.A(net908),
    .X(net655));
 sky130_fd_sc_hd__buf_8 clone39 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .X(net656));
 sky130_fd_sc_hd__clkbuf_2 rebuffer44 (.A(_0268_),
    .X(net661));
 sky130_fd_sc_hd__clkbuf_2 rebuffer45 (.A(_0268_),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer46 (.A(_0446_),
    .X(net663));
 sky130_fd_sc_hd__buf_8 clone47 (.A(net979),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer48 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ),
    .X(net665));
 sky130_fd_sc_hd__clkbuf_1 clone49 (.A(_1422_),
    .X(net666));
 sky130_fd_sc_hd__buf_6 rebuffer50 (.A(net826),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer51 (.A(_0225_),
    .X(net668));
 sky130_fd_sc_hd__buf_8 clone52 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer53 (.A(_0439_),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer59 (.A(net765),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer148 (.A(net766),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer149 (.A(net767),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer150 (.A(net768),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer151 (.A(net769),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer152 (.A(net770),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer153 (.A(net771),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer154 (.A(net772),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer155 (.A(net773),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer156 (.A(net774),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer157 (.A(net775),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer158 (.A(net776),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer159 (.A(net777),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer160 (.A(net778),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer161 (.A(net779),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer162 (.A(net780),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer163 (.A(net781),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer164 (.A(net782),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer165 (.A(net783),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer166 (.A(net784),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer167 (.A(net785),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer168 (.A(net786),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer169 (.A(net787),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer170 (.A(net788),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer171 (.A(net789),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer172 (.A(net790),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer173 (.A(net791),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer174 (.A(net792),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer175 (.A(net793),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer176 (.A(net794),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer177 (.A(net795),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer178 (.A(net796),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer179 (.A(net797),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer180 (.A(net798),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer181 (.A(net799),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer182 (.A(net800),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer183 (.A(net801),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer184 (.A(net802),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer185 (.A(net803),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer186 (.A(net804),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer187 (.A(net805),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer188 (.A(net806),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer189 (.A(net807),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer190 (.A(net808),
    .X(net807));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer191 (.A(net810),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer192 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ),
    .X(net809));
 sky130_fd_sc_hd__buf_1 rebuffer193 (.A(\Tile_X0Y1_DSP_bot.C1 ),
    .X(net810));
 sky130_fd_sc_hd__buf_6 clone194 (.A(net926),
    .X(net811));
 sky130_fd_sc_hd__buf_8 clone195 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .X(net812));
 sky130_fd_sc_hd__mux4_2 clone196 (.A0(net993),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ),
    .A2(net816),
    .A3(net814),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q ),
    .X(net813));
 sky130_fd_sc_hd__buf_6 rebuffer197 (.A(_0405_),
    .X(net814));
 sky130_fd_sc_hd__buf_6 clone198 (.A(net1020),
    .X(net815));
 sky130_fd_sc_hd__buf_6 rebuffer199 (.A(_0413_),
    .X(net816));
 sky130_fd_sc_hd__buf_8 rebuffer200 (.A(net919),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer201 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ),
    .X(net818));
 sky130_fd_sc_hd__buf_6 rebuffer202 (.A(_0237_),
    .X(net819));
 sky130_fd_sc_hd__clkbuf_2 rebuffer203 (.A(_0254_),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer204 (.A(_0217_),
    .X(net821));
 sky130_fd_sc_hd__buf_8 clone205 (.A(net1058),
    .X(net822));
 sky130_fd_sc_hd__buf_8 clone206 (.A(net1039),
    .X(net823));
 sky130_fd_sc_hd__buf_6 clone207 (.A(net1027),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_2 rebuffer208 (.A(net835),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer209 (.A(_0229_),
    .X(net826));
 sky130_fd_sc_hd__buf_6 clone211 (.A(net1049),
    .X(net828));
 sky130_fd_sc_hd__buf_8 rebuffer212 (.A(_1125_),
    .X(net829));
 sky130_fd_sc_hd__clkbuf_1 clone213 (.A(net999),
    .X(net830));
 sky130_fd_sc_hd__buf_6 clone214 (.A(net1001),
    .X(net831));
 sky130_fd_sc_hd__buf_12 rebuffer215 (.A(_1029_),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer216 (.A(_0257_),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer217 (.A(_0254_),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_2 rebuffer218 (.A(net836),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_2 rebuffer219 (.A(net837),
    .X(net836));
 sky130_fd_sc_hd__clkbuf_2 rebuffer220 (.A(net838),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_2 rebuffer221 (.A(net839),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_2 rebuffer222 (.A(net840),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_2 rebuffer223 (.A(net841),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_2 rebuffer224 (.A(net842),
    .X(net841));
 sky130_fd_sc_hd__clkbuf_2 rebuffer225 (.A(net843),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_2 rebuffer226 (.A(net844),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_2 rebuffer227 (.A(net845),
    .X(net844));
 sky130_fd_sc_hd__clkbuf_2 rebuffer228 (.A(net846),
    .X(net845));
 sky130_fd_sc_hd__clkbuf_2 rebuffer229 (.A(net847),
    .X(net846));
 sky130_fd_sc_hd__clkbuf_2 rebuffer230 (.A(net848),
    .X(net847));
 sky130_fd_sc_hd__clkbuf_2 rebuffer231 (.A(net849),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_2 rebuffer232 (.A(net850),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_2 rebuffer233 (.A(net851),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_2 rebuffer234 (.A(net852),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_2 rebuffer235 (.A(net853),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_2 rebuffer236 (.A(net854),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_2 rebuffer237 (.A(net855),
    .X(net854));
 sky130_fd_sc_hd__clkbuf_2 rebuffer238 (.A(net856),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_2 rebuffer239 (.A(net857),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_2 rebuffer240 (.A(net858),
    .X(net857));
 sky130_fd_sc_hd__clkbuf_2 rebuffer241 (.A(net859),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_2 rebuffer242 (.A(net860),
    .X(net859));
 sky130_fd_sc_hd__clkbuf_2 rebuffer243 (.A(net861),
    .X(net860));
 sky130_fd_sc_hd__clkbuf_2 rebuffer244 (.A(net862),
    .X(net861));
 sky130_fd_sc_hd__clkbuf_2 rebuffer245 (.A(net863),
    .X(net862));
 sky130_fd_sc_hd__clkbuf_2 rebuffer246 (.A(_0243_),
    .X(net863));
 sky130_fd_sc_hd__clkbuf_1 clone247 (.A(net996),
    .X(net864));
 sky130_fd_sc_hd__buf_6 clone248 (.A(net986),
    .X(net865));
 sky130_fd_sc_hd__buf_6 clone250 (.A(net1041),
    .X(net867));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer251 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .X(net868));
 sky130_fd_sc_hd__buf_6 clone252 (.A(net972),
    .X(net869));
 sky130_fd_sc_hd__buf_4 rebuffer259 (.A(net877),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer260 (.A(net878),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer261 (.A(net879),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer262 (.A(net880),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer263 (.A(net881),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer264 (.A(net882),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer265 (.A(net883),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer266 (.A(net884),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer267 (.A(net885),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer268 (.A(net886),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer269 (.A(net887),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer270 (.A(net888),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer271 (.A(net889),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer272 (.A(net890),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer273 (.A(net891),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer274 (.A(net892),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer275 (.A(net893),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer276 (.A(net894),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer277 (.A(net895),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer278 (.A(net896),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer279 (.A(net897),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer280 (.A(net898),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer281 (.A(net899),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer282 (.A(net900),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer283 (.A(net901),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer284 (.A(net902),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer285 (.A(net903),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer286 (.A(net904),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer287 (.A(net905),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer288 (.A(net906),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer289 (.A(net907),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer290 (.A(net874),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer291 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .X(net908));
 sky130_fd_sc_hd__buf_6 rebuffer292 (.A(net927),
    .X(net909));
 sky130_fd_sc_hd__clkbuf_2 rebuffer295 (.A(net911),
    .X(net912));
 sky130_fd_sc_hd__clkbuf_1 rebuffer296 (.A(net914),
    .X(net913));
 sky130_fd_sc_hd__clkbuf_1 rebuffer298 (.A(_0340_),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer301 (.A(_0413_),
    .X(net918));
 sky130_fd_sc_hd__buf_6 rebuffer303 (.A(net813),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer304 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer305 (.A(net976),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer306 (.A(net922),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer307 (.A(net976),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer308 (.A(net975),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer309 (.A(net925),
    .X(net926));
 sky130_fd_sc_hd__clkbuf_2 rebuffer310 (.A(net946),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_2 rebuffer330 (.A(net948),
    .X(net947));
 sky130_fd_sc_hd__clkbuf_2 rebuffer331 (.A(net949),
    .X(net948));
 sky130_fd_sc_hd__clkbuf_2 rebuffer332 (.A(net950),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_2 rebuffer333 (.A(net951),
    .X(net950));
 sky130_fd_sc_hd__clkbuf_2 rebuffer334 (.A(net952),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_2 rebuffer335 (.A(net953),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_2 rebuffer336 (.A(net954),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_2 rebuffer337 (.A(net955),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_2 rebuffer338 (.A(net956),
    .X(net955));
 sky130_fd_sc_hd__clkbuf_2 rebuffer339 (.A(net957),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_2 rebuffer340 (.A(net958),
    .X(net957));
 sky130_fd_sc_hd__clkbuf_2 rebuffer341 (.A(net959),
    .X(net958));
 sky130_fd_sc_hd__clkbuf_2 rebuffer342 (.A(net1276),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_2 rebuffer360 (.A(net1277),
    .X(net1276));
 sky130_fd_sc_hd__clkbuf_2 rebuffer361 (.A(net1278),
    .X(net1277));
 sky130_fd_sc_hd__clkbuf_2 rebuffer362 (.A(net1279),
    .X(net1278));
 sky130_fd_sc_hd__clkbuf_2 rebuffer363 (.A(net1280),
    .X(net1279));
 sky130_fd_sc_hd__clkbuf_2 rebuffer364 (.A(net1281),
    .X(net1280));
 sky130_fd_sc_hd__clkbuf_2 rebuffer365 (.A(net1282),
    .X(net1281));
 sky130_fd_sc_hd__clkbuf_2 rebuffer366 (.A(net1283),
    .X(net1282));
 sky130_fd_sc_hd__clkbuf_2 rebuffer367 (.A(net1284),
    .X(net1283));
 sky130_fd_sc_hd__clkbuf_2 rebuffer368 (.A(net1285),
    .X(net1284));
 sky130_fd_sc_hd__clkbuf_2 rebuffer369 (.A(net1286),
    .X(net1285));
 sky130_fd_sc_hd__clkbuf_2 rebuffer370 (.A(net1287),
    .X(net1286));
 sky130_fd_sc_hd__clkbuf_2 rebuffer371 (.A(net1288),
    .X(net1287));
 sky130_fd_sc_hd__clkbuf_2 rebuffer372 (.A(net1289),
    .X(net1288));
 sky130_fd_sc_hd__clkbuf_2 rebuffer373 (.A(net1290),
    .X(net1289));
 sky130_fd_sc_hd__clkbuf_2 rebuffer374 (.A(net1291),
    .X(net1290));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer375 (.A(net973),
    .X(net1291));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(Tile_X0Y0_E6END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(Tile_X0Y0_E6END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(Tile_X0Y0_E6END[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(Tile_X0Y0_E6END[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(Tile_X0Y0_E6END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(Tile_X0Y0_E6END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(Tile_X0Y0_E6END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(Tile_X0Y0_E6END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(Tile_X0Y0_E6END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(Tile_X0Y0_EE4END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(Tile_X0Y0_EE4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(Tile_X0Y0_EE4END[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(Tile_X0Y0_EE4END[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(Tile_X0Y0_EE4END[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(Tile_X0Y0_EE4END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(Tile_X0Y0_EE4END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(Tile_X0Y0_EE4END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(Tile_X0Y0_EE4END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(Tile_X0Y0_EE4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(Tile_X0Y0_EE4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(Tile_X0Y0_FrameData[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(Tile_X0Y0_FrameData[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(Tile_X0Y0_S4END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(Tile_X0Y0_S4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(Tile_X0Y0_S4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(Tile_X0Y0_S4END[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(Tile_X0Y0_S4END[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(Tile_X0Y0_S4END[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(Tile_X0Y0_S4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(Tile_X0Y0_S4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(Tile_X0Y0_S4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(Tile_X0Y0_W2MID[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(Tile_X0Y0_WW4END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(Tile_X0Y0_WW4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(\Tile_X0Y1_DSP_bot.A2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(\Tile_X0Y1_DSP_bot.A2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(Tile_X0Y1_E6END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(Tile_X0Y1_E6END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(Tile_X0Y1_E6END[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(Tile_X0Y1_E6END[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(Tile_X0Y1_E6END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(Tile_X0Y1_E6END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(Tile_X0Y1_E6END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(Tile_X0Y1_E6END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(Tile_X0Y1_E6END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(Tile_X0Y1_E6END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(Tile_X0Y1_EE4END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(Tile_X0Y1_EE4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(Tile_X0Y1_EE4END[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(Tile_X0Y1_EE4END[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(Tile_X0Y1_EE4END[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(Tile_X0Y1_EE4END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(Tile_X0Y1_EE4END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(Tile_X0Y1_EE4END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(Tile_X0Y1_EE4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(Tile_X0Y1_EE4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(Tile_X0Y1_FrameData[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(Tile_X0Y1_FrameData[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(Tile_X0Y1_FrameStrobe[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(Tile_X0Y1_FrameStrobe[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(Tile_X0Y1_FrameStrobe[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(Tile_X0Y1_FrameStrobe[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(Tile_X0Y1_FrameStrobe[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(Tile_X0Y1_FrameStrobe[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(Tile_X0Y1_FrameStrobe[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(Tile_X0Y1_FrameStrobe[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(Tile_X0Y1_FrameStrobe[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(Tile_X0Y1_FrameStrobe[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(Tile_X0Y1_FrameStrobe[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(Tile_X0Y1_FrameStrobe[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(Tile_X0Y1_FrameStrobe[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(Tile_X0Y1_FrameStrobe[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(Tile_X0Y1_FrameStrobe[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(Tile_X0Y1_FrameStrobe[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(Tile_X0Y1_FrameStrobe[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(Tile_X0Y1_FrameStrobe[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(Tile_X0Y1_FrameStrobe[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(Tile_X0Y1_FrameStrobe[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(Tile_X0Y1_N4END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(Tile_X0Y1_N4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(Tile_X0Y1_N4END[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(Tile_X0Y1_N4END[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(Tile_X0Y1_N4END[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(Tile_X0Y1_N4END[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(Tile_X0Y1_N4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(Tile_X0Y1_N4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(Tile_X0Y1_N4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(Tile_X0Y1_N4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(Tile_X0Y1_N4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(Tile_X0Y1_N4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(Tile_X0Y1_N4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(Tile_X0Y1_N4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(Tile_X0Y1_N4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(Tile_X0Y1_N4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(Tile_X0Y1_N4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(Tile_X0Y1_N4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(Tile_X0Y1_N4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(Tile_X0Y1_N4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(Tile_X0Y1_N4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(Tile_X0Y1_NN4END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(Tile_X0Y1_NN4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(Tile_X0Y1_NN4END[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(Tile_X0Y1_NN4END[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(Tile_X0Y1_NN4END[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(Tile_X0Y1_NN4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(Tile_X0Y1_NN4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(Tile_X0Y1_W6END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(Tile_X0Y1_WW4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(Tile_X0Y1_WW4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(_0239_));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(_1565_));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(Tile_X0Y0_W6END[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(Tile_X0Y0_W6END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(Tile_X0Y1_FrameStrobe[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(Tile_X0Y1_FrameStrobe[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(Tile_X0Y1_FrameStrobe[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(Tile_X0Y1_FrameStrobe[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(_0344_));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(_0344_));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(_0494_));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_299 (.DIODE(net1195));
 sky130_fd_sc_hd__diode_2 ANTENNA_300 (.DIODE(net1199));
 sky130_fd_sc_hd__diode_2 ANTENNA_301 (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA_302 (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA_303 (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA_304 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_305 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_306 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_307 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_308 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_309 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_310 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_311 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_312 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_313 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_314 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_315 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_316 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_317 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_318 (.DIODE(Tile_X0Y0_E6END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_319 (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA_320 (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA_321 (.DIODE(net1234));
 sky130_fd_sc_hd__diode_2 ANTENNA_322 (.DIODE(net1234));
 sky130_fd_sc_hd__diode_2 ANTENNA_323 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_324 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_325 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_326 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_327 (.DIODE(net216));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_461 ();
endmodule
