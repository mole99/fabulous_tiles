module N_term_IHP_SRAM (UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1END,
    N2END,
    N2MID,
    N4END,
    S1BEG,
    S2BEG,
    S2BEGb,
    S4BEG);
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] N1END;
 input [7:0] N2END;
 input [7:0] N2MID;
 input [15:0] N4END;
 output [3:0] S1BEG;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 output [15:0] S4BEG;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;

 sg13g2_buf_1 _00_ (.A(FrameData[0]),
    .X(net1));
 sg13g2_buf_1 _01_ (.A(FrameData[1]),
    .X(net12));
 sg13g2_buf_1 _02_ (.A(FrameData[2]),
    .X(net23));
 sg13g2_buf_1 _03_ (.A(FrameData[3]),
    .X(net26));
 sg13g2_buf_1 _04_ (.A(FrameData[4]),
    .X(net27));
 sg13g2_buf_1 _05_ (.A(FrameData[5]),
    .X(net28));
 sg13g2_buf_1 _06_ (.A(FrameData[6]),
    .X(net29));
 sg13g2_buf_1 _07_ (.A(FrameData[7]),
    .X(net30));
 sg13g2_buf_1 _08_ (.A(FrameData[8]),
    .X(net31));
 sg13g2_buf_1 _09_ (.A(FrameData[9]),
    .X(net32));
 sg13g2_buf_1 _10_ (.A(FrameData[10]),
    .X(net2));
 sg13g2_buf_1 _11_ (.A(FrameData[11]),
    .X(net3));
 sg13g2_buf_1 _12_ (.A(FrameData[12]),
    .X(net4));
 sg13g2_buf_1 _13_ (.A(FrameData[13]),
    .X(net5));
 sg13g2_buf_1 _14_ (.A(FrameData[14]),
    .X(net6));
 sg13g2_buf_1 _15_ (.A(FrameData[15]),
    .X(net7));
 sg13g2_buf_1 _16_ (.A(FrameData[16]),
    .X(net8));
 sg13g2_buf_1 _17_ (.A(FrameData[17]),
    .X(net9));
 sg13g2_buf_1 _18_ (.A(FrameData[18]),
    .X(net10));
 sg13g2_buf_1 _19_ (.A(FrameData[19]),
    .X(net11));
 sg13g2_buf_1 _20_ (.A(FrameData[20]),
    .X(net13));
 sg13g2_buf_1 _21_ (.A(FrameData[21]),
    .X(net14));
 sg13g2_buf_1 _22_ (.A(FrameData[22]),
    .X(net15));
 sg13g2_buf_1 _23_ (.A(FrameData[23]),
    .X(net16));
 sg13g2_buf_1 _24_ (.A(FrameData[24]),
    .X(net17));
 sg13g2_buf_1 _25_ (.A(FrameData[25]),
    .X(net18));
 sg13g2_buf_1 _26_ (.A(FrameData[26]),
    .X(net19));
 sg13g2_buf_1 _27_ (.A(FrameData[27]),
    .X(net20));
 sg13g2_buf_1 _28_ (.A(FrameData[28]),
    .X(net21));
 sg13g2_buf_1 _29_ (.A(FrameData[29]),
    .X(net22));
 sg13g2_buf_1 _30_ (.A(FrameData[30]),
    .X(net24));
 sg13g2_buf_1 _31_ (.A(FrameData[31]),
    .X(net25));
 sg13g2_buf_1 _32_ (.A(FrameStrobe[0]),
    .X(net33));
 sg13g2_buf_1 _33_ (.A(FrameStrobe[1]),
    .X(net44));
 sg13g2_buf_1 _34_ (.A(FrameStrobe[2]),
    .X(net45));
 sg13g2_buf_1 _35_ (.A(FrameStrobe[3]),
    .X(net46));
 sg13g2_buf_1 _36_ (.A(FrameStrobe[4]),
    .X(net47));
 sg13g2_buf_1 _37_ (.A(FrameStrobe[5]),
    .X(net48));
 sg13g2_buf_1 _38_ (.A(FrameStrobe[6]),
    .X(net49));
 sg13g2_buf_1 _39_ (.A(FrameStrobe[7]),
    .X(net50));
 sg13g2_buf_1 _40_ (.A(FrameStrobe[8]),
    .X(net51));
 sg13g2_buf_1 _41_ (.A(FrameStrobe[9]),
    .X(net52));
 sg13g2_buf_1 _42_ (.A(FrameStrobe[10]),
    .X(net34));
 sg13g2_buf_1 _43_ (.A(FrameStrobe[11]),
    .X(net35));
 sg13g2_buf_1 _44_ (.A(FrameStrobe[12]),
    .X(net36));
 sg13g2_buf_1 _45_ (.A(FrameStrobe[13]),
    .X(net37));
 sg13g2_buf_1 _46_ (.A(FrameStrobe[14]),
    .X(net38));
 sg13g2_buf_1 _47_ (.A(FrameStrobe[15]),
    .X(net39));
 sg13g2_buf_1 _48_ (.A(FrameStrobe[16]),
    .X(net40));
 sg13g2_buf_1 _49_ (.A(FrameStrobe[17]),
    .X(net41));
 sg13g2_buf_1 _50_ (.A(FrameStrobe[18]),
    .X(net42));
 sg13g2_buf_1 _51_ (.A(FrameStrobe[19]),
    .X(net43));
 sg13g2_buf_1 _52_ (.A(N1END[3]),
    .X(net53));
 sg13g2_buf_1 _53_ (.A(N1END[2]),
    .X(net54));
 sg13g2_buf_1 _54_ (.A(N1END[1]),
    .X(net55));
 sg13g2_buf_1 _55_ (.A(N1END[0]),
    .X(net56));
 sg13g2_buf_1 _56_ (.A(N2MID[7]),
    .X(net57));
 sg13g2_buf_1 _57_ (.A(N2MID[6]),
    .X(net58));
 sg13g2_buf_1 _58_ (.A(N2MID[5]),
    .X(net59));
 sg13g2_buf_1 _59_ (.A(N2MID[4]),
    .X(net60));
 sg13g2_buf_1 _60_ (.A(N2MID[3]),
    .X(net61));
 sg13g2_buf_1 _61_ (.A(N2MID[2]),
    .X(net62));
 sg13g2_buf_1 _62_ (.A(N2MID[1]),
    .X(net63));
 sg13g2_buf_1 _63_ (.A(N2MID[0]),
    .X(net64));
 sg13g2_buf_1 _64_ (.A(N2END[7]),
    .X(net65));
 sg13g2_buf_1 _65_ (.A(N2END[6]),
    .X(net66));
 sg13g2_buf_1 _66_ (.A(N2END[5]),
    .X(net67));
 sg13g2_buf_1 _67_ (.A(N2END[4]),
    .X(net68));
 sg13g2_buf_1 _68_ (.A(N2END[3]),
    .X(net69));
 sg13g2_buf_1 _69_ (.A(N2END[2]),
    .X(net70));
 sg13g2_buf_1 _70_ (.A(N2END[1]),
    .X(net71));
 sg13g2_buf_1 _71_ (.A(N2END[0]),
    .X(net72));
 sg13g2_buf_1 _72_ (.A(N4END[15]),
    .X(net73));
 sg13g2_buf_1 _73_ (.A(N4END[14]),
    .X(net80));
 sg13g2_buf_1 _74_ (.A(N4END[13]),
    .X(net81));
 sg13g2_buf_1 _75_ (.A(N4END[12]),
    .X(net82));
 sg13g2_buf_1 _76_ (.A(N4END[11]),
    .X(net83));
 sg13g2_buf_1 _77_ (.A(N4END[10]),
    .X(net84));
 sg13g2_buf_1 _78_ (.A(N4END[9]),
    .X(net85));
 sg13g2_buf_1 _79_ (.A(N4END[8]),
    .X(net86));
 sg13g2_buf_1 _80_ (.A(N4END[7]),
    .X(net87));
 sg13g2_buf_1 _81_ (.A(N4END[6]),
    .X(net88));
 sg13g2_buf_1 _82_ (.A(N4END[5]),
    .X(net74));
 sg13g2_buf_1 _83_ (.A(N4END[4]),
    .X(net75));
 sg13g2_buf_1 _84_ (.A(N4END[3]),
    .X(net76));
 sg13g2_buf_1 _85_ (.A(N4END[2]),
    .X(net77));
 sg13g2_buf_1 _86_ (.A(N4END[1]),
    .X(net78));
 sg13g2_buf_1 _87_ (.A(N4END[0]),
    .X(net79));
 sg13g2_buf_1 _88_ (.A(UserCLK),
    .X(net89));
 sg13g2_buf_1 output1 (.A(net1),
    .X(FrameData_O[0]));
 sg13g2_buf_1 output2 (.A(net2),
    .X(FrameData_O[10]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(FrameData_O[11]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(FrameData_O[12]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(FrameData_O[13]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(FrameData_O[14]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(FrameData_O[15]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(FrameData_O[16]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(FrameData_O[17]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(FrameData_O[18]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(FrameData_O[19]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(FrameData_O[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(FrameData_O[20]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(FrameData_O[21]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(FrameData_O[22]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(FrameData_O[23]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(FrameData_O[24]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(FrameData_O[25]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(FrameData_O[26]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(FrameData_O[27]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(FrameData_O[28]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(FrameData_O[29]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(FrameData_O[2]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(FrameData_O[30]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(FrameData_O[31]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(FrameData_O[3]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(FrameData_O[4]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(FrameData_O[5]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(FrameData_O[6]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(FrameData_O[7]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(FrameData_O[8]));
 sg13g2_buf_1 output32 (.A(net32),
    .X(FrameData_O[9]));
 sg13g2_buf_1 output33 (.A(net33),
    .X(FrameStrobe_O[0]));
 sg13g2_buf_1 output34 (.A(net34),
    .X(FrameStrobe_O[10]));
 sg13g2_buf_1 output35 (.A(net35),
    .X(FrameStrobe_O[11]));
 sg13g2_buf_1 output36 (.A(net36),
    .X(FrameStrobe_O[12]));
 sg13g2_buf_1 output37 (.A(net37),
    .X(FrameStrobe_O[13]));
 sg13g2_buf_1 output38 (.A(net38),
    .X(FrameStrobe_O[14]));
 sg13g2_buf_1 output39 (.A(net39),
    .X(FrameStrobe_O[15]));
 sg13g2_buf_1 output40 (.A(net40),
    .X(FrameStrobe_O[16]));
 sg13g2_buf_1 output41 (.A(net41),
    .X(FrameStrobe_O[17]));
 sg13g2_buf_1 output42 (.A(net42),
    .X(FrameStrobe_O[18]));
 sg13g2_buf_1 output43 (.A(net43),
    .X(FrameStrobe_O[19]));
 sg13g2_buf_1 output44 (.A(net44),
    .X(FrameStrobe_O[1]));
 sg13g2_buf_1 output45 (.A(net45),
    .X(FrameStrobe_O[2]));
 sg13g2_buf_1 output46 (.A(net46),
    .X(FrameStrobe_O[3]));
 sg13g2_buf_1 output47 (.A(net47),
    .X(FrameStrobe_O[4]));
 sg13g2_buf_1 output48 (.A(net48),
    .X(FrameStrobe_O[5]));
 sg13g2_buf_1 output49 (.A(net49),
    .X(FrameStrobe_O[6]));
 sg13g2_buf_1 output50 (.A(net50),
    .X(FrameStrobe_O[7]));
 sg13g2_buf_1 output51 (.A(net51),
    .X(FrameStrobe_O[8]));
 sg13g2_buf_1 output52 (.A(net52),
    .X(FrameStrobe_O[9]));
 sg13g2_buf_1 output53 (.A(net53),
    .X(S1BEG[0]));
 sg13g2_buf_1 output54 (.A(net54),
    .X(S1BEG[1]));
 sg13g2_buf_1 output55 (.A(net55),
    .X(S1BEG[2]));
 sg13g2_buf_1 output56 (.A(net56),
    .X(S1BEG[3]));
 sg13g2_buf_1 output57 (.A(net57),
    .X(S2BEG[0]));
 sg13g2_buf_1 output58 (.A(net58),
    .X(S2BEG[1]));
 sg13g2_buf_1 output59 (.A(net59),
    .X(S2BEG[2]));
 sg13g2_buf_1 output60 (.A(net60),
    .X(S2BEG[3]));
 sg13g2_buf_1 output61 (.A(net61),
    .X(S2BEG[4]));
 sg13g2_buf_1 output62 (.A(net62),
    .X(S2BEG[5]));
 sg13g2_buf_1 output63 (.A(net63),
    .X(S2BEG[6]));
 sg13g2_buf_1 output64 (.A(net64),
    .X(S2BEG[7]));
 sg13g2_buf_1 output65 (.A(net65),
    .X(S2BEGb[0]));
 sg13g2_buf_1 output66 (.A(net66),
    .X(S2BEGb[1]));
 sg13g2_buf_1 output67 (.A(net67),
    .X(S2BEGb[2]));
 sg13g2_buf_1 output68 (.A(net68),
    .X(S2BEGb[3]));
 sg13g2_buf_1 output69 (.A(net69),
    .X(S2BEGb[4]));
 sg13g2_buf_1 output70 (.A(net70),
    .X(S2BEGb[5]));
 sg13g2_buf_1 output71 (.A(net71),
    .X(S2BEGb[6]));
 sg13g2_buf_1 output72 (.A(net72),
    .X(S2BEGb[7]));
 sg13g2_buf_1 output73 (.A(net73),
    .X(S4BEG[0]));
 sg13g2_buf_1 output74 (.A(net74),
    .X(S4BEG[10]));
 sg13g2_buf_1 output75 (.A(net75),
    .X(S4BEG[11]));
 sg13g2_buf_1 output76 (.A(net76),
    .X(S4BEG[12]));
 sg13g2_buf_1 output77 (.A(net77),
    .X(S4BEG[13]));
 sg13g2_buf_1 output78 (.A(net78),
    .X(S4BEG[14]));
 sg13g2_buf_1 output79 (.A(net79),
    .X(S4BEG[15]));
 sg13g2_buf_1 output80 (.A(net80),
    .X(S4BEG[1]));
 sg13g2_buf_1 output81 (.A(net81),
    .X(S4BEG[2]));
 sg13g2_buf_1 output82 (.A(net82),
    .X(S4BEG[3]));
 sg13g2_buf_1 output83 (.A(net83),
    .X(S4BEG[4]));
 sg13g2_buf_1 output84 (.A(net84),
    .X(S4BEG[5]));
 sg13g2_buf_1 output85 (.A(net85),
    .X(S4BEG[6]));
 sg13g2_buf_1 output86 (.A(net86),
    .X(S4BEG[7]));
 sg13g2_buf_1 output87 (.A(net87),
    .X(S4BEG[8]));
 sg13g2_buf_1 output88 (.A(net88),
    .X(S4BEG[9]));
 sg13g2_buf_1 output89 (.A(net89),
    .X(UserCLKo));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_fill_2 FILLER_0_70 ();
 sg13g2_fill_1 FILLER_0_72 ();
 sg13g2_decap_8 FILLER_0_165 ();
 sg13g2_decap_4 FILLER_0_172 ();
 sg13g2_fill_1 FILLER_0_176 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_fill_2 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_17 ();
 sg13g2_decap_8 FILLER_1_24 ();
 sg13g2_decap_8 FILLER_1_31 ();
 sg13g2_decap_8 FILLER_1_38 ();
 sg13g2_decap_8 FILLER_1_45 ();
 sg13g2_decap_8 FILLER_1_52 ();
 sg13g2_decap_8 FILLER_1_59 ();
 sg13g2_decap_8 FILLER_1_66 ();
 sg13g2_decap_8 FILLER_1_73 ();
 sg13g2_fill_1 FILLER_1_80 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_fill_1 FILLER_1_147 ();
 sg13g2_decap_4 FILLER_1_156 ();
 sg13g2_decap_8 FILLER_1_172 ();
 sg13g2_decap_4 FILLER_1_179 ();
 sg13g2_fill_1 FILLER_1_183 ();
 sg13g2_fill_1 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_4 FILLER_2_7 ();
 sg13g2_fill_2 FILLER_2_11 ();
 sg13g2_decap_8 FILLER_2_17 ();
 sg13g2_decap_8 FILLER_2_24 ();
 sg13g2_decap_8 FILLER_2_31 ();
 sg13g2_decap_8 FILLER_2_38 ();
 sg13g2_decap_4 FILLER_2_45 ();
 sg13g2_fill_1 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_54 ();
 sg13g2_decap_8 FILLER_2_61 ();
 sg13g2_decap_8 FILLER_2_68 ();
 sg13g2_decap_8 FILLER_2_75 ();
 sg13g2_decap_8 FILLER_2_82 ();
 sg13g2_decap_8 FILLER_2_89 ();
 sg13g2_decap_8 FILLER_2_96 ();
 sg13g2_decap_8 FILLER_2_103 ();
 sg13g2_decap_8 FILLER_2_110 ();
 sg13g2_decap_8 FILLER_2_117 ();
 sg13g2_decap_8 FILLER_2_124 ();
 sg13g2_decap_8 FILLER_2_131 ();
 sg13g2_decap_8 FILLER_2_138 ();
 sg13g2_decap_4 FILLER_2_145 ();
 sg13g2_decap_8 FILLER_2_153 ();
 sg13g2_fill_2 FILLER_2_160 ();
 sg13g2_fill_1 FILLER_2_162 ();
 sg13g2_decap_8 FILLER_2_167 ();
 sg13g2_decap_8 FILLER_2_174 ();
 sg13g2_decap_4 FILLER_2_181 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_4 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_15 ();
 sg13g2_fill_2 FILLER_3_22 ();
 sg13g2_fill_1 FILLER_3_24 ();
 sg13g2_decap_8 FILLER_3_29 ();
 sg13g2_decap_8 FILLER_3_36 ();
 sg13g2_decap_8 FILLER_3_43 ();
 sg13g2_fill_2 FILLER_3_50 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_fill_2 FILLER_3_91 ();
 sg13g2_fill_1 FILLER_3_93 ();
 sg13g2_decap_4 FILLER_3_102 ();
 sg13g2_fill_2 FILLER_3_106 ();
 sg13g2_decap_8 FILLER_3_116 ();
 sg13g2_decap_4 FILLER_3_123 ();
 sg13g2_fill_2 FILLER_3_131 ();
 sg13g2_fill_1 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_142 ();
 sg13g2_decap_8 FILLER_3_149 ();
 sg13g2_decap_8 FILLER_3_160 ();
 sg13g2_decap_4 FILLER_3_167 ();
 sg13g2_fill_1 FILLER_3_171 ();
 sg13g2_decap_8 FILLER_3_176 ();
 sg13g2_fill_2 FILLER_3_183 ();
 sg13g2_fill_1 FILLER_3_185 ();
 sg13g2_fill_2 FILLER_3_194 ();
 sg13g2_fill_1 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_4 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_43 ();
 sg13g2_decap_8 FILLER_4_50 ();
 sg13g2_decap_8 FILLER_4_57 ();
 sg13g2_decap_8 FILLER_4_64 ();
 sg13g2_decap_8 FILLER_4_71 ();
 sg13g2_decap_8 FILLER_4_86 ();
 sg13g2_decap_8 FILLER_4_93 ();
 sg13g2_decap_8 FILLER_4_100 ();
 sg13g2_decap_8 FILLER_4_107 ();
 sg13g2_decap_8 FILLER_4_114 ();
 sg13g2_decap_8 FILLER_4_121 ();
 sg13g2_decap_8 FILLER_4_128 ();
 sg13g2_decap_8 FILLER_4_135 ();
 sg13g2_decap_8 FILLER_4_142 ();
 sg13g2_decap_8 FILLER_4_149 ();
 sg13g2_decap_8 FILLER_4_156 ();
 sg13g2_fill_2 FILLER_4_163 ();
 sg13g2_decap_8 FILLER_4_169 ();
 sg13g2_decap_4 FILLER_4_176 ();
 sg13g2_fill_2 FILLER_4_180 ();
 sg13g2_fill_2 FILLER_4_194 ();
 sg13g2_fill_1 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_7 ();
 sg13g2_fill_1 FILLER_5_12 ();
 sg13g2_decap_8 FILLER_5_17 ();
 sg13g2_decap_8 FILLER_5_24 ();
 sg13g2_decap_4 FILLER_5_31 ();
 sg13g2_fill_1 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_40 ();
 sg13g2_decap_8 FILLER_5_47 ();
 sg13g2_decap_8 FILLER_5_54 ();
 sg13g2_decap_8 FILLER_5_61 ();
 sg13g2_decap_8 FILLER_5_68 ();
 sg13g2_decap_4 FILLER_5_75 ();
 sg13g2_fill_2 FILLER_5_79 ();
 sg13g2_decap_8 FILLER_5_85 ();
 sg13g2_decap_8 FILLER_5_92 ();
 sg13g2_decap_8 FILLER_5_99 ();
 sg13g2_decap_8 FILLER_5_106 ();
 sg13g2_decap_8 FILLER_5_113 ();
 sg13g2_decap_8 FILLER_5_120 ();
 sg13g2_decap_8 FILLER_5_127 ();
 sg13g2_decap_8 FILLER_5_134 ();
 sg13g2_decap_8 FILLER_5_141 ();
 sg13g2_fill_2 FILLER_5_148 ();
 sg13g2_fill_1 FILLER_5_150 ();
 sg13g2_decap_8 FILLER_5_155 ();
 sg13g2_fill_2 FILLER_5_162 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_4 FILLER_5_175 ();
 sg13g2_fill_1 FILLER_5_179 ();
 sg13g2_fill_1 FILLER_5_188 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_13 ();
 sg13g2_decap_4 FILLER_6_20 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_4 FILLER_6_46 ();
 sg13g2_fill_2 FILLER_6_50 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_fill_2 FILLER_6_77 ();
 sg13g2_fill_1 FILLER_6_79 ();
 sg13g2_fill_1 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_89 ();
 sg13g2_decap_8 FILLER_6_96 ();
 sg13g2_decap_8 FILLER_6_103 ();
 sg13g2_decap_8 FILLER_6_110 ();
 sg13g2_decap_4 FILLER_6_117 ();
 sg13g2_decap_8 FILLER_6_125 ();
 sg13g2_decap_4 FILLER_6_132 ();
 sg13g2_fill_2 FILLER_6_136 ();
 sg13g2_decap_8 FILLER_6_142 ();
 sg13g2_decap_8 FILLER_6_149 ();
 sg13g2_decap_4 FILLER_6_156 ();
 sg13g2_fill_1 FILLER_6_160 ();
 sg13g2_decap_8 FILLER_6_169 ();
 sg13g2_decap_8 FILLER_6_176 ();
 sg13g2_decap_4 FILLER_6_183 ();
 sg13g2_fill_1 FILLER_6_187 ();
 sg13g2_fill_1 FILLER_6_192 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_13 ();
 sg13g2_decap_8 FILLER_7_20 ();
 sg13g2_decap_8 FILLER_7_27 ();
 sg13g2_decap_4 FILLER_7_34 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_fill_1 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_72 ();
 sg13g2_decap_8 FILLER_7_79 ();
 sg13g2_decap_8 FILLER_7_86 ();
 sg13g2_decap_8 FILLER_7_93 ();
 sg13g2_decap_8 FILLER_7_100 ();
 sg13g2_decap_8 FILLER_7_107 ();
 sg13g2_decap_8 FILLER_7_114 ();
 sg13g2_decap_8 FILLER_7_121 ();
 sg13g2_decap_8 FILLER_7_128 ();
 sg13g2_decap_8 FILLER_7_135 ();
 sg13g2_decap_4 FILLER_7_142 ();
 sg13g2_decap_8 FILLER_7_150 ();
 sg13g2_decap_8 FILLER_7_157 ();
 sg13g2_decap_8 FILLER_7_164 ();
 sg13g2_decap_8 FILLER_7_171 ();
 sg13g2_decap_8 FILLER_7_178 ();
 sg13g2_fill_1 FILLER_7_185 ();
 sg13g2_fill_2 FILLER_7_198 ();
 sg13g2_fill_1 FILLER_7_200 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_12 ();
 sg13g2_decap_8 FILLER_8_19 ();
 sg13g2_decap_8 FILLER_8_26 ();
 sg13g2_fill_1 FILLER_8_33 ();
 sg13g2_decap_8 FILLER_8_38 ();
 sg13g2_decap_8 FILLER_8_45 ();
 sg13g2_decap_4 FILLER_8_52 ();
 sg13g2_fill_2 FILLER_8_56 ();
 sg13g2_decap_4 FILLER_8_62 ();
 sg13g2_fill_1 FILLER_8_66 ();
 sg13g2_decap_4 FILLER_8_71 ();
 sg13g2_fill_2 FILLER_8_79 ();
 sg13g2_decap_4 FILLER_8_85 ();
 sg13g2_fill_2 FILLER_8_89 ();
 sg13g2_decap_8 FILLER_8_95 ();
 sg13g2_decap_8 FILLER_8_102 ();
 sg13g2_decap_8 FILLER_8_109 ();
 sg13g2_decap_8 FILLER_8_116 ();
 sg13g2_decap_8 FILLER_8_123 ();
 sg13g2_decap_8 FILLER_8_130 ();
 sg13g2_decap_8 FILLER_8_137 ();
 sg13g2_fill_2 FILLER_8_144 ();
 sg13g2_fill_1 FILLER_8_146 ();
 sg13g2_decap_8 FILLER_8_155 ();
 sg13g2_fill_2 FILLER_8_162 ();
 sg13g2_fill_1 FILLER_8_164 ();
 sg13g2_decap_4 FILLER_8_169 ();
 sg13g2_fill_1 FILLER_8_173 ();
 sg13g2_decap_8 FILLER_8_178 ();
 sg13g2_decap_8 FILLER_8_185 ();
 sg13g2_fill_1 FILLER_8_192 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_11 ();
 sg13g2_decap_8 FILLER_9_18 ();
 sg13g2_decap_8 FILLER_9_25 ();
 sg13g2_decap_8 FILLER_9_32 ();
 sg13g2_decap_8 FILLER_9_39 ();
 sg13g2_decap_8 FILLER_9_46 ();
 sg13g2_decap_8 FILLER_9_53 ();
 sg13g2_decap_8 FILLER_9_60 ();
 sg13g2_decap_8 FILLER_9_67 ();
 sg13g2_decap_4 FILLER_9_74 ();
 sg13g2_fill_1 FILLER_9_78 ();
 sg13g2_decap_8 FILLER_9_83 ();
 sg13g2_decap_8 FILLER_9_90 ();
 sg13g2_decap_8 FILLER_9_97 ();
 sg13g2_decap_8 FILLER_9_104 ();
 sg13g2_decap_8 FILLER_9_111 ();
 sg13g2_decap_4 FILLER_9_118 ();
 sg13g2_fill_1 FILLER_9_122 ();
 sg13g2_decap_8 FILLER_9_135 ();
 sg13g2_decap_4 FILLER_9_142 ();
 sg13g2_fill_2 FILLER_9_146 ();
 sg13g2_decap_8 FILLER_9_152 ();
 sg13g2_decap_8 FILLER_9_159 ();
 sg13g2_fill_1 FILLER_9_166 ();
 sg13g2_decap_8 FILLER_9_171 ();
 sg13g2_decap_8 FILLER_9_178 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_1 FILLER_10_11 ();
 sg13g2_decap_8 FILLER_10_16 ();
 sg13g2_decap_8 FILLER_10_23 ();
 sg13g2_decap_8 FILLER_10_30 ();
 sg13g2_decap_8 FILLER_10_37 ();
 sg13g2_decap_8 FILLER_10_44 ();
 sg13g2_decap_8 FILLER_10_51 ();
 sg13g2_decap_8 FILLER_10_58 ();
 sg13g2_decap_8 FILLER_10_65 ();
 sg13g2_decap_8 FILLER_10_72 ();
 sg13g2_decap_8 FILLER_10_79 ();
 sg13g2_decap_8 FILLER_10_86 ();
 sg13g2_decap_8 FILLER_10_93 ();
 sg13g2_fill_1 FILLER_10_100 ();
 sg13g2_decap_8 FILLER_10_109 ();
 sg13g2_decap_8 FILLER_10_116 ();
 sg13g2_decap_8 FILLER_10_123 ();
 sg13g2_fill_1 FILLER_10_130 ();
 sg13g2_fill_2 FILLER_10_139 ();
 sg13g2_fill_1 FILLER_10_141 ();
 sg13g2_decap_8 FILLER_10_146 ();
 sg13g2_decap_4 FILLER_10_153 ();
 sg13g2_fill_1 FILLER_10_157 ();
 sg13g2_decap_8 FILLER_10_162 ();
 sg13g2_fill_1 FILLER_10_169 ();
 sg13g2_fill_2 FILLER_10_174 ();
 sg13g2_fill_1 FILLER_10_196 ();
 sg13g2_decap_4 FILLER_11_4 ();
 sg13g2_fill_1 FILLER_11_8 ();
 sg13g2_decap_4 FILLER_11_13 ();
 sg13g2_fill_2 FILLER_11_17 ();
 sg13g2_decap_4 FILLER_11_23 ();
 sg13g2_fill_2 FILLER_11_27 ();
 sg13g2_decap_4 FILLER_11_33 ();
 sg13g2_fill_2 FILLER_11_37 ();
 sg13g2_decap_4 FILLER_11_43 ();
 sg13g2_fill_2 FILLER_11_47 ();
 sg13g2_decap_4 FILLER_11_53 ();
 sg13g2_fill_2 FILLER_11_57 ();
 sg13g2_decap_4 FILLER_11_63 ();
 sg13g2_fill_2 FILLER_11_67 ();
 sg13g2_decap_4 FILLER_11_73 ();
 sg13g2_fill_2 FILLER_11_77 ();
 sg13g2_decap_4 FILLER_11_83 ();
 sg13g2_fill_2 FILLER_11_87 ();
 sg13g2_decap_4 FILLER_11_93 ();
 sg13g2_fill_2 FILLER_11_97 ();
 sg13g2_decap_4 FILLER_11_103 ();
 sg13g2_fill_2 FILLER_11_107 ();
 sg13g2_decap_4 FILLER_11_113 ();
 sg13g2_fill_2 FILLER_11_117 ();
 sg13g2_decap_4 FILLER_11_123 ();
 sg13g2_fill_2 FILLER_11_127 ();
 sg13g2_decap_4 FILLER_11_133 ();
 sg13g2_fill_2 FILLER_11_137 ();
 sg13g2_decap_4 FILLER_11_143 ();
 sg13g2_fill_2 FILLER_11_147 ();
 sg13g2_decap_4 FILLER_11_153 ();
 sg13g2_fill_2 FILLER_11_157 ();
 sg13g2_decap_4 FILLER_11_163 ();
 sg13g2_fill_2 FILLER_11_167 ();
 sg13g2_fill_2 FILLER_11_173 ();
 sg13g2_fill_2 FILLER_11_183 ();
endmodule
