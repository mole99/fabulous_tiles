magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741601325
<< metal1 >>
rect 1152 45380 10656 45404
rect 1152 45340 4928 45380
rect 4968 45340 5010 45380
rect 5050 45340 5092 45380
rect 5132 45340 5174 45380
rect 5214 45340 5256 45380
rect 5296 45340 10656 45380
rect 1152 45316 10656 45340
rect 3483 45212 3525 45221
rect 3483 45172 3484 45212
rect 3524 45172 3525 45212
rect 3483 45163 3525 45172
rect 3963 45212 4005 45221
rect 3963 45172 3964 45212
rect 4004 45172 4005 45212
rect 3963 45163 4005 45172
rect 4347 45212 4389 45221
rect 4347 45172 4348 45212
rect 4388 45172 4389 45212
rect 4347 45163 4389 45172
rect 4731 45212 4773 45221
rect 4731 45172 4732 45212
rect 4772 45172 4773 45212
rect 4731 45163 4773 45172
rect 5115 45212 5157 45221
rect 5115 45172 5116 45212
rect 5156 45172 5157 45212
rect 5115 45163 5157 45172
rect 5883 45212 5925 45221
rect 5883 45172 5884 45212
rect 5924 45172 5925 45212
rect 5883 45163 5925 45172
rect 6267 45212 6309 45221
rect 6267 45172 6268 45212
rect 6308 45172 6309 45212
rect 6267 45163 6309 45172
rect 6651 45212 6693 45221
rect 6651 45172 6652 45212
rect 6692 45172 6693 45212
rect 6651 45163 6693 45172
rect 7035 45212 7077 45221
rect 7035 45172 7036 45212
rect 7076 45172 7077 45212
rect 7035 45163 7077 45172
rect 7419 45212 7461 45221
rect 7419 45172 7420 45212
rect 7460 45172 7461 45212
rect 7419 45163 7461 45172
rect 7803 45212 7845 45221
rect 7803 45172 7804 45212
rect 7844 45172 7845 45212
rect 7803 45163 7845 45172
rect 8187 45212 8229 45221
rect 8187 45172 8188 45212
rect 8228 45172 8229 45212
rect 8187 45163 8229 45172
rect 8571 45212 8613 45221
rect 8571 45172 8572 45212
rect 8612 45172 8613 45212
rect 8571 45163 8613 45172
rect 8955 45212 8997 45221
rect 8955 45172 8956 45212
rect 8996 45172 8997 45212
rect 8955 45163 8997 45172
rect 9339 45212 9381 45221
rect 9339 45172 9340 45212
rect 9380 45172 9381 45212
rect 9339 45163 9381 45172
rect 9723 45212 9765 45221
rect 9723 45172 9724 45212
rect 9764 45172 9765 45212
rect 9723 45163 9765 45172
rect 2331 45128 2373 45137
rect 2331 45088 2332 45128
rect 2372 45088 2373 45128
rect 2331 45079 2373 45088
rect 3387 45128 3429 45137
rect 3387 45088 3388 45128
rect 3428 45088 3429 45128
rect 3387 45079 3429 45088
rect 5499 45128 5541 45137
rect 5499 45088 5500 45128
rect 5540 45088 5541 45128
rect 5499 45079 5541 45088
rect 1306 45044 1364 45045
rect 1306 45004 1315 45044
rect 1355 45004 1364 45044
rect 1306 45003 1364 45004
rect 2122 45044 2180 45045
rect 2811 45044 2853 45053
rect 2122 45004 2131 45044
rect 2171 45004 2180 45044
rect 2122 45003 2180 45004
rect 2658 45035 2704 45044
rect 2658 44995 2659 45035
rect 2699 44995 2704 45035
rect 2811 45004 2812 45044
rect 2852 45004 2853 45044
rect 2811 44995 2853 45004
rect 2658 44986 2704 44995
rect 3147 44960 3189 44969
rect 3147 44920 3148 44960
rect 3188 44920 3189 44960
rect 3147 44911 3189 44920
rect 3723 44960 3765 44969
rect 3723 44920 3724 44960
rect 3764 44920 3765 44960
rect 3723 44911 3765 44920
rect 4203 44960 4245 44969
rect 4203 44920 4204 44960
rect 4244 44920 4245 44960
rect 4203 44911 4245 44920
rect 4587 44960 4629 44969
rect 4587 44920 4588 44960
rect 4628 44920 4629 44960
rect 4587 44911 4629 44920
rect 4971 44960 5013 44969
rect 4971 44920 4972 44960
rect 5012 44920 5013 44960
rect 4971 44911 5013 44920
rect 5355 44960 5397 44969
rect 5355 44920 5356 44960
rect 5396 44920 5397 44960
rect 5355 44911 5397 44920
rect 5739 44960 5781 44969
rect 5739 44920 5740 44960
rect 5780 44920 5781 44960
rect 5739 44911 5781 44920
rect 6123 44960 6165 44969
rect 6123 44920 6124 44960
rect 6164 44920 6165 44960
rect 6123 44911 6165 44920
rect 6507 44960 6549 44969
rect 6507 44920 6508 44960
rect 6548 44920 6549 44960
rect 6507 44911 6549 44920
rect 6891 44960 6933 44969
rect 6891 44920 6892 44960
rect 6932 44920 6933 44960
rect 6891 44911 6933 44920
rect 7275 44960 7317 44969
rect 7275 44920 7276 44960
rect 7316 44920 7317 44960
rect 7275 44911 7317 44920
rect 7659 44960 7701 44969
rect 7659 44920 7660 44960
rect 7700 44920 7701 44960
rect 7659 44911 7701 44920
rect 8043 44960 8085 44969
rect 8043 44920 8044 44960
rect 8084 44920 8085 44960
rect 8043 44911 8085 44920
rect 8427 44960 8469 44969
rect 8427 44920 8428 44960
rect 8468 44920 8469 44960
rect 8427 44911 8469 44920
rect 8811 44960 8853 44969
rect 8811 44920 8812 44960
rect 8852 44920 8853 44960
rect 8811 44911 8853 44920
rect 9195 44960 9237 44969
rect 9195 44920 9196 44960
rect 9236 44920 9237 44960
rect 9195 44911 9237 44920
rect 9579 44960 9621 44969
rect 9579 44920 9580 44960
rect 9620 44920 9621 44960
rect 9579 44911 9621 44920
rect 9963 44960 10005 44969
rect 9963 44920 9964 44960
rect 10004 44920 10005 44960
rect 9963 44911 10005 44920
rect 10347 44960 10389 44969
rect 10347 44920 10348 44960
rect 10388 44920 10389 44960
rect 10347 44911 10389 44920
rect 1515 44792 1557 44801
rect 1515 44752 1516 44792
rect 1556 44752 1557 44792
rect 1515 44743 1557 44752
rect 10587 44792 10629 44801
rect 10587 44752 10588 44792
rect 10628 44752 10629 44792
rect 10587 44743 10629 44752
rect 1152 44624 10656 44648
rect 1152 44584 3688 44624
rect 3728 44584 3770 44624
rect 3810 44584 3852 44624
rect 3892 44584 3934 44624
rect 3974 44584 4016 44624
rect 4056 44584 10656 44624
rect 1152 44560 10656 44584
rect 3867 44456 3909 44465
rect 3867 44416 3868 44456
rect 3908 44416 3909 44456
rect 3867 44407 3909 44416
rect 5211 44456 5253 44465
rect 5211 44416 5212 44456
rect 5252 44416 5253 44456
rect 5211 44407 5253 44416
rect 5595 44456 5637 44465
rect 5595 44416 5596 44456
rect 5636 44416 5637 44456
rect 5595 44407 5637 44416
rect 6171 44456 6213 44465
rect 6171 44416 6172 44456
rect 6212 44416 6213 44456
rect 6171 44407 6213 44416
rect 6555 44456 6597 44465
rect 6555 44416 6556 44456
rect 6596 44416 6597 44456
rect 6555 44407 6597 44416
rect 7035 44456 7077 44465
rect 7035 44416 7036 44456
rect 7076 44416 7077 44456
rect 7035 44407 7077 44416
rect 7419 44456 7461 44465
rect 7419 44416 7420 44456
rect 7460 44416 7461 44456
rect 7419 44407 7461 44416
rect 7803 44456 7845 44465
rect 7803 44416 7804 44456
rect 7844 44416 7845 44456
rect 7803 44407 7845 44416
rect 9243 44456 9285 44465
rect 9243 44416 9244 44456
rect 9284 44416 9285 44456
rect 9243 44407 9285 44416
rect 10203 44456 10245 44465
rect 10203 44416 10204 44456
rect 10244 44416 10245 44456
rect 10203 44407 10245 44416
rect 10587 44456 10629 44465
rect 10587 44416 10588 44456
rect 10628 44416 10629 44456
rect 10587 44407 10629 44416
rect 5115 44372 5157 44381
rect 5115 44332 5116 44372
rect 5156 44332 5157 44372
rect 5115 44323 5157 44332
rect 9627 44372 9669 44381
rect 9627 44332 9628 44372
rect 9668 44332 9669 44372
rect 9627 44323 9669 44332
rect 2475 44288 2517 44297
rect 2475 44248 2476 44288
rect 2516 44248 2517 44288
rect 2475 44239 2517 44248
rect 3627 44288 3669 44297
rect 3627 44248 3628 44288
rect 3668 44248 3669 44288
rect 3627 44239 3669 44248
rect 4011 44288 4053 44297
rect 4011 44248 4012 44288
rect 4052 44248 4053 44288
rect 4011 44239 4053 44248
rect 4395 44288 4437 44297
rect 4395 44248 4396 44288
rect 4436 44248 4437 44288
rect 4395 44239 4437 44248
rect 4827 44288 4869 44297
rect 4827 44248 4828 44288
rect 4868 44248 4869 44288
rect 4827 44239 4869 44248
rect 5451 44288 5493 44297
rect 5451 44248 5452 44288
rect 5492 44248 5493 44288
rect 5451 44239 5493 44248
rect 5835 44288 5877 44297
rect 5835 44248 5836 44288
rect 5876 44248 5877 44288
rect 5835 44239 5877 44248
rect 6411 44288 6453 44297
rect 6411 44248 6412 44288
rect 6452 44248 6453 44288
rect 6411 44239 6453 44248
rect 6795 44288 6837 44297
rect 6795 44248 6796 44288
rect 6836 44248 6837 44288
rect 6795 44239 6837 44248
rect 7275 44288 7317 44297
rect 7275 44248 7276 44288
rect 7316 44248 7317 44288
rect 7275 44239 7317 44248
rect 7659 44288 7701 44297
rect 7659 44248 7660 44288
rect 7700 44248 7701 44288
rect 7659 44239 7701 44248
rect 8043 44288 8085 44297
rect 8043 44248 8044 44288
rect 8084 44248 8085 44288
rect 8043 44239 8085 44248
rect 9003 44288 9045 44297
rect 9003 44248 9004 44288
rect 9044 44248 9045 44288
rect 9003 44239 9045 44248
rect 9387 44288 9429 44297
rect 9387 44248 9388 44288
rect 9428 44248 9429 44288
rect 9387 44239 9429 44248
rect 9963 44288 10005 44297
rect 9963 44248 9964 44288
rect 10004 44248 10005 44288
rect 9963 44239 10005 44248
rect 10347 44288 10389 44297
rect 10347 44248 10348 44288
rect 10388 44248 10389 44288
rect 10347 44239 10389 44248
rect 1306 44204 1364 44205
rect 1306 44164 1315 44204
rect 1355 44164 1364 44204
rect 1306 44163 1364 44164
rect 1930 44204 1988 44205
rect 1930 44164 1939 44204
rect 1979 44164 1988 44204
rect 1930 44163 1988 44164
rect 2715 44120 2757 44129
rect 2715 44080 2716 44120
rect 2756 44080 2757 44120
rect 2715 44071 2757 44080
rect 8523 44120 8565 44129
rect 8523 44080 8524 44120
rect 8564 44080 8565 44120
rect 8523 44071 8565 44080
rect 1515 44036 1557 44045
rect 1515 43996 1516 44036
rect 1556 43996 1557 44036
rect 1515 43987 1557 43996
rect 2139 44036 2181 44045
rect 2139 43996 2140 44036
rect 2180 43996 2181 44036
rect 2139 43987 2181 43996
rect 2938 44036 2996 44037
rect 2938 43996 2947 44036
rect 2987 43996 2996 44036
rect 2938 43995 2996 43996
rect 3226 44036 3284 44037
rect 3226 43996 3235 44036
rect 3275 43996 3284 44036
rect 3226 43995 3284 43996
rect 4251 44036 4293 44045
rect 4251 43996 4252 44036
rect 4292 43996 4293 44036
rect 4251 43987 4293 43996
rect 4635 44036 4677 44045
rect 4635 43996 4636 44036
rect 4676 43996 4677 44036
rect 4635 43987 4677 43996
rect 8218 44036 8276 44037
rect 8218 43996 8227 44036
rect 8267 43996 8276 44036
rect 8218 43995 8276 43996
rect 1152 43868 10656 43892
rect 1152 43828 4928 43868
rect 4968 43828 5010 43868
rect 5050 43828 5092 43868
rect 5132 43828 5174 43868
rect 5214 43828 5256 43868
rect 5296 43828 10656 43868
rect 1152 43804 10656 43828
rect 2458 43700 2516 43701
rect 2458 43660 2467 43700
rect 2507 43660 2516 43700
rect 2458 43659 2516 43660
rect 3483 43700 3525 43709
rect 3483 43660 3484 43700
rect 3524 43660 3525 43700
rect 3483 43651 3525 43660
rect 4107 43700 4149 43709
rect 4107 43660 4108 43700
rect 4148 43660 4149 43700
rect 4107 43651 4149 43660
rect 6394 43700 6452 43701
rect 6394 43660 6403 43700
rect 6443 43660 6452 43700
rect 6394 43659 6452 43660
rect 6682 43700 6740 43701
rect 6682 43660 6691 43700
rect 6731 43660 6740 43700
rect 6682 43659 6740 43660
rect 8026 43700 8084 43701
rect 8026 43660 8035 43700
rect 8075 43660 8084 43700
rect 8026 43659 8084 43660
rect 8506 43700 8564 43701
rect 8506 43660 8515 43700
rect 8555 43660 8564 43700
rect 8506 43659 8564 43660
rect 8986 43700 9044 43701
rect 8986 43660 8995 43700
rect 9035 43660 9044 43700
rect 8986 43659 9044 43660
rect 9370 43700 9428 43701
rect 9370 43660 9379 43700
rect 9419 43660 9428 43700
rect 9370 43659 9428 43660
rect 4875 43616 4917 43625
rect 4875 43576 4876 43616
rect 4916 43576 4917 43616
rect 4875 43567 4917 43576
rect 5739 43616 5781 43625
rect 5739 43576 5740 43616
rect 5780 43576 5781 43616
rect 5739 43567 5781 43576
rect 7083 43616 7125 43625
rect 7083 43576 7084 43616
rect 7124 43576 7125 43616
rect 7083 43567 7125 43576
rect 7371 43616 7413 43625
rect 7371 43576 7372 43616
rect 7412 43576 7413 43616
rect 7371 43567 7413 43576
rect 7659 43616 7701 43625
rect 7659 43576 7660 43616
rect 7700 43576 7701 43616
rect 7659 43567 7701 43576
rect 9675 43616 9717 43625
rect 9675 43576 9676 43616
rect 9716 43576 9717 43616
rect 9675 43567 9717 43576
rect 1786 43532 1844 43533
rect 1218 43523 1264 43532
rect 1218 43483 1219 43523
rect 1259 43483 1264 43523
rect 1786 43492 1795 43532
rect 1835 43492 1844 43532
rect 1786 43491 1844 43492
rect 1218 43474 1264 43483
rect 1371 43448 1413 43457
rect 1371 43408 1372 43448
rect 1412 43408 1413 43448
rect 1371 43399 1413 43408
rect 2859 43448 2901 43457
rect 2859 43408 2860 43448
rect 2900 43408 2901 43448
rect 2859 43399 2901 43408
rect 3243 43448 3285 43457
rect 3243 43408 3244 43448
rect 3284 43408 3285 43448
rect 3243 43399 3285 43408
rect 3579 43448 3621 43457
rect 3579 43408 3580 43448
rect 3620 43408 3621 43448
rect 3579 43399 3621 43408
rect 3867 43448 3909 43457
rect 3867 43408 3868 43448
rect 3908 43408 3909 43448
rect 3867 43399 3909 43408
rect 4395 43448 4437 43457
rect 4395 43408 4396 43448
rect 4436 43408 4437 43448
rect 4395 43399 4437 43408
rect 5115 43448 5157 43457
rect 5115 43408 5116 43448
rect 5156 43408 5157 43448
rect 5115 43399 5157 43408
rect 5355 43448 5397 43457
rect 5355 43408 5356 43448
rect 5396 43408 5397 43448
rect 5355 43399 5397 43408
rect 6027 43448 6069 43457
rect 6027 43408 6028 43448
rect 6068 43408 6069 43448
rect 6027 43399 6069 43408
rect 6315 43448 6357 43457
rect 6315 43408 6316 43448
rect 6356 43408 6357 43448
rect 6315 43399 6357 43408
rect 8235 43448 8277 43457
rect 8235 43408 8236 43448
rect 8276 43408 8277 43448
rect 8235 43399 8277 43408
rect 8523 43448 8565 43457
rect 8523 43408 8524 43448
rect 8564 43408 8565 43448
rect 8523 43399 8565 43408
rect 9963 43448 10005 43457
rect 9963 43408 9964 43448
rect 10004 43408 10005 43448
rect 9963 43399 10005 43408
rect 10347 43448 10389 43457
rect 10347 43408 10348 43448
rect 10388 43408 10389 43448
rect 10347 43399 10389 43408
rect 3099 43364 3141 43373
rect 3099 43324 3100 43364
rect 3140 43324 3141 43364
rect 3099 43315 3141 43324
rect 4635 43364 4677 43373
rect 4635 43324 4636 43364
rect 4676 43324 4677 43364
rect 4635 43315 4677 43324
rect 10203 43364 10245 43373
rect 10203 43324 10204 43364
rect 10244 43324 10245 43364
rect 10203 43315 10245 43324
rect 1995 43280 2037 43289
rect 1995 43240 1996 43280
rect 2036 43240 2037 43280
rect 1995 43231 2037 43240
rect 10587 43280 10629 43289
rect 10587 43240 10588 43280
rect 10628 43240 10629 43280
rect 10587 43231 10629 43240
rect 1152 43112 10656 43136
rect 1152 43072 3688 43112
rect 3728 43072 3770 43112
rect 3810 43072 3852 43112
rect 3892 43072 3934 43112
rect 3974 43072 4016 43112
rect 4056 43072 10656 43112
rect 1152 43048 10656 43072
rect 1707 42944 1749 42953
rect 1707 42904 1708 42944
rect 1748 42904 1749 42944
rect 1707 42895 1749 42904
rect 3483 42944 3525 42953
rect 3483 42904 3484 42944
rect 3524 42904 3525 42944
rect 3483 42895 3525 42904
rect 5499 42944 5541 42953
rect 5499 42904 5500 42944
rect 5540 42904 5541 42944
rect 5499 42895 5541 42904
rect 2763 42776 2805 42785
rect 2763 42736 2764 42776
rect 2804 42736 2805 42776
rect 2763 42727 2805 42736
rect 3723 42776 3765 42785
rect 3723 42736 3724 42776
rect 3764 42736 3765 42776
rect 3723 42727 3765 42736
rect 4827 42776 4869 42785
rect 4827 42736 4828 42776
rect 4868 42736 4869 42776
rect 4827 42727 4869 42736
rect 5067 42776 5109 42785
rect 5067 42736 5068 42776
rect 5108 42736 5109 42776
rect 5067 42727 5109 42736
rect 5259 42776 5301 42785
rect 5259 42736 5260 42776
rect 5300 42736 5301 42776
rect 5259 42727 5301 42736
rect 8427 42776 8469 42785
rect 8427 42736 8428 42776
rect 8468 42736 8469 42776
rect 8427 42727 8469 42736
rect 9963 42776 10005 42785
rect 9963 42736 9964 42776
rect 10004 42736 10005 42776
rect 9963 42727 10005 42736
rect 10347 42776 10389 42785
rect 10347 42736 10348 42776
rect 10388 42736 10389 42776
rect 10347 42727 10389 42736
rect 1306 42692 1364 42693
rect 1306 42652 1315 42692
rect 1355 42652 1364 42692
rect 1306 42651 1364 42652
rect 2074 42692 2132 42693
rect 2074 42652 2083 42692
rect 2123 42652 2132 42692
rect 2074 42651 2132 42652
rect 3865 42692 3923 42693
rect 3865 42652 3874 42692
rect 3914 42652 3923 42692
rect 3865 42651 3923 42652
rect 4345 42692 4403 42693
rect 4345 42652 4354 42692
rect 4394 42652 4403 42692
rect 4345 42651 4403 42652
rect 6795 42692 6837 42701
rect 6795 42652 6796 42692
rect 6836 42652 6837 42692
rect 6795 42643 6837 42652
rect 8715 42692 8757 42701
rect 8715 42652 8716 42692
rect 8756 42652 8757 42692
rect 8715 42643 8757 42652
rect 9387 42692 9429 42701
rect 9387 42652 9388 42692
rect 9428 42652 9429 42692
rect 9387 42643 9429 42652
rect 6507 42608 6549 42617
rect 6507 42568 6508 42608
rect 6548 42568 6549 42608
rect 6507 42559 6549 42568
rect 7083 42608 7125 42617
rect 7083 42568 7084 42608
rect 7124 42568 7125 42608
rect 7083 42559 7125 42568
rect 7947 42608 7989 42617
rect 7947 42568 7948 42608
rect 7988 42568 7989 42608
rect 7947 42559 7989 42568
rect 9675 42608 9717 42617
rect 9675 42568 9676 42608
rect 9716 42568 9717 42608
rect 9675 42559 9717 42568
rect 10203 42608 10245 42617
rect 10203 42568 10204 42608
rect 10244 42568 10245 42608
rect 10203 42559 10245 42568
rect 2283 42524 2325 42533
rect 2283 42484 2284 42524
rect 2324 42484 2325 42524
rect 2283 42475 2325 42484
rect 3003 42524 3045 42533
rect 3003 42484 3004 42524
rect 3044 42484 3045 42524
rect 3003 42475 3045 42484
rect 3322 42524 3380 42525
rect 3322 42484 3331 42524
rect 3371 42484 3380 42524
rect 3322 42483 3380 42484
rect 4059 42524 4101 42533
rect 4059 42484 4060 42524
rect 4100 42484 4101 42524
rect 4059 42475 4101 42484
rect 4539 42524 4581 42533
rect 4539 42484 4540 42524
rect 4580 42484 4581 42524
rect 4539 42475 4581 42484
rect 5722 42524 5780 42525
rect 5722 42484 5731 42524
rect 5771 42484 5780 42524
rect 5722 42483 5780 42484
rect 5914 42524 5972 42525
rect 5914 42484 5923 42524
rect 5963 42484 5972 42524
rect 5914 42483 5972 42484
rect 6298 42524 6356 42525
rect 6298 42484 6307 42524
rect 6347 42484 6356 42524
rect 6298 42483 6356 42484
rect 7354 42524 7412 42525
rect 7354 42484 7363 42524
rect 7403 42484 7412 42524
rect 7354 42483 7412 42484
rect 7642 42524 7700 42525
rect 7642 42484 7651 42524
rect 7691 42484 7700 42524
rect 7642 42483 7700 42484
rect 8986 42524 9044 42525
rect 8986 42484 8995 42524
rect 9035 42484 9044 42524
rect 8986 42483 9044 42484
rect 9466 42524 9524 42525
rect 9466 42484 9475 42524
rect 9515 42484 9524 42524
rect 9466 42483 9524 42484
rect 10587 42524 10629 42533
rect 10587 42484 10588 42524
rect 10628 42484 10629 42524
rect 10587 42475 10629 42484
rect 1152 42356 10656 42380
rect 1152 42316 4928 42356
rect 4968 42316 5010 42356
rect 5050 42316 5092 42356
rect 5132 42316 5174 42356
rect 5214 42316 5256 42356
rect 5296 42316 10656 42356
rect 1152 42292 10656 42316
rect 2283 42188 2325 42197
rect 2283 42148 2284 42188
rect 2324 42148 2325 42188
rect 2283 42139 2325 42148
rect 4731 42188 4773 42197
rect 4731 42148 4732 42188
rect 4772 42148 4773 42188
rect 4731 42139 4773 42148
rect 7995 42188 8037 42197
rect 7995 42148 7996 42188
rect 8036 42148 8037 42188
rect 7995 42139 8037 42148
rect 8410 42188 8468 42189
rect 8410 42148 8419 42188
rect 8459 42148 8468 42188
rect 8410 42147 8468 42148
rect 9627 42188 9669 42197
rect 9627 42148 9628 42188
rect 9668 42148 9669 42188
rect 9627 42139 9669 42148
rect 1707 42104 1749 42113
rect 1707 42064 1708 42104
rect 1748 42064 1749 42104
rect 1707 42055 1749 42064
rect 3675 42104 3717 42113
rect 3675 42064 3676 42104
rect 3716 42064 3717 42104
rect 3675 42055 3717 42064
rect 4875 42104 4917 42113
rect 4875 42064 4876 42104
rect 4916 42064 4917 42104
rect 4875 42055 4917 42064
rect 5931 42104 5973 42113
rect 5931 42064 5932 42104
rect 5972 42064 5973 42104
rect 5931 42055 5973 42064
rect 8715 42104 8757 42113
rect 8715 42064 8716 42104
rect 8756 42064 8757 42104
rect 8715 42055 8757 42064
rect 9003 42104 9045 42113
rect 9003 42064 9004 42104
rect 9044 42064 9045 42104
rect 9003 42055 9045 42064
rect 1306 42020 1364 42021
rect 1306 41980 1315 42020
rect 1355 41980 1364 42020
rect 1306 41979 1364 41980
rect 2074 42020 2132 42021
rect 2074 41980 2083 42020
rect 2123 41980 2132 42020
rect 2074 41979 2132 41980
rect 2842 42020 2900 42021
rect 5643 42020 5685 42029
rect 2842 41980 2851 42020
rect 2891 41980 2900 42020
rect 2842 41979 2900 41980
rect 3522 42011 3568 42020
rect 3522 41971 3523 42011
rect 3563 41971 3568 42011
rect 3522 41962 3568 41971
rect 4002 42011 4048 42020
rect 4002 41971 4003 42011
rect 4043 41971 4048 42011
rect 4002 41962 4048 41971
rect 5154 42011 5200 42020
rect 5154 41971 5155 42011
rect 5195 41971 5200 42011
rect 5643 41980 5644 42020
rect 5684 41980 5685 42020
rect 5643 41971 5685 41980
rect 6411 42020 6453 42029
rect 10059 42020 10101 42029
rect 6411 41980 6412 42020
rect 6452 41980 6453 42020
rect 6411 41971 6453 41980
rect 7659 42011 7701 42020
rect 7659 41971 7660 42011
rect 7700 41971 7701 42011
rect 10059 41980 10060 42020
rect 10100 41980 10101 42020
rect 10059 41971 10101 41980
rect 5154 41962 5200 41971
rect 7659 41962 7701 41971
rect 4155 41936 4197 41945
rect 4155 41896 4156 41936
rect 4196 41896 4197 41936
rect 4155 41887 4197 41896
rect 4491 41936 4533 41945
rect 4491 41896 4492 41936
rect 4532 41896 4533 41936
rect 4491 41887 4533 41896
rect 5307 41936 5349 41945
rect 5307 41896 5308 41936
rect 5348 41896 5349 41936
rect 5307 41887 5349 41896
rect 8235 41936 8277 41945
rect 8235 41896 8236 41936
rect 8276 41896 8277 41936
rect 8235 41887 8277 41896
rect 9291 41936 9333 41945
rect 9291 41896 9292 41936
rect 9332 41896 9333 41936
rect 9291 41887 9333 41896
rect 9867 41936 9909 41945
rect 9867 41896 9868 41936
rect 9908 41896 9909 41936
rect 9867 41887 9909 41896
rect 10347 41936 10389 41945
rect 10347 41896 10348 41936
rect 10388 41896 10389 41936
rect 10347 41887 10389 41896
rect 10587 41936 10629 41945
rect 10587 41896 10588 41936
rect 10628 41896 10629 41936
rect 10587 41887 10629 41896
rect 3051 41852 3093 41861
rect 3051 41812 3052 41852
rect 3092 41812 3093 41852
rect 3051 41803 3093 41812
rect 7851 41852 7893 41861
rect 7851 41812 7852 41852
rect 7892 41812 7893 41852
rect 7851 41803 7893 41812
rect 9531 41852 9573 41861
rect 9531 41812 9532 41852
rect 9572 41812 9573 41852
rect 9531 41803 9573 41812
rect 1152 41600 10656 41624
rect 1152 41560 3688 41600
rect 3728 41560 3770 41600
rect 3810 41560 3852 41600
rect 3892 41560 3934 41600
rect 3974 41560 4016 41600
rect 4056 41560 10656 41600
rect 1152 41536 10656 41560
rect 1227 41264 1269 41273
rect 1227 41224 1228 41264
rect 1268 41224 1269 41264
rect 1227 41215 1269 41224
rect 3339 41264 3381 41273
rect 3339 41224 3340 41264
rect 3380 41224 3381 41264
rect 3339 41215 3381 41224
rect 6123 41264 6165 41273
rect 6123 41224 6124 41264
rect 6164 41224 6165 41264
rect 6123 41215 6165 41224
rect 9963 41264 10005 41273
rect 9963 41224 9964 41264
rect 10004 41224 10005 41264
rect 9963 41215 10005 41224
rect 10347 41264 10389 41273
rect 10347 41224 10348 41264
rect 10388 41224 10389 41264
rect 10347 41215 10389 41224
rect 1611 41180 1653 41189
rect 1611 41140 1612 41180
rect 1652 41140 1653 41180
rect 1611 41131 1653 41140
rect 2851 41180 2909 41181
rect 2851 41140 2860 41180
rect 2900 41140 2909 41180
rect 2851 41139 2909 41140
rect 3819 41180 3861 41189
rect 3819 41140 3820 41180
rect 3860 41140 3861 41180
rect 3819 41131 3861 41140
rect 5063 41180 5121 41181
rect 5063 41140 5072 41180
rect 5112 41140 5121 41180
rect 5063 41139 5121 41140
rect 5593 41180 5651 41181
rect 5593 41140 5602 41180
rect 5642 41140 5651 41180
rect 5593 41139 5651 41140
rect 6411 41180 6453 41189
rect 6411 41140 6412 41180
rect 6452 41140 6453 41180
rect 6411 41131 6453 41140
rect 7651 41180 7709 41181
rect 7651 41140 7660 41180
rect 7700 41140 7709 41180
rect 7651 41139 7709 41140
rect 8043 41180 8085 41189
rect 8043 41140 8044 41180
rect 8084 41140 8085 41180
rect 8043 41131 8085 41140
rect 9283 41180 9341 41181
rect 9283 41140 9292 41180
rect 9332 41140 9341 41180
rect 9283 41139 9341 41140
rect 10203 41096 10245 41105
rect 10203 41056 10204 41096
rect 10244 41056 10245 41096
rect 10203 41047 10245 41056
rect 1467 41012 1509 41021
rect 1467 40972 1468 41012
rect 1508 40972 1509 41012
rect 1467 40963 1509 40972
rect 3051 41012 3093 41021
rect 3051 40972 3052 41012
rect 3092 40972 3093 41012
rect 3051 40963 3093 40972
rect 3322 41012 3380 41013
rect 3322 40972 3331 41012
rect 3371 40972 3380 41012
rect 3322 40971 3380 40972
rect 3610 41012 3668 41013
rect 3610 40972 3619 41012
rect 3659 40972 3668 41012
rect 3610 40971 3668 40972
rect 5259 41012 5301 41021
rect 5259 40972 5260 41012
rect 5300 40972 5301 41012
rect 5259 40963 5301 40972
rect 5787 41012 5829 41021
rect 5787 40972 5788 41012
rect 5828 40972 5829 41012
rect 5787 40963 5829 40972
rect 6202 41012 6260 41013
rect 6202 40972 6211 41012
rect 6251 40972 6260 41012
rect 6202 40971 6260 40972
rect 7851 41012 7893 41021
rect 7851 40972 7852 41012
rect 7892 40972 7893 41012
rect 7851 40963 7893 40972
rect 9483 41012 9525 41021
rect 9483 40972 9484 41012
rect 9524 40972 9525 41012
rect 9483 40963 9525 40972
rect 9754 41012 9812 41013
rect 9754 40972 9763 41012
rect 9803 40972 9812 41012
rect 9754 40971 9812 40972
rect 10587 41012 10629 41021
rect 10587 40972 10588 41012
rect 10628 40972 10629 41012
rect 10587 40963 10629 40972
rect 1152 40844 10656 40868
rect 1152 40804 4928 40844
rect 4968 40804 5010 40844
rect 5050 40804 5092 40844
rect 5132 40804 5174 40844
rect 5214 40804 5256 40844
rect 5296 40804 10656 40844
rect 1152 40780 10656 40804
rect 5547 40676 5589 40685
rect 5547 40636 5548 40676
rect 5588 40636 5589 40676
rect 5547 40627 5589 40636
rect 5979 40676 6021 40685
rect 5979 40636 5980 40676
rect 6020 40636 6021 40676
rect 5979 40627 6021 40636
rect 9579 40676 9621 40685
rect 9579 40636 9580 40676
rect 9620 40636 9621 40676
rect 9579 40627 9621 40636
rect 3531 40592 3573 40601
rect 3531 40552 3532 40592
rect 3572 40552 3573 40592
rect 3531 40543 3573 40552
rect 7563 40592 7605 40601
rect 7563 40552 7564 40592
rect 7604 40552 7605 40592
rect 7563 40543 7605 40552
rect 1306 40508 1364 40509
rect 1306 40468 1315 40508
rect 1355 40468 1364 40508
rect 1306 40467 1364 40468
rect 2091 40508 2133 40517
rect 3802 40508 3860 40509
rect 2091 40468 2092 40508
rect 2132 40468 2133 40508
rect 2091 40459 2133 40468
rect 3339 40499 3381 40508
rect 3339 40459 3340 40499
rect 3380 40459 3381 40499
rect 3802 40468 3811 40508
rect 3851 40468 3860 40508
rect 3802 40467 3860 40468
rect 3915 40508 3957 40517
rect 3915 40468 3916 40508
rect 3956 40468 3957 40508
rect 3915 40459 3957 40468
rect 4299 40508 4341 40517
rect 6123 40508 6165 40517
rect 7834 40508 7892 40509
rect 4299 40468 4300 40508
rect 4340 40468 4341 40508
rect 4299 40459 4341 40468
rect 4875 40499 4917 40508
rect 4875 40459 4876 40499
rect 4916 40459 4917 40499
rect 3339 40450 3381 40459
rect 4875 40450 4917 40459
rect 5355 40499 5397 40508
rect 5355 40459 5356 40499
rect 5396 40459 5397 40499
rect 6123 40468 6124 40508
rect 6164 40468 6165 40508
rect 6123 40459 6165 40468
rect 7371 40499 7413 40508
rect 7371 40459 7372 40499
rect 7412 40459 7413 40499
rect 7834 40468 7843 40508
rect 7883 40468 7892 40508
rect 7834 40467 7892 40468
rect 7947 40508 7989 40517
rect 7947 40468 7948 40508
rect 7988 40468 7989 40508
rect 7947 40459 7989 40468
rect 8331 40508 8373 40517
rect 8331 40468 8332 40508
rect 8372 40468 8373 40508
rect 8331 40459 8373 40468
rect 8907 40499 8949 40508
rect 8907 40459 8908 40499
rect 8948 40459 8949 40499
rect 5355 40450 5397 40459
rect 7371 40450 7413 40459
rect 8907 40450 8949 40459
rect 9387 40499 9429 40508
rect 9387 40459 9388 40499
rect 9428 40459 9429 40499
rect 9387 40450 9429 40459
rect 10242 40499 10288 40508
rect 10242 40459 10243 40499
rect 10283 40459 10288 40499
rect 10242 40450 10288 40459
rect 4395 40424 4437 40433
rect 4395 40384 4396 40424
rect 4436 40384 4437 40424
rect 4395 40375 4437 40384
rect 5739 40424 5781 40433
rect 5739 40384 5740 40424
rect 5780 40384 5781 40424
rect 5739 40375 5781 40384
rect 8427 40424 8469 40433
rect 8427 40384 8428 40424
rect 8468 40384 8469 40424
rect 8427 40375 8469 40384
rect 9963 40424 10005 40433
rect 9963 40384 9964 40424
rect 10004 40384 10005 40424
rect 9963 40375 10005 40384
rect 10395 40424 10437 40433
rect 10395 40384 10396 40424
rect 10436 40384 10437 40424
rect 10395 40375 10437 40384
rect 1515 40340 1557 40349
rect 1515 40300 1516 40340
rect 1556 40300 1557 40340
rect 1515 40291 1557 40300
rect 1152 40088 10656 40112
rect 1152 40048 3688 40088
rect 3728 40048 3770 40088
rect 3810 40048 3852 40088
rect 3892 40048 3934 40088
rect 3974 40048 4016 40088
rect 4056 40048 10656 40088
rect 1152 40024 10656 40048
rect 6267 39836 6309 39845
rect 6267 39796 6268 39836
rect 6308 39796 6309 39836
rect 6267 39787 6309 39796
rect 3723 39752 3765 39761
rect 3723 39712 3724 39752
rect 3764 39712 3765 39752
rect 3723 39703 3765 39712
rect 5163 39752 5205 39761
rect 5163 39712 5164 39752
rect 5204 39712 5205 39752
rect 5163 39703 5205 39712
rect 5691 39752 5733 39761
rect 5691 39712 5692 39752
rect 5732 39712 5733 39752
rect 5691 39703 5733 39712
rect 6027 39752 6069 39761
rect 6027 39712 6028 39752
rect 6068 39712 6069 39752
rect 6027 39703 6069 39712
rect 6603 39752 6645 39761
rect 6603 39712 6604 39752
rect 6644 39712 6645 39752
rect 6603 39703 6645 39712
rect 8427 39752 8469 39761
rect 8427 39712 8428 39752
rect 8468 39712 8469 39752
rect 8427 39703 8469 39712
rect 9867 39752 9909 39761
rect 9867 39712 9868 39752
rect 9908 39712 9909 39752
rect 9867 39703 9909 39712
rect 1419 39668 1461 39677
rect 1419 39628 1420 39668
rect 1460 39628 1461 39668
rect 1419 39619 1461 39628
rect 2659 39668 2717 39669
rect 2659 39628 2668 39668
rect 2708 39628 2717 39668
rect 2659 39627 2717 39628
rect 3226 39668 3284 39669
rect 3226 39628 3235 39668
rect 3275 39628 3284 39668
rect 3226 39627 3284 39628
rect 3339 39668 3381 39677
rect 3339 39628 3340 39668
rect 3380 39628 3381 39668
rect 3339 39619 3381 39628
rect 3819 39668 3861 39677
rect 3819 39628 3820 39668
rect 3860 39628 3861 39668
rect 3819 39619 3861 39628
rect 4291 39668 4349 39669
rect 4291 39628 4300 39668
rect 4340 39628 4349 39668
rect 4291 39627 4349 39628
rect 4779 39668 4837 39669
rect 4779 39628 4788 39668
rect 4828 39628 4837 39668
rect 4779 39627 4837 39628
rect 5527 39668 5585 39669
rect 5527 39628 5536 39668
rect 5576 39628 5585 39668
rect 5527 39627 5585 39628
rect 7917 39668 7959 39677
rect 7917 39628 7918 39668
rect 7958 39628 7959 39668
rect 7917 39619 7959 39628
rect 8032 39668 8090 39669
rect 8032 39628 8041 39668
rect 8081 39628 8090 39668
rect 8032 39627 8090 39628
rect 8523 39668 8565 39677
rect 8523 39628 8524 39668
rect 8564 39628 8565 39668
rect 8523 39619 8565 39628
rect 8995 39668 9053 39669
rect 8995 39628 9004 39668
rect 9044 39628 9053 39668
rect 8995 39627 9053 39628
rect 9483 39668 9541 39669
rect 9483 39628 9492 39668
rect 9532 39628 9541 39668
rect 9483 39627 9541 39628
rect 10186 39668 10244 39669
rect 10186 39628 10195 39668
rect 10235 39628 10244 39668
rect 10186 39627 10244 39628
rect 5403 39584 5445 39593
rect 5403 39544 5404 39584
rect 5444 39544 5445 39584
rect 5403 39535 5445 39544
rect 2859 39500 2901 39509
rect 2859 39460 2860 39500
rect 2900 39460 2901 39500
rect 2859 39451 2901 39460
rect 4971 39500 5013 39509
rect 4971 39460 4972 39500
rect 5012 39460 5013 39500
rect 4971 39451 5013 39460
rect 6363 39500 6405 39509
rect 6363 39460 6364 39500
rect 6404 39460 6405 39500
rect 6363 39451 6405 39460
rect 6874 39500 6932 39501
rect 6874 39460 6883 39500
rect 6923 39460 6932 39500
rect 6874 39459 6932 39460
rect 7066 39500 7124 39501
rect 7066 39460 7075 39500
rect 7115 39460 7124 39500
rect 7066 39459 7124 39460
rect 7354 39500 7412 39501
rect 7354 39460 7363 39500
rect 7403 39460 7412 39500
rect 7354 39459 7412 39460
rect 9675 39500 9717 39509
rect 9675 39460 9676 39500
rect 9716 39460 9717 39500
rect 9675 39451 9717 39460
rect 10107 39500 10149 39509
rect 10107 39460 10108 39500
rect 10148 39460 10149 39500
rect 10107 39451 10149 39460
rect 10395 39500 10437 39509
rect 10395 39460 10396 39500
rect 10436 39460 10437 39500
rect 10395 39451 10437 39460
rect 1152 39332 10656 39356
rect 1152 39292 4928 39332
rect 4968 39292 5010 39332
rect 5050 39292 5092 39332
rect 5132 39292 5174 39332
rect 5214 39292 5256 39332
rect 5296 39292 10656 39332
rect 1152 39268 10656 39292
rect 3195 39164 3237 39173
rect 3195 39124 3196 39164
rect 3236 39124 3237 39164
rect 3195 39115 3237 39124
rect 5451 39164 5493 39173
rect 5451 39124 5452 39164
rect 5492 39124 5493 39164
rect 5451 39115 5493 39124
rect 9963 39164 10005 39173
rect 9963 39124 9964 39164
rect 10004 39124 10005 39164
rect 9963 39115 10005 39124
rect 2859 39080 2901 39089
rect 2859 39040 2860 39080
rect 2900 39040 2901 39080
rect 2859 39031 2901 39040
rect 1419 38996 1461 39005
rect 4011 38996 4053 39005
rect 6123 38996 6165 39005
rect 8214 38996 8272 38997
rect 1419 38956 1420 38996
rect 1460 38956 1461 38996
rect 1419 38947 1461 38956
rect 2667 38987 2709 38996
rect 2667 38947 2668 38987
rect 2708 38947 2709 38987
rect 2667 38938 2709 38947
rect 3042 38987 3088 38996
rect 3042 38947 3043 38987
rect 3083 38947 3088 38987
rect 3042 38938 3088 38947
rect 3522 38987 3568 38996
rect 3522 38947 3523 38987
rect 3563 38947 3568 38987
rect 4011 38956 4012 38996
rect 4052 38956 4053 38996
rect 4011 38947 4053 38956
rect 5259 38987 5301 38996
rect 5259 38947 5260 38987
rect 5300 38947 5301 38987
rect 3522 38938 3568 38947
rect 5259 38938 5301 38947
rect 5634 38987 5680 38996
rect 5634 38947 5635 38987
rect 5675 38947 5680 38987
rect 6123 38956 6124 38996
rect 6164 38956 6165 38996
rect 6123 38947 6165 38956
rect 7371 38987 7413 38996
rect 7371 38947 7372 38987
rect 7412 38947 7413 38987
rect 8214 38956 8223 38996
rect 8263 38956 8272 38996
rect 8214 38955 8272 38956
rect 8331 38996 8373 39005
rect 8331 38956 8332 38996
rect 8372 38956 8373 38996
rect 8331 38947 8373 38956
rect 8715 38996 8757 39005
rect 8715 38956 8716 38996
rect 8756 38956 8757 38996
rect 8715 38947 8757 38956
rect 9291 38987 9333 38996
rect 9291 38947 9292 38987
rect 9332 38947 9333 38987
rect 5634 38938 5680 38947
rect 7371 38938 7413 38947
rect 9291 38938 9333 38947
rect 9771 38987 9813 38996
rect 9771 38947 9772 38987
rect 9812 38947 9813 38987
rect 9771 38938 9813 38947
rect 10146 38987 10192 38996
rect 10146 38947 10147 38987
rect 10187 38947 10192 38987
rect 10146 38938 10192 38947
rect 3675 38912 3717 38921
rect 3675 38872 3676 38912
rect 3716 38872 3717 38912
rect 3675 38863 3717 38872
rect 5787 38912 5829 38921
rect 5787 38872 5788 38912
rect 5828 38872 5829 38912
rect 5787 38863 5829 38872
rect 7755 38912 7797 38921
rect 7755 38872 7756 38912
rect 7796 38872 7797 38912
rect 7755 38863 7797 38872
rect 8811 38912 8853 38921
rect 8811 38872 8812 38912
rect 8852 38872 8853 38912
rect 8811 38863 8853 38872
rect 10299 38912 10341 38921
rect 10299 38872 10300 38912
rect 10340 38872 10341 38912
rect 10299 38863 10341 38872
rect 7563 38744 7605 38753
rect 7563 38704 7564 38744
rect 7604 38704 7605 38744
rect 7563 38695 7605 38704
rect 7995 38744 8037 38753
rect 7995 38704 7996 38744
rect 8036 38704 8037 38744
rect 7995 38695 8037 38704
rect 1152 38576 10656 38600
rect 1152 38536 3688 38576
rect 3728 38536 3770 38576
rect 3810 38536 3852 38576
rect 3892 38536 3934 38576
rect 3974 38536 4016 38576
rect 4056 38536 10656 38576
rect 1152 38512 10656 38536
rect 8427 38408 8469 38417
rect 8427 38368 8428 38408
rect 8468 38368 8469 38408
rect 8427 38359 8469 38368
rect 10251 38408 10293 38417
rect 10251 38368 10252 38408
rect 10292 38368 10293 38408
rect 10251 38359 10293 38368
rect 2235 38324 2277 38333
rect 2235 38284 2236 38324
rect 2276 38284 2277 38324
rect 2235 38275 2277 38284
rect 1995 38240 2037 38249
rect 1995 38200 1996 38240
rect 2036 38200 2037 38240
rect 1995 38191 2037 38200
rect 10443 38240 10485 38249
rect 10443 38200 10444 38240
rect 10484 38200 10485 38240
rect 10443 38191 10485 38200
rect 1306 38156 1364 38157
rect 1306 38116 1315 38156
rect 1355 38116 1364 38156
rect 1306 38115 1364 38116
rect 2379 38156 2421 38165
rect 2379 38116 2380 38156
rect 2420 38116 2421 38156
rect 2379 38107 2421 38116
rect 3619 38156 3677 38157
rect 3619 38116 3628 38156
rect 3668 38116 3677 38156
rect 3619 38115 3677 38116
rect 4203 38156 4245 38165
rect 4203 38116 4204 38156
rect 4244 38116 4245 38156
rect 4203 38107 4245 38116
rect 5443 38156 5501 38157
rect 5443 38116 5452 38156
rect 5492 38116 5501 38156
rect 5443 38115 5501 38116
rect 5866 38156 5924 38157
rect 5866 38116 5875 38156
rect 5915 38116 5924 38156
rect 5866 38115 5924 38116
rect 6361 38156 6419 38157
rect 6361 38116 6370 38156
rect 6410 38116 6419 38156
rect 6361 38115 6419 38116
rect 6987 38156 7029 38165
rect 6987 38116 6988 38156
rect 7028 38116 7029 38156
rect 6987 38107 7029 38116
rect 8227 38156 8285 38157
rect 8227 38116 8236 38156
rect 8276 38116 8285 38156
rect 8227 38115 8285 38116
rect 8811 38156 8853 38165
rect 8811 38116 8812 38156
rect 8852 38116 8853 38156
rect 8811 38107 8853 38116
rect 10051 38156 10109 38157
rect 10051 38116 10060 38156
rect 10100 38116 10109 38156
rect 10051 38115 10109 38116
rect 1594 38072 1652 38073
rect 1594 38032 1603 38072
rect 1643 38032 1652 38072
rect 1594 38031 1652 38032
rect 6555 38072 6597 38081
rect 6555 38032 6556 38072
rect 6596 38032 6597 38072
rect 6555 38023 6597 38032
rect 3819 37988 3861 37997
rect 3819 37948 3820 37988
rect 3860 37948 3861 37988
rect 3819 37939 3861 37948
rect 5643 37988 5685 37997
rect 5643 37948 5644 37988
rect 5684 37948 5685 37988
rect 5643 37939 5685 37948
rect 6075 37988 6117 37997
rect 6075 37948 6076 37988
rect 6116 37948 6117 37988
rect 6075 37939 6117 37948
rect 1152 37820 10656 37844
rect 1152 37780 4928 37820
rect 4968 37780 5010 37820
rect 5050 37780 5092 37820
rect 5132 37780 5174 37820
rect 5214 37780 5256 37820
rect 5296 37780 10656 37820
rect 1152 37756 10656 37780
rect 3562 37652 3620 37653
rect 3562 37612 3571 37652
rect 3611 37612 3620 37652
rect 3562 37611 3620 37612
rect 5739 37652 5781 37661
rect 5739 37612 5740 37652
rect 5780 37612 5781 37652
rect 5739 37603 5781 37612
rect 8218 37652 8276 37653
rect 8218 37612 8227 37652
rect 8267 37612 8276 37652
rect 8218 37611 8276 37612
rect 3099 37568 3141 37577
rect 3099 37528 3100 37568
rect 3140 37528 3141 37568
rect 3099 37519 3141 37528
rect 1306 37484 1364 37485
rect 2139 37484 2181 37493
rect 2619 37484 2661 37493
rect 3757 37484 3815 37485
rect 1306 37444 1315 37484
rect 1355 37444 1364 37484
rect 1306 37443 1364 37444
rect 1986 37475 2032 37484
rect 1986 37435 1987 37475
rect 2027 37435 2032 37475
rect 2139 37444 2140 37484
rect 2180 37444 2181 37484
rect 2139 37435 2181 37444
rect 2466 37475 2512 37484
rect 2466 37435 2467 37475
rect 2507 37435 2512 37475
rect 2619 37444 2620 37484
rect 2660 37444 2661 37484
rect 2619 37435 2661 37444
rect 2946 37475 2992 37484
rect 2946 37435 2947 37475
rect 2987 37435 2992 37475
rect 3757 37444 3766 37484
rect 3806 37444 3815 37484
rect 3757 37443 3815 37444
rect 3994 37484 4052 37485
rect 3994 37444 4003 37484
rect 4043 37444 4052 37484
rect 3994 37443 4052 37444
rect 4107 37484 4149 37493
rect 4107 37444 4108 37484
rect 4148 37444 4149 37484
rect 4107 37435 4149 37444
rect 4491 37484 4533 37493
rect 6123 37484 6165 37493
rect 7899 37484 7941 37493
rect 10347 37484 10389 37493
rect 4491 37444 4492 37484
rect 4532 37444 4533 37484
rect 4491 37435 4533 37444
rect 5067 37475 5109 37484
rect 5067 37435 5068 37475
rect 5108 37435 5109 37475
rect 1986 37426 2032 37435
rect 2466 37426 2512 37435
rect 2946 37426 2992 37435
rect 5067 37426 5109 37435
rect 5547 37475 5589 37484
rect 5547 37435 5548 37475
rect 5588 37435 5589 37475
rect 6123 37444 6124 37484
rect 6164 37444 6165 37484
rect 6123 37435 6165 37444
rect 7371 37475 7413 37484
rect 7371 37435 7372 37475
rect 7412 37435 7413 37475
rect 5547 37426 5589 37435
rect 7371 37426 7413 37435
rect 7746 37475 7792 37484
rect 7746 37435 7747 37475
rect 7787 37435 7792 37475
rect 7899 37444 7900 37484
rect 7940 37444 7941 37484
rect 7899 37435 7941 37444
rect 9095 37475 9137 37484
rect 9095 37435 9096 37475
rect 9136 37435 9137 37475
rect 10347 37444 10348 37484
rect 10388 37444 10389 37484
rect 10347 37435 10389 37444
rect 7746 37426 7792 37435
rect 9095 37426 9137 37435
rect 4587 37400 4629 37409
rect 4587 37360 4588 37400
rect 4628 37360 4629 37400
rect 4587 37351 4629 37360
rect 8523 37400 8565 37409
rect 8523 37360 8524 37400
rect 8564 37360 8565 37400
rect 8523 37351 8565 37360
rect 8763 37316 8805 37325
rect 8763 37276 8764 37316
rect 8804 37276 8805 37316
rect 8763 37267 8805 37276
rect 1515 37232 1557 37241
rect 1515 37192 1516 37232
rect 1556 37192 1557 37232
rect 1515 37183 1557 37192
rect 7563 37232 7605 37241
rect 7563 37192 7564 37232
rect 7604 37192 7605 37232
rect 7563 37183 7605 37192
rect 8907 37232 8949 37241
rect 8907 37192 8908 37232
rect 8948 37192 8949 37232
rect 8907 37183 8949 37192
rect 1152 37064 10656 37088
rect 1152 37024 3688 37064
rect 3728 37024 3770 37064
rect 3810 37024 3852 37064
rect 3892 37024 3934 37064
rect 3974 37024 4016 37064
rect 4056 37024 10656 37064
rect 1152 37000 10656 37024
rect 3531 36728 3573 36737
rect 3531 36688 3532 36728
rect 3572 36688 3573 36728
rect 3531 36679 3573 36688
rect 5643 36728 5685 36737
rect 5643 36688 5644 36728
rect 5684 36688 5685 36728
rect 5643 36679 5685 36688
rect 7755 36728 7797 36737
rect 7755 36688 7756 36728
rect 7796 36688 7797 36728
rect 7755 36679 7797 36688
rect 9963 36728 10005 36737
rect 9963 36688 9964 36728
rect 10004 36688 10005 36728
rect 9963 36679 10005 36688
rect 10347 36728 10389 36737
rect 10347 36688 10348 36728
rect 10388 36688 10389 36728
rect 10347 36679 10389 36688
rect 1323 36644 1365 36653
rect 1323 36604 1324 36644
rect 1364 36604 1365 36644
rect 1323 36595 1365 36604
rect 2563 36644 2621 36645
rect 2563 36604 2572 36644
rect 2612 36604 2621 36644
rect 2563 36603 2621 36604
rect 3034 36644 3092 36645
rect 3034 36604 3043 36644
rect 3083 36604 3092 36644
rect 3034 36603 3092 36604
rect 3147 36644 3189 36653
rect 3147 36604 3148 36644
rect 3188 36604 3189 36644
rect 3147 36595 3189 36604
rect 3627 36644 3669 36653
rect 3627 36604 3628 36644
rect 3668 36604 3669 36644
rect 3627 36595 3669 36604
rect 4099 36644 4157 36645
rect 4099 36604 4108 36644
rect 4148 36604 4157 36644
rect 4099 36603 4157 36604
rect 4587 36644 4645 36645
rect 4587 36604 4596 36644
rect 4636 36604 4645 36644
rect 4587 36603 4645 36604
rect 5146 36644 5204 36645
rect 5146 36604 5155 36644
rect 5195 36604 5204 36644
rect 5146 36603 5204 36604
rect 5259 36644 5301 36653
rect 5259 36604 5260 36644
rect 5300 36604 5301 36644
rect 5259 36595 5301 36604
rect 5739 36644 5781 36653
rect 5739 36604 5740 36644
rect 5780 36604 5781 36644
rect 5739 36595 5781 36604
rect 6211 36644 6269 36645
rect 6211 36604 6220 36644
rect 6260 36604 6269 36644
rect 6211 36603 6269 36604
rect 6730 36644 6788 36645
rect 6730 36604 6739 36644
rect 6779 36604 6788 36644
rect 6730 36603 6788 36604
rect 7258 36644 7316 36645
rect 7258 36604 7267 36644
rect 7307 36604 7316 36644
rect 7258 36603 7316 36604
rect 7371 36644 7413 36653
rect 7371 36604 7372 36644
rect 7412 36604 7413 36644
rect 7371 36595 7413 36604
rect 7851 36644 7893 36653
rect 7851 36604 7852 36644
rect 7892 36604 7893 36644
rect 7851 36595 7893 36604
rect 8323 36644 8381 36645
rect 8323 36604 8332 36644
rect 8372 36604 8381 36644
rect 8323 36603 8381 36604
rect 8811 36644 8869 36645
rect 8811 36604 8820 36644
rect 8860 36604 8869 36644
rect 8811 36603 8869 36604
rect 9226 36644 9284 36645
rect 9226 36604 9235 36644
rect 9275 36604 9284 36644
rect 9226 36603 9284 36604
rect 2763 36560 2805 36569
rect 2763 36520 2764 36560
rect 2804 36520 2805 36560
rect 2763 36511 2805 36520
rect 10203 36560 10245 36569
rect 10203 36520 10204 36560
rect 10244 36520 10245 36560
rect 10203 36511 10245 36520
rect 4779 36476 4821 36485
rect 4779 36436 4780 36476
rect 4820 36436 4821 36476
rect 4779 36427 4821 36436
rect 6891 36476 6933 36485
rect 6891 36436 6892 36476
rect 6932 36436 6933 36476
rect 6891 36427 6933 36436
rect 9003 36476 9045 36485
rect 9003 36436 9004 36476
rect 9044 36436 9045 36476
rect 9003 36427 9045 36436
rect 9435 36476 9477 36485
rect 9435 36436 9436 36476
rect 9476 36436 9477 36476
rect 9435 36427 9477 36436
rect 10587 36476 10629 36485
rect 10587 36436 10588 36476
rect 10628 36436 10629 36476
rect 10587 36427 10629 36436
rect 1152 36308 10656 36332
rect 1152 36268 4928 36308
rect 4968 36268 5010 36308
rect 5050 36268 5092 36308
rect 5132 36268 5174 36308
rect 5214 36268 5256 36308
rect 5296 36268 10656 36308
rect 1152 36244 10656 36268
rect 1851 36140 1893 36149
rect 1851 36100 1852 36140
rect 1892 36100 1893 36140
rect 1851 36091 1893 36100
rect 4378 36140 4436 36141
rect 4378 36100 4387 36140
rect 4427 36100 4436 36140
rect 4378 36099 4436 36100
rect 8619 36140 8661 36149
rect 8619 36100 8620 36140
rect 8660 36100 8661 36140
rect 8619 36091 8661 36100
rect 10522 36140 10580 36141
rect 10522 36100 10531 36140
rect 10571 36100 10580 36140
rect 10522 36099 10580 36100
rect 1371 36056 1413 36065
rect 1371 36016 1372 36056
rect 1412 36016 1413 36056
rect 1371 36007 1413 36016
rect 2667 35972 2709 35981
rect 4666 35972 4724 35973
rect 1218 35963 1264 35972
rect 1218 35923 1219 35963
rect 1259 35923 1264 35963
rect 1218 35914 1264 35923
rect 1698 35963 1744 35972
rect 1698 35923 1699 35963
rect 1739 35923 1744 35963
rect 1698 35914 1744 35923
rect 2178 35963 2224 35972
rect 2178 35923 2179 35963
rect 2219 35923 2224 35963
rect 2667 35932 2668 35972
rect 2708 35932 2709 35972
rect 2667 35923 2709 35932
rect 3915 35963 3957 35972
rect 3915 35923 3916 35963
rect 3956 35923 3957 35963
rect 4666 35932 4675 35972
rect 4715 35932 4724 35972
rect 4666 35931 4724 35932
rect 4779 35972 4821 35981
rect 4779 35932 4780 35972
rect 4820 35932 4821 35972
rect 4779 35923 4821 35932
rect 5163 35972 5205 35981
rect 6442 35972 6500 35973
rect 7179 35972 7221 35981
rect 10251 35972 10293 35981
rect 5163 35932 5164 35972
rect 5204 35932 5205 35972
rect 5163 35923 5205 35932
rect 5739 35963 5781 35972
rect 5739 35923 5740 35963
rect 5780 35923 5781 35963
rect 2178 35914 2224 35923
rect 3915 35914 3957 35923
rect 5739 35914 5781 35923
rect 6219 35963 6261 35972
rect 6219 35923 6220 35963
rect 6260 35923 6261 35963
rect 6442 35932 6451 35972
rect 6491 35932 6500 35972
rect 6442 35931 6500 35932
rect 6594 35963 6640 35972
rect 6219 35914 6261 35923
rect 6594 35923 6595 35963
rect 6635 35923 6640 35963
rect 7179 35932 7180 35972
rect 7220 35932 7221 35972
rect 7179 35923 7221 35932
rect 8427 35963 8469 35972
rect 8427 35923 8428 35963
rect 8468 35923 8469 35963
rect 6594 35914 6640 35923
rect 8427 35914 8469 35923
rect 9003 35963 9045 35972
rect 9003 35923 9004 35963
rect 9044 35923 9045 35963
rect 10251 35932 10252 35972
rect 10292 35932 10293 35972
rect 10251 35923 10293 35932
rect 9003 35914 9045 35923
rect 2331 35888 2373 35897
rect 2331 35848 2332 35888
rect 2372 35848 2373 35888
rect 2331 35839 2373 35848
rect 5259 35888 5301 35897
rect 5259 35848 5260 35888
rect 5300 35848 5301 35888
rect 5259 35839 5301 35848
rect 6747 35888 6789 35897
rect 6747 35848 6748 35888
rect 6788 35848 6789 35888
rect 6747 35839 6789 35848
rect 4107 35804 4149 35813
rect 4107 35764 4108 35804
rect 4148 35764 4149 35804
rect 4107 35755 4149 35764
rect 8811 35804 8853 35813
rect 8811 35764 8812 35804
rect 8852 35764 8853 35804
rect 8811 35755 8853 35764
rect 1152 35552 10656 35576
rect 1152 35512 3688 35552
rect 3728 35512 3770 35552
rect 3810 35512 3852 35552
rect 3892 35512 3934 35552
rect 3974 35512 4016 35552
rect 4056 35512 10656 35552
rect 1152 35488 10656 35512
rect 1467 35384 1509 35393
rect 1467 35344 1468 35384
rect 1508 35344 1509 35384
rect 1467 35335 1509 35344
rect 3051 35384 3093 35393
rect 3051 35344 3052 35384
rect 3092 35344 3093 35384
rect 3051 35335 3093 35344
rect 5451 35384 5493 35393
rect 5451 35344 5452 35384
rect 5492 35344 5493 35384
rect 5451 35335 5493 35344
rect 5883 35300 5925 35309
rect 5883 35260 5884 35300
rect 5924 35260 5925 35300
rect 5883 35251 5925 35260
rect 1227 35216 1269 35225
rect 1227 35176 1228 35216
rect 1268 35176 1269 35216
rect 1227 35167 1269 35176
rect 5643 35216 5685 35225
rect 5643 35176 5644 35216
rect 5684 35176 5685 35216
rect 5643 35167 5685 35176
rect 6027 35216 6069 35225
rect 6027 35176 6028 35216
rect 6068 35176 6069 35216
rect 6027 35167 6069 35176
rect 6267 35216 6309 35225
rect 6267 35176 6268 35216
rect 6308 35176 6309 35216
rect 6267 35167 6309 35176
rect 10347 35216 10389 35225
rect 10347 35176 10348 35216
rect 10388 35176 10389 35216
rect 10347 35167 10389 35176
rect 1611 35132 1653 35141
rect 1611 35092 1612 35132
rect 1652 35092 1653 35132
rect 1611 35083 1653 35092
rect 2851 35132 2909 35133
rect 2851 35092 2860 35132
rect 2900 35092 2909 35132
rect 2851 35091 2909 35092
rect 3178 35132 3236 35133
rect 3178 35092 3187 35132
rect 3227 35092 3236 35132
rect 3178 35091 3236 35092
rect 4011 35132 4053 35141
rect 4011 35092 4012 35132
rect 4052 35092 4053 35132
rect 4011 35083 4053 35092
rect 5251 35132 5309 35133
rect 5251 35092 5260 35132
rect 5300 35092 5309 35132
rect 5251 35091 5309 35092
rect 6411 35132 6453 35141
rect 6411 35092 6412 35132
rect 6452 35092 6453 35132
rect 6411 35083 6453 35092
rect 7651 35132 7709 35133
rect 7651 35092 7660 35132
rect 7700 35092 7709 35132
rect 7651 35091 7709 35092
rect 8527 35132 8585 35133
rect 8527 35092 8536 35132
rect 8576 35092 8585 35132
rect 8527 35091 8585 35092
rect 8715 35132 8757 35141
rect 8715 35092 8716 35132
rect 8756 35092 8757 35132
rect 8715 35083 8757 35092
rect 9955 35132 10013 35133
rect 9955 35092 9964 35132
rect 10004 35092 10013 35132
rect 9955 35091 10013 35092
rect 8362 35048 8420 35049
rect 8362 35008 8371 35048
rect 8411 35008 8420 35048
rect 8362 35007 8420 35008
rect 3387 34964 3429 34973
rect 3387 34924 3388 34964
rect 3428 34924 3429 34964
rect 3387 34915 3429 34924
rect 3802 34964 3860 34965
rect 3802 34924 3811 34964
rect 3851 34924 3860 34964
rect 3802 34923 3860 34924
rect 7851 34964 7893 34973
rect 7851 34924 7852 34964
rect 7892 34924 7893 34964
rect 7851 34915 7893 34924
rect 10155 34964 10197 34973
rect 10155 34924 10156 34964
rect 10196 34924 10197 34964
rect 10155 34915 10197 34924
rect 10587 34964 10629 34973
rect 10587 34924 10588 34964
rect 10628 34924 10629 34964
rect 10587 34915 10629 34924
rect 1152 34796 10656 34820
rect 1152 34756 4928 34796
rect 4968 34756 5010 34796
rect 5050 34756 5092 34796
rect 5132 34756 5174 34796
rect 5214 34756 5256 34796
rect 5296 34756 10656 34796
rect 1152 34732 10656 34756
rect 7515 34628 7557 34637
rect 7515 34588 7516 34628
rect 7556 34588 7557 34628
rect 7515 34579 7557 34588
rect 10522 34628 10580 34629
rect 10522 34588 10531 34628
rect 10571 34588 10580 34628
rect 10522 34587 10580 34588
rect 7371 34544 7413 34553
rect 7371 34504 7372 34544
rect 7412 34504 7413 34544
rect 7371 34495 7413 34504
rect 1995 34460 2037 34469
rect 3915 34460 3957 34469
rect 5931 34460 5973 34469
rect 8026 34460 8084 34461
rect 1218 34451 1264 34460
rect 1218 34411 1219 34451
rect 1259 34411 1264 34451
rect 1995 34420 1996 34460
rect 2036 34420 2037 34460
rect 1995 34411 2037 34420
rect 3243 34451 3285 34460
rect 3243 34411 3244 34451
rect 3284 34411 3285 34451
rect 3915 34420 3916 34460
rect 3956 34420 3957 34460
rect 3915 34411 3957 34420
rect 5163 34451 5205 34460
rect 5163 34411 5164 34451
rect 5204 34411 5205 34451
rect 5931 34420 5932 34460
rect 5972 34420 5973 34460
rect 5931 34411 5973 34420
rect 7179 34451 7221 34460
rect 7179 34411 7180 34451
rect 7220 34411 7221 34451
rect 8026 34420 8035 34460
rect 8075 34420 8084 34460
rect 8026 34419 8084 34420
rect 8139 34460 8181 34469
rect 8139 34420 8140 34460
rect 8180 34420 8181 34460
rect 8139 34411 8181 34420
rect 8523 34460 8565 34469
rect 9802 34460 9860 34461
rect 8523 34420 8524 34460
rect 8564 34420 8565 34460
rect 8523 34411 8565 34420
rect 9099 34451 9141 34460
rect 9099 34411 9100 34451
rect 9140 34411 9141 34451
rect 1218 34402 1264 34411
rect 3243 34402 3285 34411
rect 5163 34402 5205 34411
rect 7179 34402 7221 34411
rect 9099 34402 9141 34411
rect 9579 34451 9621 34460
rect 9579 34411 9580 34451
rect 9620 34411 9621 34451
rect 9802 34420 9811 34460
rect 9851 34420 9860 34460
rect 9802 34419 9860 34420
rect 9954 34451 10000 34460
rect 9579 34402 9621 34411
rect 9954 34411 9955 34451
rect 9995 34411 10000 34451
rect 9954 34402 10000 34411
rect 1371 34376 1413 34385
rect 1371 34336 1372 34376
rect 1412 34336 1413 34376
rect 1371 34327 1413 34336
rect 1803 34376 1845 34385
rect 1803 34336 1804 34376
rect 1844 34336 1845 34376
rect 1803 34327 1845 34336
rect 3627 34376 3669 34385
rect 3627 34336 3628 34376
rect 3668 34336 3669 34376
rect 3627 34327 3669 34336
rect 5547 34376 5589 34385
rect 5547 34336 5548 34376
rect 5588 34336 5589 34376
rect 5547 34327 5589 34336
rect 7755 34376 7797 34385
rect 7755 34336 7756 34376
rect 7796 34336 7797 34376
rect 7755 34327 7797 34336
rect 8619 34376 8661 34385
rect 8619 34336 8620 34376
rect 8660 34336 8661 34376
rect 8619 34327 8661 34336
rect 10107 34376 10149 34385
rect 10107 34336 10108 34376
rect 10148 34336 10149 34376
rect 10107 34327 10149 34336
rect 3435 34208 3477 34217
rect 3435 34168 3436 34208
rect 3476 34168 3477 34208
rect 3435 34159 3477 34168
rect 5355 34208 5397 34217
rect 5355 34168 5356 34208
rect 5396 34168 5397 34208
rect 5355 34159 5397 34168
rect 5787 34208 5829 34217
rect 5787 34168 5788 34208
rect 5828 34168 5829 34208
rect 5787 34159 5829 34168
rect 1152 34040 10656 34064
rect 1152 34000 3688 34040
rect 3728 34000 3770 34040
rect 3810 34000 3852 34040
rect 3892 34000 3934 34040
rect 3974 34000 4016 34040
rect 4056 34000 10656 34040
rect 1152 33976 10656 34000
rect 3963 33704 4005 33713
rect 3963 33664 3964 33704
rect 4004 33664 4005 33704
rect 3963 33655 4005 33664
rect 4443 33704 4485 33713
rect 4443 33664 4444 33704
rect 4484 33664 4485 33704
rect 4443 33655 4485 33664
rect 6411 33704 6453 33713
rect 6411 33664 6412 33704
rect 6452 33664 6453 33704
rect 6411 33655 6453 33664
rect 6747 33704 6789 33713
rect 6747 33664 6748 33704
rect 6788 33664 6789 33704
rect 6747 33655 6789 33664
rect 6987 33704 7029 33713
rect 6987 33664 6988 33704
rect 7028 33664 7029 33704
rect 6987 33655 7029 33664
rect 7179 33704 7221 33713
rect 7179 33664 7180 33704
rect 7220 33664 7221 33704
rect 7179 33655 7221 33664
rect 7851 33704 7893 33713
rect 7851 33664 7852 33704
rect 7892 33664 7893 33704
rect 7851 33655 7893 33664
rect 8715 33704 8757 33713
rect 8715 33664 8716 33704
rect 8756 33664 8757 33704
rect 8715 33655 8757 33664
rect 1162 33620 1220 33621
rect 1162 33580 1171 33620
rect 1211 33580 1220 33620
rect 1162 33579 1220 33580
rect 1707 33620 1749 33629
rect 1707 33580 1708 33620
rect 1748 33580 1749 33620
rect 1707 33571 1749 33580
rect 2947 33620 3005 33621
rect 2947 33580 2956 33620
rect 2996 33580 3005 33620
rect 2947 33579 3005 33580
rect 3319 33620 3377 33621
rect 3319 33580 3328 33620
rect 3368 33580 3377 33620
rect 3319 33579 3377 33580
rect 3769 33620 3827 33621
rect 3769 33580 3778 33620
rect 3818 33580 3827 33620
rect 3769 33579 3827 33580
rect 4279 33620 4337 33621
rect 4279 33580 4288 33620
rect 4328 33580 4337 33620
rect 4279 33579 4337 33580
rect 4779 33620 4821 33629
rect 4779 33580 4780 33620
rect 4820 33580 4821 33620
rect 4779 33571 4821 33580
rect 6019 33620 6077 33621
rect 6019 33580 6028 33620
rect 6068 33580 6077 33620
rect 6019 33579 6077 33580
rect 7467 33620 7509 33629
rect 7467 33580 7468 33620
rect 7508 33580 7509 33620
rect 7467 33571 7509 33580
rect 8218 33620 8276 33621
rect 8218 33580 8227 33620
rect 8267 33580 8276 33620
rect 8218 33579 8276 33580
rect 8331 33620 8373 33629
rect 8331 33580 8332 33620
rect 8372 33580 8373 33620
rect 8331 33571 8373 33580
rect 8811 33620 8853 33629
rect 8811 33580 8812 33620
rect 8852 33580 8853 33620
rect 8811 33571 8853 33580
rect 9283 33620 9341 33621
rect 9283 33580 9292 33620
rect 9332 33580 9341 33620
rect 9283 33579 9341 33580
rect 9802 33620 9860 33621
rect 9802 33580 9811 33620
rect 9851 33580 9860 33620
rect 9802 33579 9860 33580
rect 10090 33620 10148 33621
rect 10090 33580 10099 33620
rect 10139 33580 10148 33620
rect 10090 33579 10148 33580
rect 6651 33536 6693 33545
rect 6651 33496 6652 33536
rect 6692 33496 6693 33536
rect 6651 33487 6693 33496
rect 1371 33452 1413 33461
rect 1371 33412 1372 33452
rect 1412 33412 1413 33452
rect 1371 33403 1413 33412
rect 3147 33452 3189 33461
rect 3147 33412 3148 33452
rect 3188 33412 3189 33452
rect 3147 33403 3189 33412
rect 3483 33452 3525 33461
rect 3483 33412 3484 33452
rect 3524 33412 3525 33452
rect 3483 33403 3525 33412
rect 6219 33452 6261 33461
rect 6219 33412 6220 33452
rect 6260 33412 6261 33452
rect 6219 33403 6261 33412
rect 7258 33452 7316 33453
rect 7258 33412 7267 33452
rect 7307 33412 7316 33452
rect 7258 33411 7316 33412
rect 9963 33452 10005 33461
rect 9963 33412 9964 33452
rect 10004 33412 10005 33452
rect 9963 33403 10005 33412
rect 10299 33452 10341 33461
rect 10299 33412 10300 33452
rect 10340 33412 10341 33452
rect 10299 33403 10341 33412
rect 1152 33284 10656 33308
rect 1152 33244 4928 33284
rect 4968 33244 5010 33284
rect 5050 33244 5092 33284
rect 5132 33244 5174 33284
rect 5214 33244 5256 33284
rect 5296 33244 10656 33284
rect 1152 33220 10656 33244
rect 1515 33116 1557 33125
rect 1515 33076 1516 33116
rect 1556 33076 1557 33116
rect 1515 33067 1557 33076
rect 5451 33116 5493 33125
rect 5451 33076 5452 33116
rect 5492 33076 5493 33116
rect 5451 33067 5493 33076
rect 9771 33116 9813 33125
rect 9771 33076 9772 33116
rect 9812 33076 9813 33116
rect 9771 33067 9813 33076
rect 10522 33116 10580 33117
rect 10522 33076 10531 33116
rect 10571 33076 10580 33116
rect 10522 33075 10580 33076
rect 7755 33032 7797 33041
rect 7755 32992 7756 33032
rect 7796 32992 7797 33032
rect 7755 32983 7797 32992
rect 1306 32948 1364 32949
rect 1306 32908 1315 32948
rect 1355 32908 1364 32948
rect 1306 32907 1364 32908
rect 1995 32948 2037 32957
rect 3706 32948 3764 32949
rect 1995 32908 1996 32948
rect 2036 32908 2037 32948
rect 1995 32899 2037 32908
rect 3243 32939 3285 32948
rect 3243 32899 3244 32939
rect 3284 32899 3285 32939
rect 3706 32908 3715 32948
rect 3755 32908 3764 32948
rect 3706 32907 3764 32908
rect 3819 32948 3861 32957
rect 3819 32908 3820 32948
rect 3860 32908 3861 32948
rect 3819 32899 3861 32908
rect 4203 32948 4245 32957
rect 6315 32948 6357 32957
rect 8026 32948 8084 32949
rect 4203 32908 4204 32948
rect 4244 32908 4245 32948
rect 4203 32899 4245 32908
rect 4779 32939 4821 32948
rect 4779 32899 4780 32939
rect 4820 32899 4821 32939
rect 3243 32890 3285 32899
rect 4779 32890 4821 32899
rect 5259 32939 5301 32948
rect 5259 32899 5260 32939
rect 5300 32899 5301 32939
rect 5259 32890 5301 32899
rect 5634 32939 5680 32948
rect 5634 32899 5635 32939
rect 5675 32899 5680 32939
rect 6315 32908 6316 32948
rect 6356 32908 6357 32948
rect 6315 32899 6357 32908
rect 7563 32939 7605 32948
rect 7563 32899 7564 32939
rect 7604 32899 7605 32939
rect 8026 32908 8035 32948
rect 8075 32908 8084 32948
rect 8026 32907 8084 32908
rect 8139 32948 8181 32957
rect 8139 32908 8140 32948
rect 8180 32908 8181 32948
rect 8139 32899 8181 32908
rect 8527 32948 8569 32957
rect 8527 32908 8528 32948
rect 8568 32908 8569 32948
rect 8527 32899 8569 32908
rect 9099 32939 9141 32948
rect 9099 32899 9100 32939
rect 9140 32899 9141 32939
rect 5634 32890 5680 32899
rect 7563 32890 7605 32899
rect 9099 32890 9141 32899
rect 9579 32939 9621 32948
rect 9579 32899 9580 32939
rect 9620 32899 9621 32939
rect 9579 32890 9621 32899
rect 9954 32939 10000 32948
rect 9954 32899 9955 32939
rect 9995 32899 10000 32939
rect 9954 32890 10000 32899
rect 4299 32864 4341 32873
rect 4299 32824 4300 32864
rect 4340 32824 4341 32864
rect 4299 32815 4341 32824
rect 5787 32864 5829 32873
rect 5787 32824 5788 32864
rect 5828 32824 5829 32864
rect 5787 32815 5829 32824
rect 8619 32864 8661 32873
rect 8619 32824 8620 32864
rect 8660 32824 8661 32864
rect 8619 32815 8661 32824
rect 10107 32864 10149 32873
rect 10107 32824 10108 32864
rect 10148 32824 10149 32864
rect 10107 32815 10149 32824
rect 1515 32696 1557 32705
rect 1515 32656 1516 32696
rect 1556 32656 1557 32696
rect 1515 32647 1557 32656
rect 3435 32696 3477 32705
rect 3435 32656 3436 32696
rect 3476 32656 3477 32696
rect 3435 32647 3477 32656
rect 1152 32528 10656 32552
rect 1152 32488 3688 32528
rect 3728 32488 3770 32528
rect 3810 32488 3852 32528
rect 3892 32488 3934 32528
rect 3974 32488 4016 32528
rect 4056 32488 10656 32528
rect 1152 32464 10656 32488
rect 7851 32360 7893 32369
rect 7851 32320 7852 32360
rect 7892 32320 7893 32360
rect 7851 32311 7893 32320
rect 9819 32276 9861 32285
rect 9819 32236 9820 32276
rect 9860 32236 9861 32276
rect 9819 32227 9861 32236
rect 3435 32192 3477 32201
rect 3435 32152 3436 32192
rect 3476 32152 3477 32192
rect 3435 32143 3477 32152
rect 8170 32192 8228 32193
rect 8170 32152 8179 32192
rect 8219 32152 8228 32192
rect 8170 32151 8228 32152
rect 9003 32192 9045 32201
rect 9003 32152 9004 32192
rect 9044 32152 9045 32192
rect 9003 32143 9045 32152
rect 9291 32192 9333 32201
rect 9291 32152 9292 32192
rect 9332 32152 9333 32192
rect 9291 32143 9333 32152
rect 9579 32192 9621 32201
rect 9579 32152 9580 32192
rect 9620 32152 9621 32192
rect 9579 32143 9621 32152
rect 9963 32192 10005 32201
rect 9963 32152 9964 32192
rect 10004 32152 10005 32192
rect 9963 32143 10005 32152
rect 10347 32192 10389 32201
rect 10347 32152 10348 32192
rect 10388 32152 10389 32192
rect 10347 32143 10389 32152
rect 1227 32108 1269 32117
rect 1227 32068 1228 32108
rect 1268 32068 1269 32108
rect 1227 32059 1269 32068
rect 2467 32108 2525 32109
rect 2467 32068 2476 32108
rect 2516 32068 2525 32108
rect 2467 32067 2525 32068
rect 2938 32108 2996 32109
rect 2938 32068 2947 32108
rect 2987 32068 2996 32108
rect 2938 32067 2996 32068
rect 3051 32108 3093 32117
rect 3051 32068 3052 32108
rect 3092 32068 3093 32108
rect 3051 32059 3093 32068
rect 3531 32108 3573 32117
rect 3531 32068 3532 32108
rect 3572 32068 3573 32108
rect 3531 32059 3573 32068
rect 4003 32108 4061 32109
rect 4003 32068 4012 32108
rect 4052 32068 4061 32108
rect 4003 32067 4061 32068
rect 4491 32108 4549 32109
rect 4491 32068 4500 32108
rect 4540 32068 4549 32108
rect 4491 32067 4549 32068
rect 4810 32108 4868 32109
rect 4810 32068 4819 32108
rect 4859 32068 4868 32108
rect 4810 32067 4868 32068
rect 5305 32108 5363 32109
rect 5305 32068 5314 32108
rect 5354 32068 5363 32108
rect 5305 32067 5363 32068
rect 5835 32108 5877 32117
rect 5835 32068 5836 32108
rect 5876 32068 5877 32108
rect 5835 32059 5877 32068
rect 6411 32108 6453 32117
rect 6411 32068 6412 32108
rect 6452 32068 6453 32108
rect 6411 32059 6453 32068
rect 7651 32108 7709 32109
rect 7651 32068 7660 32108
rect 7700 32068 7709 32108
rect 7651 32067 7709 32068
rect 8335 32108 8393 32109
rect 8335 32068 8344 32108
rect 8384 32068 8393 32108
rect 8335 32067 8393 32068
rect 8523 32108 8565 32117
rect 8523 32068 8524 32108
rect 8564 32068 8565 32108
rect 8523 32059 8565 32068
rect 2667 32024 2709 32033
rect 2667 31984 2668 32024
rect 2708 31984 2709 32024
rect 2667 31975 2709 31984
rect 10203 32024 10245 32033
rect 10203 31984 10204 32024
rect 10244 31984 10245 32024
rect 10203 31975 10245 31984
rect 4683 31940 4725 31949
rect 4683 31900 4684 31940
rect 4724 31900 4725 31940
rect 4683 31891 4725 31900
rect 5019 31940 5061 31949
rect 5019 31900 5020 31940
rect 5060 31900 5061 31940
rect 5019 31891 5061 31900
rect 5499 31940 5541 31949
rect 5499 31900 5500 31940
rect 5540 31900 5541 31940
rect 5499 31891 5541 31900
rect 6106 31940 6164 31941
rect 6106 31900 6115 31940
rect 6155 31900 6164 31940
rect 6106 31899 6164 31900
rect 9082 31940 9140 31941
rect 9082 31900 9091 31940
rect 9131 31900 9140 31940
rect 9082 31899 9140 31900
rect 10587 31940 10629 31949
rect 10587 31900 10588 31940
rect 10628 31900 10629 31940
rect 10587 31891 10629 31900
rect 1152 31772 10656 31796
rect 1152 31732 4928 31772
rect 4968 31732 5010 31772
rect 5050 31732 5092 31772
rect 5132 31732 5174 31772
rect 5214 31732 5256 31772
rect 5296 31732 10656 31772
rect 1152 31708 10656 31732
rect 2619 31604 2661 31613
rect 2619 31564 2620 31604
rect 2660 31564 2661 31604
rect 2619 31555 2661 31564
rect 3195 31604 3237 31613
rect 3195 31564 3196 31604
rect 3236 31564 3237 31604
rect 3195 31555 3237 31564
rect 5163 31604 5205 31613
rect 5163 31564 5164 31604
rect 5204 31564 5205 31604
rect 5163 31555 5205 31564
rect 7066 31604 7124 31605
rect 7066 31564 7075 31604
rect 7115 31564 7124 31604
rect 7066 31563 7124 31564
rect 8170 31604 8228 31605
rect 8170 31564 8179 31604
rect 8219 31564 8228 31604
rect 8170 31563 8228 31564
rect 6219 31520 6261 31529
rect 6219 31480 6220 31520
rect 6260 31480 6261 31520
rect 6219 31471 6261 31480
rect 7275 31520 7317 31529
rect 7275 31480 7276 31520
rect 7316 31480 7317 31520
rect 7275 31471 7317 31480
rect 7707 31520 7749 31529
rect 7707 31480 7708 31520
rect 7748 31480 7749 31520
rect 7707 31471 7749 31480
rect 1306 31436 1364 31437
rect 3418 31436 3476 31437
rect 1306 31396 1315 31436
rect 1355 31396 1364 31436
rect 1306 31395 1364 31396
rect 1986 31427 2032 31436
rect 1986 31387 1987 31427
rect 2027 31387 2032 31427
rect 1986 31378 2032 31387
rect 2466 31427 2512 31436
rect 2466 31387 2467 31427
rect 2507 31387 2512 31427
rect 3418 31396 3427 31436
rect 3467 31396 3476 31436
rect 3418 31395 3476 31396
rect 3531 31436 3573 31445
rect 3531 31396 3532 31436
rect 3572 31396 3573 31436
rect 3531 31387 3573 31396
rect 3915 31436 3957 31445
rect 6507 31436 6549 31445
rect 8602 31436 8660 31437
rect 3915 31396 3916 31436
rect 3956 31396 3957 31436
rect 3915 31387 3957 31396
rect 4491 31427 4533 31436
rect 4491 31387 4492 31427
rect 4532 31387 4533 31427
rect 2466 31378 2512 31387
rect 4491 31378 4533 31387
rect 4971 31427 5013 31436
rect 4971 31387 4972 31427
rect 5012 31387 5013 31427
rect 4971 31378 5013 31387
rect 5346 31427 5392 31436
rect 5346 31387 5347 31427
rect 5387 31387 5392 31427
rect 6507 31396 6508 31436
rect 6548 31396 6549 31436
rect 6507 31387 6549 31396
rect 7554 31427 7600 31436
rect 7554 31387 7555 31427
rect 7595 31387 7600 31427
rect 8602 31396 8611 31436
rect 8651 31396 8660 31436
rect 8602 31395 8660 31396
rect 8715 31436 8757 31445
rect 8715 31396 8716 31436
rect 8756 31396 8757 31436
rect 5346 31378 5392 31387
rect 7554 31378 7600 31387
rect 8362 31394 8420 31395
rect 2139 31352 2181 31361
rect 2139 31312 2140 31352
rect 2180 31312 2181 31352
rect 2139 31303 2181 31312
rect 2955 31352 2997 31361
rect 2955 31312 2956 31352
rect 2996 31312 2997 31352
rect 2955 31303 2997 31312
rect 4011 31352 4053 31361
rect 4011 31312 4012 31352
rect 4052 31312 4053 31352
rect 4011 31303 4053 31312
rect 5499 31352 5541 31361
rect 5499 31312 5500 31352
rect 5540 31312 5541 31352
rect 5499 31303 5541 31312
rect 5835 31352 5877 31361
rect 8362 31354 8371 31394
rect 8411 31354 8420 31394
rect 8715 31387 8757 31396
rect 9099 31436 9141 31445
rect 9099 31396 9100 31436
rect 9140 31396 9141 31436
rect 9099 31387 9141 31396
rect 9675 31427 9717 31436
rect 9675 31387 9676 31427
rect 9716 31387 9717 31427
rect 9675 31378 9717 31387
rect 10155 31427 10197 31436
rect 10155 31387 10156 31427
rect 10196 31387 10197 31427
rect 10155 31378 10197 31387
rect 8362 31353 8420 31354
rect 5835 31312 5836 31352
rect 5876 31312 5877 31352
rect 5835 31303 5877 31312
rect 9195 31352 9237 31361
rect 9195 31312 9196 31352
rect 9236 31312 9237 31352
rect 9195 31303 9237 31312
rect 1515 31184 1557 31193
rect 1515 31144 1516 31184
rect 1556 31144 1557 31184
rect 1515 31135 1557 31144
rect 6075 31184 6117 31193
rect 6075 31144 6076 31184
rect 6116 31144 6117 31184
rect 6075 31135 6117 31144
rect 10378 31184 10436 31185
rect 10378 31144 10387 31184
rect 10427 31144 10436 31184
rect 10378 31143 10436 31144
rect 1152 31016 10656 31040
rect 1152 30976 3688 31016
rect 3728 30976 3770 31016
rect 3810 30976 3852 31016
rect 3892 30976 3934 31016
rect 3974 30976 4016 31016
rect 4056 30976 10656 31016
rect 1152 30952 10656 30976
rect 9291 30848 9333 30857
rect 9291 30808 9292 30848
rect 9332 30808 9333 30848
rect 9291 30799 9333 30808
rect 10395 30848 10437 30857
rect 10395 30808 10396 30848
rect 10436 30808 10437 30848
rect 10395 30799 10437 30808
rect 3867 30680 3909 30689
rect 3867 30640 3868 30680
rect 3908 30640 3909 30680
rect 3867 30631 3909 30640
rect 10155 30680 10197 30689
rect 10155 30640 10156 30680
rect 10196 30640 10197 30680
rect 9994 30638 10052 30639
rect 1419 30596 1461 30605
rect 1419 30556 1420 30596
rect 1460 30556 1461 30596
rect 1419 30547 1461 30556
rect 2659 30596 2717 30597
rect 2659 30556 2668 30596
rect 2708 30556 2717 30596
rect 2659 30555 2717 30556
rect 3339 30596 3381 30605
rect 3339 30556 3340 30596
rect 3380 30556 3381 30596
rect 3339 30547 3381 30556
rect 3458 30596 3500 30605
rect 3458 30556 3459 30596
rect 3499 30556 3500 30596
rect 3458 30547 3500 30556
rect 3568 30596 3626 30597
rect 3568 30556 3577 30596
rect 3617 30556 3626 30596
rect 3568 30555 3626 30556
rect 3703 30596 3761 30597
rect 3703 30556 3712 30596
rect 3752 30556 3761 30596
rect 3703 30555 3761 30556
rect 4203 30596 4245 30605
rect 4203 30556 4204 30596
rect 4244 30556 4245 30596
rect 4203 30547 4245 30556
rect 4395 30596 4437 30605
rect 4395 30556 4396 30596
rect 4436 30556 4437 30596
rect 4395 30547 4437 30556
rect 4587 30596 4629 30605
rect 4587 30556 4588 30596
rect 4628 30556 4629 30596
rect 4587 30547 4629 30556
rect 5827 30596 5885 30597
rect 5827 30556 5836 30596
rect 5876 30556 5885 30596
rect 5827 30555 5885 30556
rect 6219 30596 6261 30605
rect 6219 30556 6220 30596
rect 6260 30556 6261 30596
rect 6219 30547 6261 30556
rect 7459 30596 7517 30597
rect 7459 30556 7468 30596
rect 7508 30556 7517 30596
rect 7459 30555 7517 30556
rect 7851 30596 7893 30605
rect 9994 30598 10003 30638
rect 10043 30598 10052 30638
rect 10155 30631 10197 30640
rect 9994 30597 10052 30598
rect 7851 30556 7852 30596
rect 7892 30556 7893 30596
rect 7851 30547 7893 30556
rect 9091 30596 9149 30597
rect 9091 30556 9100 30596
rect 9140 30556 9149 30596
rect 9091 30555 9149 30556
rect 2859 30428 2901 30437
rect 2859 30388 2860 30428
rect 2900 30388 2901 30428
rect 2859 30379 2901 30388
rect 3243 30428 3285 30437
rect 3243 30388 3244 30428
rect 3284 30388 3285 30428
rect 3243 30379 3285 30388
rect 4299 30428 4341 30437
rect 4299 30388 4300 30428
rect 4340 30388 4341 30428
rect 4299 30379 4341 30388
rect 6027 30428 6069 30437
rect 6027 30388 6028 30428
rect 6068 30388 6069 30428
rect 6027 30379 6069 30388
rect 7659 30428 7701 30437
rect 7659 30388 7660 30428
rect 7700 30388 7701 30428
rect 7659 30379 7701 30388
rect 9802 30428 9860 30429
rect 9802 30388 9811 30428
rect 9851 30388 9860 30428
rect 9802 30387 9860 30388
rect 1152 30260 10656 30284
rect 1152 30220 4928 30260
rect 4968 30220 5010 30260
rect 5050 30220 5092 30260
rect 5132 30220 5174 30260
rect 5214 30220 5256 30260
rect 5296 30220 10656 30260
rect 1152 30196 10656 30220
rect 2667 30092 2709 30101
rect 2667 30052 2668 30092
rect 2708 30052 2709 30092
rect 2667 30043 2709 30052
rect 5211 30092 5253 30101
rect 5211 30052 5212 30092
rect 5252 30052 5253 30092
rect 4378 30050 4436 30051
rect 4378 30010 4387 30050
rect 4427 30010 4436 30050
rect 5211 30043 5253 30052
rect 7851 30092 7893 30101
rect 7851 30052 7852 30092
rect 7892 30052 7893 30092
rect 7851 30043 7893 30052
rect 10539 30092 10581 30101
rect 10539 30052 10540 30092
rect 10580 30052 10581 30092
rect 10539 30043 10581 30052
rect 4378 30009 4436 30010
rect 1227 29924 1269 29933
rect 3095 29924 3153 29925
rect 1227 29884 1228 29924
rect 1268 29884 1269 29924
rect 1227 29875 1269 29884
rect 2475 29915 2517 29924
rect 2475 29875 2476 29915
rect 2516 29875 2517 29915
rect 2475 29866 2517 29875
rect 2986 29906 3028 29915
rect 2986 29866 2987 29906
rect 3027 29866 3028 29906
rect 3095 29884 3104 29924
rect 3144 29884 3153 29924
rect 3095 29883 3153 29884
rect 3217 29924 3275 29925
rect 3217 29884 3226 29924
rect 3266 29884 3275 29924
rect 3217 29883 3275 29884
rect 3435 29924 3477 29933
rect 3435 29884 3436 29924
rect 3476 29884 3477 29924
rect 3435 29875 3477 29884
rect 3723 29924 3765 29933
rect 3723 29884 3724 29924
rect 3764 29884 3765 29924
rect 3723 29875 3765 29884
rect 4155 29924 4197 29933
rect 4155 29884 4156 29924
rect 4196 29884 4197 29924
rect 4155 29875 4197 29884
rect 4456 29924 4498 29933
rect 4456 29884 4457 29924
rect 4497 29884 4498 29924
rect 4456 29875 4498 29884
rect 4610 29924 4652 29933
rect 6106 29924 6164 29925
rect 4610 29884 4611 29924
rect 4651 29884 4652 29924
rect 4610 29875 4652 29884
rect 4770 29915 4816 29924
rect 4770 29875 4771 29915
rect 4811 29875 4816 29915
rect 6106 29884 6115 29924
rect 6155 29884 6164 29924
rect 6106 29883 6164 29884
rect 6224 29924 6266 29933
rect 6224 29884 6225 29924
rect 6265 29884 6266 29924
rect 6224 29875 6266 29884
rect 6603 29924 6645 29933
rect 9099 29924 9141 29933
rect 6603 29884 6604 29924
rect 6644 29884 6645 29924
rect 6603 29875 6645 29884
rect 7179 29915 7221 29924
rect 7179 29875 7180 29915
rect 7220 29875 7221 29915
rect 4770 29866 4816 29875
rect 7179 29866 7221 29875
rect 7659 29915 7701 29924
rect 7659 29875 7660 29915
rect 7700 29875 7701 29915
rect 7659 29866 7701 29875
rect 8034 29915 8080 29924
rect 8034 29875 8035 29915
rect 8075 29875 8080 29915
rect 9099 29884 9100 29924
rect 9140 29884 9141 29924
rect 9099 29875 9141 29884
rect 10347 29915 10389 29924
rect 10347 29875 10348 29915
rect 10388 29875 10389 29915
rect 8034 29866 8080 29875
rect 10347 29866 10389 29875
rect 2986 29857 3028 29866
rect 4299 29840 4341 29849
rect 4299 29800 4300 29840
rect 4340 29800 4341 29840
rect 4299 29791 4341 29800
rect 4923 29840 4965 29849
rect 4923 29800 4924 29840
rect 4964 29800 4965 29840
rect 4923 29791 4965 29800
rect 5451 29840 5493 29849
rect 5451 29800 5452 29840
rect 5492 29800 5493 29840
rect 5451 29791 5493 29800
rect 5835 29840 5877 29849
rect 5835 29800 5836 29840
rect 5876 29800 5877 29840
rect 5835 29791 5877 29800
rect 6699 29840 6741 29849
rect 6699 29800 6700 29840
rect 6740 29800 6741 29840
rect 6699 29791 6741 29800
rect 8187 29840 8229 29849
rect 8187 29800 8188 29840
rect 8228 29800 8229 29840
rect 8187 29791 8229 29800
rect 8715 29840 8757 29849
rect 8715 29800 8716 29840
rect 8756 29800 8757 29840
rect 8715 29791 8757 29800
rect 3147 29672 3189 29681
rect 3147 29632 3148 29672
rect 3188 29632 3189 29672
rect 3147 29623 3189 29632
rect 3915 29672 3957 29681
rect 3915 29632 3916 29672
rect 3956 29632 3957 29672
rect 3915 29623 3957 29632
rect 5595 29672 5637 29681
rect 5595 29632 5596 29672
rect 5636 29632 5637 29672
rect 5595 29623 5637 29632
rect 8955 29672 8997 29681
rect 8955 29632 8956 29672
rect 8996 29632 8997 29672
rect 8955 29623 8997 29632
rect 1152 29504 10656 29528
rect 1152 29464 3688 29504
rect 3728 29464 3770 29504
rect 3810 29464 3852 29504
rect 3892 29464 3934 29504
rect 3974 29464 4016 29504
rect 4056 29464 10656 29504
rect 1152 29440 10656 29464
rect 3130 29336 3188 29337
rect 3130 29296 3139 29336
rect 3179 29296 3188 29336
rect 3130 29295 3188 29296
rect 4203 29336 4245 29345
rect 4203 29296 4204 29336
rect 4244 29296 4245 29336
rect 4203 29287 4245 29296
rect 2410 29168 2468 29169
rect 2410 29128 2419 29168
rect 2459 29128 2468 29168
rect 2410 29127 2468 29128
rect 2763 29168 2805 29177
rect 2763 29128 2764 29168
rect 2804 29128 2805 29168
rect 2763 29119 2805 29128
rect 5163 29168 5205 29177
rect 5163 29128 5164 29168
rect 5204 29128 5205 29168
rect 5163 29119 5205 29128
rect 7083 29168 7125 29177
rect 7083 29128 7084 29168
rect 7124 29128 7125 29168
rect 7083 29119 7125 29128
rect 9291 29168 9333 29177
rect 9291 29128 9292 29168
rect 9332 29128 9333 29168
rect 9291 29119 9333 29128
rect 10347 29168 10389 29177
rect 10347 29128 10348 29168
rect 10388 29128 10389 29168
rect 10347 29119 10389 29128
rect 1162 29084 1220 29085
rect 1162 29044 1171 29084
rect 1211 29044 1220 29084
rect 1162 29043 1220 29044
rect 1657 29084 1715 29085
rect 1657 29044 1666 29084
rect 1706 29044 1715 29084
rect 1657 29043 1715 29044
rect 2575 29084 2633 29085
rect 2575 29044 2584 29084
rect 2624 29044 2633 29084
rect 2575 29043 2633 29044
rect 3130 29084 3188 29085
rect 3130 29044 3139 29084
rect 3179 29044 3188 29084
rect 3130 29043 3188 29044
rect 3248 29084 3306 29085
rect 3248 29044 3257 29084
rect 3297 29044 3306 29084
rect 3248 29043 3306 29044
rect 3380 29084 3438 29085
rect 3380 29044 3389 29084
rect 3429 29044 3438 29084
rect 3380 29043 3438 29044
rect 3514 29084 3572 29085
rect 3514 29044 3523 29084
rect 3563 29044 3572 29084
rect 3514 29043 3572 29044
rect 3691 29084 3749 29085
rect 3691 29044 3700 29084
rect 3740 29044 3749 29084
rect 3691 29043 3749 29044
rect 3898 29084 3956 29085
rect 3898 29044 3907 29084
rect 3947 29044 3956 29084
rect 3898 29043 3956 29044
rect 4203 29084 4245 29093
rect 4203 29044 4204 29084
rect 4244 29044 4245 29084
rect 4203 29035 4245 29044
rect 4666 29084 4724 29085
rect 4666 29044 4675 29084
rect 4715 29044 4724 29084
rect 4666 29043 4724 29044
rect 4779 29084 4821 29093
rect 4779 29044 4780 29084
rect 4820 29044 4821 29084
rect 4779 29035 4821 29044
rect 5259 29084 5301 29093
rect 5259 29044 5260 29084
rect 5300 29044 5301 29084
rect 5259 29035 5301 29044
rect 5731 29084 5789 29085
rect 5731 29044 5740 29084
rect 5780 29044 5789 29084
rect 5731 29043 5789 29044
rect 6219 29084 6277 29085
rect 6219 29044 6228 29084
rect 6268 29044 6277 29084
rect 6219 29043 6277 29044
rect 6442 29084 6500 29085
rect 6442 29044 6451 29084
rect 6491 29044 6500 29084
rect 6442 29043 6500 29044
rect 6538 29084 6596 29085
rect 6538 29044 6547 29084
rect 6587 29044 6596 29084
rect 6538 29043 6596 29044
rect 7563 29084 7605 29093
rect 7563 29044 7564 29084
rect 7604 29044 7605 29084
rect 7563 29035 7605 29044
rect 8803 29084 8861 29085
rect 8803 29044 8812 29084
rect 8852 29044 8861 29084
rect 8803 29043 8861 29044
rect 9997 29084 10055 29085
rect 9997 29044 10006 29084
rect 10046 29044 10055 29084
rect 9997 29043 10055 29044
rect 1851 29000 1893 29009
rect 1851 28960 1852 29000
rect 1892 28960 1893 29000
rect 1851 28951 1893 28960
rect 3003 29000 3045 29009
rect 3003 28960 3004 29000
rect 3044 28960 3045 29000
rect 3003 28951 3045 28960
rect 1371 28916 1413 28925
rect 1371 28876 1372 28916
rect 1412 28876 1413 28916
rect 1371 28867 1413 28876
rect 6747 28916 6789 28925
rect 6747 28876 6748 28916
rect 6788 28876 6789 28916
rect 6747 28867 6789 28876
rect 7066 28916 7124 28917
rect 7066 28876 7075 28916
rect 7115 28876 7124 28916
rect 7066 28875 7124 28876
rect 9003 28916 9045 28925
rect 9003 28876 9004 28916
rect 9044 28876 9045 28916
rect 9003 28867 9045 28876
rect 9531 28916 9573 28925
rect 9531 28876 9532 28916
rect 9572 28876 9573 28916
rect 9531 28867 9573 28876
rect 9802 28916 9860 28917
rect 9802 28876 9811 28916
rect 9851 28876 9860 28916
rect 9802 28875 9860 28876
rect 10587 28916 10629 28925
rect 10587 28876 10588 28916
rect 10628 28876 10629 28916
rect 10587 28867 10629 28876
rect 1152 28748 10656 28772
rect 1152 28708 4928 28748
rect 4968 28708 5010 28748
rect 5050 28708 5092 28748
rect 5132 28708 5174 28748
rect 5214 28708 5256 28748
rect 5296 28708 10656 28748
rect 1152 28684 10656 28708
rect 2859 28580 2901 28589
rect 2859 28540 2860 28580
rect 2900 28540 2901 28580
rect 2859 28531 2901 28540
rect 3723 28580 3765 28589
rect 3723 28540 3724 28580
rect 3764 28540 3765 28580
rect 3723 28531 3765 28540
rect 6219 28580 6261 28589
rect 6219 28540 6220 28580
rect 6260 28540 6261 28580
rect 6219 28531 6261 28540
rect 6874 28580 6932 28581
rect 6874 28540 6883 28580
rect 6923 28540 6932 28580
rect 6874 28539 6932 28540
rect 7162 28580 7220 28581
rect 7162 28540 7171 28580
rect 7211 28540 7220 28580
rect 7162 28539 7220 28540
rect 7546 28580 7604 28581
rect 7546 28540 7555 28580
rect 7595 28540 7604 28580
rect 7546 28539 7604 28540
rect 7930 28580 7988 28581
rect 7930 28540 7939 28580
rect 7979 28540 7988 28580
rect 7930 28539 7988 28540
rect 10251 28580 10293 28589
rect 10251 28540 10252 28580
rect 10292 28540 10293 28580
rect 10251 28531 10293 28540
rect 10522 28580 10580 28581
rect 10522 28540 10531 28580
rect 10571 28540 10580 28580
rect 10522 28539 10580 28540
rect 3178 28496 3236 28497
rect 3178 28456 3187 28496
rect 3227 28456 3236 28496
rect 3178 28455 3236 28456
rect 3627 28496 3669 28505
rect 3627 28456 3628 28496
rect 3668 28456 3669 28496
rect 3627 28447 3669 28456
rect 3833 28496 3875 28505
rect 3833 28456 3834 28496
rect 3874 28456 3875 28496
rect 3833 28447 3875 28456
rect 4107 28496 4149 28505
rect 4107 28456 4108 28496
rect 4148 28456 4149 28496
rect 4107 28447 4149 28456
rect 10443 28496 10485 28505
rect 10443 28456 10444 28496
rect 10484 28456 10485 28496
rect 10443 28447 10485 28456
rect 1419 28412 1461 28421
rect 3343 28412 3401 28413
rect 1419 28372 1420 28412
rect 1460 28372 1461 28412
rect 1419 28363 1461 28372
rect 2667 28403 2709 28412
rect 2667 28363 2668 28403
rect 2708 28363 2709 28403
rect 3343 28372 3352 28412
rect 3392 28372 3401 28412
rect 3343 28371 3401 28372
rect 3514 28412 3572 28413
rect 3514 28372 3523 28412
rect 3563 28372 3572 28412
rect 3514 28371 3572 28372
rect 4011 28412 4053 28421
rect 4011 28372 4012 28412
rect 4052 28372 4053 28412
rect 4011 28363 4053 28372
rect 4186 28412 4244 28413
rect 4186 28372 4195 28412
rect 4235 28372 4244 28412
rect 4186 28371 4244 28372
rect 4474 28412 4532 28413
rect 4474 28372 4483 28412
rect 4523 28372 4532 28412
rect 4474 28371 4532 28372
rect 4587 28412 4629 28421
rect 4587 28372 4588 28412
rect 4628 28372 4629 28412
rect 4587 28363 4629 28372
rect 4971 28412 5013 28421
rect 8506 28412 8564 28413
rect 4971 28372 4972 28412
rect 5012 28372 5013 28412
rect 4971 28363 5013 28372
rect 5547 28403 5589 28412
rect 5547 28363 5548 28403
rect 5588 28363 5589 28403
rect 2667 28354 2709 28363
rect 5547 28354 5589 28363
rect 6027 28403 6069 28412
rect 6027 28363 6028 28403
rect 6068 28363 6069 28403
rect 6027 28354 6069 28363
rect 6402 28403 6448 28412
rect 6402 28363 6403 28403
rect 6443 28363 6448 28403
rect 8506 28372 8515 28412
rect 8555 28372 8564 28412
rect 8506 28371 8564 28372
rect 8619 28412 8661 28421
rect 8619 28372 8620 28412
rect 8660 28372 8661 28412
rect 8619 28363 8661 28372
rect 9003 28412 9045 28421
rect 9003 28372 9004 28412
rect 9044 28372 9045 28412
rect 9003 28363 9045 28372
rect 9579 28403 9621 28412
rect 9579 28363 9580 28403
rect 9620 28363 9621 28403
rect 6402 28354 6448 28363
rect 9579 28354 9621 28363
rect 10059 28403 10101 28412
rect 10059 28363 10060 28403
rect 10100 28363 10101 28403
rect 10059 28354 10101 28363
rect 5067 28328 5109 28337
rect 5067 28288 5068 28328
rect 5108 28288 5109 28328
rect 5067 28279 5109 28288
rect 6555 28328 6597 28337
rect 6555 28288 6556 28328
rect 6596 28288 6597 28328
rect 6555 28279 6597 28288
rect 7851 28328 7893 28337
rect 7851 28288 7852 28328
rect 7892 28288 7893 28328
rect 7851 28279 7893 28288
rect 8139 28328 8181 28337
rect 8139 28288 8140 28328
rect 8180 28288 8181 28328
rect 8139 28279 8181 28288
rect 9099 28328 9141 28337
rect 9099 28288 9100 28328
rect 9140 28288 9141 28328
rect 9099 28279 9141 28288
rect 1152 27992 10656 28016
rect 1152 27952 3688 27992
rect 3728 27952 3770 27992
rect 3810 27952 3852 27992
rect 3892 27952 3934 27992
rect 3974 27952 4016 27992
rect 4056 27952 10656 27992
rect 1152 27928 10656 27952
rect 3915 27824 3957 27833
rect 3915 27784 3916 27824
rect 3956 27784 3957 27824
rect 3915 27775 3957 27784
rect 5931 27824 5973 27833
rect 5931 27784 5932 27824
rect 5972 27784 5973 27824
rect 5931 27775 5973 27784
rect 10347 27824 10389 27833
rect 10347 27784 10348 27824
rect 10388 27784 10389 27824
rect 10347 27775 10389 27784
rect 4347 27740 4389 27749
rect 4347 27700 4348 27740
rect 4388 27700 4389 27740
rect 4347 27691 4389 27700
rect 2122 27656 2180 27657
rect 2122 27616 2131 27656
rect 2171 27616 2180 27656
rect 2122 27615 2180 27616
rect 4107 27656 4149 27665
rect 4107 27616 4108 27656
rect 4148 27616 4149 27656
rect 4107 27607 4149 27616
rect 8139 27656 8181 27665
rect 8139 27616 8140 27656
rect 8180 27616 8181 27656
rect 8139 27607 8181 27616
rect 1162 27572 1220 27573
rect 1162 27532 1171 27572
rect 1211 27532 1220 27572
rect 1162 27531 1220 27532
rect 2317 27572 2375 27573
rect 2317 27532 2326 27572
rect 2366 27532 2375 27572
rect 2317 27531 2375 27532
rect 2475 27572 2517 27581
rect 2475 27532 2476 27572
rect 2516 27532 2517 27572
rect 2475 27523 2517 27532
rect 3715 27572 3773 27573
rect 3715 27532 3724 27572
rect 3764 27532 3773 27572
rect 3715 27531 3773 27532
rect 4491 27572 4533 27581
rect 4491 27532 4492 27572
rect 4532 27532 4533 27572
rect 4491 27523 4533 27532
rect 5731 27572 5789 27573
rect 5731 27532 5740 27572
rect 5780 27532 5789 27572
rect 5731 27531 5789 27532
rect 6219 27572 6261 27581
rect 6219 27532 6220 27572
rect 6260 27532 6261 27572
rect 6219 27523 6261 27532
rect 7459 27572 7517 27573
rect 7459 27532 7468 27572
rect 7508 27532 7517 27572
rect 7459 27531 7517 27532
rect 8362 27572 8420 27573
rect 8362 27532 8371 27572
rect 8411 27532 8420 27572
rect 8362 27531 8420 27532
rect 8907 27572 8949 27581
rect 8907 27532 8908 27572
rect 8948 27532 8949 27572
rect 8907 27523 8949 27532
rect 10147 27572 10205 27573
rect 10147 27532 10156 27572
rect 10196 27532 10205 27572
rect 10147 27531 10205 27532
rect 7659 27488 7701 27497
rect 7659 27448 7660 27488
rect 7700 27448 7701 27488
rect 7659 27439 7701 27448
rect 1371 27404 1413 27413
rect 1371 27364 1372 27404
rect 1412 27364 1413 27404
rect 1371 27355 1413 27364
rect 1786 27404 1844 27405
rect 1786 27364 1795 27404
rect 1835 27364 1844 27404
rect 1786 27363 1844 27364
rect 7930 27404 7988 27405
rect 7930 27364 7939 27404
rect 7979 27364 7988 27404
rect 7930 27363 7988 27364
rect 8218 27404 8276 27405
rect 8218 27364 8227 27404
rect 8267 27364 8276 27404
rect 8218 27363 8276 27364
rect 8571 27404 8613 27413
rect 8571 27364 8572 27404
rect 8612 27364 8613 27404
rect 8571 27355 8613 27364
rect 1152 27236 10656 27260
rect 1152 27196 4928 27236
rect 4968 27196 5010 27236
rect 5050 27196 5092 27236
rect 5132 27196 5174 27236
rect 5214 27196 5256 27236
rect 5296 27196 10656 27236
rect 1152 27172 10656 27196
rect 1707 27068 1749 27077
rect 1707 27028 1708 27068
rect 1748 27028 1749 27068
rect 1707 27019 1749 27028
rect 2139 27068 2181 27077
rect 2139 27028 2140 27068
rect 2180 27028 2181 27068
rect 2139 27019 2181 27028
rect 3099 27068 3141 27077
rect 3099 27028 3100 27068
rect 3140 27028 3141 27068
rect 3099 27019 3141 27028
rect 4683 27068 4725 27077
rect 4683 27028 4684 27068
rect 4724 27028 4725 27068
rect 4683 27019 4725 27028
rect 8331 27068 8373 27077
rect 8331 27028 8332 27068
rect 8372 27028 8373 27068
rect 8331 27019 8373 27028
rect 2619 26984 2661 26993
rect 2619 26944 2620 26984
rect 2660 26944 2661 26984
rect 2619 26935 2661 26944
rect 6315 26984 6357 26993
rect 6315 26944 6316 26984
rect 6356 26944 6357 26984
rect 6315 26935 6357 26944
rect 2955 26900 2997 26909
rect 1218 26891 1264 26900
rect 1218 26851 1219 26891
rect 1259 26851 1264 26891
rect 1218 26842 1264 26851
rect 1986 26891 2032 26900
rect 1986 26851 1987 26891
rect 2027 26851 2032 26891
rect 1986 26842 2032 26851
rect 2466 26891 2512 26900
rect 2466 26851 2467 26891
rect 2507 26851 2512 26891
rect 2955 26860 2956 26900
rect 2996 26860 2997 26900
rect 2955 26851 2997 26860
rect 3243 26900 3285 26909
rect 4875 26900 4917 26909
rect 6586 26900 6644 26901
rect 3243 26860 3244 26900
rect 3284 26860 3285 26900
rect 3243 26851 3285 26860
rect 4491 26891 4533 26900
rect 4491 26851 4492 26891
rect 4532 26851 4533 26891
rect 4875 26860 4876 26900
rect 4916 26860 4917 26900
rect 4875 26851 4917 26860
rect 6123 26891 6165 26900
rect 6123 26851 6124 26891
rect 6164 26851 6165 26891
rect 6586 26860 6595 26900
rect 6635 26860 6644 26900
rect 6586 26859 6644 26860
rect 6699 26900 6741 26909
rect 6699 26860 6700 26900
rect 6740 26860 6741 26900
rect 6699 26851 6741 26860
rect 7083 26900 7125 26909
rect 9099 26900 9141 26909
rect 7083 26860 7084 26900
rect 7124 26860 7125 26900
rect 7083 26851 7125 26860
rect 7659 26891 7701 26900
rect 7659 26851 7660 26891
rect 7700 26851 7701 26891
rect 2466 26842 2512 26851
rect 4491 26842 4533 26851
rect 6123 26842 6165 26851
rect 7659 26842 7701 26851
rect 8139 26891 8181 26900
rect 8139 26851 8140 26891
rect 8180 26851 8181 26891
rect 8139 26842 8181 26851
rect 8514 26891 8560 26900
rect 8514 26851 8515 26891
rect 8555 26851 8560 26891
rect 9099 26860 9100 26900
rect 9140 26860 9141 26900
rect 9099 26851 9141 26860
rect 10347 26891 10389 26900
rect 10347 26851 10348 26891
rect 10388 26851 10389 26891
rect 8514 26842 8560 26851
rect 10347 26842 10389 26851
rect 1371 26816 1413 26825
rect 1371 26776 1372 26816
rect 1412 26776 1413 26816
rect 1371 26767 1413 26776
rect 7179 26816 7221 26825
rect 7179 26776 7180 26816
rect 7220 26776 7221 26816
rect 7179 26767 7221 26776
rect 8667 26816 8709 26825
rect 8667 26776 8668 26816
rect 8708 26776 8709 26816
rect 8667 26767 8709 26776
rect 10539 26648 10581 26657
rect 10539 26608 10540 26648
rect 10580 26608 10581 26648
rect 10539 26599 10581 26608
rect 1152 26480 10656 26504
rect 1152 26440 3688 26480
rect 3728 26440 3770 26480
rect 3810 26440 3852 26480
rect 3892 26440 3934 26480
rect 3974 26440 4016 26480
rect 4056 26440 10656 26480
rect 1152 26416 10656 26440
rect 4635 26312 4677 26321
rect 4635 26272 4636 26312
rect 4676 26272 4677 26312
rect 4635 26263 4677 26272
rect 5019 26312 5061 26321
rect 5019 26272 5020 26312
rect 5060 26272 5061 26312
rect 5019 26263 5061 26272
rect 9627 26312 9669 26321
rect 9627 26272 9628 26312
rect 9668 26272 9669 26312
rect 9627 26263 9669 26272
rect 10203 26228 10245 26237
rect 10203 26188 10204 26228
rect 10244 26188 10245 26228
rect 10203 26179 10245 26188
rect 1371 26144 1413 26153
rect 1371 26104 1372 26144
rect 1412 26104 1413 26144
rect 1371 26095 1413 26104
rect 3675 26144 3717 26153
rect 3675 26104 3676 26144
rect 3716 26104 3717 26144
rect 3675 26095 3717 26104
rect 4395 26144 4437 26153
rect 4395 26104 4396 26144
rect 4436 26104 4437 26144
rect 4395 26095 4437 26104
rect 4779 26144 4821 26153
rect 4779 26104 4780 26144
rect 4820 26104 4821 26144
rect 4779 26095 4821 26104
rect 5451 26144 5493 26153
rect 5451 26104 5452 26144
rect 5492 26104 5493 26144
rect 5451 26095 5493 26104
rect 6315 26144 6357 26153
rect 6315 26104 6316 26144
rect 6356 26104 6357 26144
rect 6315 26095 6357 26104
rect 6891 26144 6933 26153
rect 6891 26104 6892 26144
rect 6932 26104 6933 26144
rect 6891 26095 6933 26104
rect 9387 26144 9429 26153
rect 9387 26104 9388 26144
rect 9428 26104 9429 26144
rect 9387 26095 9429 26104
rect 9963 26144 10005 26153
rect 9963 26104 9964 26144
rect 10004 26104 10005 26144
rect 9963 26095 10005 26104
rect 10347 26144 10389 26153
rect 10347 26104 10348 26144
rect 10388 26104 10389 26144
rect 10347 26095 10389 26104
rect 1162 26060 1220 26061
rect 1162 26020 1171 26060
rect 1211 26020 1220 26060
rect 1162 26019 1220 26020
rect 1803 26060 1845 26069
rect 1803 26020 1804 26060
rect 1844 26020 1845 26060
rect 1803 26011 1845 26020
rect 3043 26060 3101 26061
rect 3043 26020 3052 26060
rect 3092 26020 3101 26060
rect 3043 26019 3101 26020
rect 3466 26060 3524 26061
rect 3466 26020 3475 26060
rect 3515 26020 3524 26060
rect 3466 26019 3524 26020
rect 4011 26060 4053 26069
rect 4011 26020 4012 26060
rect 4052 26020 4053 26060
rect 4011 26011 4053 26020
rect 4186 26060 4244 26061
rect 4186 26020 4195 26060
rect 4235 26020 4244 26060
rect 4186 26019 4244 26020
rect 7755 26060 7797 26069
rect 7755 26020 7756 26060
rect 7796 26020 7797 26060
rect 7755 26011 7797 26020
rect 8995 26060 9053 26061
rect 8995 26020 9004 26060
rect 9044 26020 9053 26060
rect 8995 26019 9053 26020
rect 10587 25976 10629 25985
rect 10587 25936 10588 25976
rect 10628 25936 10629 25976
rect 10587 25927 10629 25936
rect 3243 25892 3285 25901
rect 3243 25852 3244 25892
rect 3284 25852 3285 25892
rect 3243 25843 3285 25852
rect 4107 25892 4149 25901
rect 4107 25852 4108 25892
rect 4148 25852 4149 25892
rect 4107 25843 4149 25852
rect 5242 25892 5300 25893
rect 5242 25852 5251 25892
rect 5291 25852 5300 25892
rect 5242 25851 5300 25852
rect 5722 25892 5780 25893
rect 5722 25852 5731 25892
rect 5771 25852 5780 25892
rect 5722 25851 5780 25852
rect 6106 25892 6164 25893
rect 6106 25852 6115 25892
rect 6155 25852 6164 25892
rect 6106 25851 6164 25852
rect 6682 25892 6740 25893
rect 6682 25852 6691 25892
rect 6731 25852 6740 25892
rect 6682 25851 6740 25852
rect 7258 25892 7316 25893
rect 7258 25852 7267 25892
rect 7307 25852 7316 25892
rect 7258 25851 7316 25852
rect 7546 25892 7604 25893
rect 7546 25852 7555 25892
rect 7595 25852 7604 25892
rect 7546 25851 7604 25852
rect 9195 25892 9237 25901
rect 9195 25852 9196 25892
rect 9236 25852 9237 25892
rect 9195 25843 9237 25852
rect 1152 25724 10656 25748
rect 1152 25684 4928 25724
rect 4968 25684 5010 25724
rect 5050 25684 5092 25724
rect 5132 25684 5174 25724
rect 5214 25684 5256 25724
rect 5296 25684 10656 25724
rect 1152 25660 10656 25684
rect 4731 25556 4773 25565
rect 4731 25516 4732 25556
rect 4772 25516 4773 25556
rect 4731 25507 4773 25516
rect 4829 25556 4887 25557
rect 4829 25516 4838 25556
rect 4878 25516 4887 25556
rect 4829 25515 4887 25516
rect 9675 25556 9717 25565
rect 9675 25516 9676 25556
rect 9716 25516 9717 25556
rect 9675 25507 9717 25516
rect 3147 25472 3189 25481
rect 3147 25432 3148 25472
rect 3188 25432 3189 25472
rect 3147 25423 3189 25432
rect 4395 25472 4437 25481
rect 4395 25432 4396 25472
rect 4436 25432 4437 25472
rect 4395 25423 4437 25432
rect 7467 25472 7509 25481
rect 7467 25432 7468 25472
rect 7508 25432 7509 25472
rect 7467 25423 7509 25432
rect 1227 25388 1269 25397
rect 2938 25388 2996 25389
rect 1227 25348 1228 25388
rect 1268 25348 1269 25388
rect 1227 25339 1269 25348
rect 2475 25379 2517 25388
rect 2475 25339 2476 25379
rect 2516 25339 2517 25379
rect 2938 25348 2947 25388
rect 2987 25348 2996 25388
rect 2938 25347 2996 25348
rect 3243 25388 3285 25397
rect 3243 25348 3244 25388
rect 3284 25348 3285 25388
rect 3243 25339 3285 25348
rect 3435 25388 3477 25397
rect 3435 25348 3436 25388
rect 3476 25348 3477 25388
rect 3435 25339 3477 25348
rect 3552 25388 3610 25389
rect 3552 25348 3561 25388
rect 3601 25348 3610 25388
rect 3552 25347 3610 25348
rect 3723 25388 3765 25397
rect 3723 25348 3724 25388
rect 3764 25348 3765 25388
rect 3723 25339 3765 25348
rect 4011 25388 4053 25397
rect 4011 25348 4012 25388
rect 4052 25348 4053 25388
rect 4011 25339 4053 25348
rect 4282 25388 4340 25389
rect 4282 25348 4291 25388
rect 4331 25348 4340 25388
rect 4282 25347 4340 25348
rect 4954 25388 5012 25389
rect 5499 25388 5541 25397
rect 4954 25348 4963 25388
rect 5003 25348 5012 25388
rect 4954 25347 5012 25348
rect 5067 25379 5109 25388
rect 5067 25339 5068 25379
rect 5108 25339 5109 25379
rect 5499 25348 5500 25388
rect 5540 25348 5541 25388
rect 5499 25339 5541 25348
rect 5643 25388 5685 25397
rect 5643 25348 5644 25388
rect 5684 25348 5685 25388
rect 5643 25339 5685 25348
rect 6027 25388 6069 25397
rect 7930 25388 7988 25389
rect 6027 25348 6028 25388
rect 6068 25348 6069 25388
rect 6027 25339 6069 25348
rect 7275 25379 7317 25388
rect 7275 25339 7276 25379
rect 7316 25339 7317 25379
rect 7930 25348 7939 25388
rect 7979 25348 7988 25388
rect 7930 25347 7988 25348
rect 8043 25388 8085 25397
rect 8043 25348 8044 25388
rect 8084 25348 8085 25388
rect 8043 25339 8085 25348
rect 8427 25388 8469 25397
rect 10011 25388 10053 25397
rect 8427 25348 8428 25388
rect 8468 25348 8469 25388
rect 8427 25339 8469 25348
rect 9003 25379 9045 25388
rect 9003 25339 9004 25379
rect 9044 25339 9045 25379
rect 2475 25330 2517 25339
rect 5067 25330 5109 25339
rect 7275 25330 7317 25339
rect 9003 25330 9045 25339
rect 9483 25379 9525 25388
rect 9483 25339 9484 25379
rect 9524 25339 9525 25379
rect 9483 25330 9525 25339
rect 9858 25379 9904 25388
rect 9858 25339 9859 25379
rect 9899 25339 9904 25379
rect 10011 25348 10012 25388
rect 10052 25348 10053 25388
rect 10011 25339 10053 25348
rect 9858 25330 9904 25339
rect 8523 25304 8565 25313
rect 8523 25264 8524 25304
rect 8564 25264 8565 25304
rect 8523 25255 8565 25264
rect 10347 25304 10389 25313
rect 10347 25264 10348 25304
rect 10388 25264 10389 25304
rect 10347 25255 10389 25264
rect 2667 25220 2709 25229
rect 2667 25180 2668 25220
rect 2708 25180 2709 25220
rect 2667 25171 2709 25180
rect 3435 25136 3477 25145
rect 3435 25096 3436 25136
rect 3476 25096 3477 25136
rect 3435 25087 3477 25096
rect 5355 25136 5397 25145
rect 5355 25096 5356 25136
rect 5396 25096 5397 25136
rect 5355 25087 5397 25096
rect 10587 25136 10629 25145
rect 10587 25096 10588 25136
rect 10628 25096 10629 25136
rect 10587 25087 10629 25096
rect 1152 24968 10656 24992
rect 1152 24928 3688 24968
rect 3728 24928 3770 24968
rect 3810 24928 3852 24968
rect 3892 24928 3934 24968
rect 3974 24928 4016 24968
rect 4056 24928 10656 24968
rect 1152 24904 10656 24928
rect 2667 24800 2709 24809
rect 2667 24760 2668 24800
rect 2708 24760 2709 24800
rect 2667 24751 2709 24760
rect 6027 24716 6069 24725
rect 6027 24676 6028 24716
rect 6068 24676 6069 24716
rect 6027 24667 6069 24676
rect 10539 24716 10581 24725
rect 10539 24676 10540 24716
rect 10580 24676 10581 24716
rect 10539 24667 10581 24676
rect 3610 24632 3668 24633
rect 3610 24592 3619 24632
rect 3659 24592 3668 24632
rect 3610 24591 3668 24592
rect 3819 24632 3861 24641
rect 3819 24592 3820 24632
rect 3860 24592 3861 24632
rect 3819 24583 3861 24592
rect 4322 24632 4364 24641
rect 4322 24592 4323 24632
rect 4363 24592 4364 24632
rect 4322 24583 4364 24592
rect 6795 24632 6837 24641
rect 6795 24592 6796 24632
rect 6836 24592 6837 24632
rect 6795 24583 6837 24592
rect 8379 24632 8421 24641
rect 8379 24592 8380 24632
rect 8420 24592 8421 24632
rect 8379 24583 8421 24592
rect 1227 24548 1269 24557
rect 1227 24508 1228 24548
rect 1268 24508 1269 24548
rect 1227 24499 1269 24508
rect 2467 24548 2525 24549
rect 2467 24508 2476 24548
rect 2516 24508 2525 24548
rect 2467 24507 2525 24508
rect 3051 24548 3093 24557
rect 3051 24508 3052 24548
rect 3092 24508 3093 24548
rect 3051 24499 3093 24508
rect 3185 24548 3243 24549
rect 3185 24508 3194 24548
rect 3234 24508 3243 24548
rect 3185 24507 3243 24508
rect 3495 24548 3537 24557
rect 3495 24508 3496 24548
rect 3536 24508 3537 24548
rect 3495 24499 3537 24508
rect 3723 24548 3765 24557
rect 3723 24508 3724 24548
rect 3764 24508 3765 24548
rect 3723 24499 3765 24508
rect 4203 24548 4245 24557
rect 4203 24508 4204 24548
rect 4244 24508 4245 24548
rect 4203 24499 4245 24508
rect 4420 24548 4462 24557
rect 4420 24508 4421 24548
rect 4461 24508 4462 24548
rect 4420 24499 4462 24508
rect 4627 24548 4669 24557
rect 4627 24508 4628 24548
rect 4668 24508 4669 24548
rect 4627 24499 4669 24508
rect 5827 24548 5885 24549
rect 5827 24508 5836 24548
rect 5876 24508 5885 24548
rect 5827 24507 5885 24508
rect 6298 24548 6356 24549
rect 6298 24508 6307 24548
rect 6347 24508 6356 24548
rect 6298 24507 6356 24508
rect 6411 24548 6453 24557
rect 6411 24508 6412 24548
rect 6452 24508 6453 24548
rect 6411 24499 6453 24508
rect 6891 24548 6933 24557
rect 6891 24508 6892 24548
rect 6932 24508 6933 24548
rect 6891 24499 6933 24508
rect 7363 24548 7421 24549
rect 7363 24508 7372 24548
rect 7412 24508 7421 24548
rect 7363 24507 7421 24508
rect 7851 24548 7909 24549
rect 7851 24508 7860 24548
rect 7900 24508 7909 24548
rect 7851 24507 7909 24508
rect 8074 24548 8132 24549
rect 8074 24508 8083 24548
rect 8123 24508 8132 24548
rect 8074 24507 8132 24508
rect 8170 24548 8228 24549
rect 8170 24508 8179 24548
rect 8219 24508 8228 24548
rect 8170 24507 8228 24508
rect 9099 24548 9141 24557
rect 9099 24508 9100 24548
rect 9140 24508 9141 24548
rect 9099 24499 9141 24508
rect 10339 24548 10397 24549
rect 10339 24508 10348 24548
rect 10388 24508 10397 24548
rect 10339 24507 10397 24508
rect 8715 24464 8757 24473
rect 8715 24424 8716 24464
rect 8756 24424 8757 24464
rect 8715 24415 8757 24424
rect 2667 24380 2709 24389
rect 2667 24340 2668 24380
rect 2708 24340 2709 24380
rect 2667 24331 2709 24340
rect 3339 24380 3381 24389
rect 3339 24340 3340 24380
rect 3380 24340 3381 24380
rect 3339 24331 3381 24340
rect 4107 24380 4149 24389
rect 4107 24340 4108 24380
rect 4148 24340 4149 24380
rect 4107 24331 4149 24340
rect 1152 24212 10656 24236
rect 1152 24172 4928 24212
rect 4968 24172 5010 24212
rect 5050 24172 5092 24212
rect 5132 24172 5174 24212
rect 5214 24172 5256 24212
rect 5296 24172 10656 24212
rect 1152 24148 10656 24172
rect 4011 24044 4053 24053
rect 4011 24004 4012 24044
rect 4052 24004 4053 24044
rect 4011 23995 4053 24004
rect 4779 24044 4821 24053
rect 4779 24004 4780 24044
rect 4820 24004 4821 24044
rect 4779 23995 4821 24004
rect 5146 24044 5204 24045
rect 5146 24004 5155 24044
rect 5195 24004 5204 24044
rect 5146 24003 5204 24004
rect 5722 24044 5780 24045
rect 5722 24004 5731 24044
rect 5771 24004 5780 24044
rect 5722 24003 5780 24004
rect 7371 24044 7413 24053
rect 7371 24004 7372 24044
rect 7412 24004 7413 24044
rect 7371 23995 7413 24004
rect 8410 24044 8468 24045
rect 8410 24004 8419 24044
rect 8459 24004 8468 24044
rect 8410 24003 8468 24004
rect 1707 23960 1749 23969
rect 1707 23920 1708 23960
rect 1748 23920 1749 23960
rect 1707 23911 1749 23920
rect 4347 23960 4389 23969
rect 4347 23920 4348 23960
rect 4388 23920 4389 23960
rect 4347 23911 4389 23920
rect 7563 23960 7605 23969
rect 7563 23920 7564 23960
rect 7604 23920 7605 23960
rect 7563 23911 7605 23920
rect 7851 23960 7893 23969
rect 7851 23920 7852 23960
rect 7892 23920 7893 23960
rect 7851 23911 7893 23920
rect 8619 23960 8661 23969
rect 8619 23920 8620 23960
rect 8660 23920 8661 23960
rect 8619 23911 8661 23920
rect 1323 23876 1365 23885
rect 1323 23836 1324 23876
rect 1364 23836 1365 23876
rect 1323 23827 1365 23836
rect 1594 23876 1652 23877
rect 1594 23836 1603 23876
rect 1643 23836 1652 23876
rect 1594 23835 1652 23836
rect 2266 23876 2324 23877
rect 2266 23836 2275 23876
rect 2315 23836 2324 23876
rect 2266 23835 2324 23836
rect 2379 23876 2421 23885
rect 2379 23836 2380 23876
rect 2420 23836 2421 23876
rect 2379 23827 2421 23836
rect 2763 23876 2805 23885
rect 4683 23876 4725 23885
rect 2763 23836 2764 23876
rect 2804 23836 2805 23876
rect 2763 23827 2805 23836
rect 3338 23867 3380 23876
rect 3338 23827 3339 23867
rect 3379 23827 3380 23867
rect 3338 23818 3380 23827
rect 3819 23867 3861 23876
rect 3819 23827 3820 23867
rect 3860 23827 3861 23867
rect 3819 23818 3861 23827
rect 4194 23867 4240 23876
rect 4194 23827 4195 23867
rect 4235 23827 4240 23867
rect 4683 23836 4684 23876
rect 4724 23836 4725 23876
rect 4683 23827 4725 23836
rect 4875 23876 4917 23885
rect 4875 23836 4876 23876
rect 4916 23836 4917 23876
rect 4875 23827 4917 23836
rect 5931 23876 5973 23885
rect 10347 23876 10389 23885
rect 5931 23836 5932 23876
rect 5972 23836 5973 23876
rect 5931 23827 5973 23836
rect 7179 23867 7221 23876
rect 7179 23827 7180 23867
rect 7220 23827 7221 23867
rect 4194 23818 4240 23827
rect 7179 23818 7221 23827
rect 9099 23867 9141 23876
rect 9099 23827 9100 23867
rect 9140 23827 9141 23867
rect 10347 23836 10348 23876
rect 10388 23836 10389 23876
rect 10347 23827 10389 23836
rect 9099 23818 9141 23827
rect 2859 23792 2901 23801
rect 2859 23752 2860 23792
rect 2900 23752 2901 23792
rect 2859 23743 2901 23752
rect 5355 23792 5397 23801
rect 5355 23752 5356 23792
rect 5396 23752 5397 23792
rect 5355 23743 5397 23752
rect 8331 23792 8373 23801
rect 8331 23752 8332 23792
rect 8372 23752 8373 23792
rect 8331 23743 8373 23752
rect 1995 23708 2037 23717
rect 1995 23668 1996 23708
rect 2036 23668 2037 23708
rect 1995 23659 2037 23668
rect 8907 23624 8949 23633
rect 8907 23584 8908 23624
rect 8948 23584 8949 23624
rect 8907 23575 8949 23584
rect 1152 23456 10656 23480
rect 1152 23416 3688 23456
rect 3728 23416 3770 23456
rect 3810 23416 3852 23456
rect 3892 23416 3934 23456
rect 3974 23416 4016 23456
rect 4056 23416 10656 23456
rect 1152 23392 10656 23416
rect 3435 23288 3477 23297
rect 3435 23248 3436 23288
rect 3476 23248 3477 23288
rect 3435 23239 3477 23248
rect 5787 23288 5829 23297
rect 5787 23248 5788 23288
rect 5828 23248 5829 23288
rect 5787 23239 5829 23248
rect 5067 23204 5109 23213
rect 5067 23164 5068 23204
rect 5108 23164 5109 23204
rect 5067 23155 5109 23164
rect 6123 23120 6165 23129
rect 6123 23080 6124 23120
rect 6164 23080 6165 23120
rect 6123 23071 6165 23080
rect 6603 23120 6645 23129
rect 6603 23080 6604 23120
rect 6644 23080 6645 23120
rect 6603 23071 6645 23080
rect 8523 23120 8565 23129
rect 8523 23080 8524 23120
rect 8564 23080 8565 23120
rect 8523 23071 8565 23080
rect 1162 23036 1220 23037
rect 1162 22996 1171 23036
rect 1211 22996 1220 23036
rect 1162 22995 1220 22996
rect 1657 23036 1715 23037
rect 1657 22996 1666 23036
rect 1706 22996 1715 23036
rect 1657 22995 1715 22996
rect 2137 23036 2195 23037
rect 2137 22996 2146 23036
rect 2186 22996 2195 23036
rect 2137 22995 2195 22996
rect 2763 23036 2805 23045
rect 2763 22996 2764 23036
rect 2804 22996 2805 23036
rect 2763 22987 2805 22996
rect 3034 23036 3092 23037
rect 3034 22996 3043 23036
rect 3083 22996 3092 23036
rect 3034 22995 3092 22996
rect 3577 23036 3635 23037
rect 3577 22996 3586 23036
rect 3626 22996 3635 23036
rect 3577 22995 3635 22996
rect 4057 23036 4115 23037
rect 4057 22996 4066 23036
rect 4106 22996 4115 23036
rect 4057 22995 4115 22996
rect 4587 23036 4629 23045
rect 4587 22996 4588 23036
rect 4628 22996 4629 23036
rect 4587 22987 4629 22996
rect 4875 23036 4917 23045
rect 4875 22996 4876 23036
rect 4916 22996 4917 23036
rect 4875 22987 4917 22996
rect 5067 23036 5109 23045
rect 5067 22996 5068 23036
rect 5108 22996 5109 23036
rect 5067 22987 5109 22996
rect 5259 23036 5301 23045
rect 5259 22996 5260 23036
rect 5300 22996 5301 23036
rect 5259 22987 5301 22996
rect 5643 23036 5685 23045
rect 5643 22996 5644 23036
rect 5684 22996 5685 23036
rect 5643 22987 5685 22996
rect 6967 23036 7025 23037
rect 6967 22996 6976 23036
rect 7016 22996 7025 23036
rect 6967 22995 7025 22996
rect 7131 23036 7173 23045
rect 7131 22996 7132 23036
rect 7172 22996 7173 23036
rect 7131 22987 7173 22996
rect 8026 23036 8084 23037
rect 8026 22996 8035 23036
rect 8075 22996 8084 23036
rect 8026 22995 8084 22996
rect 8139 23036 8181 23045
rect 8139 22996 8140 23036
rect 8180 22996 8181 23036
rect 8139 22987 8181 22996
rect 8619 23036 8661 23045
rect 8619 22996 8620 23036
rect 8660 22996 8661 23036
rect 8619 22987 8661 22996
rect 9091 23036 9149 23037
rect 9091 22996 9100 23036
rect 9140 22996 9149 23036
rect 9091 22995 9149 22996
rect 9610 23036 9668 23037
rect 9610 22996 9619 23036
rect 9659 22996 9668 23036
rect 9610 22995 9668 22996
rect 9898 23036 9956 23037
rect 9898 22996 9907 23036
rect 9947 22996 9956 23036
rect 9898 22995 9956 22996
rect 10443 23036 10485 23045
rect 10443 22996 10444 23036
rect 10484 22996 10485 23036
rect 10443 22987 10485 22996
rect 2331 22952 2373 22961
rect 2331 22912 2332 22952
rect 2372 22912 2373 22952
rect 2331 22903 2373 22912
rect 3147 22952 3189 22961
rect 3147 22912 3148 22952
rect 3188 22912 3189 22952
rect 3147 22903 3189 22912
rect 1371 22868 1413 22877
rect 1371 22828 1372 22868
rect 1412 22828 1413 22868
rect 1371 22819 1413 22828
rect 1851 22868 1893 22877
rect 1851 22828 1852 22868
rect 1892 22828 1893 22868
rect 1851 22819 1893 22828
rect 3771 22868 3813 22877
rect 3771 22828 3772 22868
rect 3812 22828 3813 22868
rect 3771 22819 3813 22828
rect 4251 22868 4293 22877
rect 4251 22828 4252 22868
rect 4292 22828 4293 22868
rect 4251 22819 4293 22828
rect 4666 22868 4724 22869
rect 4666 22828 4675 22868
rect 4715 22828 4724 22868
rect 4666 22827 4724 22828
rect 5883 22868 5925 22877
rect 5883 22828 5884 22868
rect 5924 22828 5925 22868
rect 5883 22819 5925 22828
rect 6394 22868 6452 22869
rect 6394 22828 6403 22868
rect 6443 22828 6452 22868
rect 6394 22827 6452 22828
rect 7546 22868 7604 22869
rect 7546 22828 7555 22868
rect 7595 22828 7604 22868
rect 7546 22827 7604 22828
rect 9771 22868 9813 22877
rect 9771 22828 9772 22868
rect 9812 22828 9813 22868
rect 9771 22819 9813 22828
rect 10107 22868 10149 22877
rect 10107 22828 10108 22868
rect 10148 22828 10149 22868
rect 10107 22819 10149 22828
rect 1152 22700 10656 22724
rect 1152 22660 4928 22700
rect 4968 22660 5010 22700
rect 5050 22660 5092 22700
rect 5132 22660 5174 22700
rect 5214 22660 5256 22700
rect 5296 22660 10656 22700
rect 1152 22636 10656 22660
rect 5739 22532 5781 22541
rect 5739 22492 5740 22532
rect 5780 22492 5781 22532
rect 5739 22483 5781 22492
rect 7738 22532 7796 22533
rect 7738 22492 7747 22532
rect 7787 22492 7796 22532
rect 7738 22491 7796 22492
rect 8026 22532 8084 22533
rect 8026 22492 8035 22532
rect 8075 22492 8084 22532
rect 8026 22491 8084 22492
rect 9867 22532 9909 22541
rect 9867 22492 9868 22532
rect 9908 22492 9909 22532
rect 9867 22483 9909 22492
rect 10587 22532 10629 22541
rect 10587 22492 10588 22532
rect 10628 22492 10629 22532
rect 10587 22483 10629 22492
rect 2667 22448 2709 22457
rect 2667 22408 2668 22448
rect 2708 22408 2709 22448
rect 2667 22399 2709 22408
rect 1227 22364 1269 22373
rect 3147 22364 3189 22373
rect 1227 22324 1228 22364
rect 1268 22324 1269 22364
rect 1227 22315 1269 22324
rect 2475 22355 2517 22364
rect 2475 22315 2476 22355
rect 2516 22315 2517 22355
rect 3147 22324 3148 22364
rect 3188 22324 3189 22364
rect 3147 22315 3189 22324
rect 3248 22364 3306 22365
rect 3248 22324 3257 22364
rect 3297 22324 3306 22364
rect 3248 22323 3306 22324
rect 3531 22364 3573 22373
rect 3531 22324 3532 22364
rect 3572 22324 3573 22364
rect 3531 22315 3573 22324
rect 3994 22364 4052 22365
rect 3994 22324 4003 22364
rect 4043 22324 4052 22364
rect 3994 22323 4052 22324
rect 4107 22364 4149 22373
rect 4107 22324 4108 22364
rect 4148 22324 4149 22364
rect 4107 22315 4149 22324
rect 4491 22364 4533 22373
rect 7563 22364 7605 22373
rect 4491 22324 4492 22364
rect 4532 22324 4533 22364
rect 4491 22315 4533 22324
rect 5067 22355 5109 22364
rect 5067 22315 5068 22355
rect 5108 22315 5109 22355
rect 2475 22306 2517 22315
rect 5067 22306 5109 22315
rect 5547 22355 5589 22364
rect 5547 22315 5548 22355
rect 5588 22315 5589 22355
rect 5547 22306 5589 22315
rect 6315 22355 6357 22364
rect 6315 22315 6316 22355
rect 6356 22315 6357 22355
rect 7563 22324 7564 22364
rect 7604 22324 7605 22364
rect 7563 22315 7605 22324
rect 8427 22364 8469 22373
rect 8427 22324 8428 22364
rect 8468 22324 8469 22364
rect 8427 22315 8469 22324
rect 9675 22355 9717 22364
rect 9675 22315 9676 22355
rect 9716 22315 9717 22355
rect 6315 22306 6357 22315
rect 9675 22306 9717 22315
rect 4587 22280 4629 22289
rect 4587 22240 4588 22280
rect 4628 22240 4629 22280
rect 4587 22231 4629 22240
rect 6106 22280 6164 22281
rect 6106 22240 6115 22280
rect 6155 22240 6164 22280
rect 6106 22239 6164 22240
rect 10059 22280 10101 22289
rect 10059 22240 10060 22280
rect 10100 22240 10101 22280
rect 10059 22231 10101 22240
rect 10347 22280 10389 22289
rect 10347 22240 10348 22280
rect 10388 22240 10389 22280
rect 10347 22231 10389 22240
rect 2859 22196 2901 22205
rect 2859 22156 2860 22196
rect 2900 22156 2901 22196
rect 2859 22147 2901 22156
rect 1152 21944 10656 21968
rect 1152 21904 3688 21944
rect 3728 21904 3770 21944
rect 3810 21904 3852 21944
rect 3892 21904 3934 21944
rect 3974 21904 4016 21944
rect 4056 21904 10656 21944
rect 1152 21880 10656 21904
rect 2667 21776 2709 21785
rect 2667 21736 2668 21776
rect 2708 21736 2709 21776
rect 2667 21727 2709 21736
rect 8715 21776 8757 21785
rect 8715 21736 8716 21776
rect 8756 21736 8757 21776
rect 8715 21727 8757 21736
rect 10587 21776 10629 21785
rect 10587 21736 10588 21776
rect 10628 21736 10629 21776
rect 10587 21727 10629 21736
rect 1371 21608 1413 21617
rect 1371 21568 1372 21608
rect 1412 21568 1413 21608
rect 1371 21559 1413 21568
rect 3435 21608 3477 21617
rect 3435 21568 3436 21608
rect 3476 21568 3477 21608
rect 3435 21559 3477 21568
rect 6682 21608 6740 21609
rect 6682 21568 6691 21608
rect 6731 21568 6740 21608
rect 6682 21567 6740 21568
rect 8331 21608 8373 21617
rect 8331 21568 8332 21608
rect 8372 21568 8373 21608
rect 6027 21557 6069 21566
rect 8331 21559 8373 21568
rect 10347 21608 10389 21617
rect 10347 21568 10348 21608
rect 10388 21568 10389 21608
rect 10347 21559 10389 21568
rect 1162 21524 1220 21525
rect 1162 21484 1171 21524
rect 1211 21484 1220 21524
rect 1162 21483 1220 21484
rect 1995 21524 2037 21533
rect 1995 21484 1996 21524
rect 2036 21484 2037 21524
rect 1995 21475 2037 21484
rect 2266 21524 2324 21525
rect 2266 21484 2275 21524
rect 2315 21484 2324 21524
rect 2266 21483 2324 21484
rect 2938 21524 2996 21525
rect 2938 21484 2947 21524
rect 2987 21484 2996 21524
rect 2938 21483 2996 21484
rect 3051 21524 3093 21533
rect 3051 21484 3052 21524
rect 3092 21484 3093 21524
rect 3051 21475 3093 21484
rect 3531 21524 3573 21533
rect 3531 21484 3532 21524
rect 3572 21484 3573 21524
rect 3531 21475 3573 21484
rect 4003 21524 4061 21525
rect 4003 21484 4012 21524
rect 4052 21484 4061 21524
rect 4003 21483 4061 21484
rect 4491 21524 4549 21525
rect 4491 21484 4500 21524
rect 4540 21484 4549 21524
rect 4491 21483 4549 21484
rect 4971 21524 5013 21533
rect 4971 21484 4972 21524
rect 5012 21484 5013 21524
rect 4971 21475 5013 21484
rect 5218 21524 5276 21525
rect 5218 21484 5227 21524
rect 5267 21484 5276 21524
rect 5218 21483 5276 21484
rect 5338 21524 5396 21525
rect 5338 21484 5347 21524
rect 5387 21484 5396 21524
rect 5338 21483 5396 21484
rect 5914 21524 5972 21525
rect 5914 21484 5923 21524
rect 5963 21484 5972 21524
rect 6027 21517 6028 21557
rect 6068 21517 6069 21557
rect 6027 21508 6069 21517
rect 6883 21524 6941 21525
rect 5914 21483 5972 21484
rect 6883 21484 6892 21524
rect 6932 21484 6941 21524
rect 6883 21483 6941 21484
rect 8139 21524 8181 21533
rect 8139 21484 8140 21524
rect 8180 21484 8181 21524
rect 8139 21475 8181 21484
rect 8899 21524 8957 21525
rect 8899 21484 8908 21524
rect 8948 21484 8957 21524
rect 8899 21483 8957 21484
rect 10155 21524 10197 21533
rect 10155 21484 10156 21524
rect 10196 21484 10197 21524
rect 10155 21475 10197 21484
rect 2379 21440 2421 21449
rect 2379 21400 2380 21440
rect 2420 21400 2421 21440
rect 2379 21391 2421 21400
rect 6346 21440 6404 21441
rect 6346 21400 6355 21440
rect 6395 21400 6404 21440
rect 6346 21399 6404 21400
rect 4683 21356 4725 21365
rect 4683 21316 4684 21356
rect 4724 21316 4725 21356
rect 4683 21307 4725 21316
rect 5691 21356 5733 21365
rect 8571 21356 8613 21365
rect 5691 21316 5692 21356
rect 5732 21316 5733 21356
rect 5691 21307 5733 21316
rect 5826 21347 5872 21356
rect 5826 21307 5827 21347
rect 5867 21307 5872 21347
rect 8571 21316 8572 21356
rect 8612 21316 8613 21356
rect 8571 21307 8613 21316
rect 5826 21298 5872 21307
rect 1152 21188 10656 21212
rect 1152 21148 4928 21188
rect 4968 21148 5010 21188
rect 5050 21148 5092 21188
rect 5132 21148 5174 21188
rect 5214 21148 5256 21188
rect 5296 21148 10656 21188
rect 1152 21124 10656 21148
rect 1371 21020 1413 21029
rect 1371 20980 1372 21020
rect 1412 20980 1413 21020
rect 1371 20971 1413 20980
rect 5547 21020 5589 21029
rect 5547 20980 5548 21020
rect 5588 20980 5589 21020
rect 5547 20971 5589 20980
rect 6490 21020 6548 21021
rect 6490 20980 6499 21020
rect 6539 20980 6548 21020
rect 6490 20979 6548 20980
rect 7066 21020 7124 21021
rect 7066 20980 7075 21020
rect 7115 20980 7124 21020
rect 7066 20979 7124 20980
rect 2283 20936 2325 20945
rect 2283 20896 2284 20936
rect 2324 20896 2325 20936
rect 2283 20887 2325 20896
rect 3243 20936 3285 20945
rect 3243 20896 3244 20936
rect 3284 20896 3285 20936
rect 3243 20887 3285 20896
rect 7275 20936 7317 20945
rect 7275 20896 7276 20936
rect 7316 20896 7317 20936
rect 7275 20887 7317 20896
rect 1899 20852 1941 20861
rect 1218 20843 1264 20852
rect 1218 20803 1219 20843
rect 1259 20803 1264 20843
rect 1899 20812 1900 20852
rect 1940 20812 1941 20852
rect 1899 20803 1941 20812
rect 2170 20852 2228 20853
rect 2170 20812 2179 20852
rect 2219 20812 2228 20852
rect 2170 20811 2228 20812
rect 2859 20852 2901 20861
rect 2859 20812 2860 20852
rect 2900 20812 2901 20852
rect 2859 20803 2901 20812
rect 3130 20852 3188 20853
rect 3130 20812 3139 20852
rect 3179 20812 3188 20852
rect 3130 20811 3188 20812
rect 3802 20852 3860 20853
rect 3802 20812 3811 20852
rect 3851 20812 3860 20852
rect 3802 20811 3860 20812
rect 3915 20852 3957 20861
rect 3915 20812 3916 20852
rect 3956 20812 3957 20852
rect 3915 20803 3957 20812
rect 4299 20852 4341 20861
rect 5686 20852 5728 20861
rect 4299 20812 4300 20852
rect 4340 20812 4341 20852
rect 4299 20803 4341 20812
rect 4875 20843 4917 20852
rect 4875 20803 4876 20843
rect 4916 20803 4917 20843
rect 1218 20794 1264 20803
rect 4875 20794 4917 20803
rect 5355 20843 5397 20852
rect 5355 20803 5356 20843
rect 5396 20803 5397 20843
rect 5686 20812 5687 20852
rect 5727 20812 5728 20852
rect 5686 20803 5728 20812
rect 5931 20852 5973 20861
rect 5931 20812 5932 20852
rect 5972 20812 5973 20852
rect 5931 20803 5973 20812
rect 6166 20852 6208 20861
rect 6166 20812 6167 20852
rect 6207 20812 6208 20852
rect 6166 20803 6208 20812
rect 6411 20852 6453 20861
rect 8715 20852 8757 20861
rect 10347 20852 10389 20861
rect 6411 20812 6412 20852
rect 6452 20812 6453 20852
rect 6411 20803 6453 20812
rect 7467 20843 7509 20852
rect 7467 20803 7468 20843
rect 7508 20803 7509 20843
rect 8715 20812 8716 20852
rect 8756 20812 8757 20852
rect 8715 20803 8757 20812
rect 9099 20843 9141 20852
rect 9099 20803 9100 20843
rect 9140 20803 9141 20843
rect 10347 20812 10348 20852
rect 10388 20812 10389 20852
rect 10347 20803 10389 20812
rect 5355 20794 5397 20803
rect 7467 20794 7509 20803
rect 9099 20794 9141 20803
rect 4395 20768 4437 20777
rect 4395 20728 4396 20768
rect 4436 20728 4437 20768
rect 4395 20719 4437 20728
rect 5818 20768 5876 20769
rect 5818 20728 5827 20768
rect 5867 20728 5876 20768
rect 5818 20727 5876 20728
rect 6027 20768 6069 20777
rect 6027 20728 6028 20768
rect 6068 20728 6069 20768
rect 6027 20719 6069 20728
rect 6298 20768 6356 20769
rect 6298 20728 6307 20768
rect 6347 20728 6356 20768
rect 6298 20727 6356 20728
rect 6699 20768 6741 20777
rect 6699 20728 6700 20768
rect 6740 20728 6741 20768
rect 6699 20719 6741 20728
rect 8907 20684 8949 20693
rect 8907 20644 8908 20684
rect 8948 20644 8949 20684
rect 8907 20635 8949 20644
rect 2571 20600 2613 20609
rect 2571 20560 2572 20600
rect 2612 20560 2613 20600
rect 2571 20551 2613 20560
rect 3531 20600 3573 20609
rect 3531 20560 3532 20600
rect 3572 20560 3573 20600
rect 3531 20551 3573 20560
rect 1152 20432 10656 20456
rect 1152 20392 3688 20432
rect 3728 20392 3770 20432
rect 3810 20392 3852 20432
rect 3892 20392 3934 20432
rect 3974 20392 4016 20432
rect 4056 20392 10656 20432
rect 1152 20368 10656 20392
rect 5931 20264 5973 20273
rect 5931 20224 5932 20264
rect 5972 20224 5973 20264
rect 5931 20215 5973 20224
rect 2763 20180 2805 20189
rect 2763 20140 2764 20180
rect 2804 20140 2805 20180
rect 2763 20131 2805 20140
rect 5163 20180 5205 20189
rect 5163 20140 5164 20180
rect 5204 20140 5205 20180
rect 5163 20131 5205 20140
rect 8763 20180 8805 20189
rect 8763 20140 8764 20180
rect 8804 20140 8805 20180
rect 8763 20131 8805 20140
rect 3531 20096 3573 20105
rect 3531 20056 3532 20096
rect 3572 20056 3573 20096
rect 3531 20047 3573 20056
rect 8523 20096 8565 20105
rect 8523 20056 8524 20096
rect 8564 20056 8565 20096
rect 8523 20047 8565 20056
rect 1162 20012 1220 20013
rect 1162 19972 1171 20012
rect 1211 19972 1220 20012
rect 1162 19971 1220 19972
rect 1803 20012 1845 20021
rect 1803 19972 1804 20012
rect 1844 19972 1845 20012
rect 1803 19963 1845 19972
rect 2091 20012 2133 20021
rect 2091 19972 2092 20012
rect 2132 19972 2133 20012
rect 2091 19963 2133 19972
rect 2362 20012 2420 20013
rect 3147 20012 3189 20021
rect 2362 19972 2371 20012
rect 2411 19972 2420 20012
rect 2362 19971 2420 19972
rect 3034 20011 3092 20012
rect 3034 19971 3043 20011
rect 3083 19971 3092 20011
rect 3034 19970 3092 19971
rect 3147 19972 3148 20012
rect 3188 19972 3189 20012
rect 3147 19963 3189 19972
rect 3627 20012 3669 20021
rect 3627 19972 3628 20012
rect 3668 19972 3669 20012
rect 3627 19963 3669 19972
rect 4099 20012 4157 20013
rect 4099 19972 4108 20012
rect 4148 19972 4157 20012
rect 4099 19971 4157 19972
rect 4618 20012 4676 20013
rect 4618 19972 4627 20012
rect 4667 19972 4676 20012
rect 4618 19971 4676 19972
rect 4971 20012 5013 20021
rect 4971 19972 4972 20012
rect 5012 19972 5013 20012
rect 4971 19963 5013 19972
rect 5088 20012 5146 20013
rect 5088 19972 5097 20012
rect 5137 19972 5146 20012
rect 5088 19971 5146 19972
rect 5259 20012 5301 20021
rect 5259 19972 5260 20012
rect 5300 19972 5301 20012
rect 5259 19963 5301 19972
rect 5595 20012 5637 20021
rect 5595 19972 5596 20012
rect 5636 19972 5637 20012
rect 5595 19963 5637 19972
rect 5739 20012 5781 20021
rect 5739 19972 5740 20012
rect 5780 19972 5781 20012
rect 5739 19963 5781 19972
rect 5931 20012 5973 20021
rect 5931 19972 5932 20012
rect 5972 19972 5973 20012
rect 5931 19963 5973 19972
rect 6123 20012 6165 20021
rect 6123 19972 6124 20012
rect 6164 19972 6165 20012
rect 6123 19963 6165 19972
rect 6603 20012 6645 20021
rect 6603 19972 6604 20012
rect 6644 19972 6645 20012
rect 6603 19963 6645 19972
rect 7843 20012 7901 20013
rect 7843 19972 7852 20012
rect 7892 19972 7901 20012
rect 7843 19971 7901 19972
rect 8907 20012 8949 20021
rect 8907 19972 8908 20012
rect 8948 19972 8949 20012
rect 8907 19963 8949 19972
rect 10147 20012 10205 20013
rect 10147 19972 10156 20012
rect 10196 19972 10205 20012
rect 10147 19971 10205 19972
rect 2475 19928 2517 19937
rect 2475 19888 2476 19928
rect 2516 19888 2517 19928
rect 2475 19879 2517 19888
rect 8235 19928 8277 19937
rect 8235 19888 8236 19928
rect 8276 19888 8277 19928
rect 8235 19879 8277 19888
rect 1371 19844 1413 19853
rect 1371 19804 1372 19844
rect 1412 19804 1413 19844
rect 1371 19795 1413 19804
rect 4779 19844 4821 19853
rect 4779 19804 4780 19844
rect 4820 19804 4821 19844
rect 4779 19795 4821 19804
rect 5434 19844 5492 19845
rect 5434 19804 5443 19844
rect 5483 19804 5492 19844
rect 5434 19803 5492 19804
rect 6394 19844 6452 19845
rect 6394 19804 6403 19844
rect 6443 19804 6452 19844
rect 6394 19803 6452 19804
rect 8043 19844 8085 19853
rect 8043 19804 8044 19844
rect 8084 19804 8085 19844
rect 8043 19795 8085 19804
rect 10347 19844 10389 19853
rect 10347 19804 10348 19844
rect 10388 19804 10389 19844
rect 10347 19795 10389 19804
rect 1152 19676 10656 19700
rect 1152 19636 4928 19676
rect 4968 19636 5010 19676
rect 5050 19636 5092 19676
rect 5132 19636 5174 19676
rect 5214 19636 5256 19676
rect 5296 19636 10656 19676
rect 1152 19612 10656 19636
rect 3195 19508 3237 19517
rect 3195 19468 3196 19508
rect 3236 19468 3237 19508
rect 3195 19459 3237 19468
rect 3675 19508 3717 19517
rect 3675 19468 3676 19508
rect 3716 19468 3717 19508
rect 3675 19459 3717 19468
rect 8619 19508 8661 19517
rect 8619 19468 8620 19508
rect 8660 19468 8661 19508
rect 8619 19459 8661 19468
rect 2571 19424 2613 19433
rect 2571 19384 2572 19424
rect 2612 19384 2613 19424
rect 2571 19375 2613 19384
rect 4635 19424 4677 19433
rect 4635 19384 4636 19424
rect 4676 19384 4677 19424
rect 4635 19375 4677 19384
rect 6603 19424 6645 19433
rect 6603 19384 6604 19424
rect 6644 19384 6645 19424
rect 6603 19375 6645 19384
rect 1371 19340 1413 19349
rect 1218 19331 1264 19340
rect 1218 19291 1219 19331
rect 1259 19291 1264 19331
rect 1371 19300 1372 19340
rect 1412 19300 1413 19340
rect 1371 19291 1413 19300
rect 2139 19340 2181 19349
rect 2139 19300 2140 19340
rect 2180 19300 2181 19340
rect 2139 19291 2181 19300
rect 2458 19340 2516 19341
rect 5163 19340 5205 19349
rect 6874 19340 6932 19341
rect 2458 19300 2467 19340
rect 2507 19300 2516 19340
rect 2458 19299 2516 19300
rect 3042 19331 3088 19340
rect 3042 19291 3043 19331
rect 3083 19291 3088 19331
rect 1218 19282 1264 19291
rect 3042 19282 3088 19291
rect 3522 19331 3568 19340
rect 3522 19291 3523 19331
rect 3563 19291 3568 19331
rect 3522 19282 3568 19291
rect 4002 19331 4048 19340
rect 4002 19291 4003 19331
rect 4043 19291 4048 19331
rect 4002 19282 4048 19291
rect 4482 19331 4528 19340
rect 4482 19291 4483 19331
rect 4523 19291 4528 19331
rect 5163 19300 5164 19340
rect 5204 19300 5205 19340
rect 5163 19291 5205 19300
rect 6411 19331 6453 19340
rect 6411 19291 6412 19331
rect 6452 19291 6453 19331
rect 6874 19300 6883 19340
rect 6923 19300 6932 19340
rect 6874 19299 6932 19300
rect 6987 19340 7029 19349
rect 6987 19300 6988 19340
rect 7028 19300 7029 19340
rect 6987 19291 7029 19300
rect 7371 19340 7413 19349
rect 10539 19340 10581 19349
rect 7371 19300 7372 19340
rect 7412 19300 7413 19340
rect 7371 19291 7413 19300
rect 7947 19331 7989 19340
rect 7947 19291 7948 19331
rect 7988 19291 7989 19331
rect 4482 19282 4528 19291
rect 6411 19282 6453 19291
rect 7947 19282 7989 19291
rect 8427 19331 8469 19340
rect 8427 19291 8428 19331
rect 8468 19291 8469 19331
rect 8427 19282 8469 19291
rect 9291 19331 9333 19340
rect 9291 19291 9292 19331
rect 9332 19291 9333 19331
rect 10539 19300 10540 19340
rect 10580 19300 10581 19340
rect 10539 19291 10581 19300
rect 9291 19282 9333 19291
rect 1707 19256 1749 19265
rect 1707 19216 1708 19256
rect 1748 19216 1749 19256
rect 1707 19207 1749 19216
rect 4155 19256 4197 19265
rect 4155 19216 4156 19256
rect 4196 19216 4197 19256
rect 4155 19207 4197 19216
rect 7467 19256 7509 19265
rect 7467 19216 7468 19256
rect 7508 19216 7509 19256
rect 7467 19207 7509 19216
rect 8811 19256 8853 19265
rect 8811 19216 8812 19256
rect 8852 19216 8853 19256
rect 8811 19207 8853 19216
rect 2859 19172 2901 19181
rect 2859 19132 2860 19172
rect 2900 19132 2901 19172
rect 2859 19123 2901 19132
rect 1947 19088 1989 19097
rect 1947 19048 1948 19088
rect 1988 19048 1989 19088
rect 1947 19039 1989 19048
rect 9099 19088 9141 19097
rect 9099 19048 9100 19088
rect 9140 19048 9141 19088
rect 9099 19039 9141 19048
rect 1152 18920 10656 18944
rect 1152 18880 3688 18920
rect 3728 18880 3770 18920
rect 3810 18880 3852 18920
rect 3892 18880 3934 18920
rect 3974 18880 4016 18920
rect 4056 18880 10656 18920
rect 1152 18856 10656 18880
rect 7323 18752 7365 18761
rect 7323 18712 7324 18752
rect 7364 18712 7365 18752
rect 7323 18703 7365 18712
rect 4347 18668 4389 18677
rect 4347 18628 4348 18668
rect 4388 18628 4389 18668
rect 4347 18619 4389 18628
rect 1371 18584 1413 18593
rect 1371 18544 1372 18584
rect 1412 18544 1413 18584
rect 1371 18535 1413 18544
rect 2475 18584 2517 18593
rect 2475 18544 2476 18584
rect 2516 18544 2517 18584
rect 2475 18535 2517 18544
rect 4059 18584 4101 18593
rect 4059 18544 4060 18584
rect 4100 18544 4101 18584
rect 3906 18533 3952 18542
rect 4059 18535 4101 18544
rect 4587 18584 4629 18593
rect 4587 18544 4588 18584
rect 4628 18544 4629 18584
rect 4587 18535 4629 18544
rect 4971 18584 5013 18593
rect 4971 18544 4972 18584
rect 5012 18544 5013 18584
rect 4971 18535 5013 18544
rect 7083 18584 7125 18593
rect 7083 18544 7084 18584
rect 7124 18544 7125 18584
rect 7083 18535 7125 18544
rect 7467 18584 7509 18593
rect 7467 18544 7468 18584
rect 7508 18544 7509 18584
rect 7467 18535 7509 18544
rect 8523 18584 8565 18593
rect 8523 18544 8524 18584
rect 8564 18544 8565 18584
rect 8523 18535 8565 18544
rect 1162 18500 1220 18501
rect 1162 18460 1171 18500
rect 1211 18460 1220 18500
rect 1162 18459 1220 18460
rect 1978 18500 2036 18501
rect 1978 18460 1987 18500
rect 2027 18460 2036 18500
rect 1978 18459 2036 18460
rect 2091 18500 2133 18509
rect 2091 18460 2092 18500
rect 2132 18460 2133 18500
rect 2091 18451 2133 18460
rect 2571 18500 2613 18509
rect 2571 18460 2572 18500
rect 2612 18460 2613 18500
rect 2571 18451 2613 18460
rect 3043 18500 3101 18501
rect 3043 18460 3052 18500
rect 3092 18460 3101 18500
rect 3043 18459 3101 18460
rect 3531 18500 3589 18501
rect 3531 18460 3540 18500
rect 3580 18460 3589 18500
rect 3906 18493 3907 18533
rect 3947 18493 3952 18533
rect 3906 18484 3952 18493
rect 5451 18500 5493 18509
rect 3531 18459 3589 18460
rect 5451 18460 5452 18500
rect 5492 18460 5493 18500
rect 5451 18451 5493 18460
rect 6691 18500 6749 18501
rect 6691 18460 6700 18500
rect 6740 18460 6749 18500
rect 6691 18459 6749 18460
rect 8026 18500 8084 18501
rect 8026 18460 8035 18500
rect 8075 18460 8084 18500
rect 8026 18459 8084 18460
rect 8139 18500 8181 18509
rect 8139 18460 8140 18500
rect 8180 18460 8181 18500
rect 8139 18451 8181 18460
rect 8619 18500 8661 18509
rect 8619 18460 8620 18500
rect 8660 18460 8661 18500
rect 8619 18451 8661 18460
rect 9091 18500 9149 18501
rect 9091 18460 9100 18500
rect 9140 18460 9149 18500
rect 9091 18459 9149 18460
rect 9610 18500 9668 18501
rect 9610 18460 9619 18500
rect 9659 18460 9668 18500
rect 9610 18459 9668 18460
rect 9898 18500 9956 18501
rect 9898 18460 9907 18500
rect 9947 18460 9956 18500
rect 9898 18459 9956 18460
rect 3723 18332 3765 18341
rect 3723 18292 3724 18332
rect 3764 18292 3765 18332
rect 3723 18283 3765 18292
rect 4731 18332 4773 18341
rect 4731 18292 4732 18332
rect 4772 18292 4773 18332
rect 4731 18283 4773 18292
rect 5242 18332 5300 18333
rect 5242 18292 5251 18332
rect 5291 18292 5300 18332
rect 5242 18291 5300 18292
rect 6891 18332 6933 18341
rect 6891 18292 6892 18332
rect 6932 18292 6933 18332
rect 6891 18283 6933 18292
rect 7450 18332 7508 18333
rect 7450 18292 7459 18332
rect 7499 18292 7508 18332
rect 7450 18291 7508 18292
rect 9771 18332 9813 18341
rect 9771 18292 9772 18332
rect 9812 18292 9813 18332
rect 9771 18283 9813 18292
rect 10107 18332 10149 18341
rect 10107 18292 10108 18332
rect 10148 18292 10149 18332
rect 10107 18283 10149 18292
rect 1152 18164 10656 18188
rect 1152 18124 4928 18164
rect 4968 18124 5010 18164
rect 5050 18124 5092 18164
rect 5132 18124 5174 18164
rect 5214 18124 5256 18164
rect 5296 18124 10656 18164
rect 1152 18100 10656 18124
rect 3627 17996 3669 18005
rect 3627 17956 3628 17996
rect 3668 17956 3669 17996
rect 3627 17947 3669 17956
rect 6219 17996 6261 18005
rect 6219 17956 6220 17996
rect 6260 17956 6261 17996
rect 6219 17947 6261 17956
rect 9483 17996 9525 18005
rect 9483 17956 9484 17996
rect 9524 17956 9525 17996
rect 9483 17947 9525 17956
rect 10587 17996 10629 18005
rect 10587 17956 10588 17996
rect 10628 17956 10629 17996
rect 10587 17947 10629 17956
rect 1371 17912 1413 17921
rect 1371 17872 1372 17912
rect 1412 17872 1413 17912
rect 1371 17863 1413 17872
rect 1882 17828 1940 17829
rect 1218 17819 1264 17828
rect 1218 17779 1219 17819
rect 1259 17779 1264 17819
rect 1882 17788 1891 17828
rect 1931 17788 1940 17828
rect 1882 17787 1940 17788
rect 1995 17828 2037 17837
rect 1995 17788 1996 17828
rect 2036 17788 2037 17828
rect 1995 17779 2037 17788
rect 2379 17828 2421 17837
rect 3915 17828 3957 17837
rect 2379 17788 2380 17828
rect 2420 17788 2421 17828
rect 2379 17779 2421 17788
rect 2955 17819 2997 17828
rect 2955 17779 2956 17819
rect 2996 17779 2997 17819
rect 1218 17770 1264 17779
rect 2955 17770 2997 17779
rect 3435 17819 3477 17828
rect 3435 17779 3436 17819
rect 3476 17779 3477 17819
rect 3915 17788 3916 17828
rect 3956 17788 3957 17828
rect 3915 17779 3957 17788
rect 4090 17828 4148 17829
rect 4090 17788 4099 17828
rect 4139 17788 4148 17828
rect 4090 17787 4148 17788
rect 4203 17828 4245 17837
rect 4203 17788 4204 17828
rect 4244 17788 4245 17828
rect 4203 17779 4245 17788
rect 4474 17828 4532 17829
rect 4474 17788 4483 17828
rect 4523 17788 4532 17828
rect 4474 17787 4532 17788
rect 4587 17828 4629 17837
rect 4587 17788 4588 17828
rect 4628 17788 4629 17828
rect 4587 17779 4629 17788
rect 4971 17828 5013 17837
rect 7738 17828 7796 17829
rect 4971 17788 4972 17828
rect 5012 17788 5013 17828
rect 4971 17779 5013 17788
rect 5547 17819 5589 17828
rect 5547 17779 5548 17819
rect 5588 17779 5589 17819
rect 3435 17770 3477 17779
rect 5547 17770 5589 17779
rect 6027 17819 6069 17828
rect 6027 17779 6028 17819
rect 6068 17779 6069 17819
rect 7738 17788 7747 17828
rect 7787 17788 7796 17828
rect 7738 17787 7796 17788
rect 7851 17828 7893 17837
rect 7851 17788 7852 17828
rect 7892 17788 7893 17828
rect 7851 17779 7893 17788
rect 8235 17828 8277 17837
rect 8235 17788 8236 17828
rect 8276 17788 8277 17828
rect 8235 17779 8277 17788
rect 8811 17819 8853 17828
rect 8811 17779 8812 17819
rect 8852 17779 8853 17819
rect 6027 17770 6069 17779
rect 8811 17770 8853 17779
rect 9291 17819 9333 17828
rect 9291 17779 9292 17819
rect 9332 17779 9333 17819
rect 9291 17770 9333 17779
rect 2475 17744 2517 17753
rect 2475 17704 2476 17744
rect 2516 17704 2517 17744
rect 2475 17695 2517 17704
rect 5067 17744 5109 17753
rect 5067 17704 5068 17744
rect 5108 17704 5109 17744
rect 5067 17695 5109 17704
rect 6411 17744 6453 17753
rect 6411 17704 6412 17744
rect 6452 17704 6453 17744
rect 6411 17695 6453 17704
rect 8331 17744 8373 17753
rect 8331 17704 8332 17744
rect 8372 17704 8373 17744
rect 8331 17695 8373 17704
rect 9867 17744 9909 17753
rect 9867 17704 9868 17744
rect 9908 17704 9909 17744
rect 9867 17695 9909 17704
rect 10347 17744 10389 17753
rect 10347 17704 10348 17744
rect 10388 17704 10389 17744
rect 10347 17695 10389 17704
rect 4203 17576 4245 17585
rect 4203 17536 4204 17576
rect 4244 17536 4245 17576
rect 4203 17527 4245 17536
rect 9627 17576 9669 17585
rect 9627 17536 9628 17576
rect 9668 17536 9669 17576
rect 9627 17527 9669 17536
rect 1152 17408 10656 17432
rect 1152 17368 3688 17408
rect 3728 17368 3770 17408
rect 3810 17368 3852 17408
rect 3892 17368 3934 17408
rect 3974 17368 4016 17408
rect 4056 17368 10656 17408
rect 1152 17344 10656 17368
rect 5242 17240 5300 17241
rect 5242 17200 5251 17240
rect 5291 17200 5300 17240
rect 5242 17199 5300 17200
rect 9291 17240 9333 17249
rect 9291 17200 9292 17240
rect 9332 17200 9333 17240
rect 9291 17191 9333 17200
rect 10587 17240 10629 17249
rect 10587 17200 10588 17240
rect 10628 17200 10629 17240
rect 10587 17191 10629 17200
rect 3147 17156 3189 17165
rect 3147 17116 3148 17156
rect 3188 17116 3189 17156
rect 3147 17107 3189 17116
rect 4587 17156 4629 17165
rect 4587 17116 4588 17156
rect 4628 17116 4629 17156
rect 4587 17107 4629 17116
rect 3898 17072 3956 17073
rect 3898 17032 3907 17072
rect 3947 17032 3956 17072
rect 3898 17031 3956 17032
rect 4107 17072 4149 17081
rect 4107 17032 4108 17072
rect 4148 17032 4149 17072
rect 4107 17023 4149 17032
rect 6507 17072 6549 17081
rect 6507 17032 6508 17072
rect 6548 17032 6549 17072
rect 6507 17023 6549 17032
rect 10155 17072 10197 17081
rect 10155 17032 10156 17072
rect 10196 17032 10197 17072
rect 10155 17023 10197 17032
rect 10347 17072 10389 17081
rect 10347 17032 10348 17072
rect 10388 17032 10389 17072
rect 10347 17023 10389 17032
rect 1162 16988 1220 16989
rect 1162 16948 1171 16988
rect 1211 16948 1220 16988
rect 1162 16947 1220 16948
rect 1707 16988 1749 16997
rect 1707 16948 1708 16988
rect 1748 16948 1749 16988
rect 1707 16939 1749 16948
rect 2947 16988 3005 16989
rect 2947 16948 2956 16988
rect 2996 16948 3005 16988
rect 2947 16947 3005 16948
rect 3286 16988 3328 16997
rect 3286 16948 3287 16988
rect 3327 16948 3328 16988
rect 3286 16939 3328 16948
rect 3418 16988 3476 16989
rect 3418 16948 3427 16988
rect 3467 16948 3476 16988
rect 3418 16947 3476 16948
rect 3531 16988 3573 16997
rect 3531 16948 3532 16988
rect 3572 16948 3573 16988
rect 3531 16939 3573 16948
rect 3766 16988 3808 16997
rect 3766 16948 3767 16988
rect 3807 16948 3808 16988
rect 3766 16939 3808 16948
rect 4011 16988 4053 16997
rect 4011 16948 4012 16988
rect 4052 16948 4053 16988
rect 4011 16939 4053 16948
rect 4282 16988 4340 16989
rect 4282 16948 4291 16988
rect 4331 16948 4340 16988
rect 4282 16947 4340 16948
rect 4587 16988 4629 16997
rect 4587 16948 4588 16988
rect 4628 16948 4629 16988
rect 4587 16939 4629 16948
rect 4779 16988 4821 16997
rect 4779 16948 4780 16988
rect 4820 16948 4821 16988
rect 4779 16939 4821 16948
rect 4893 16988 4951 16989
rect 4893 16948 4902 16988
rect 4942 16948 4951 16988
rect 4893 16947 4951 16948
rect 5020 16988 5078 16989
rect 5020 16948 5029 16988
rect 5069 16948 5078 16988
rect 5020 16947 5078 16948
rect 5245 16988 5287 16997
rect 5245 16948 5246 16988
rect 5286 16948 5287 16988
rect 5245 16939 5287 16948
rect 5539 16988 5597 16989
rect 5539 16948 5548 16988
rect 5588 16948 5597 16988
rect 5539 16947 5597 16948
rect 5770 16988 5828 16989
rect 5770 16948 5779 16988
rect 5819 16948 5828 16988
rect 5770 16947 5828 16948
rect 5873 16988 5931 16989
rect 5873 16948 5882 16988
rect 5922 16948 5931 16988
rect 5873 16947 5931 16948
rect 7183 16988 7241 16989
rect 7183 16948 7192 16988
rect 7232 16948 7241 16988
rect 7183 16947 7241 16948
rect 7321 16988 7379 16989
rect 7321 16948 7330 16988
rect 7370 16948 7379 16988
rect 7321 16947 7379 16948
rect 7851 16988 7893 16997
rect 7851 16948 7852 16988
rect 7892 16948 7893 16988
rect 7851 16939 7893 16948
rect 9091 16988 9149 16989
rect 9091 16948 9100 16988
rect 9140 16948 9149 16988
rect 9091 16947 9149 16948
rect 9418 16988 9476 16989
rect 9418 16948 9427 16988
rect 9467 16948 9476 16988
rect 9418 16947 9476 16948
rect 6267 16904 6309 16913
rect 6267 16864 6268 16904
rect 6308 16864 6309 16904
rect 6267 16855 6309 16864
rect 9627 16904 9669 16913
rect 9627 16864 9628 16904
rect 9668 16864 9669 16904
rect 9627 16855 9669 16864
rect 1371 16820 1413 16829
rect 1371 16780 1372 16820
rect 1412 16780 1413 16820
rect 1371 16771 1413 16780
rect 3610 16820 3668 16821
rect 3610 16780 3619 16820
rect 3659 16780 3668 16820
rect 3610 16779 3668 16780
rect 5067 16820 5109 16829
rect 5067 16780 5068 16820
rect 5108 16780 5109 16820
rect 5067 16771 5109 16780
rect 5451 16820 5493 16829
rect 5451 16780 5452 16820
rect 5492 16780 5493 16820
rect 5451 16771 5493 16780
rect 6027 16820 6069 16829
rect 6027 16780 6028 16820
rect 6068 16780 6069 16820
rect 6027 16771 6069 16780
rect 7018 16820 7076 16821
rect 7018 16780 7027 16820
rect 7067 16780 7076 16820
rect 7018 16779 7076 16780
rect 7515 16820 7557 16829
rect 7515 16780 7516 16820
rect 7556 16780 7557 16820
rect 7515 16771 7557 16780
rect 9915 16820 9957 16829
rect 9915 16780 9916 16820
rect 9956 16780 9957 16820
rect 9915 16771 9957 16780
rect 1152 16652 10656 16676
rect 1152 16612 4928 16652
rect 4968 16612 5010 16652
rect 5050 16612 5092 16652
rect 5132 16612 5174 16652
rect 5214 16612 5256 16652
rect 5296 16612 10656 16652
rect 1152 16588 10656 16612
rect 4090 16484 4148 16485
rect 4090 16444 4099 16484
rect 4139 16444 4148 16484
rect 4090 16443 4148 16444
rect 5050 16484 5108 16485
rect 5050 16444 5059 16484
rect 5099 16444 5108 16484
rect 5050 16443 5108 16444
rect 5451 16484 5493 16493
rect 5451 16444 5452 16484
rect 5492 16444 5493 16484
rect 5451 16435 5493 16444
rect 9579 16484 9621 16493
rect 9579 16444 9580 16484
rect 9620 16444 9621 16484
rect 9579 16435 9621 16444
rect 3243 16400 3285 16409
rect 3243 16360 3244 16400
rect 3284 16360 3285 16400
rect 3243 16351 3285 16360
rect 9850 16400 9908 16401
rect 9850 16360 9859 16400
rect 9899 16360 9908 16400
rect 9850 16359 9908 16360
rect 1803 16316 1845 16325
rect 3915 16316 3957 16325
rect 1218 16307 1264 16316
rect 1218 16267 1219 16307
rect 1259 16267 1264 16307
rect 1803 16276 1804 16316
rect 1844 16276 1845 16316
rect 1803 16267 1845 16276
rect 3051 16307 3093 16316
rect 3051 16267 3052 16307
rect 3092 16267 3093 16307
rect 3915 16276 3916 16316
rect 3956 16276 3957 16316
rect 3915 16267 3957 16276
rect 4106 16316 4148 16325
rect 4106 16276 4107 16316
rect 4147 16276 4148 16316
rect 4106 16267 4148 16276
rect 4258 16316 4316 16317
rect 4258 16276 4267 16316
rect 4307 16276 4316 16316
rect 4258 16275 4316 16276
rect 4491 16316 4533 16325
rect 4491 16276 4492 16316
rect 4532 16276 4533 16316
rect 4491 16267 4533 16276
rect 4731 16316 4773 16325
rect 4731 16276 4732 16316
rect 4772 16276 4773 16316
rect 4731 16267 4773 16276
rect 4858 16316 4916 16317
rect 4858 16276 4867 16316
rect 4907 16276 4916 16316
rect 4858 16275 4916 16276
rect 4971 16316 5013 16325
rect 6891 16316 6933 16325
rect 4971 16276 4972 16316
rect 5012 16276 5013 16316
rect 4971 16267 5013 16276
rect 5643 16307 5685 16316
rect 5643 16267 5644 16307
rect 5684 16267 5685 16307
rect 6891 16276 6892 16316
rect 6932 16276 6933 16316
rect 6891 16267 6933 16276
rect 7834 16316 7892 16317
rect 7834 16276 7843 16316
rect 7883 16276 7892 16316
rect 7834 16275 7892 16276
rect 7947 16316 7989 16325
rect 7947 16276 7948 16316
rect 7988 16276 7989 16316
rect 7947 16267 7989 16276
rect 8331 16316 8373 16325
rect 10251 16316 10293 16325
rect 8331 16276 8332 16316
rect 8372 16276 8373 16316
rect 8331 16267 8373 16276
rect 8907 16307 8949 16316
rect 8907 16267 8908 16307
rect 8948 16267 8949 16307
rect 1218 16258 1264 16267
rect 3051 16258 3093 16267
rect 5643 16258 5685 16267
rect 8907 16258 8949 16267
rect 9387 16307 9429 16316
rect 9387 16267 9388 16307
rect 9428 16267 9429 16307
rect 10251 16276 10252 16316
rect 10292 16276 10293 16316
rect 10251 16267 10293 16276
rect 9387 16258 9429 16267
rect 1371 16232 1413 16241
rect 1371 16192 1372 16232
rect 1412 16192 1413 16232
rect 1371 16183 1413 16192
rect 3627 16232 3669 16241
rect 3627 16192 3628 16232
rect 3668 16192 3669 16232
rect 3627 16183 3669 16192
rect 4378 16232 4436 16233
rect 4378 16192 4387 16232
rect 4427 16192 4436 16232
rect 4378 16191 4436 16192
rect 4587 16232 4629 16241
rect 4587 16192 4588 16232
rect 4628 16192 4629 16232
rect 4587 16183 4629 16192
rect 8427 16232 8469 16241
rect 8427 16192 8428 16232
rect 8468 16192 8469 16232
rect 8427 16183 8469 16192
rect 3387 16148 3429 16157
rect 3387 16108 3388 16148
rect 3428 16108 3429 16148
rect 3387 16099 3429 16108
rect 1152 15896 10656 15920
rect 1152 15856 3688 15896
rect 3728 15856 3770 15896
rect 3810 15856 3852 15896
rect 3892 15856 3934 15896
rect 3974 15856 4016 15896
rect 4056 15856 10656 15896
rect 1152 15832 10656 15856
rect 2667 15728 2709 15737
rect 2667 15688 2668 15728
rect 2708 15688 2709 15728
rect 2667 15679 2709 15688
rect 3195 15728 3237 15737
rect 3195 15688 3196 15728
rect 3236 15688 3237 15728
rect 3195 15679 3237 15688
rect 7563 15728 7605 15737
rect 7563 15688 7564 15728
rect 7604 15688 7605 15728
rect 7563 15679 7605 15688
rect 9771 15728 9813 15737
rect 9771 15688 9772 15728
rect 9812 15688 9813 15728
rect 9771 15679 9813 15688
rect 10587 15728 10629 15737
rect 10587 15688 10588 15728
rect 10628 15688 10629 15728
rect 10587 15679 10629 15688
rect 2811 15644 2853 15653
rect 2811 15604 2812 15644
rect 2852 15604 2853 15644
rect 2811 15595 2853 15604
rect 4731 15644 4773 15653
rect 4731 15604 4732 15644
rect 4772 15604 4773 15644
rect 4731 15595 4773 15604
rect 3051 15560 3093 15569
rect 3051 15520 3052 15560
rect 3092 15520 3093 15560
rect 3051 15511 3093 15520
rect 3435 15560 3477 15569
rect 3435 15520 3436 15560
rect 3476 15520 3477 15560
rect 3435 15511 3477 15520
rect 3819 15560 3861 15569
rect 3819 15520 3820 15560
rect 3860 15520 3861 15560
rect 3819 15511 3861 15520
rect 4203 15560 4245 15569
rect 4203 15520 4204 15560
rect 4244 15520 4245 15560
rect 4203 15511 4245 15520
rect 4587 15560 4629 15569
rect 4587 15520 4588 15560
rect 4628 15520 4629 15560
rect 4587 15511 4629 15520
rect 4971 15560 5013 15569
rect 4971 15520 4972 15560
rect 5012 15520 5013 15560
rect 4971 15511 5013 15520
rect 10155 15560 10197 15569
rect 10155 15520 10156 15560
rect 10196 15520 10197 15560
rect 10155 15511 10197 15520
rect 10347 15560 10389 15569
rect 10347 15520 10348 15560
rect 10388 15520 10389 15560
rect 10347 15511 10389 15520
rect 1227 15476 1269 15485
rect 1227 15436 1228 15476
rect 1268 15436 1269 15476
rect 1227 15427 1269 15436
rect 2467 15476 2525 15477
rect 2467 15436 2476 15476
rect 2516 15436 2525 15476
rect 2467 15435 2525 15436
rect 5259 15476 5301 15485
rect 5259 15436 5260 15476
rect 5300 15436 5301 15476
rect 5259 15427 5301 15436
rect 6123 15476 6165 15485
rect 6123 15436 6124 15476
rect 6164 15436 6165 15476
rect 6123 15427 6165 15436
rect 7363 15476 7421 15477
rect 7363 15436 7372 15476
rect 7412 15436 7421 15476
rect 7363 15435 7421 15436
rect 8331 15476 8373 15485
rect 8331 15436 8332 15476
rect 8372 15436 8373 15476
rect 8331 15427 8373 15436
rect 9571 15476 9629 15477
rect 9571 15436 9580 15476
rect 9620 15436 9629 15476
rect 9571 15435 9629 15436
rect 3579 15392 3621 15401
rect 3579 15352 3580 15392
rect 3620 15352 3621 15392
rect 3579 15343 3621 15352
rect 3963 15308 4005 15317
rect 3963 15268 3964 15308
rect 4004 15268 4005 15308
rect 3963 15259 4005 15268
rect 4347 15308 4389 15317
rect 4347 15268 4348 15308
rect 4388 15268 4389 15308
rect 4347 15259 4389 15268
rect 5115 15308 5157 15317
rect 5115 15268 5116 15308
rect 5156 15268 5157 15308
rect 5115 15259 5157 15268
rect 9915 15308 9957 15317
rect 9915 15268 9916 15308
rect 9956 15268 9957 15308
rect 9915 15259 9957 15268
rect 1152 15140 10656 15164
rect 1152 15100 4928 15140
rect 4968 15100 5010 15140
rect 5050 15100 5092 15140
rect 5132 15100 5174 15140
rect 5214 15100 5256 15140
rect 5296 15100 10656 15140
rect 1152 15076 10656 15100
rect 1563 14972 1605 14981
rect 1563 14932 1564 14972
rect 1604 14932 1605 14972
rect 1563 14923 1605 14932
rect 4203 14972 4245 14981
rect 4203 14932 4204 14972
rect 4244 14932 4245 14972
rect 4203 14923 4245 14932
rect 4491 14972 4533 14981
rect 4491 14932 4492 14972
rect 4532 14932 4533 14972
rect 4491 14923 4533 14932
rect 10587 14972 10629 14981
rect 10587 14932 10588 14972
rect 10628 14932 10629 14972
rect 10587 14923 10629 14932
rect 1947 14888 1989 14897
rect 1947 14848 1948 14888
rect 1988 14848 1989 14888
rect 1947 14839 1989 14848
rect 7563 14888 7605 14897
rect 7563 14848 7564 14888
rect 7604 14848 7605 14888
rect 7563 14839 7605 14848
rect 2458 14804 2516 14805
rect 2458 14764 2467 14804
rect 2507 14764 2516 14804
rect 2458 14763 2516 14764
rect 2571 14804 2613 14813
rect 2571 14764 2572 14804
rect 2612 14764 2613 14804
rect 2571 14755 2613 14764
rect 2955 14804 2997 14813
rect 5931 14804 5973 14813
rect 2955 14764 2956 14804
rect 2996 14764 2997 14804
rect 2955 14755 2997 14764
rect 3531 14795 3573 14804
rect 3531 14755 3532 14795
rect 3572 14755 3573 14795
rect 3531 14746 3573 14755
rect 4011 14795 4053 14804
rect 4011 14755 4012 14795
rect 4052 14755 4053 14795
rect 4011 14746 4053 14755
rect 4683 14795 4725 14804
rect 4683 14755 4684 14795
rect 4724 14755 4725 14795
rect 5931 14764 5932 14804
rect 5972 14764 5973 14804
rect 5931 14755 5973 14764
rect 6123 14804 6165 14813
rect 7834 14804 7892 14805
rect 6123 14764 6124 14804
rect 6164 14764 6165 14804
rect 6123 14755 6165 14764
rect 7371 14795 7413 14804
rect 7371 14755 7372 14795
rect 7412 14755 7413 14795
rect 7834 14764 7843 14804
rect 7883 14764 7892 14804
rect 7834 14763 7892 14764
rect 7947 14804 7989 14813
rect 7947 14764 7948 14804
rect 7988 14764 7989 14804
rect 7947 14755 7989 14764
rect 8331 14804 8373 14813
rect 8331 14764 8332 14804
rect 8372 14764 8373 14804
rect 8331 14755 8373 14764
rect 8907 14795 8949 14804
rect 8907 14755 8908 14795
rect 8948 14755 8949 14795
rect 4683 14746 4725 14755
rect 7371 14746 7413 14755
rect 8907 14746 8949 14755
rect 9387 14795 9429 14804
rect 9387 14755 9388 14795
rect 9428 14755 9429 14795
rect 9387 14746 9429 14755
rect 1227 14720 1269 14729
rect 1227 14680 1228 14720
rect 1268 14680 1269 14720
rect 1227 14671 1269 14680
rect 1803 14720 1845 14729
rect 1803 14680 1804 14720
rect 1844 14680 1845 14720
rect 1803 14671 1845 14680
rect 2187 14720 2229 14729
rect 2187 14680 2188 14720
rect 2228 14680 2229 14720
rect 2187 14671 2229 14680
rect 3051 14720 3093 14729
rect 3051 14680 3052 14720
rect 3092 14680 3093 14720
rect 3051 14671 3093 14680
rect 8427 14720 8469 14729
rect 8427 14680 8428 14720
rect 8468 14680 8469 14720
rect 8427 14671 8469 14680
rect 9610 14720 9668 14721
rect 9610 14680 9619 14720
rect 9659 14680 9668 14720
rect 9610 14679 9668 14680
rect 9963 14720 10005 14729
rect 9963 14680 9964 14720
rect 10004 14680 10005 14720
rect 9963 14671 10005 14680
rect 10347 14720 10389 14729
rect 10347 14680 10348 14720
rect 10388 14680 10389 14720
rect 10347 14671 10389 14680
rect 1467 14552 1509 14561
rect 1467 14512 1468 14552
rect 1508 14512 1509 14552
rect 1467 14503 1509 14512
rect 9723 14552 9765 14561
rect 9723 14512 9724 14552
rect 9764 14512 9765 14552
rect 9723 14503 9765 14512
rect 1152 14384 10656 14408
rect 1152 14344 3688 14384
rect 3728 14344 3770 14384
rect 3810 14344 3852 14384
rect 3892 14344 3934 14384
rect 3974 14344 4016 14384
rect 4056 14344 10656 14384
rect 1152 14320 10656 14344
rect 4827 14216 4869 14225
rect 4827 14176 4828 14216
rect 4868 14176 4869 14216
rect 4827 14167 4869 14176
rect 5787 14216 5829 14225
rect 5787 14176 5788 14216
rect 5828 14176 5829 14216
rect 5787 14167 5829 14176
rect 9195 14216 9237 14225
rect 9195 14176 9196 14216
rect 9236 14176 9237 14216
rect 9195 14167 9237 14176
rect 10587 14216 10629 14225
rect 10587 14176 10588 14216
rect 10628 14176 10629 14216
rect 10587 14167 10629 14176
rect 1179 14132 1221 14141
rect 1179 14092 1180 14132
rect 1220 14092 1221 14132
rect 1179 14083 1221 14092
rect 6267 14132 6309 14141
rect 6267 14092 6268 14132
rect 6308 14092 6309 14132
rect 6267 14083 6309 14092
rect 10203 14132 10245 14141
rect 10203 14092 10204 14132
rect 10244 14092 10245 14132
rect 10203 14083 10245 14092
rect 1419 14048 1461 14057
rect 1419 14008 1420 14048
rect 1460 14008 1461 14048
rect 1419 13999 1461 14008
rect 1803 14048 1845 14057
rect 1803 14008 1804 14048
rect 1844 14008 1845 14048
rect 1803 13999 1845 14008
rect 2187 14048 2229 14057
rect 2187 14008 2188 14048
rect 2228 14008 2229 14048
rect 2187 13999 2229 14008
rect 3051 14048 3093 14057
rect 3051 14008 3052 14048
rect 3092 14008 3093 14048
rect 3051 13999 3093 14008
rect 4330 14048 4388 14049
rect 4330 14008 4339 14048
rect 4379 14008 4388 14048
rect 4330 14007 4388 14008
rect 4683 14048 4725 14057
rect 4683 14008 4684 14048
rect 4724 14008 4725 14048
rect 4683 13999 4725 14008
rect 5067 14048 5109 14057
rect 5067 14008 5068 14048
rect 5108 14008 5109 14048
rect 5067 13999 5109 14008
rect 5547 14048 5589 14057
rect 5547 14008 5548 14048
rect 5588 14008 5589 14048
rect 5547 13999 5589 14008
rect 6027 14048 6069 14057
rect 6027 14008 6028 14048
rect 6068 14008 6069 14048
rect 6027 13999 6069 14008
rect 9531 14048 9573 14057
rect 9531 14008 9532 14048
rect 9572 14008 9573 14048
rect 9531 13999 9573 14008
rect 9963 14048 10005 14057
rect 9963 14008 9964 14048
rect 10004 14008 10005 14048
rect 9963 13999 10005 14008
rect 10347 14048 10389 14057
rect 10347 14008 10348 14048
rect 10388 14008 10389 14048
rect 10347 13999 10389 14008
rect 2554 13964 2612 13965
rect 2554 13924 2563 13964
rect 2603 13924 2612 13964
rect 2554 13923 2612 13924
rect 2667 13964 2709 13973
rect 2667 13924 2668 13964
rect 2708 13924 2709 13964
rect 2667 13915 2709 13924
rect 3147 13964 3189 13973
rect 3147 13924 3148 13964
rect 3188 13924 3189 13964
rect 3147 13915 3189 13924
rect 3619 13964 3677 13965
rect 3619 13924 3628 13964
rect 3668 13924 3677 13964
rect 3619 13923 3677 13924
rect 4138 13964 4196 13965
rect 4138 13924 4147 13964
rect 4187 13924 4196 13964
rect 4138 13923 4196 13924
rect 7210 13964 7268 13965
rect 7210 13924 7219 13964
rect 7259 13924 7268 13964
rect 7210 13923 7268 13924
rect 7755 13964 7797 13973
rect 7755 13924 7756 13964
rect 7796 13924 7797 13964
rect 7755 13915 7797 13924
rect 8995 13964 9053 13965
rect 8995 13924 9004 13964
rect 9044 13924 9053 13964
rect 8995 13923 9053 13924
rect 9367 13964 9425 13965
rect 9367 13924 9376 13964
rect 9416 13924 9425 13964
rect 9367 13923 9425 13924
rect 1947 13880 1989 13889
rect 1947 13840 1948 13880
rect 1988 13840 1989 13880
rect 1947 13831 1989 13840
rect 1563 13796 1605 13805
rect 1563 13756 1564 13796
rect 1604 13756 1605 13796
rect 1563 13747 1605 13756
rect 4443 13796 4485 13805
rect 4443 13756 4444 13796
rect 4484 13756 4485 13796
rect 4443 13747 4485 13756
rect 7419 13796 7461 13805
rect 7419 13756 7420 13796
rect 7460 13756 7461 13796
rect 7419 13747 7461 13756
rect 1152 13628 10656 13652
rect 1152 13588 4928 13628
rect 4968 13588 5010 13628
rect 5050 13588 5092 13628
rect 5132 13588 5174 13628
rect 5214 13588 5256 13628
rect 5296 13588 10656 13628
rect 1152 13564 10656 13588
rect 2859 13460 2901 13469
rect 2859 13420 2860 13460
rect 2900 13420 2901 13460
rect 2859 13411 2901 13420
rect 4491 13460 4533 13469
rect 4491 13420 4492 13460
rect 4532 13420 4533 13460
rect 4491 13411 4533 13420
rect 6123 13376 6165 13385
rect 6123 13336 6124 13376
rect 6164 13336 6165 13376
rect 6123 13327 6165 13336
rect 7371 13376 7413 13385
rect 7371 13336 7372 13376
rect 7412 13336 7413 13376
rect 7371 13327 7413 13336
rect 10251 13376 10293 13385
rect 10251 13336 10252 13376
rect 10292 13336 10293 13376
rect 10251 13327 10293 13336
rect 1419 13292 1461 13301
rect 3051 13292 3093 13301
rect 4683 13292 4725 13301
rect 6987 13292 7029 13301
rect 1419 13252 1420 13292
rect 1460 13252 1461 13292
rect 1419 13243 1461 13252
rect 2667 13283 2709 13292
rect 2667 13243 2668 13283
rect 2708 13243 2709 13283
rect 3051 13252 3052 13292
rect 3092 13252 3093 13292
rect 3051 13243 3093 13252
rect 4299 13283 4341 13292
rect 4299 13243 4300 13283
rect 4340 13243 4341 13283
rect 4683 13252 4684 13292
rect 4724 13252 4725 13292
rect 4683 13243 4725 13252
rect 5931 13283 5973 13292
rect 5931 13243 5932 13283
rect 5972 13243 5973 13283
rect 6987 13252 6988 13292
rect 7028 13252 7029 13292
rect 6987 13243 7029 13252
rect 7258 13292 7316 13293
rect 7258 13252 7267 13292
rect 7307 13252 7316 13292
rect 7258 13251 7316 13252
rect 8811 13292 8853 13301
rect 8811 13252 8812 13292
rect 8852 13252 8853 13292
rect 8811 13243 8853 13252
rect 10059 13283 10101 13292
rect 10059 13243 10060 13283
rect 10100 13243 10101 13283
rect 2667 13234 2709 13243
rect 4299 13234 4341 13243
rect 5931 13234 5973 13243
rect 10059 13234 10101 13243
rect 8043 13208 8085 13217
rect 8043 13168 8044 13208
rect 8084 13168 8085 13208
rect 8043 13159 8085 13168
rect 8427 13208 8469 13217
rect 8427 13168 8428 13208
rect 8468 13168 8469 13208
rect 8427 13159 8469 13168
rect 7803 13124 7845 13133
rect 7803 13084 7804 13124
rect 7844 13084 7845 13124
rect 7803 13075 7845 13084
rect 8667 13124 8709 13133
rect 8667 13084 8668 13124
rect 8708 13084 8709 13124
rect 8667 13075 8709 13084
rect 7659 13040 7701 13049
rect 7659 13000 7660 13040
rect 7700 13000 7701 13040
rect 7659 12991 7701 13000
rect 1152 12872 10656 12896
rect 1152 12832 3688 12872
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 4056 12832 10656 12872
rect 1152 12808 10656 12832
rect 2859 12704 2901 12713
rect 2859 12664 2860 12704
rect 2900 12664 2901 12704
rect 2859 12655 2901 12664
rect 6075 12704 6117 12713
rect 6075 12664 6076 12704
rect 6116 12664 6117 12704
rect 6075 12655 6117 12664
rect 9099 12704 9141 12713
rect 9099 12664 9100 12704
rect 9140 12664 9141 12704
rect 9099 12655 9141 12664
rect 2667 12620 2709 12629
rect 2667 12580 2668 12620
rect 2708 12580 2709 12620
rect 2667 12571 2709 12580
rect 8907 12620 8949 12629
rect 8907 12580 8908 12620
rect 8948 12580 8949 12620
rect 8907 12571 8949 12580
rect 4683 12536 4725 12545
rect 4683 12496 4684 12536
rect 4724 12496 4725 12536
rect 4683 12487 4725 12496
rect 5067 12536 5109 12545
rect 5067 12496 5068 12536
rect 5108 12496 5109 12536
rect 5067 12487 5109 12496
rect 5451 12536 5493 12545
rect 5451 12496 5452 12536
rect 5492 12496 5493 12536
rect 5451 12487 5493 12496
rect 6315 12536 6357 12545
rect 6315 12496 6316 12536
rect 6356 12496 6357 12536
rect 6315 12487 6357 12496
rect 1227 12452 1269 12461
rect 1227 12412 1228 12452
rect 1268 12412 1269 12452
rect 1227 12403 1269 12412
rect 2467 12452 2525 12453
rect 2467 12412 2476 12452
rect 2516 12412 2525 12452
rect 2467 12411 2525 12412
rect 3043 12452 3101 12453
rect 3043 12412 3052 12452
rect 3092 12412 3101 12452
rect 3043 12411 3101 12412
rect 4299 12452 4341 12461
rect 4299 12412 4300 12452
rect 4340 12412 4341 12452
rect 4299 12403 4341 12412
rect 7213 12452 7271 12453
rect 7213 12412 7222 12452
rect 7262 12412 7271 12452
rect 7213 12411 7271 12412
rect 8074 12452 8132 12453
rect 8074 12412 8083 12452
rect 8123 12412 8132 12452
rect 8074 12411 8132 12412
rect 9283 12452 9341 12453
rect 9283 12412 9292 12452
rect 9332 12412 9341 12452
rect 9283 12411 9341 12412
rect 10539 12452 10581 12461
rect 10539 12412 10540 12452
rect 10580 12412 10581 12452
rect 10539 12403 10581 12412
rect 5211 12368 5253 12377
rect 5211 12328 5212 12368
rect 5252 12328 5253 12368
rect 5211 12319 5253 12328
rect 4443 12284 4485 12293
rect 4443 12244 4444 12284
rect 4484 12244 4485 12284
rect 4443 12235 4485 12244
rect 4827 12284 4869 12293
rect 4827 12244 4828 12284
rect 4868 12244 4869 12284
rect 4827 12235 4869 12244
rect 7018 12284 7076 12285
rect 7018 12244 7027 12284
rect 7067 12244 7076 12284
rect 7018 12243 7076 12244
rect 8283 12284 8325 12293
rect 8283 12244 8284 12284
rect 8324 12244 8325 12284
rect 8283 12235 8325 12244
rect 1152 12116 10656 12140
rect 1152 12076 4928 12116
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 5296 12076 10656 12116
rect 1152 12052 10656 12076
rect 2955 11948 2997 11957
rect 2955 11908 2956 11948
rect 2996 11908 2997 11948
rect 2955 11899 2997 11908
rect 3579 11948 3621 11957
rect 3579 11908 3580 11948
rect 3620 11908 3621 11948
rect 3579 11899 3621 11908
rect 5931 11948 5973 11957
rect 5931 11908 5932 11948
rect 5972 11908 5973 11948
rect 5931 11899 5973 11908
rect 7803 11948 7845 11957
rect 7803 11908 7804 11948
rect 7844 11908 7845 11948
rect 7803 11899 7845 11908
rect 10539 11948 10581 11957
rect 10539 11908 10540 11948
rect 10580 11908 10581 11948
rect 10539 11899 10581 11908
rect 1515 11780 1557 11789
rect 3469 11780 3527 11781
rect 1515 11740 1516 11780
rect 1556 11740 1557 11780
rect 1515 11731 1557 11740
rect 2763 11771 2805 11780
rect 2763 11731 2764 11771
rect 2804 11731 2805 11771
rect 3469 11740 3478 11780
rect 3518 11740 3527 11780
rect 3469 11739 3527 11740
rect 4173 11780 4215 11789
rect 4173 11740 4174 11780
rect 4214 11740 4215 11780
rect 4173 11731 4215 11740
rect 4299 11780 4341 11789
rect 4299 11740 4300 11780
rect 4340 11740 4341 11780
rect 4299 11731 4341 11740
rect 4683 11780 4725 11789
rect 6219 11780 6261 11789
rect 8602 11780 8660 11781
rect 4683 11740 4684 11780
rect 4724 11740 4725 11780
rect 4683 11731 4725 11740
rect 5259 11771 5301 11780
rect 5259 11731 5260 11771
rect 5300 11731 5301 11771
rect 2763 11722 2805 11731
rect 5259 11722 5301 11731
rect 5739 11771 5781 11780
rect 5739 11731 5740 11771
rect 5780 11731 5781 11771
rect 6219 11740 6220 11780
rect 6260 11740 6261 11780
rect 6219 11731 6261 11740
rect 7467 11771 7509 11780
rect 7467 11731 7468 11771
rect 7508 11731 7509 11771
rect 8602 11740 8611 11780
rect 8651 11740 8660 11780
rect 8602 11739 8660 11740
rect 5739 11722 5781 11731
rect 7467 11722 7509 11731
rect 3274 11696 3332 11697
rect 3274 11656 3283 11696
rect 3323 11656 3332 11696
rect 3274 11655 3332 11656
rect 3819 11696 3861 11705
rect 3819 11656 3820 11696
rect 3860 11656 3861 11696
rect 3819 11647 3861 11656
rect 4779 11696 4821 11705
rect 4779 11656 4780 11696
rect 4820 11656 4821 11696
rect 4779 11647 4821 11656
rect 8043 11696 8085 11705
rect 8043 11656 8044 11696
rect 8084 11656 8085 11696
rect 8043 11647 8085 11656
rect 8235 11696 8277 11705
rect 8235 11656 8236 11696
rect 8276 11656 8277 11696
rect 8235 11647 8277 11656
rect 7659 11528 7701 11537
rect 7659 11488 7660 11528
rect 7700 11488 7701 11528
rect 7659 11479 7701 11488
rect 1152 11360 10656 11384
rect 1152 11320 3688 11360
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 4056 11320 10656 11360
rect 1152 11296 10656 11320
rect 1179 11192 1221 11201
rect 1179 11152 1180 11192
rect 1220 11152 1221 11192
rect 1179 11143 1221 11152
rect 1563 11192 1605 11201
rect 1563 11152 1564 11192
rect 1604 11152 1605 11192
rect 1563 11143 1605 11152
rect 3627 11192 3669 11201
rect 3627 11152 3628 11192
rect 3668 11152 3669 11192
rect 3627 11143 3669 11152
rect 5835 11192 5877 11201
rect 5835 11152 5836 11192
rect 5876 11152 5877 11192
rect 5835 11143 5877 11152
rect 10539 11192 10581 11201
rect 10539 11152 10540 11192
rect 10580 11152 10581 11192
rect 10539 11143 10581 11152
rect 1419 11024 1461 11033
rect 1419 10984 1420 11024
rect 1460 10984 1461 11024
rect 1419 10975 1461 10984
rect 1803 11024 1845 11033
rect 1803 10984 1804 11024
rect 1844 10984 1845 11024
rect 1803 10975 1845 10984
rect 3819 11024 3861 11033
rect 3819 10984 3820 11024
rect 3860 10984 3861 11024
rect 3819 10975 3861 10984
rect 4059 11024 4101 11033
rect 4059 10984 4060 11024
rect 4100 10984 4101 11024
rect 4059 10975 4101 10984
rect 6699 11024 6741 11033
rect 6699 10984 6700 11024
rect 6740 10984 6741 11024
rect 6699 10975 6741 10984
rect 2187 10940 2229 10949
rect 2187 10900 2188 10940
rect 2228 10900 2229 10940
rect 2187 10891 2229 10900
rect 3427 10940 3485 10941
rect 3427 10900 3436 10940
rect 3476 10900 3485 10940
rect 3427 10899 3485 10900
rect 4395 10940 4437 10949
rect 4395 10900 4396 10940
rect 4436 10900 4437 10940
rect 4395 10891 4437 10900
rect 5635 10940 5693 10941
rect 5635 10900 5644 10940
rect 5684 10900 5693 10940
rect 5635 10899 5693 10900
rect 6202 10940 6260 10941
rect 6202 10900 6211 10940
rect 6251 10900 6260 10940
rect 6202 10899 6260 10900
rect 6315 10940 6357 10949
rect 6315 10900 6316 10940
rect 6356 10900 6357 10940
rect 6315 10891 6357 10900
rect 6795 10940 6837 10949
rect 6795 10900 6796 10940
rect 6836 10900 6837 10940
rect 6795 10891 6837 10900
rect 7267 10940 7325 10941
rect 7267 10900 7276 10940
rect 7316 10900 7325 10940
rect 7267 10899 7325 10900
rect 7755 10940 7813 10941
rect 7755 10900 7764 10940
rect 7804 10900 7813 10940
rect 7755 10899 7813 10900
rect 8602 10940 8660 10941
rect 8602 10900 8611 10940
rect 8651 10900 8660 10940
rect 8602 10899 8660 10900
rect 8218 10856 8276 10857
rect 8218 10816 8227 10856
rect 8267 10816 8276 10856
rect 8218 10815 8276 10816
rect 7947 10772 7989 10781
rect 7947 10732 7948 10772
rect 7988 10732 7989 10772
rect 7947 10723 7989 10732
rect 1152 10604 10656 10628
rect 1152 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 10656 10604
rect 1152 10540 10656 10564
rect 1179 10436 1221 10445
rect 1179 10396 1180 10436
rect 1220 10396 1221 10436
rect 1179 10387 1221 10396
rect 3723 10436 3765 10445
rect 3723 10396 3724 10436
rect 3764 10396 3765 10436
rect 3723 10387 3765 10396
rect 8379 10436 8421 10445
rect 8379 10396 8380 10436
rect 8420 10396 8421 10436
rect 8379 10387 8421 10396
rect 10203 10436 10245 10445
rect 10203 10396 10204 10436
rect 10244 10396 10245 10436
rect 10203 10387 10245 10396
rect 10587 10436 10629 10445
rect 10587 10396 10588 10436
rect 10628 10396 10629 10436
rect 10587 10387 10629 10396
rect 1563 10352 1605 10361
rect 1563 10312 1564 10352
rect 1604 10312 1605 10352
rect 1563 10303 1605 10312
rect 2283 10268 2325 10277
rect 4282 10268 4340 10269
rect 2283 10228 2284 10268
rect 2324 10228 2325 10268
rect 2283 10219 2325 10228
rect 3531 10259 3573 10268
rect 3531 10219 3532 10259
rect 3572 10219 3573 10259
rect 4282 10228 4291 10268
rect 4331 10228 4340 10268
rect 4282 10227 4340 10228
rect 4395 10268 4437 10277
rect 4395 10228 4396 10268
rect 4436 10228 4437 10268
rect 4395 10219 4437 10228
rect 4779 10268 4821 10277
rect 4779 10228 4780 10268
rect 4820 10228 4821 10268
rect 4779 10219 4821 10228
rect 5355 10259 5397 10268
rect 5355 10219 5356 10259
rect 5396 10219 5397 10259
rect 3531 10210 3573 10219
rect 5355 10210 5397 10219
rect 5835 10259 5877 10268
rect 5835 10219 5836 10259
rect 5876 10219 5877 10259
rect 5835 10210 5877 10219
rect 1419 10184 1461 10193
rect 1419 10144 1420 10184
rect 1460 10144 1461 10184
rect 1419 10135 1461 10144
rect 1803 10184 1845 10193
rect 1803 10144 1804 10184
rect 1844 10144 1845 10184
rect 1803 10135 1845 10144
rect 4875 10184 4917 10193
rect 4875 10144 4876 10184
rect 4916 10144 4917 10184
rect 4875 10135 4917 10144
rect 6058 10184 6116 10185
rect 6058 10144 6067 10184
rect 6107 10144 6116 10184
rect 6058 10143 6116 10144
rect 6411 10184 6453 10193
rect 6411 10144 6412 10184
rect 6452 10144 6453 10184
rect 6411 10135 6453 10144
rect 6795 10184 6837 10193
rect 6795 10144 6796 10184
rect 6836 10144 6837 10184
rect 6795 10135 6837 10144
rect 8235 10184 8277 10193
rect 8235 10144 8236 10184
rect 8276 10144 8277 10184
rect 8235 10135 8277 10144
rect 8619 10184 8661 10193
rect 8619 10144 8620 10184
rect 8660 10144 8661 10184
rect 8619 10135 8661 10144
rect 8907 10184 8949 10193
rect 8907 10144 8908 10184
rect 8948 10144 8949 10184
rect 8907 10135 8949 10144
rect 9147 10184 9189 10193
rect 9147 10144 9148 10184
rect 9188 10144 9189 10184
rect 9147 10135 9189 10144
rect 9963 10184 10005 10193
rect 9963 10144 9964 10184
rect 10004 10144 10005 10184
rect 9963 10135 10005 10144
rect 10347 10184 10389 10193
rect 10347 10144 10348 10184
rect 10388 10144 10389 10184
rect 10347 10135 10389 10144
rect 6171 10100 6213 10109
rect 6171 10060 6172 10100
rect 6212 10060 6213 10100
rect 6171 10051 6213 10060
rect 7995 10100 8037 10109
rect 7995 10060 7996 10100
rect 8036 10060 8037 10100
rect 7995 10051 8037 10060
rect 9291 10100 9333 10109
rect 9291 10060 9292 10100
rect 9332 10060 9333 10100
rect 9291 10051 9333 10060
rect 6555 10016 6597 10025
rect 6555 9976 6556 10016
rect 6596 9976 6597 10016
rect 6555 9967 6597 9976
rect 1152 9848 10656 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 10656 9848
rect 1152 9784 10656 9808
rect 3435 9680 3477 9689
rect 3435 9640 3436 9680
rect 3476 9640 3477 9680
rect 3435 9631 3477 9640
rect 5451 9680 5493 9689
rect 5451 9640 5452 9680
rect 5492 9640 5493 9680
rect 5451 9631 5493 9640
rect 8170 9680 8228 9681
rect 8170 9640 8179 9680
rect 8219 9640 8228 9680
rect 8170 9639 8228 9640
rect 1179 9596 1221 9605
rect 1179 9556 1180 9596
rect 1220 9556 1221 9596
rect 1179 9547 1221 9556
rect 1563 9596 1605 9605
rect 1563 9556 1564 9596
rect 1604 9556 1605 9596
rect 1563 9547 1605 9556
rect 3579 9596 3621 9605
rect 3579 9556 3580 9596
rect 3620 9556 3621 9596
rect 3579 9547 3621 9556
rect 8331 9596 8373 9605
rect 8331 9556 8332 9596
rect 8372 9556 8373 9596
rect 8331 9547 8373 9556
rect 1419 9512 1461 9521
rect 1419 9472 1420 9512
rect 1460 9472 1461 9512
rect 1419 9463 1461 9472
rect 1803 9512 1845 9521
rect 1803 9472 1804 9512
rect 1844 9472 1845 9512
rect 1803 9463 1845 9472
rect 3819 9512 3861 9521
rect 3819 9472 3820 9512
rect 3860 9472 3861 9512
rect 3819 9463 3861 9472
rect 6123 9512 6165 9521
rect 6123 9472 6124 9512
rect 6164 9472 6165 9512
rect 6123 9463 6165 9472
rect 6891 9512 6933 9521
rect 6891 9472 6892 9512
rect 6932 9472 6933 9512
rect 6891 9463 6933 9472
rect 10090 9512 10148 9513
rect 10090 9472 10099 9512
rect 10139 9472 10148 9512
rect 10090 9471 10148 9472
rect 1995 9428 2037 9437
rect 1995 9388 1996 9428
rect 2036 9388 2037 9428
rect 1995 9379 2037 9388
rect 3235 9428 3293 9429
rect 3235 9388 3244 9428
rect 3284 9388 3293 9428
rect 3235 9387 3293 9388
rect 4011 9428 4053 9437
rect 4011 9388 4012 9428
rect 4052 9388 4053 9428
rect 4011 9379 4053 9388
rect 5251 9428 5309 9429
rect 5251 9388 5260 9428
rect 5300 9388 5309 9428
rect 5251 9387 5309 9388
rect 6394 9428 6452 9429
rect 6394 9388 6403 9428
rect 6443 9388 6452 9428
rect 6394 9387 6452 9388
rect 6507 9428 6549 9437
rect 6507 9388 6508 9428
rect 6548 9388 6549 9428
rect 6507 9379 6549 9388
rect 6987 9428 7029 9437
rect 6987 9388 6988 9428
rect 7028 9388 7029 9428
rect 6987 9379 7029 9388
rect 7459 9428 7517 9429
rect 7459 9388 7468 9428
rect 7508 9388 7517 9428
rect 7459 9387 7517 9388
rect 7978 9428 8036 9429
rect 7978 9388 7987 9428
rect 8027 9388 8036 9428
rect 7978 9387 8036 9388
rect 8515 9428 8573 9429
rect 8515 9388 8524 9428
rect 8564 9388 8573 9428
rect 8515 9387 8573 9388
rect 9771 9428 9813 9437
rect 9771 9388 9772 9428
rect 9812 9388 9813 9428
rect 9771 9379 9813 9388
rect 10285 9428 10343 9429
rect 10285 9388 10294 9428
rect 10334 9388 10343 9428
rect 10285 9387 10343 9388
rect 5883 9260 5925 9269
rect 5883 9220 5884 9260
rect 5924 9220 5925 9260
rect 5883 9211 5925 9220
rect 1152 9092 10656 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 10656 9092
rect 1152 9028 10656 9052
rect 1467 8924 1509 8933
rect 1467 8884 1468 8924
rect 1508 8884 1509 8924
rect 1467 8875 1509 8884
rect 3723 8924 3765 8933
rect 3723 8884 3724 8924
rect 3764 8884 3765 8924
rect 3723 8875 3765 8884
rect 6651 8924 6693 8933
rect 6651 8884 6652 8924
rect 6692 8884 6693 8924
rect 6651 8875 6693 8884
rect 8427 8924 8469 8933
rect 8427 8884 8428 8924
rect 8468 8884 8469 8924
rect 8427 8875 8469 8884
rect 5451 8840 5493 8849
rect 5451 8800 5452 8840
rect 5492 8800 5493 8840
rect 5451 8791 5493 8800
rect 6315 8840 6357 8849
rect 6315 8800 6316 8840
rect 6356 8800 6357 8840
rect 6315 8791 6357 8800
rect 2283 8756 2325 8765
rect 4011 8756 4053 8765
rect 5931 8756 5973 8765
rect 1314 8747 1360 8756
rect 1314 8707 1315 8747
rect 1355 8707 1360 8747
rect 1314 8698 1360 8707
rect 1794 8747 1840 8756
rect 1794 8707 1795 8747
rect 1835 8707 1840 8747
rect 2283 8716 2284 8756
rect 2324 8716 2325 8756
rect 2283 8707 2325 8716
rect 3531 8747 3573 8756
rect 3531 8707 3532 8747
rect 3572 8707 3573 8747
rect 4011 8716 4012 8756
rect 4052 8716 4053 8756
rect 4011 8707 4053 8716
rect 5259 8747 5301 8756
rect 5259 8707 5260 8747
rect 5300 8707 5301 8747
rect 5931 8716 5932 8756
rect 5972 8716 5973 8756
rect 5931 8707 5973 8716
rect 6202 8756 6260 8757
rect 6202 8716 6211 8756
rect 6251 8716 6260 8756
rect 6202 8715 6260 8716
rect 6987 8756 7029 8765
rect 9099 8756 9141 8765
rect 6987 8716 6988 8756
rect 7028 8716 7029 8756
rect 6987 8707 7029 8716
rect 8235 8747 8277 8756
rect 8235 8707 8236 8747
rect 8276 8707 8277 8747
rect 9099 8716 9100 8756
rect 9140 8716 9141 8756
rect 9099 8707 9141 8716
rect 10347 8747 10389 8756
rect 10347 8707 10348 8747
rect 10388 8707 10389 8747
rect 1794 8698 1840 8707
rect 3531 8698 3573 8707
rect 5259 8698 5301 8707
rect 8235 8698 8277 8707
rect 10347 8698 10389 8707
rect 1947 8672 1989 8681
rect 1947 8632 1948 8672
rect 1988 8632 1989 8672
rect 1947 8623 1989 8632
rect 8715 8672 8757 8681
rect 8715 8632 8716 8672
rect 8756 8632 8757 8672
rect 8715 8623 8757 8632
rect 8955 8672 8997 8681
rect 8955 8632 8956 8672
rect 8996 8632 8997 8672
rect 8955 8623 8997 8632
rect 10539 8504 10581 8513
rect 10539 8464 10540 8504
rect 10580 8464 10581 8504
rect 10539 8455 10581 8464
rect 1152 8336 10656 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 10656 8336
rect 1152 8272 10656 8296
rect 2955 8168 2997 8177
rect 2955 8128 2956 8168
rect 2996 8128 2997 8168
rect 2955 8119 2997 8128
rect 6171 8168 6213 8177
rect 6171 8128 6172 8168
rect 6212 8128 6213 8168
rect 6171 8119 6213 8128
rect 9003 8168 9045 8177
rect 9003 8128 9004 8168
rect 9044 8128 9045 8168
rect 9003 8119 9045 8128
rect 5643 8084 5685 8093
rect 5643 8044 5644 8084
rect 5684 8044 5685 8084
rect 5643 8035 5685 8044
rect 8427 8084 8469 8093
rect 8427 8044 8428 8084
rect 8468 8044 8469 8084
rect 8427 8035 8469 8044
rect 1227 8000 1269 8009
rect 1227 7960 1228 8000
rect 1268 7960 1269 8000
rect 1227 7951 1269 7960
rect 6027 8000 6069 8009
rect 6027 7960 6028 8000
rect 6068 7960 6069 8000
rect 6027 7951 6069 7960
rect 6411 8000 6453 8009
rect 6411 7960 6412 8000
rect 6452 7960 6453 8000
rect 6411 7951 6453 7960
rect 6555 8000 6597 8009
rect 6555 7960 6556 8000
rect 6596 7960 6597 8000
rect 6555 7951 6597 7960
rect 6795 8000 6837 8009
rect 6795 7960 6796 8000
rect 6836 7960 6837 8000
rect 6795 7951 6837 7960
rect 1515 7916 1557 7925
rect 1515 7876 1516 7916
rect 1556 7876 1557 7916
rect 1515 7867 1557 7876
rect 2755 7916 2813 7917
rect 2755 7876 2764 7916
rect 2804 7876 2813 7916
rect 2755 7875 2813 7876
rect 3147 7916 3189 7925
rect 3147 7876 3148 7916
rect 3188 7876 3189 7916
rect 3147 7867 3189 7876
rect 4387 7916 4445 7917
rect 4387 7876 4396 7916
rect 4436 7876 4445 7916
rect 4387 7875 4445 7876
rect 4971 7916 5013 7925
rect 4971 7876 4972 7916
rect 5012 7876 5013 7916
rect 4971 7867 5013 7876
rect 5242 7916 5300 7917
rect 5242 7876 5251 7916
rect 5291 7876 5300 7916
rect 5242 7875 5300 7876
rect 7755 7916 7797 7925
rect 7755 7876 7756 7916
rect 7796 7876 7797 7916
rect 7755 7867 7797 7876
rect 8026 7916 8084 7917
rect 8026 7876 8035 7916
rect 8075 7876 8084 7916
rect 8026 7875 8084 7876
rect 9187 7916 9245 7917
rect 9187 7876 9196 7916
rect 9236 7876 9245 7916
rect 9187 7875 9245 7876
rect 10443 7916 10485 7925
rect 10443 7876 10444 7916
rect 10484 7876 10485 7916
rect 10443 7867 10485 7876
rect 4587 7832 4629 7841
rect 4587 7792 4588 7832
rect 4628 7792 4629 7832
rect 4587 7783 4629 7792
rect 5355 7832 5397 7841
rect 5355 7792 5356 7832
rect 5396 7792 5397 7832
rect 5355 7783 5397 7792
rect 8139 7832 8181 7841
rect 8139 7792 8140 7832
rect 8180 7792 8181 7832
rect 8139 7783 8181 7792
rect 5787 7748 5829 7757
rect 5787 7708 5788 7748
rect 5828 7708 5829 7748
rect 5787 7699 5829 7708
rect 1152 7580 10656 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 10656 7580
rect 1152 7516 10656 7540
rect 3003 7412 3045 7421
rect 3003 7372 3004 7412
rect 3044 7372 3045 7412
rect 3003 7363 3045 7372
rect 7563 7412 7605 7421
rect 7563 7372 7564 7412
rect 7604 7372 7605 7412
rect 7563 7363 7605 7372
rect 1227 7244 1269 7253
rect 4299 7244 4341 7253
rect 6123 7244 6165 7253
rect 8523 7244 8565 7253
rect 1227 7204 1228 7244
rect 1268 7204 1269 7244
rect 1227 7195 1269 7204
rect 2475 7235 2517 7244
rect 2475 7195 2476 7235
rect 2516 7195 2517 7235
rect 2475 7186 2517 7195
rect 2850 7235 2896 7244
rect 2850 7195 2851 7235
rect 2891 7195 2896 7235
rect 4299 7204 4300 7244
rect 4340 7204 4341 7244
rect 4299 7195 4341 7204
rect 5547 7235 5589 7244
rect 5547 7195 5548 7235
rect 5588 7195 5589 7235
rect 6123 7204 6124 7244
rect 6164 7204 6165 7244
rect 6123 7195 6165 7204
rect 7371 7235 7413 7244
rect 7371 7195 7372 7235
rect 7412 7195 7413 7235
rect 8523 7204 8524 7244
rect 8564 7204 8565 7244
rect 8523 7195 8565 7204
rect 9771 7235 9813 7244
rect 9771 7195 9772 7235
rect 9812 7195 9813 7235
rect 2850 7186 2896 7195
rect 5547 7186 5589 7195
rect 7371 7186 7413 7195
rect 9771 7186 9813 7195
rect 3531 7160 3573 7169
rect 3531 7120 3532 7160
rect 3572 7120 3573 7160
rect 3531 7111 3573 7120
rect 3915 7160 3957 7169
rect 3915 7120 3916 7160
rect 3956 7120 3957 7160
rect 3915 7111 3957 7120
rect 8331 7160 8373 7169
rect 8331 7120 8332 7160
rect 8372 7120 8373 7160
rect 8331 7111 8373 7120
rect 10347 7160 10389 7169
rect 10347 7120 10348 7160
rect 10388 7120 10389 7160
rect 10347 7111 10389 7120
rect 2667 7076 2709 7085
rect 2667 7036 2668 7076
rect 2708 7036 2709 7076
rect 2667 7027 2709 7036
rect 3291 7076 3333 7085
rect 3291 7036 3292 7076
rect 3332 7036 3333 7076
rect 3291 7027 3333 7036
rect 9963 7076 10005 7085
rect 9963 7036 9964 7076
rect 10004 7036 10005 7076
rect 9963 7027 10005 7036
rect 10587 7076 10629 7085
rect 10587 7036 10588 7076
rect 10628 7036 10629 7076
rect 10587 7027 10629 7036
rect 3675 6992 3717 7001
rect 3675 6952 3676 6992
rect 3716 6952 3717 6992
rect 3675 6943 3717 6952
rect 5739 6992 5781 7001
rect 5739 6952 5740 6992
rect 5780 6952 5781 6992
rect 5739 6943 5781 6952
rect 8091 6992 8133 7001
rect 8091 6952 8092 6992
rect 8132 6952 8133 6992
rect 8091 6943 8133 6952
rect 1152 6824 10656 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 10656 6824
rect 1152 6760 10656 6784
rect 1371 6656 1413 6665
rect 1371 6616 1372 6656
rect 1412 6616 1413 6656
rect 1371 6607 1413 6616
rect 10587 6656 10629 6665
rect 10587 6616 10588 6656
rect 10628 6616 10629 6656
rect 10587 6607 10629 6616
rect 7755 6572 7797 6581
rect 7755 6532 7756 6572
rect 7796 6532 7797 6572
rect 7755 6523 7797 6532
rect 1611 6488 1653 6497
rect 1611 6448 1612 6488
rect 1652 6448 1653 6488
rect 1611 6439 1653 6448
rect 4587 6488 4629 6497
rect 4587 6448 4588 6488
rect 4628 6448 4629 6488
rect 4587 6439 4629 6448
rect 9963 6488 10005 6497
rect 9963 6448 9964 6488
rect 10004 6448 10005 6488
rect 9963 6439 10005 6448
rect 10347 6488 10389 6497
rect 10347 6448 10348 6488
rect 10388 6448 10389 6488
rect 10347 6439 10389 6448
rect 1803 6404 1845 6413
rect 1803 6364 1804 6404
rect 1844 6364 1845 6404
rect 1803 6355 1845 6364
rect 3043 6404 3101 6405
rect 3043 6364 3052 6404
rect 3092 6364 3101 6404
rect 3043 6363 3101 6364
rect 4090 6404 4148 6405
rect 4090 6364 4099 6404
rect 4139 6364 4148 6404
rect 4090 6363 4148 6364
rect 4203 6404 4245 6413
rect 4203 6364 4204 6404
rect 4244 6364 4245 6404
rect 4203 6355 4245 6364
rect 4683 6404 4725 6413
rect 4683 6364 4684 6404
rect 4724 6364 4725 6404
rect 4683 6355 4725 6364
rect 5155 6404 5213 6405
rect 5155 6364 5164 6404
rect 5204 6364 5213 6404
rect 5155 6363 5213 6364
rect 5674 6404 5732 6405
rect 5674 6364 5683 6404
rect 5723 6364 5732 6404
rect 5674 6363 5732 6364
rect 6315 6404 6357 6413
rect 6315 6364 6316 6404
rect 6356 6364 6357 6404
rect 6315 6355 6357 6364
rect 7555 6404 7613 6405
rect 7555 6364 7564 6404
rect 7604 6364 7613 6404
rect 7555 6363 7613 6364
rect 3243 6320 3285 6329
rect 3243 6280 3244 6320
rect 3284 6280 3285 6320
rect 3243 6271 3285 6280
rect 10203 6320 10245 6329
rect 10203 6280 10204 6320
rect 10244 6280 10245 6320
rect 10203 6271 10245 6280
rect 3514 6236 3572 6237
rect 3514 6196 3523 6236
rect 3563 6196 3572 6236
rect 3514 6195 3572 6196
rect 3802 6236 3860 6237
rect 3802 6196 3811 6236
rect 3851 6196 3860 6236
rect 3802 6195 3860 6196
rect 5835 6236 5877 6245
rect 5835 6196 5836 6236
rect 5876 6196 5877 6236
rect 5835 6187 5877 6196
rect 6106 6236 6164 6237
rect 6106 6196 6115 6236
rect 6155 6196 6164 6236
rect 6106 6195 6164 6196
rect 1152 6068 10656 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 10656 6068
rect 1152 6004 10656 6028
rect 6202 5900 6260 5901
rect 6202 5860 6211 5900
rect 6251 5860 6260 5900
rect 6202 5859 6260 5860
rect 8427 5900 8469 5909
rect 8427 5860 8428 5900
rect 8468 5860 8469 5900
rect 8427 5851 8469 5860
rect 2859 5816 2901 5825
rect 2859 5776 2860 5816
rect 2900 5776 2901 5816
rect 2859 5767 2901 5776
rect 1419 5732 1461 5741
rect 3130 5732 3188 5733
rect 1419 5692 1420 5732
rect 1460 5692 1461 5732
rect 1419 5683 1461 5692
rect 2667 5723 2709 5732
rect 2667 5683 2668 5723
rect 2708 5683 2709 5723
rect 3130 5692 3139 5732
rect 3179 5692 3188 5732
rect 3130 5691 3188 5692
rect 3243 5732 3285 5741
rect 3243 5692 3244 5732
rect 3284 5692 3285 5732
rect 3243 5683 3285 5692
rect 3627 5732 3669 5741
rect 6682 5732 6740 5733
rect 3627 5692 3628 5732
rect 3668 5692 3669 5732
rect 3627 5683 3669 5692
rect 4203 5723 4245 5732
rect 4203 5683 4204 5723
rect 4244 5683 4245 5723
rect 2667 5674 2709 5683
rect 4203 5674 4245 5683
rect 4683 5723 4725 5732
rect 4683 5683 4684 5723
rect 4724 5683 4725 5723
rect 6682 5692 6691 5732
rect 6731 5692 6740 5732
rect 6682 5691 6740 5692
rect 6795 5732 6837 5741
rect 6795 5692 6796 5732
rect 6836 5692 6837 5732
rect 6795 5683 6837 5692
rect 7179 5732 7221 5741
rect 8763 5732 8805 5741
rect 7179 5692 7180 5732
rect 7220 5692 7221 5732
rect 7179 5683 7221 5692
rect 7755 5723 7797 5732
rect 7755 5683 7756 5723
rect 7796 5683 7797 5723
rect 4683 5674 4725 5683
rect 7755 5674 7797 5683
rect 8235 5723 8277 5732
rect 8235 5683 8236 5723
rect 8276 5683 8277 5723
rect 8235 5674 8277 5683
rect 8610 5723 8656 5732
rect 8610 5683 8611 5723
rect 8651 5683 8656 5723
rect 8763 5692 8764 5732
rect 8804 5692 8805 5732
rect 8763 5683 8805 5692
rect 8610 5674 8656 5683
rect 3723 5648 3765 5657
rect 3723 5608 3724 5648
rect 3764 5608 3765 5648
rect 3723 5599 3765 5608
rect 4906 5648 4964 5649
rect 4906 5608 4915 5648
rect 4955 5608 4964 5648
rect 4906 5607 4964 5608
rect 5259 5648 5301 5657
rect 5259 5608 5260 5648
rect 5300 5608 5301 5648
rect 5259 5599 5301 5608
rect 5643 5648 5685 5657
rect 5643 5608 5644 5648
rect 5684 5608 5685 5648
rect 5643 5599 5685 5608
rect 5835 5648 5877 5657
rect 5835 5608 5836 5648
rect 5876 5608 5877 5648
rect 5835 5599 5877 5608
rect 7275 5648 7317 5657
rect 7275 5608 7276 5648
rect 7316 5608 7317 5648
rect 7275 5599 7317 5608
rect 9291 5648 9333 5657
rect 9291 5608 9292 5648
rect 9332 5608 9333 5648
rect 9291 5599 9333 5608
rect 10347 5648 10389 5657
rect 10347 5608 10348 5648
rect 10388 5608 10389 5648
rect 10347 5599 10389 5608
rect 6075 5564 6117 5573
rect 6075 5524 6076 5564
rect 6116 5524 6117 5564
rect 6075 5515 6117 5524
rect 9051 5564 9093 5573
rect 9051 5524 9052 5564
rect 9092 5524 9093 5564
rect 9051 5515 9093 5524
rect 5019 5480 5061 5489
rect 5019 5440 5020 5480
rect 5060 5440 5061 5480
rect 5019 5431 5061 5440
rect 5403 5480 5445 5489
rect 5403 5440 5404 5480
rect 5444 5440 5445 5480
rect 5403 5431 5445 5440
rect 10587 5480 10629 5489
rect 10587 5440 10588 5480
rect 10628 5440 10629 5480
rect 10587 5431 10629 5440
rect 1152 5312 10656 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 10656 5312
rect 1152 5248 10656 5272
rect 4011 5144 4053 5153
rect 4011 5104 4012 5144
rect 4052 5104 4053 5144
rect 4011 5095 4053 5104
rect 8427 5144 8469 5153
rect 8427 5104 8428 5144
rect 8468 5104 8469 5144
rect 8427 5095 8469 5104
rect 4875 4976 4917 4985
rect 4875 4936 4876 4976
rect 4916 4936 4917 4976
rect 4875 4927 4917 4936
rect 6154 4976 6212 4977
rect 6154 4936 6163 4976
rect 6203 4936 6212 4976
rect 6154 4935 6212 4936
rect 6507 4976 6549 4985
rect 6507 4936 6508 4976
rect 6548 4936 6549 4976
rect 6507 4927 6549 4936
rect 1711 4892 1769 4893
rect 1711 4852 1720 4892
rect 1760 4852 1769 4892
rect 1711 4851 1769 4852
rect 1879 4892 1937 4893
rect 1879 4852 1888 4892
rect 1928 4852 1937 4892
rect 1879 4851 1937 4852
rect 2571 4892 2613 4901
rect 2571 4852 2572 4892
rect 2612 4852 2613 4892
rect 2571 4843 2613 4852
rect 3811 4892 3869 4893
rect 3811 4852 3820 4892
rect 3860 4852 3869 4892
rect 3811 4851 3869 4852
rect 4365 4892 4407 4901
rect 4365 4852 4366 4892
rect 4406 4852 4407 4892
rect 4365 4843 4407 4852
rect 4480 4892 4538 4893
rect 4480 4852 4489 4892
rect 4529 4852 4538 4892
rect 4480 4851 4538 4852
rect 4971 4892 5013 4901
rect 4971 4852 4972 4892
rect 5012 4852 5013 4892
rect 4971 4843 5013 4852
rect 5443 4892 5501 4893
rect 5443 4852 5452 4892
rect 5492 4852 5501 4892
rect 5443 4851 5501 4852
rect 5931 4892 5989 4893
rect 5931 4852 5940 4892
rect 5980 4852 5989 4892
rect 5931 4851 5989 4852
rect 6987 4892 7029 4901
rect 6987 4852 6988 4892
rect 7028 4852 7029 4892
rect 6987 4843 7029 4852
rect 8227 4892 8285 4893
rect 8227 4852 8236 4892
rect 8276 4852 8285 4892
rect 8227 4851 8285 4852
rect 1546 4808 1604 4809
rect 1546 4768 1555 4808
rect 1595 4768 1604 4808
rect 1546 4767 1604 4768
rect 2043 4724 2085 4733
rect 2043 4684 2044 4724
rect 2084 4684 2085 4724
rect 2043 4675 2085 4684
rect 6267 4724 6309 4733
rect 6267 4684 6268 4724
rect 6308 4684 6309 4724
rect 6267 4675 6309 4684
rect 6682 4724 6740 4725
rect 6682 4684 6691 4724
rect 6731 4684 6740 4724
rect 6682 4683 6740 4684
rect 1152 4556 10656 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 10656 4556
rect 1152 4492 10656 4516
rect 1210 4388 1268 4389
rect 1210 4348 1219 4388
rect 1259 4348 1268 4388
rect 1210 4347 1268 4348
rect 3627 4388 3669 4397
rect 3627 4348 3628 4388
rect 3668 4348 3669 4388
rect 3627 4339 3669 4348
rect 7179 4388 7221 4397
rect 7179 4348 7180 4388
rect 7220 4348 7221 4388
rect 7179 4339 7221 4348
rect 7354 4388 7412 4389
rect 7354 4348 7363 4388
rect 7403 4348 7412 4388
rect 7354 4347 7412 4348
rect 1851 4304 1893 4313
rect 1851 4264 1852 4304
rect 1892 4264 1893 4304
rect 1851 4255 1893 4264
rect 5451 4304 5493 4313
rect 5451 4264 5452 4304
rect 5492 4264 5493 4304
rect 5451 4255 5493 4264
rect 10042 4304 10100 4305
rect 10042 4264 10051 4304
rect 10091 4264 10100 4304
rect 10042 4263 10100 4264
rect 2187 4220 2229 4229
rect 4011 4220 4053 4229
rect 1698 4211 1744 4220
rect 1698 4171 1699 4211
rect 1739 4171 1744 4211
rect 2187 4180 2188 4220
rect 2228 4180 2229 4220
rect 2187 4171 2229 4180
rect 3435 4211 3477 4220
rect 3435 4171 3436 4211
rect 3476 4171 3477 4211
rect 4011 4180 4012 4220
rect 4052 4180 4053 4220
rect 4011 4171 4053 4180
rect 5259 4220 5317 4221
rect 5259 4180 5268 4220
rect 5308 4180 5317 4220
rect 5259 4179 5317 4180
rect 5739 4220 5781 4229
rect 10443 4220 10485 4229
rect 5739 4180 5740 4220
rect 5780 4180 5781 4220
rect 5739 4171 5781 4180
rect 6987 4211 7029 4220
rect 6987 4171 6988 4211
rect 7028 4171 7029 4211
rect 10443 4180 10444 4220
rect 10484 4180 10485 4220
rect 10443 4171 10485 4180
rect 1698 4162 1744 4171
rect 3435 4162 3477 4171
rect 6987 4162 7029 4171
rect 1152 3800 10656 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 10656 3800
rect 1152 3736 10656 3760
rect 3099 3632 3141 3641
rect 3099 3592 3100 3632
rect 3140 3592 3141 3632
rect 3099 3583 3141 3592
rect 3483 3632 3525 3641
rect 3483 3592 3484 3632
rect 3524 3592 3525 3632
rect 3483 3583 3525 3592
rect 1563 3548 1605 3557
rect 1563 3508 1564 3548
rect 1604 3508 1605 3548
rect 1563 3499 1605 3508
rect 1947 3548 1989 3557
rect 1947 3508 1948 3548
rect 1988 3508 1989 3548
rect 1947 3499 1989 3508
rect 1803 3464 1845 3473
rect 1803 3424 1804 3464
rect 1844 3424 1845 3464
rect 1803 3415 1845 3424
rect 2187 3464 2229 3473
rect 2187 3424 2188 3464
rect 2228 3424 2229 3464
rect 2187 3415 2229 3424
rect 2331 3464 2373 3473
rect 2331 3424 2332 3464
rect 2372 3424 2373 3464
rect 2331 3415 2373 3424
rect 2571 3464 2613 3473
rect 2571 3424 2572 3464
rect 2612 3424 2613 3464
rect 2571 3415 2613 3424
rect 2955 3464 2997 3473
rect 2955 3424 2956 3464
rect 2996 3424 2997 3464
rect 2955 3415 2997 3424
rect 3339 3464 3381 3473
rect 3339 3424 3340 3464
rect 3380 3424 3381 3464
rect 3339 3415 3381 3424
rect 3723 3464 3765 3473
rect 3723 3424 3724 3464
rect 3764 3424 3765 3464
rect 3723 3415 3765 3424
rect 3915 3464 3957 3473
rect 3915 3424 3916 3464
rect 3956 3424 3957 3464
rect 3915 3415 3957 3424
rect 4491 3464 4533 3473
rect 4491 3424 4492 3464
rect 4532 3424 4533 3464
rect 4491 3415 4533 3424
rect 4779 3464 4821 3473
rect 4779 3424 4780 3464
rect 4820 3424 4821 3464
rect 4779 3415 4821 3424
rect 5643 3464 5685 3473
rect 5643 3424 5644 3464
rect 5684 3424 5685 3464
rect 5643 3415 5685 3424
rect 5931 3464 5973 3473
rect 5931 3424 5932 3464
rect 5972 3424 5973 3464
rect 5931 3415 5973 3424
rect 6507 3464 6549 3473
rect 6507 3424 6508 3464
rect 6548 3424 6549 3464
rect 6507 3415 6549 3424
rect 6795 3464 6837 3473
rect 6795 3424 6796 3464
rect 6836 3424 6837 3464
rect 6795 3415 6837 3424
rect 7083 3464 7125 3473
rect 7083 3424 7084 3464
rect 7124 3424 7125 3464
rect 7083 3415 7125 3424
rect 10347 3464 10389 3473
rect 10347 3424 10348 3464
rect 10388 3424 10389 3464
rect 10347 3415 10389 3424
rect 2715 3296 2757 3305
rect 2715 3256 2716 3296
rect 2756 3256 2757 3296
rect 2715 3247 2757 3256
rect 1306 3212 1364 3213
rect 1306 3172 1315 3212
rect 1355 3172 1364 3212
rect 1306 3171 1364 3172
rect 3898 3212 3956 3213
rect 3898 3172 3907 3212
rect 3947 3172 3956 3212
rect 3898 3171 3956 3172
rect 4282 3212 4340 3213
rect 4282 3172 4291 3212
rect 4331 3172 4340 3212
rect 4282 3171 4340 3172
rect 5146 3212 5204 3213
rect 5146 3172 5155 3212
rect 5195 3172 5204 3212
rect 5146 3171 5204 3172
rect 5434 3212 5492 3213
rect 5434 3172 5443 3212
rect 5483 3172 5492 3212
rect 5434 3171 5492 3172
rect 6298 3212 6356 3213
rect 6298 3172 6307 3212
rect 6347 3172 6356 3212
rect 6298 3171 6356 3172
rect 6778 3212 6836 3213
rect 6778 3172 6787 3212
rect 6827 3172 6836 3212
rect 6778 3171 6836 3172
rect 10587 3212 10629 3221
rect 10587 3172 10588 3212
rect 10628 3172 10629 3212
rect 10587 3163 10629 3172
rect 1152 3044 10656 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 10656 3044
rect 1152 2980 10656 3004
rect 1179 2876 1221 2885
rect 1179 2836 1180 2876
rect 1220 2836 1221 2876
rect 1179 2827 1221 2836
rect 2715 2876 2757 2885
rect 2715 2836 2716 2876
rect 2756 2836 2757 2876
rect 2715 2827 2757 2836
rect 3610 2876 3668 2877
rect 3610 2836 3619 2876
rect 3659 2836 3668 2876
rect 3610 2835 3668 2836
rect 3898 2876 3956 2877
rect 3898 2836 3907 2876
rect 3947 2836 3956 2876
rect 3898 2835 3956 2836
rect 5050 2876 5108 2877
rect 5050 2836 5059 2876
rect 5099 2836 5108 2876
rect 5050 2835 5108 2836
rect 5818 2876 5876 2877
rect 5818 2836 5827 2876
rect 5867 2836 5876 2876
rect 5818 2835 5876 2836
rect 2331 2792 2373 2801
rect 2331 2752 2332 2792
rect 2372 2752 2373 2792
rect 2331 2743 2373 2752
rect 4395 2792 4437 2801
rect 4395 2752 4396 2792
rect 4436 2752 4437 2792
rect 4395 2743 4437 2752
rect 4683 2792 4725 2801
rect 4683 2752 4684 2792
rect 4724 2752 4725 2792
rect 4683 2743 4725 2752
rect 5259 2792 5301 2801
rect 5259 2752 5260 2792
rect 5300 2752 5301 2792
rect 5259 2743 5301 2752
rect 5547 2792 5589 2801
rect 5547 2752 5548 2792
rect 5588 2752 5589 2792
rect 5547 2743 5589 2752
rect 6123 2792 6165 2801
rect 6123 2752 6124 2792
rect 6164 2752 6165 2792
rect 6123 2743 6165 2752
rect 6411 2792 6453 2801
rect 6411 2752 6412 2792
rect 6452 2752 6453 2792
rect 6411 2743 6453 2752
rect 1611 2708 1653 2717
rect 1611 2668 1612 2708
rect 1652 2668 1653 2708
rect 1611 2659 1653 2668
rect 1419 2624 1461 2633
rect 1419 2584 1420 2624
rect 1460 2584 1461 2624
rect 1419 2575 1461 2584
rect 1947 2624 1989 2633
rect 1947 2584 1948 2624
rect 1988 2584 1989 2624
rect 1947 2575 1989 2584
rect 2187 2624 2229 2633
rect 2187 2584 2188 2624
rect 2228 2584 2229 2624
rect 2187 2575 2229 2584
rect 2571 2624 2613 2633
rect 2571 2584 2572 2624
rect 2612 2584 2613 2624
rect 2571 2575 2613 2584
rect 2955 2624 2997 2633
rect 2955 2584 2956 2624
rect 2996 2584 2997 2624
rect 2955 2575 2997 2584
rect 3339 2624 3381 2633
rect 3339 2584 3340 2624
rect 3380 2584 3381 2624
rect 3339 2575 3381 2584
rect 4395 2624 4437 2633
rect 4395 2584 4396 2624
rect 4436 2584 4437 2624
rect 4395 2575 4437 2584
rect 10347 2624 10389 2633
rect 10347 2584 10348 2624
rect 10388 2584 10389 2624
rect 10347 2575 10389 2584
rect 3099 2456 3141 2465
rect 3099 2416 3100 2456
rect 3140 2416 3141 2456
rect 3099 2407 3141 2416
rect 10587 2456 10629 2465
rect 10587 2416 10588 2456
rect 10628 2416 10629 2456
rect 10587 2407 10629 2416
rect 1152 2288 10656 2312
rect 1152 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 10656 2288
rect 1152 2224 10656 2248
rect 1179 2120 1221 2129
rect 1179 2080 1180 2120
rect 1220 2080 1221 2120
rect 1179 2071 1221 2080
rect 2331 2120 2373 2129
rect 2331 2080 2332 2120
rect 2372 2080 2373 2120
rect 2331 2071 2373 2080
rect 2715 2120 2757 2129
rect 2715 2080 2716 2120
rect 2756 2080 2757 2120
rect 2715 2071 2757 2080
rect 10042 2120 10100 2121
rect 10042 2080 10051 2120
rect 10091 2080 10100 2120
rect 10042 2079 10100 2080
rect 1563 2036 1605 2045
rect 1563 1996 1564 2036
rect 1604 1996 1605 2036
rect 1563 1987 1605 1996
rect 1419 1952 1461 1961
rect 1419 1912 1420 1952
rect 1460 1912 1461 1952
rect 1419 1903 1461 1912
rect 1803 1952 1845 1961
rect 1803 1912 1804 1952
rect 1844 1912 1845 1952
rect 1803 1903 1845 1912
rect 2187 1952 2229 1961
rect 2187 1912 2188 1952
rect 2228 1912 2229 1952
rect 2187 1903 2229 1912
rect 2571 1952 2613 1961
rect 2571 1912 2572 1952
rect 2612 1912 2613 1952
rect 2571 1903 2613 1912
rect 2955 1952 2997 1961
rect 2955 1912 2956 1952
rect 2996 1912 2997 1952
rect 2955 1903 2997 1912
rect 3339 1952 3381 1961
rect 3339 1912 3340 1952
rect 3380 1912 3381 1952
rect 3339 1903 3381 1912
rect 3723 1952 3765 1961
rect 3723 1912 3724 1952
rect 3764 1912 3765 1952
rect 3723 1903 3765 1912
rect 4299 1952 4341 1961
rect 4299 1912 4300 1952
rect 4340 1912 4341 1952
rect 4299 1903 4341 1912
rect 4587 1952 4629 1961
rect 4587 1912 4588 1952
rect 4628 1912 4629 1952
rect 4587 1903 4629 1912
rect 5451 1952 5493 1961
rect 5451 1912 5452 1952
rect 5492 1912 5493 1952
rect 5451 1903 5493 1912
rect 5163 1868 5205 1877
rect 5163 1828 5164 1868
rect 5204 1828 5205 1868
rect 5163 1819 5205 1828
rect 10443 1868 10485 1877
rect 10443 1828 10444 1868
rect 10484 1828 10485 1868
rect 10443 1819 10485 1828
rect 1947 1784 1989 1793
rect 1947 1744 1948 1784
rect 1988 1744 1989 1784
rect 1947 1735 1989 1744
rect 3099 1784 3141 1793
rect 3099 1744 3100 1784
rect 3140 1744 3141 1784
rect 3099 1735 3141 1744
rect 4011 1784 4053 1793
rect 4011 1744 4012 1784
rect 4052 1744 4053 1784
rect 4011 1735 4053 1744
rect 5739 1784 5781 1793
rect 5739 1744 5740 1784
rect 5780 1744 5781 1784
rect 5739 1735 5781 1744
rect 6027 1784 6069 1793
rect 6027 1744 6028 1784
rect 6068 1744 6069 1784
rect 6027 1735 6069 1744
rect 3483 1700 3525 1709
rect 3483 1660 3484 1700
rect 3524 1660 3525 1700
rect 3483 1651 3525 1660
rect 4858 1700 4916 1701
rect 4858 1660 4867 1700
rect 4907 1660 4916 1700
rect 4858 1659 4916 1660
rect 1152 1532 10656 1556
rect 1152 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 10656 1532
rect 1152 1468 10656 1492
<< via1 >>
rect 4928 45340 4968 45380
rect 5010 45340 5050 45380
rect 5092 45340 5132 45380
rect 5174 45340 5214 45380
rect 5256 45340 5296 45380
rect 3484 45172 3524 45212
rect 3964 45172 4004 45212
rect 4348 45172 4388 45212
rect 4732 45172 4772 45212
rect 5116 45172 5156 45212
rect 5884 45172 5924 45212
rect 6268 45172 6308 45212
rect 6652 45172 6692 45212
rect 7036 45172 7076 45212
rect 7420 45172 7460 45212
rect 7804 45172 7844 45212
rect 8188 45172 8228 45212
rect 8572 45172 8612 45212
rect 8956 45172 8996 45212
rect 9340 45172 9380 45212
rect 9724 45172 9764 45212
rect 2332 45088 2372 45128
rect 3388 45088 3428 45128
rect 5500 45088 5540 45128
rect 1315 45004 1355 45044
rect 2131 45004 2171 45044
rect 2659 44995 2699 45035
rect 2812 45004 2852 45044
rect 3148 44920 3188 44960
rect 3724 44920 3764 44960
rect 4204 44920 4244 44960
rect 4588 44920 4628 44960
rect 4972 44920 5012 44960
rect 5356 44920 5396 44960
rect 5740 44920 5780 44960
rect 6124 44920 6164 44960
rect 6508 44920 6548 44960
rect 6892 44920 6932 44960
rect 7276 44920 7316 44960
rect 7660 44920 7700 44960
rect 8044 44920 8084 44960
rect 8428 44920 8468 44960
rect 8812 44920 8852 44960
rect 9196 44920 9236 44960
rect 9580 44920 9620 44960
rect 9964 44920 10004 44960
rect 10348 44920 10388 44960
rect 1516 44752 1556 44792
rect 10588 44752 10628 44792
rect 3688 44584 3728 44624
rect 3770 44584 3810 44624
rect 3852 44584 3892 44624
rect 3934 44584 3974 44624
rect 4016 44584 4056 44624
rect 3868 44416 3908 44456
rect 5212 44416 5252 44456
rect 5596 44416 5636 44456
rect 6172 44416 6212 44456
rect 6556 44416 6596 44456
rect 7036 44416 7076 44456
rect 7420 44416 7460 44456
rect 7804 44416 7844 44456
rect 9244 44416 9284 44456
rect 10204 44416 10244 44456
rect 10588 44416 10628 44456
rect 5116 44332 5156 44372
rect 9628 44332 9668 44372
rect 2476 44248 2516 44288
rect 3628 44248 3668 44288
rect 4012 44248 4052 44288
rect 4396 44248 4436 44288
rect 4828 44248 4868 44288
rect 5452 44248 5492 44288
rect 5836 44248 5876 44288
rect 6412 44248 6452 44288
rect 6796 44248 6836 44288
rect 7276 44248 7316 44288
rect 7660 44248 7700 44288
rect 8044 44248 8084 44288
rect 9004 44248 9044 44288
rect 9388 44248 9428 44288
rect 9964 44248 10004 44288
rect 10348 44248 10388 44288
rect 1315 44164 1355 44204
rect 1939 44164 1979 44204
rect 2716 44080 2756 44120
rect 8524 44080 8564 44120
rect 1516 43996 1556 44036
rect 2140 43996 2180 44036
rect 2947 43996 2987 44036
rect 3235 43996 3275 44036
rect 4252 43996 4292 44036
rect 4636 43996 4676 44036
rect 8227 43996 8267 44036
rect 4928 43828 4968 43868
rect 5010 43828 5050 43868
rect 5092 43828 5132 43868
rect 5174 43828 5214 43868
rect 5256 43828 5296 43868
rect 2467 43660 2507 43700
rect 3484 43660 3524 43700
rect 4108 43660 4148 43700
rect 6403 43660 6443 43700
rect 6691 43660 6731 43700
rect 8035 43660 8075 43700
rect 8515 43660 8555 43700
rect 8995 43660 9035 43700
rect 9379 43660 9419 43700
rect 4876 43576 4916 43616
rect 5740 43576 5780 43616
rect 7084 43576 7124 43616
rect 7372 43576 7412 43616
rect 7660 43576 7700 43616
rect 9676 43576 9716 43616
rect 1219 43483 1259 43523
rect 1795 43492 1835 43532
rect 1372 43408 1412 43448
rect 2860 43408 2900 43448
rect 3244 43408 3284 43448
rect 3580 43408 3620 43448
rect 3868 43408 3908 43448
rect 4396 43408 4436 43448
rect 5116 43408 5156 43448
rect 5356 43408 5396 43448
rect 6028 43408 6068 43448
rect 6316 43408 6356 43448
rect 8236 43408 8276 43448
rect 8524 43408 8564 43448
rect 9964 43408 10004 43448
rect 10348 43408 10388 43448
rect 3100 43324 3140 43364
rect 4636 43324 4676 43364
rect 10204 43324 10244 43364
rect 1996 43240 2036 43280
rect 10588 43240 10628 43280
rect 3688 43072 3728 43112
rect 3770 43072 3810 43112
rect 3852 43072 3892 43112
rect 3934 43072 3974 43112
rect 4016 43072 4056 43112
rect 1708 42904 1748 42944
rect 3484 42904 3524 42944
rect 5500 42904 5540 42944
rect 2764 42736 2804 42776
rect 3724 42736 3764 42776
rect 4828 42736 4868 42776
rect 5068 42736 5108 42776
rect 5260 42736 5300 42776
rect 8428 42736 8468 42776
rect 9964 42736 10004 42776
rect 10348 42736 10388 42776
rect 1315 42652 1355 42692
rect 2083 42652 2123 42692
rect 3874 42652 3914 42692
rect 4354 42652 4394 42692
rect 6796 42652 6836 42692
rect 8716 42652 8756 42692
rect 9388 42652 9428 42692
rect 6508 42568 6548 42608
rect 7084 42568 7124 42608
rect 7948 42568 7988 42608
rect 9676 42568 9716 42608
rect 10204 42568 10244 42608
rect 2284 42484 2324 42524
rect 3004 42484 3044 42524
rect 3331 42484 3371 42524
rect 4060 42484 4100 42524
rect 4540 42484 4580 42524
rect 5731 42484 5771 42524
rect 5923 42484 5963 42524
rect 6307 42484 6347 42524
rect 7363 42484 7403 42524
rect 7651 42484 7691 42524
rect 8995 42484 9035 42524
rect 9475 42484 9515 42524
rect 10588 42484 10628 42524
rect 4928 42316 4968 42356
rect 5010 42316 5050 42356
rect 5092 42316 5132 42356
rect 5174 42316 5214 42356
rect 5256 42316 5296 42356
rect 2284 42148 2324 42188
rect 4732 42148 4772 42188
rect 7996 42148 8036 42188
rect 8419 42148 8459 42188
rect 9628 42148 9668 42188
rect 1708 42064 1748 42104
rect 3676 42064 3716 42104
rect 4876 42064 4916 42104
rect 5932 42064 5972 42104
rect 8716 42064 8756 42104
rect 9004 42064 9044 42104
rect 1315 41980 1355 42020
rect 2083 41980 2123 42020
rect 2851 41980 2891 42020
rect 3523 41971 3563 42011
rect 4003 41971 4043 42011
rect 5155 41971 5195 42011
rect 5644 41980 5684 42020
rect 6412 41980 6452 42020
rect 7660 41971 7700 42011
rect 10060 41980 10100 42020
rect 4156 41896 4196 41936
rect 4492 41896 4532 41936
rect 5308 41896 5348 41936
rect 8236 41896 8276 41936
rect 9292 41896 9332 41936
rect 9868 41896 9908 41936
rect 10348 41896 10388 41936
rect 10588 41896 10628 41936
rect 3052 41812 3092 41852
rect 7852 41812 7892 41852
rect 9532 41812 9572 41852
rect 3688 41560 3728 41600
rect 3770 41560 3810 41600
rect 3852 41560 3892 41600
rect 3934 41560 3974 41600
rect 4016 41560 4056 41600
rect 1228 41224 1268 41264
rect 3340 41224 3380 41264
rect 6124 41224 6164 41264
rect 9964 41224 10004 41264
rect 10348 41224 10388 41264
rect 1612 41140 1652 41180
rect 2860 41140 2900 41180
rect 3820 41140 3860 41180
rect 5072 41140 5112 41180
rect 5602 41140 5642 41180
rect 6412 41140 6452 41180
rect 7660 41140 7700 41180
rect 8044 41140 8084 41180
rect 9292 41140 9332 41180
rect 10204 41056 10244 41096
rect 1468 40972 1508 41012
rect 3052 40972 3092 41012
rect 3331 40972 3371 41012
rect 3619 40972 3659 41012
rect 5260 40972 5300 41012
rect 5788 40972 5828 41012
rect 6211 40972 6251 41012
rect 7852 40972 7892 41012
rect 9484 40972 9524 41012
rect 9763 40972 9803 41012
rect 10588 40972 10628 41012
rect 4928 40804 4968 40844
rect 5010 40804 5050 40844
rect 5092 40804 5132 40844
rect 5174 40804 5214 40844
rect 5256 40804 5296 40844
rect 5548 40636 5588 40676
rect 5980 40636 6020 40676
rect 9580 40636 9620 40676
rect 3532 40552 3572 40592
rect 7564 40552 7604 40592
rect 1315 40468 1355 40508
rect 2092 40468 2132 40508
rect 3340 40459 3380 40499
rect 3811 40468 3851 40508
rect 3916 40468 3956 40508
rect 4300 40468 4340 40508
rect 4876 40459 4916 40499
rect 5356 40459 5396 40499
rect 6124 40468 6164 40508
rect 7372 40459 7412 40499
rect 7843 40468 7883 40508
rect 7948 40468 7988 40508
rect 8332 40468 8372 40508
rect 8908 40459 8948 40499
rect 9388 40459 9428 40499
rect 10243 40459 10283 40499
rect 4396 40384 4436 40424
rect 5740 40384 5780 40424
rect 8428 40384 8468 40424
rect 9964 40384 10004 40424
rect 10396 40384 10436 40424
rect 1516 40300 1556 40340
rect 3688 40048 3728 40088
rect 3770 40048 3810 40088
rect 3852 40048 3892 40088
rect 3934 40048 3974 40088
rect 4016 40048 4056 40088
rect 6268 39796 6308 39836
rect 3724 39712 3764 39752
rect 5164 39712 5204 39752
rect 5692 39712 5732 39752
rect 6028 39712 6068 39752
rect 6604 39712 6644 39752
rect 8428 39712 8468 39752
rect 9868 39712 9908 39752
rect 1420 39628 1460 39668
rect 2668 39628 2708 39668
rect 3235 39628 3275 39668
rect 3340 39628 3380 39668
rect 3820 39628 3860 39668
rect 4300 39628 4340 39668
rect 4788 39628 4828 39668
rect 5536 39628 5576 39668
rect 7918 39628 7958 39668
rect 8041 39628 8081 39668
rect 8524 39628 8564 39668
rect 9004 39628 9044 39668
rect 9492 39628 9532 39668
rect 10195 39628 10235 39668
rect 5404 39544 5444 39584
rect 2860 39460 2900 39500
rect 4972 39460 5012 39500
rect 6364 39460 6404 39500
rect 6883 39460 6923 39500
rect 7075 39460 7115 39500
rect 7363 39460 7403 39500
rect 9676 39460 9716 39500
rect 10108 39460 10148 39500
rect 10396 39460 10436 39500
rect 4928 39292 4968 39332
rect 5010 39292 5050 39332
rect 5092 39292 5132 39332
rect 5174 39292 5214 39332
rect 5256 39292 5296 39332
rect 3196 39124 3236 39164
rect 5452 39124 5492 39164
rect 9964 39124 10004 39164
rect 2860 39040 2900 39080
rect 1420 38956 1460 38996
rect 2668 38947 2708 38987
rect 3043 38947 3083 38987
rect 3523 38947 3563 38987
rect 4012 38956 4052 38996
rect 5260 38947 5300 38987
rect 5635 38947 5675 38987
rect 6124 38956 6164 38996
rect 7372 38947 7412 38987
rect 8223 38956 8263 38996
rect 8332 38956 8372 38996
rect 8716 38956 8756 38996
rect 9292 38947 9332 38987
rect 9772 38947 9812 38987
rect 10147 38947 10187 38987
rect 3676 38872 3716 38912
rect 5788 38872 5828 38912
rect 7756 38872 7796 38912
rect 8812 38872 8852 38912
rect 10300 38872 10340 38912
rect 7564 38704 7604 38744
rect 7996 38704 8036 38744
rect 3688 38536 3728 38576
rect 3770 38536 3810 38576
rect 3852 38536 3892 38576
rect 3934 38536 3974 38576
rect 4016 38536 4056 38576
rect 8428 38368 8468 38408
rect 10252 38368 10292 38408
rect 2236 38284 2276 38324
rect 1996 38200 2036 38240
rect 10444 38200 10484 38240
rect 1315 38116 1355 38156
rect 2380 38116 2420 38156
rect 3628 38116 3668 38156
rect 4204 38116 4244 38156
rect 5452 38116 5492 38156
rect 5875 38116 5915 38156
rect 6370 38116 6410 38156
rect 6988 38116 7028 38156
rect 8236 38116 8276 38156
rect 8812 38116 8852 38156
rect 10060 38116 10100 38156
rect 1603 38032 1643 38072
rect 6556 38032 6596 38072
rect 3820 37948 3860 37988
rect 5644 37948 5684 37988
rect 6076 37948 6116 37988
rect 4928 37780 4968 37820
rect 5010 37780 5050 37820
rect 5092 37780 5132 37820
rect 5174 37780 5214 37820
rect 5256 37780 5296 37820
rect 3571 37612 3611 37652
rect 5740 37612 5780 37652
rect 8227 37612 8267 37652
rect 3100 37528 3140 37568
rect 1315 37444 1355 37484
rect 1987 37435 2027 37475
rect 2140 37444 2180 37484
rect 2467 37435 2507 37475
rect 2620 37444 2660 37484
rect 2947 37435 2987 37475
rect 3766 37444 3806 37484
rect 4003 37444 4043 37484
rect 4108 37444 4148 37484
rect 4492 37444 4532 37484
rect 5068 37435 5108 37475
rect 5548 37435 5588 37475
rect 6124 37444 6164 37484
rect 7372 37435 7412 37475
rect 7747 37435 7787 37475
rect 7900 37444 7940 37484
rect 9096 37435 9136 37475
rect 10348 37444 10388 37484
rect 4588 37360 4628 37400
rect 8524 37360 8564 37400
rect 8764 37276 8804 37316
rect 1516 37192 1556 37232
rect 7564 37192 7604 37232
rect 8908 37192 8948 37232
rect 3688 37024 3728 37064
rect 3770 37024 3810 37064
rect 3852 37024 3892 37064
rect 3934 37024 3974 37064
rect 4016 37024 4056 37064
rect 3532 36688 3572 36728
rect 5644 36688 5684 36728
rect 7756 36688 7796 36728
rect 9964 36688 10004 36728
rect 10348 36688 10388 36728
rect 1324 36604 1364 36644
rect 2572 36604 2612 36644
rect 3043 36604 3083 36644
rect 3148 36604 3188 36644
rect 3628 36604 3668 36644
rect 4108 36604 4148 36644
rect 4596 36604 4636 36644
rect 5155 36604 5195 36644
rect 5260 36604 5300 36644
rect 5740 36604 5780 36644
rect 6220 36604 6260 36644
rect 6739 36604 6779 36644
rect 7267 36604 7307 36644
rect 7372 36604 7412 36644
rect 7852 36604 7892 36644
rect 8332 36604 8372 36644
rect 8820 36604 8860 36644
rect 9235 36604 9275 36644
rect 2764 36520 2804 36560
rect 10204 36520 10244 36560
rect 4780 36436 4820 36476
rect 6892 36436 6932 36476
rect 9004 36436 9044 36476
rect 9436 36436 9476 36476
rect 10588 36436 10628 36476
rect 4928 36268 4968 36308
rect 5010 36268 5050 36308
rect 5092 36268 5132 36308
rect 5174 36268 5214 36308
rect 5256 36268 5296 36308
rect 1852 36100 1892 36140
rect 4387 36100 4427 36140
rect 8620 36100 8660 36140
rect 10531 36100 10571 36140
rect 1372 36016 1412 36056
rect 1219 35923 1259 35963
rect 1699 35923 1739 35963
rect 2179 35923 2219 35963
rect 2668 35932 2708 35972
rect 3916 35923 3956 35963
rect 4675 35932 4715 35972
rect 4780 35932 4820 35972
rect 5164 35932 5204 35972
rect 5740 35923 5780 35963
rect 6220 35923 6260 35963
rect 6451 35932 6491 35972
rect 6595 35923 6635 35963
rect 7180 35932 7220 35972
rect 8428 35923 8468 35963
rect 9004 35923 9044 35963
rect 10252 35932 10292 35972
rect 2332 35848 2372 35888
rect 5260 35848 5300 35888
rect 6748 35848 6788 35888
rect 4108 35764 4148 35804
rect 8812 35764 8852 35804
rect 3688 35512 3728 35552
rect 3770 35512 3810 35552
rect 3852 35512 3892 35552
rect 3934 35512 3974 35552
rect 4016 35512 4056 35552
rect 1468 35344 1508 35384
rect 3052 35344 3092 35384
rect 5452 35344 5492 35384
rect 5884 35260 5924 35300
rect 1228 35176 1268 35216
rect 5644 35176 5684 35216
rect 6028 35176 6068 35216
rect 6268 35176 6308 35216
rect 10348 35176 10388 35216
rect 1612 35092 1652 35132
rect 2860 35092 2900 35132
rect 3187 35092 3227 35132
rect 4012 35092 4052 35132
rect 5260 35092 5300 35132
rect 6412 35092 6452 35132
rect 7660 35092 7700 35132
rect 8536 35092 8576 35132
rect 8716 35092 8756 35132
rect 9964 35092 10004 35132
rect 8371 35008 8411 35048
rect 3388 34924 3428 34964
rect 3811 34924 3851 34964
rect 7852 34924 7892 34964
rect 10156 34924 10196 34964
rect 10588 34924 10628 34964
rect 4928 34756 4968 34796
rect 5010 34756 5050 34796
rect 5092 34756 5132 34796
rect 5174 34756 5214 34796
rect 5256 34756 5296 34796
rect 7516 34588 7556 34628
rect 10531 34588 10571 34628
rect 7372 34504 7412 34544
rect 1219 34411 1259 34451
rect 1996 34420 2036 34460
rect 3244 34411 3284 34451
rect 3916 34420 3956 34460
rect 5164 34411 5204 34451
rect 5932 34420 5972 34460
rect 7180 34411 7220 34451
rect 8035 34420 8075 34460
rect 8140 34420 8180 34460
rect 8524 34420 8564 34460
rect 9100 34411 9140 34451
rect 9580 34411 9620 34451
rect 9811 34420 9851 34460
rect 9955 34411 9995 34451
rect 1372 34336 1412 34376
rect 1804 34336 1844 34376
rect 3628 34336 3668 34376
rect 5548 34336 5588 34376
rect 7756 34336 7796 34376
rect 8620 34336 8660 34376
rect 10108 34336 10148 34376
rect 3436 34168 3476 34208
rect 5356 34168 5396 34208
rect 5788 34168 5828 34208
rect 3688 34000 3728 34040
rect 3770 34000 3810 34040
rect 3852 34000 3892 34040
rect 3934 34000 3974 34040
rect 4016 34000 4056 34040
rect 3964 33664 4004 33704
rect 4444 33664 4484 33704
rect 6412 33664 6452 33704
rect 6748 33664 6788 33704
rect 6988 33664 7028 33704
rect 7180 33664 7220 33704
rect 7852 33664 7892 33704
rect 8716 33664 8756 33704
rect 1171 33580 1211 33620
rect 1708 33580 1748 33620
rect 2956 33580 2996 33620
rect 3328 33580 3368 33620
rect 3778 33580 3818 33620
rect 4288 33580 4328 33620
rect 4780 33580 4820 33620
rect 6028 33580 6068 33620
rect 7468 33580 7508 33620
rect 8227 33580 8267 33620
rect 8332 33580 8372 33620
rect 8812 33580 8852 33620
rect 9292 33580 9332 33620
rect 9811 33580 9851 33620
rect 10099 33580 10139 33620
rect 6652 33496 6692 33536
rect 1372 33412 1412 33452
rect 3148 33412 3188 33452
rect 3484 33412 3524 33452
rect 6220 33412 6260 33452
rect 7267 33412 7307 33452
rect 9964 33412 10004 33452
rect 10300 33412 10340 33452
rect 4928 33244 4968 33284
rect 5010 33244 5050 33284
rect 5092 33244 5132 33284
rect 5174 33244 5214 33284
rect 5256 33244 5296 33284
rect 1516 33076 1556 33116
rect 5452 33076 5492 33116
rect 9772 33076 9812 33116
rect 10531 33076 10571 33116
rect 7756 32992 7796 33032
rect 1315 32908 1355 32948
rect 1996 32908 2036 32948
rect 3244 32899 3284 32939
rect 3715 32908 3755 32948
rect 3820 32908 3860 32948
rect 4204 32908 4244 32948
rect 4780 32899 4820 32939
rect 5260 32899 5300 32939
rect 5635 32899 5675 32939
rect 6316 32908 6356 32948
rect 7564 32899 7604 32939
rect 8035 32908 8075 32948
rect 8140 32908 8180 32948
rect 8528 32908 8568 32948
rect 9100 32899 9140 32939
rect 9580 32899 9620 32939
rect 9955 32899 9995 32939
rect 4300 32824 4340 32864
rect 5788 32824 5828 32864
rect 8620 32824 8660 32864
rect 10108 32824 10148 32864
rect 1516 32656 1556 32696
rect 3436 32656 3476 32696
rect 3688 32488 3728 32528
rect 3770 32488 3810 32528
rect 3852 32488 3892 32528
rect 3934 32488 3974 32528
rect 4016 32488 4056 32528
rect 7852 32320 7892 32360
rect 9820 32236 9860 32276
rect 3436 32152 3476 32192
rect 8179 32152 8219 32192
rect 9004 32152 9044 32192
rect 9292 32152 9332 32192
rect 9580 32152 9620 32192
rect 9964 32152 10004 32192
rect 10348 32152 10388 32192
rect 1228 32068 1268 32108
rect 2476 32068 2516 32108
rect 2947 32068 2987 32108
rect 3052 32068 3092 32108
rect 3532 32068 3572 32108
rect 4012 32068 4052 32108
rect 4500 32068 4540 32108
rect 4819 32068 4859 32108
rect 5314 32068 5354 32108
rect 5836 32068 5876 32108
rect 6412 32068 6452 32108
rect 7660 32068 7700 32108
rect 8344 32068 8384 32108
rect 8524 32068 8564 32108
rect 2668 31984 2708 32024
rect 10204 31984 10244 32024
rect 4684 31900 4724 31940
rect 5020 31900 5060 31940
rect 5500 31900 5540 31940
rect 6115 31900 6155 31940
rect 9091 31900 9131 31940
rect 10588 31900 10628 31940
rect 4928 31732 4968 31772
rect 5010 31732 5050 31772
rect 5092 31732 5132 31772
rect 5174 31732 5214 31772
rect 5256 31732 5296 31772
rect 2620 31564 2660 31604
rect 3196 31564 3236 31604
rect 5164 31564 5204 31604
rect 7075 31564 7115 31604
rect 8179 31564 8219 31604
rect 6220 31480 6260 31520
rect 7276 31480 7316 31520
rect 7708 31480 7748 31520
rect 1315 31396 1355 31436
rect 1987 31387 2027 31427
rect 2467 31387 2507 31427
rect 3427 31396 3467 31436
rect 3532 31396 3572 31436
rect 3916 31396 3956 31436
rect 4492 31387 4532 31427
rect 4972 31387 5012 31427
rect 5347 31387 5387 31427
rect 6508 31396 6548 31436
rect 7555 31387 7595 31427
rect 8611 31396 8651 31436
rect 8716 31396 8756 31436
rect 2140 31312 2180 31352
rect 2956 31312 2996 31352
rect 4012 31312 4052 31352
rect 5500 31312 5540 31352
rect 8371 31354 8411 31394
rect 9100 31396 9140 31436
rect 9676 31387 9716 31427
rect 10156 31387 10196 31427
rect 5836 31312 5876 31352
rect 9196 31312 9236 31352
rect 1516 31144 1556 31184
rect 6076 31144 6116 31184
rect 10387 31144 10427 31184
rect 3688 30976 3728 31016
rect 3770 30976 3810 31016
rect 3852 30976 3892 31016
rect 3934 30976 3974 31016
rect 4016 30976 4056 31016
rect 9292 30808 9332 30848
rect 10396 30808 10436 30848
rect 3868 30640 3908 30680
rect 10156 30640 10196 30680
rect 1420 30556 1460 30596
rect 2668 30556 2708 30596
rect 3340 30556 3380 30596
rect 3459 30556 3499 30596
rect 3577 30556 3617 30596
rect 3712 30556 3752 30596
rect 4204 30556 4244 30596
rect 4396 30556 4436 30596
rect 4588 30556 4628 30596
rect 5836 30556 5876 30596
rect 6220 30556 6260 30596
rect 7468 30556 7508 30596
rect 10003 30598 10043 30638
rect 7852 30556 7892 30596
rect 9100 30556 9140 30596
rect 2860 30388 2900 30428
rect 3244 30388 3284 30428
rect 4300 30388 4340 30428
rect 6028 30388 6068 30428
rect 7660 30388 7700 30428
rect 9811 30388 9851 30428
rect 4928 30220 4968 30260
rect 5010 30220 5050 30260
rect 5092 30220 5132 30260
rect 5174 30220 5214 30260
rect 5256 30220 5296 30260
rect 2668 30052 2708 30092
rect 5212 30052 5252 30092
rect 4387 30010 4427 30050
rect 7852 30052 7892 30092
rect 10540 30052 10580 30092
rect 1228 29884 1268 29924
rect 2476 29875 2516 29915
rect 2987 29866 3027 29906
rect 3104 29884 3144 29924
rect 3226 29884 3266 29924
rect 3436 29884 3476 29924
rect 3724 29884 3764 29924
rect 4156 29884 4196 29924
rect 4457 29884 4497 29924
rect 4611 29884 4651 29924
rect 4771 29875 4811 29915
rect 6115 29884 6155 29924
rect 6225 29884 6265 29924
rect 6604 29884 6644 29924
rect 7180 29875 7220 29915
rect 7660 29875 7700 29915
rect 8035 29875 8075 29915
rect 9100 29884 9140 29924
rect 10348 29875 10388 29915
rect 4300 29800 4340 29840
rect 4924 29800 4964 29840
rect 5452 29800 5492 29840
rect 5836 29800 5876 29840
rect 6700 29800 6740 29840
rect 8188 29800 8228 29840
rect 8716 29800 8756 29840
rect 3148 29632 3188 29672
rect 3916 29632 3956 29672
rect 5596 29632 5636 29672
rect 8956 29632 8996 29672
rect 3688 29464 3728 29504
rect 3770 29464 3810 29504
rect 3852 29464 3892 29504
rect 3934 29464 3974 29504
rect 4016 29464 4056 29504
rect 3139 29296 3179 29336
rect 4204 29296 4244 29336
rect 2419 29128 2459 29168
rect 2764 29128 2804 29168
rect 5164 29128 5204 29168
rect 7084 29128 7124 29168
rect 9292 29128 9332 29168
rect 10348 29128 10388 29168
rect 1171 29044 1211 29084
rect 1666 29044 1706 29084
rect 2584 29044 2624 29084
rect 3139 29044 3179 29084
rect 3257 29044 3297 29084
rect 3389 29044 3429 29084
rect 3523 29044 3563 29084
rect 3700 29044 3740 29084
rect 3907 29044 3947 29084
rect 4204 29044 4244 29084
rect 4675 29044 4715 29084
rect 4780 29044 4820 29084
rect 5260 29044 5300 29084
rect 5740 29044 5780 29084
rect 6228 29044 6268 29084
rect 6451 29044 6491 29084
rect 6547 29044 6587 29084
rect 7564 29044 7604 29084
rect 8812 29044 8852 29084
rect 10006 29044 10046 29084
rect 1852 28960 1892 29000
rect 3004 28960 3044 29000
rect 1372 28876 1412 28916
rect 6748 28876 6788 28916
rect 7075 28876 7115 28916
rect 9004 28876 9044 28916
rect 9532 28876 9572 28916
rect 9811 28876 9851 28916
rect 10588 28876 10628 28916
rect 4928 28708 4968 28748
rect 5010 28708 5050 28748
rect 5092 28708 5132 28748
rect 5174 28708 5214 28748
rect 5256 28708 5296 28748
rect 2860 28540 2900 28580
rect 3724 28540 3764 28580
rect 6220 28540 6260 28580
rect 6883 28540 6923 28580
rect 7171 28540 7211 28580
rect 7555 28540 7595 28580
rect 7939 28540 7979 28580
rect 10252 28540 10292 28580
rect 10531 28540 10571 28580
rect 3187 28456 3227 28496
rect 3628 28456 3668 28496
rect 3834 28456 3874 28496
rect 4108 28456 4148 28496
rect 10444 28456 10484 28496
rect 1420 28372 1460 28412
rect 2668 28363 2708 28403
rect 3352 28372 3392 28412
rect 3523 28372 3563 28412
rect 4012 28372 4052 28412
rect 4195 28372 4235 28412
rect 4483 28372 4523 28412
rect 4588 28372 4628 28412
rect 4972 28372 5012 28412
rect 5548 28363 5588 28403
rect 6028 28363 6068 28403
rect 6403 28363 6443 28403
rect 8515 28372 8555 28412
rect 8620 28372 8660 28412
rect 9004 28372 9044 28412
rect 9580 28363 9620 28403
rect 10060 28363 10100 28403
rect 5068 28288 5108 28328
rect 6556 28288 6596 28328
rect 7852 28288 7892 28328
rect 8140 28288 8180 28328
rect 9100 28288 9140 28328
rect 3688 27952 3728 27992
rect 3770 27952 3810 27992
rect 3852 27952 3892 27992
rect 3934 27952 3974 27992
rect 4016 27952 4056 27992
rect 3916 27784 3956 27824
rect 5932 27784 5972 27824
rect 10348 27784 10388 27824
rect 4348 27700 4388 27740
rect 2131 27616 2171 27656
rect 4108 27616 4148 27656
rect 8140 27616 8180 27656
rect 1171 27532 1211 27572
rect 2326 27532 2366 27572
rect 2476 27532 2516 27572
rect 3724 27532 3764 27572
rect 4492 27532 4532 27572
rect 5740 27532 5780 27572
rect 6220 27532 6260 27572
rect 7468 27532 7508 27572
rect 8371 27532 8411 27572
rect 8908 27532 8948 27572
rect 10156 27532 10196 27572
rect 7660 27448 7700 27488
rect 1372 27364 1412 27404
rect 1795 27364 1835 27404
rect 7939 27364 7979 27404
rect 8227 27364 8267 27404
rect 8572 27364 8612 27404
rect 4928 27196 4968 27236
rect 5010 27196 5050 27236
rect 5092 27196 5132 27236
rect 5174 27196 5214 27236
rect 5256 27196 5296 27236
rect 1708 27028 1748 27068
rect 2140 27028 2180 27068
rect 3100 27028 3140 27068
rect 4684 27028 4724 27068
rect 8332 27028 8372 27068
rect 2620 26944 2660 26984
rect 6316 26944 6356 26984
rect 1219 26851 1259 26891
rect 1987 26851 2027 26891
rect 2467 26851 2507 26891
rect 2956 26860 2996 26900
rect 3244 26860 3284 26900
rect 4492 26851 4532 26891
rect 4876 26860 4916 26900
rect 6124 26851 6164 26891
rect 6595 26860 6635 26900
rect 6700 26860 6740 26900
rect 7084 26860 7124 26900
rect 7660 26851 7700 26891
rect 8140 26851 8180 26891
rect 8515 26851 8555 26891
rect 9100 26860 9140 26900
rect 10348 26851 10388 26891
rect 1372 26776 1412 26816
rect 7180 26776 7220 26816
rect 8668 26776 8708 26816
rect 10540 26608 10580 26648
rect 3688 26440 3728 26480
rect 3770 26440 3810 26480
rect 3852 26440 3892 26480
rect 3934 26440 3974 26480
rect 4016 26440 4056 26480
rect 4636 26272 4676 26312
rect 5020 26272 5060 26312
rect 9628 26272 9668 26312
rect 10204 26188 10244 26228
rect 1372 26104 1412 26144
rect 3676 26104 3716 26144
rect 4396 26104 4436 26144
rect 4780 26104 4820 26144
rect 5452 26104 5492 26144
rect 6316 26104 6356 26144
rect 6892 26104 6932 26144
rect 9388 26104 9428 26144
rect 9964 26104 10004 26144
rect 10348 26104 10388 26144
rect 1171 26020 1211 26060
rect 1804 26020 1844 26060
rect 3052 26020 3092 26060
rect 3475 26020 3515 26060
rect 4012 26020 4052 26060
rect 4195 26020 4235 26060
rect 7756 26020 7796 26060
rect 9004 26020 9044 26060
rect 10588 25936 10628 25976
rect 3244 25852 3284 25892
rect 4108 25852 4148 25892
rect 5251 25852 5291 25892
rect 5731 25852 5771 25892
rect 6115 25852 6155 25892
rect 6691 25852 6731 25892
rect 7267 25852 7307 25892
rect 7555 25852 7595 25892
rect 9196 25852 9236 25892
rect 4928 25684 4968 25724
rect 5010 25684 5050 25724
rect 5092 25684 5132 25724
rect 5174 25684 5214 25724
rect 5256 25684 5296 25724
rect 4732 25516 4772 25556
rect 4838 25516 4878 25556
rect 9676 25516 9716 25556
rect 3148 25432 3188 25472
rect 4396 25432 4436 25472
rect 7468 25432 7508 25472
rect 1228 25348 1268 25388
rect 2476 25339 2516 25379
rect 2947 25348 2987 25388
rect 3244 25348 3284 25388
rect 3436 25348 3476 25388
rect 3561 25348 3601 25388
rect 3724 25348 3764 25388
rect 4012 25348 4052 25388
rect 4291 25348 4331 25388
rect 4963 25348 5003 25388
rect 5068 25339 5108 25379
rect 5500 25348 5540 25388
rect 5644 25348 5684 25388
rect 6028 25348 6068 25388
rect 7276 25339 7316 25379
rect 7939 25348 7979 25388
rect 8044 25348 8084 25388
rect 8428 25348 8468 25388
rect 9004 25339 9044 25379
rect 9484 25339 9524 25379
rect 9859 25339 9899 25379
rect 10012 25348 10052 25388
rect 8524 25264 8564 25304
rect 10348 25264 10388 25304
rect 2668 25180 2708 25220
rect 3436 25096 3476 25136
rect 5356 25096 5396 25136
rect 10588 25096 10628 25136
rect 3688 24928 3728 24968
rect 3770 24928 3810 24968
rect 3852 24928 3892 24968
rect 3934 24928 3974 24968
rect 4016 24928 4056 24968
rect 2668 24760 2708 24800
rect 6028 24676 6068 24716
rect 10540 24676 10580 24716
rect 3619 24592 3659 24632
rect 3820 24592 3860 24632
rect 4323 24592 4363 24632
rect 6796 24592 6836 24632
rect 8380 24592 8420 24632
rect 1228 24508 1268 24548
rect 2476 24508 2516 24548
rect 3052 24508 3092 24548
rect 3194 24508 3234 24548
rect 3496 24508 3536 24548
rect 3724 24508 3764 24548
rect 4204 24508 4244 24548
rect 4421 24508 4461 24548
rect 4628 24508 4668 24548
rect 5836 24508 5876 24548
rect 6307 24508 6347 24548
rect 6412 24508 6452 24548
rect 6892 24508 6932 24548
rect 7372 24508 7412 24548
rect 7860 24508 7900 24548
rect 8083 24508 8123 24548
rect 8179 24508 8219 24548
rect 9100 24508 9140 24548
rect 10348 24508 10388 24548
rect 8716 24424 8756 24464
rect 2668 24340 2708 24380
rect 3340 24340 3380 24380
rect 4108 24340 4148 24380
rect 4928 24172 4968 24212
rect 5010 24172 5050 24212
rect 5092 24172 5132 24212
rect 5174 24172 5214 24212
rect 5256 24172 5296 24212
rect 4012 24004 4052 24044
rect 4780 24004 4820 24044
rect 5155 24004 5195 24044
rect 5731 24004 5771 24044
rect 7372 24004 7412 24044
rect 8419 24004 8459 24044
rect 1708 23920 1748 23960
rect 4348 23920 4388 23960
rect 7564 23920 7604 23960
rect 7852 23920 7892 23960
rect 8620 23920 8660 23960
rect 1324 23836 1364 23876
rect 1603 23836 1643 23876
rect 2275 23836 2315 23876
rect 2380 23836 2420 23876
rect 2764 23836 2804 23876
rect 3339 23827 3379 23867
rect 3820 23827 3860 23867
rect 4195 23827 4235 23867
rect 4684 23836 4724 23876
rect 4876 23836 4916 23876
rect 5932 23836 5972 23876
rect 7180 23827 7220 23867
rect 9100 23827 9140 23867
rect 10348 23836 10388 23876
rect 2860 23752 2900 23792
rect 5356 23752 5396 23792
rect 8332 23752 8372 23792
rect 1996 23668 2036 23708
rect 8908 23584 8948 23624
rect 3688 23416 3728 23456
rect 3770 23416 3810 23456
rect 3852 23416 3892 23456
rect 3934 23416 3974 23456
rect 4016 23416 4056 23456
rect 3436 23248 3476 23288
rect 5788 23248 5828 23288
rect 5068 23164 5108 23204
rect 6124 23080 6164 23120
rect 6604 23080 6644 23120
rect 8524 23080 8564 23120
rect 1171 22996 1211 23036
rect 1666 22996 1706 23036
rect 2146 22996 2186 23036
rect 2764 22996 2804 23036
rect 3043 22996 3083 23036
rect 3586 22996 3626 23036
rect 4066 22996 4106 23036
rect 4588 22996 4628 23036
rect 4876 22996 4916 23036
rect 5068 22996 5108 23036
rect 5260 22996 5300 23036
rect 5644 22996 5684 23036
rect 6976 22996 7016 23036
rect 7132 22996 7172 23036
rect 8035 22996 8075 23036
rect 8140 22996 8180 23036
rect 8620 22996 8660 23036
rect 9100 22996 9140 23036
rect 9619 22996 9659 23036
rect 9907 22996 9947 23036
rect 10444 22996 10484 23036
rect 2332 22912 2372 22952
rect 3148 22912 3188 22952
rect 1372 22828 1412 22868
rect 1852 22828 1892 22868
rect 3772 22828 3812 22868
rect 4252 22828 4292 22868
rect 4675 22828 4715 22868
rect 5884 22828 5924 22868
rect 6403 22828 6443 22868
rect 7555 22828 7595 22868
rect 9772 22828 9812 22868
rect 10108 22828 10148 22868
rect 4928 22660 4968 22700
rect 5010 22660 5050 22700
rect 5092 22660 5132 22700
rect 5174 22660 5214 22700
rect 5256 22660 5296 22700
rect 5740 22492 5780 22532
rect 7747 22492 7787 22532
rect 8035 22492 8075 22532
rect 9868 22492 9908 22532
rect 10588 22492 10628 22532
rect 2668 22408 2708 22448
rect 1228 22324 1268 22364
rect 2476 22315 2516 22355
rect 3148 22324 3188 22364
rect 3257 22324 3297 22364
rect 3532 22324 3572 22364
rect 4003 22324 4043 22364
rect 4108 22324 4148 22364
rect 4492 22324 4532 22364
rect 5068 22315 5108 22355
rect 5548 22315 5588 22355
rect 6316 22315 6356 22355
rect 7564 22324 7604 22364
rect 8428 22324 8468 22364
rect 9676 22315 9716 22355
rect 4588 22240 4628 22280
rect 6115 22240 6155 22280
rect 10060 22240 10100 22280
rect 10348 22240 10388 22280
rect 2860 22156 2900 22196
rect 3688 21904 3728 21944
rect 3770 21904 3810 21944
rect 3852 21904 3892 21944
rect 3934 21904 3974 21944
rect 4016 21904 4056 21944
rect 2668 21736 2708 21776
rect 8716 21736 8756 21776
rect 10588 21736 10628 21776
rect 1372 21568 1412 21608
rect 3436 21568 3476 21608
rect 6691 21568 6731 21608
rect 8332 21568 8372 21608
rect 10348 21568 10388 21608
rect 1171 21484 1211 21524
rect 1996 21484 2036 21524
rect 2275 21484 2315 21524
rect 2947 21484 2987 21524
rect 3052 21484 3092 21524
rect 3532 21484 3572 21524
rect 4012 21484 4052 21524
rect 4500 21484 4540 21524
rect 4972 21484 5012 21524
rect 5227 21484 5267 21524
rect 5347 21484 5387 21524
rect 5923 21484 5963 21524
rect 6028 21517 6068 21557
rect 6892 21484 6932 21524
rect 8140 21484 8180 21524
rect 8908 21484 8948 21524
rect 10156 21484 10196 21524
rect 2380 21400 2420 21440
rect 6355 21400 6395 21440
rect 4684 21316 4724 21356
rect 5692 21316 5732 21356
rect 5827 21307 5867 21347
rect 8572 21316 8612 21356
rect 4928 21148 4968 21188
rect 5010 21148 5050 21188
rect 5092 21148 5132 21188
rect 5174 21148 5214 21188
rect 5256 21148 5296 21188
rect 1372 20980 1412 21020
rect 5548 20980 5588 21020
rect 6499 20980 6539 21020
rect 7075 20980 7115 21020
rect 2284 20896 2324 20936
rect 3244 20896 3284 20936
rect 7276 20896 7316 20936
rect 1219 20803 1259 20843
rect 1900 20812 1940 20852
rect 2179 20812 2219 20852
rect 2860 20812 2900 20852
rect 3139 20812 3179 20852
rect 3811 20812 3851 20852
rect 3916 20812 3956 20852
rect 4300 20812 4340 20852
rect 4876 20803 4916 20843
rect 5356 20803 5396 20843
rect 5687 20812 5727 20852
rect 5932 20812 5972 20852
rect 6167 20812 6207 20852
rect 6412 20812 6452 20852
rect 7468 20803 7508 20843
rect 8716 20812 8756 20852
rect 9100 20803 9140 20843
rect 10348 20812 10388 20852
rect 4396 20728 4436 20768
rect 5827 20728 5867 20768
rect 6028 20728 6068 20768
rect 6307 20728 6347 20768
rect 6700 20728 6740 20768
rect 8908 20644 8948 20684
rect 2572 20560 2612 20600
rect 3532 20560 3572 20600
rect 3688 20392 3728 20432
rect 3770 20392 3810 20432
rect 3852 20392 3892 20432
rect 3934 20392 3974 20432
rect 4016 20392 4056 20432
rect 5932 20224 5972 20264
rect 2764 20140 2804 20180
rect 5164 20140 5204 20180
rect 8764 20140 8804 20180
rect 3532 20056 3572 20096
rect 8524 20056 8564 20096
rect 1171 19972 1211 20012
rect 1804 19972 1844 20012
rect 2092 19972 2132 20012
rect 2371 19972 2411 20012
rect 3043 19971 3083 20011
rect 3148 19972 3188 20012
rect 3628 19972 3668 20012
rect 4108 19972 4148 20012
rect 4627 19972 4667 20012
rect 4972 19972 5012 20012
rect 5097 19972 5137 20012
rect 5260 19972 5300 20012
rect 5596 19972 5636 20012
rect 5740 19972 5780 20012
rect 5932 19972 5972 20012
rect 6124 19972 6164 20012
rect 6604 19972 6644 20012
rect 7852 19972 7892 20012
rect 8908 19972 8948 20012
rect 10156 19972 10196 20012
rect 2476 19888 2516 19928
rect 8236 19888 8276 19928
rect 1372 19804 1412 19844
rect 4780 19804 4820 19844
rect 5443 19804 5483 19844
rect 6403 19804 6443 19844
rect 8044 19804 8084 19844
rect 10348 19804 10388 19844
rect 4928 19636 4968 19676
rect 5010 19636 5050 19676
rect 5092 19636 5132 19676
rect 5174 19636 5214 19676
rect 5256 19636 5296 19676
rect 3196 19468 3236 19508
rect 3676 19468 3716 19508
rect 8620 19468 8660 19508
rect 2572 19384 2612 19424
rect 4636 19384 4676 19424
rect 6604 19384 6644 19424
rect 1219 19291 1259 19331
rect 1372 19300 1412 19340
rect 2140 19300 2180 19340
rect 2467 19300 2507 19340
rect 3043 19291 3083 19331
rect 3523 19291 3563 19331
rect 4003 19291 4043 19331
rect 4483 19291 4523 19331
rect 5164 19300 5204 19340
rect 6412 19291 6452 19331
rect 6883 19300 6923 19340
rect 6988 19300 7028 19340
rect 7372 19300 7412 19340
rect 7948 19291 7988 19331
rect 8428 19291 8468 19331
rect 9292 19291 9332 19331
rect 10540 19300 10580 19340
rect 1708 19216 1748 19256
rect 4156 19216 4196 19256
rect 7468 19216 7508 19256
rect 8812 19216 8852 19256
rect 2860 19132 2900 19172
rect 1948 19048 1988 19088
rect 9100 19048 9140 19088
rect 3688 18880 3728 18920
rect 3770 18880 3810 18920
rect 3852 18880 3892 18920
rect 3934 18880 3974 18920
rect 4016 18880 4056 18920
rect 7324 18712 7364 18752
rect 4348 18628 4388 18668
rect 1372 18544 1412 18584
rect 2476 18544 2516 18584
rect 4060 18544 4100 18584
rect 4588 18544 4628 18584
rect 4972 18544 5012 18584
rect 7084 18544 7124 18584
rect 7468 18544 7508 18584
rect 8524 18544 8564 18584
rect 1171 18460 1211 18500
rect 1987 18460 2027 18500
rect 2092 18460 2132 18500
rect 2572 18460 2612 18500
rect 3052 18460 3092 18500
rect 3540 18460 3580 18500
rect 3907 18493 3947 18533
rect 5452 18460 5492 18500
rect 6700 18460 6740 18500
rect 8035 18460 8075 18500
rect 8140 18460 8180 18500
rect 8620 18460 8660 18500
rect 9100 18460 9140 18500
rect 9619 18460 9659 18500
rect 9907 18460 9947 18500
rect 3724 18292 3764 18332
rect 4732 18292 4772 18332
rect 5251 18292 5291 18332
rect 6892 18292 6932 18332
rect 7459 18292 7499 18332
rect 9772 18292 9812 18332
rect 10108 18292 10148 18332
rect 4928 18124 4968 18164
rect 5010 18124 5050 18164
rect 5092 18124 5132 18164
rect 5174 18124 5214 18164
rect 5256 18124 5296 18164
rect 3628 17956 3668 17996
rect 6220 17956 6260 17996
rect 9484 17956 9524 17996
rect 10588 17956 10628 17996
rect 1372 17872 1412 17912
rect 1219 17779 1259 17819
rect 1891 17788 1931 17828
rect 1996 17788 2036 17828
rect 2380 17788 2420 17828
rect 2956 17779 2996 17819
rect 3436 17779 3476 17819
rect 3916 17788 3956 17828
rect 4099 17788 4139 17828
rect 4204 17788 4244 17828
rect 4483 17788 4523 17828
rect 4588 17788 4628 17828
rect 4972 17788 5012 17828
rect 5548 17779 5588 17819
rect 6028 17779 6068 17819
rect 7747 17788 7787 17828
rect 7852 17788 7892 17828
rect 8236 17788 8276 17828
rect 8812 17779 8852 17819
rect 9292 17779 9332 17819
rect 2476 17704 2516 17744
rect 5068 17704 5108 17744
rect 6412 17704 6452 17744
rect 8332 17704 8372 17744
rect 9868 17704 9908 17744
rect 10348 17704 10388 17744
rect 4204 17536 4244 17576
rect 9628 17536 9668 17576
rect 3688 17368 3728 17408
rect 3770 17368 3810 17408
rect 3852 17368 3892 17408
rect 3934 17368 3974 17408
rect 4016 17368 4056 17408
rect 5251 17200 5291 17240
rect 9292 17200 9332 17240
rect 10588 17200 10628 17240
rect 3148 17116 3188 17156
rect 4588 17116 4628 17156
rect 3907 17032 3947 17072
rect 4108 17032 4148 17072
rect 6508 17032 6548 17072
rect 10156 17032 10196 17072
rect 10348 17032 10388 17072
rect 1171 16948 1211 16988
rect 1708 16948 1748 16988
rect 2956 16948 2996 16988
rect 3287 16948 3327 16988
rect 3427 16948 3467 16988
rect 3532 16948 3572 16988
rect 3767 16948 3807 16988
rect 4012 16948 4052 16988
rect 4291 16948 4331 16988
rect 4588 16948 4628 16988
rect 4780 16948 4820 16988
rect 4902 16948 4942 16988
rect 5029 16948 5069 16988
rect 5246 16948 5286 16988
rect 5548 16948 5588 16988
rect 5779 16948 5819 16988
rect 5882 16948 5922 16988
rect 7192 16948 7232 16988
rect 7330 16948 7370 16988
rect 7852 16948 7892 16988
rect 9100 16948 9140 16988
rect 9427 16948 9467 16988
rect 6268 16864 6308 16904
rect 9628 16864 9668 16904
rect 1372 16780 1412 16820
rect 3619 16780 3659 16820
rect 5068 16780 5108 16820
rect 5452 16780 5492 16820
rect 6028 16780 6068 16820
rect 7027 16780 7067 16820
rect 7516 16780 7556 16820
rect 9916 16780 9956 16820
rect 4928 16612 4968 16652
rect 5010 16612 5050 16652
rect 5092 16612 5132 16652
rect 5174 16612 5214 16652
rect 5256 16612 5296 16652
rect 4099 16444 4139 16484
rect 5059 16444 5099 16484
rect 5452 16444 5492 16484
rect 9580 16444 9620 16484
rect 3244 16360 3284 16400
rect 9859 16360 9899 16400
rect 1219 16267 1259 16307
rect 1804 16276 1844 16316
rect 3052 16267 3092 16307
rect 3916 16276 3956 16316
rect 4107 16276 4147 16316
rect 4267 16276 4307 16316
rect 4492 16276 4532 16316
rect 4732 16276 4772 16316
rect 4867 16276 4907 16316
rect 4972 16276 5012 16316
rect 5644 16267 5684 16307
rect 6892 16276 6932 16316
rect 7843 16276 7883 16316
rect 7948 16276 7988 16316
rect 8332 16276 8372 16316
rect 8908 16267 8948 16307
rect 9388 16267 9428 16307
rect 10252 16276 10292 16316
rect 1372 16192 1412 16232
rect 3628 16192 3668 16232
rect 4387 16192 4427 16232
rect 4588 16192 4628 16232
rect 8428 16192 8468 16232
rect 3388 16108 3428 16148
rect 3688 15856 3728 15896
rect 3770 15856 3810 15896
rect 3852 15856 3892 15896
rect 3934 15856 3974 15896
rect 4016 15856 4056 15896
rect 2668 15688 2708 15728
rect 3196 15688 3236 15728
rect 7564 15688 7604 15728
rect 9772 15688 9812 15728
rect 10588 15688 10628 15728
rect 2812 15604 2852 15644
rect 4732 15604 4772 15644
rect 3052 15520 3092 15560
rect 3436 15520 3476 15560
rect 3820 15520 3860 15560
rect 4204 15520 4244 15560
rect 4588 15520 4628 15560
rect 4972 15520 5012 15560
rect 10156 15520 10196 15560
rect 10348 15520 10388 15560
rect 1228 15436 1268 15476
rect 2476 15436 2516 15476
rect 5260 15436 5300 15476
rect 6124 15436 6164 15476
rect 7372 15436 7412 15476
rect 8332 15436 8372 15476
rect 9580 15436 9620 15476
rect 3580 15352 3620 15392
rect 3964 15268 4004 15308
rect 4348 15268 4388 15308
rect 5116 15268 5156 15308
rect 9916 15268 9956 15308
rect 4928 15100 4968 15140
rect 5010 15100 5050 15140
rect 5092 15100 5132 15140
rect 5174 15100 5214 15140
rect 5256 15100 5296 15140
rect 1564 14932 1604 14972
rect 4204 14932 4244 14972
rect 4492 14932 4532 14972
rect 10588 14932 10628 14972
rect 1948 14848 1988 14888
rect 7564 14848 7604 14888
rect 2467 14764 2507 14804
rect 2572 14764 2612 14804
rect 2956 14764 2996 14804
rect 3532 14755 3572 14795
rect 4012 14755 4052 14795
rect 4684 14755 4724 14795
rect 5932 14764 5972 14804
rect 6124 14764 6164 14804
rect 7372 14755 7412 14795
rect 7843 14764 7883 14804
rect 7948 14764 7988 14804
rect 8332 14764 8372 14804
rect 8908 14755 8948 14795
rect 9388 14755 9428 14795
rect 1228 14680 1268 14720
rect 1804 14680 1844 14720
rect 2188 14680 2228 14720
rect 3052 14680 3092 14720
rect 8428 14680 8468 14720
rect 9619 14680 9659 14720
rect 9964 14680 10004 14720
rect 10348 14680 10388 14720
rect 1468 14512 1508 14552
rect 9724 14512 9764 14552
rect 3688 14344 3728 14384
rect 3770 14344 3810 14384
rect 3852 14344 3892 14384
rect 3934 14344 3974 14384
rect 4016 14344 4056 14384
rect 4828 14176 4868 14216
rect 5788 14176 5828 14216
rect 9196 14176 9236 14216
rect 10588 14176 10628 14216
rect 1180 14092 1220 14132
rect 6268 14092 6308 14132
rect 10204 14092 10244 14132
rect 1420 14008 1460 14048
rect 1804 14008 1844 14048
rect 2188 14008 2228 14048
rect 3052 14008 3092 14048
rect 4339 14008 4379 14048
rect 4684 14008 4724 14048
rect 5068 14008 5108 14048
rect 5548 14008 5588 14048
rect 6028 14008 6068 14048
rect 9532 14008 9572 14048
rect 9964 14008 10004 14048
rect 10348 14008 10388 14048
rect 2563 13924 2603 13964
rect 2668 13924 2708 13964
rect 3148 13924 3188 13964
rect 3628 13924 3668 13964
rect 4147 13924 4187 13964
rect 7219 13924 7259 13964
rect 7756 13924 7796 13964
rect 9004 13924 9044 13964
rect 9376 13924 9416 13964
rect 1948 13840 1988 13880
rect 1564 13756 1604 13796
rect 4444 13756 4484 13796
rect 7420 13756 7460 13796
rect 4928 13588 4968 13628
rect 5010 13588 5050 13628
rect 5092 13588 5132 13628
rect 5174 13588 5214 13628
rect 5256 13588 5296 13628
rect 2860 13420 2900 13460
rect 4492 13420 4532 13460
rect 6124 13336 6164 13376
rect 7372 13336 7412 13376
rect 10252 13336 10292 13376
rect 1420 13252 1460 13292
rect 2668 13243 2708 13283
rect 3052 13252 3092 13292
rect 4300 13243 4340 13283
rect 4684 13252 4724 13292
rect 5932 13243 5972 13283
rect 6988 13252 7028 13292
rect 7267 13252 7307 13292
rect 8812 13252 8852 13292
rect 10060 13243 10100 13283
rect 8044 13168 8084 13208
rect 8428 13168 8468 13208
rect 7804 13084 7844 13124
rect 8668 13084 8708 13124
rect 7660 13000 7700 13040
rect 3688 12832 3728 12872
rect 3770 12832 3810 12872
rect 3852 12832 3892 12872
rect 3934 12832 3974 12872
rect 4016 12832 4056 12872
rect 2860 12664 2900 12704
rect 6076 12664 6116 12704
rect 9100 12664 9140 12704
rect 2668 12580 2708 12620
rect 8908 12580 8948 12620
rect 4684 12496 4724 12536
rect 5068 12496 5108 12536
rect 5452 12496 5492 12536
rect 6316 12496 6356 12536
rect 1228 12412 1268 12452
rect 2476 12412 2516 12452
rect 3052 12412 3092 12452
rect 4300 12412 4340 12452
rect 7222 12412 7262 12452
rect 8083 12412 8123 12452
rect 9292 12412 9332 12452
rect 10540 12412 10580 12452
rect 5212 12328 5252 12368
rect 4444 12244 4484 12284
rect 4828 12244 4868 12284
rect 7027 12244 7067 12284
rect 8284 12244 8324 12284
rect 4928 12076 4968 12116
rect 5010 12076 5050 12116
rect 5092 12076 5132 12116
rect 5174 12076 5214 12116
rect 5256 12076 5296 12116
rect 2956 11908 2996 11948
rect 3580 11908 3620 11948
rect 5932 11908 5972 11948
rect 7804 11908 7844 11948
rect 10540 11908 10580 11948
rect 1516 11740 1556 11780
rect 2764 11731 2804 11771
rect 3478 11740 3518 11780
rect 4174 11740 4214 11780
rect 4300 11740 4340 11780
rect 4684 11740 4724 11780
rect 5260 11731 5300 11771
rect 5740 11731 5780 11771
rect 6220 11740 6260 11780
rect 7468 11731 7508 11771
rect 8611 11740 8651 11780
rect 3283 11656 3323 11696
rect 3820 11656 3860 11696
rect 4780 11656 4820 11696
rect 8044 11656 8084 11696
rect 8236 11656 8276 11696
rect 7660 11488 7700 11528
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 1180 11152 1220 11192
rect 1564 11152 1604 11192
rect 3628 11152 3668 11192
rect 5836 11152 5876 11192
rect 10540 11152 10580 11192
rect 1420 10984 1460 11024
rect 1804 10984 1844 11024
rect 3820 10984 3860 11024
rect 4060 10984 4100 11024
rect 6700 10984 6740 11024
rect 2188 10900 2228 10940
rect 3436 10900 3476 10940
rect 4396 10900 4436 10940
rect 5644 10900 5684 10940
rect 6211 10900 6251 10940
rect 6316 10900 6356 10940
rect 6796 10900 6836 10940
rect 7276 10900 7316 10940
rect 7764 10900 7804 10940
rect 8611 10900 8651 10940
rect 8227 10816 8267 10856
rect 7948 10732 7988 10772
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 1180 10396 1220 10436
rect 3724 10396 3764 10436
rect 8380 10396 8420 10436
rect 10204 10396 10244 10436
rect 10588 10396 10628 10436
rect 1564 10312 1604 10352
rect 2284 10228 2324 10268
rect 3532 10219 3572 10259
rect 4291 10228 4331 10268
rect 4396 10228 4436 10268
rect 4780 10228 4820 10268
rect 5356 10219 5396 10259
rect 5836 10219 5876 10259
rect 1420 10144 1460 10184
rect 1804 10144 1844 10184
rect 4876 10144 4916 10184
rect 6067 10144 6107 10184
rect 6412 10144 6452 10184
rect 6796 10144 6836 10184
rect 8236 10144 8276 10184
rect 8620 10144 8660 10184
rect 8908 10144 8948 10184
rect 9148 10144 9188 10184
rect 9964 10144 10004 10184
rect 10348 10144 10388 10184
rect 6172 10060 6212 10100
rect 7996 10060 8036 10100
rect 9292 10060 9332 10100
rect 6556 9976 6596 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 3436 9640 3476 9680
rect 5452 9640 5492 9680
rect 8179 9640 8219 9680
rect 1180 9556 1220 9596
rect 1564 9556 1604 9596
rect 3580 9556 3620 9596
rect 8332 9556 8372 9596
rect 1420 9472 1460 9512
rect 1804 9472 1844 9512
rect 3820 9472 3860 9512
rect 6124 9472 6164 9512
rect 6892 9472 6932 9512
rect 10099 9472 10139 9512
rect 1996 9388 2036 9428
rect 3244 9388 3284 9428
rect 4012 9388 4052 9428
rect 5260 9388 5300 9428
rect 6403 9388 6443 9428
rect 6508 9388 6548 9428
rect 6988 9388 7028 9428
rect 7468 9388 7508 9428
rect 7987 9388 8027 9428
rect 8524 9388 8564 9428
rect 9772 9388 9812 9428
rect 10294 9388 10334 9428
rect 5884 9220 5924 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 1468 8884 1508 8924
rect 3724 8884 3764 8924
rect 6652 8884 6692 8924
rect 8428 8884 8468 8924
rect 5452 8800 5492 8840
rect 6316 8800 6356 8840
rect 1315 8707 1355 8747
rect 1795 8707 1835 8747
rect 2284 8716 2324 8756
rect 3532 8707 3572 8747
rect 4012 8716 4052 8756
rect 5260 8707 5300 8747
rect 5932 8716 5972 8756
rect 6211 8716 6251 8756
rect 6988 8716 7028 8756
rect 8236 8707 8276 8747
rect 9100 8716 9140 8756
rect 10348 8707 10388 8747
rect 1948 8632 1988 8672
rect 8716 8632 8756 8672
rect 8956 8632 8996 8672
rect 10540 8464 10580 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 2956 8128 2996 8168
rect 6172 8128 6212 8168
rect 9004 8128 9044 8168
rect 5644 8044 5684 8084
rect 8428 8044 8468 8084
rect 1228 7960 1268 8000
rect 6028 7960 6068 8000
rect 6412 7960 6452 8000
rect 6556 7960 6596 8000
rect 6796 7960 6836 8000
rect 1516 7876 1556 7916
rect 2764 7876 2804 7916
rect 3148 7876 3188 7916
rect 4396 7876 4436 7916
rect 4972 7876 5012 7916
rect 5251 7876 5291 7916
rect 7756 7876 7796 7916
rect 8035 7876 8075 7916
rect 9196 7876 9236 7916
rect 10444 7876 10484 7916
rect 4588 7792 4628 7832
rect 5356 7792 5396 7832
rect 8140 7792 8180 7832
rect 5788 7708 5828 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 3004 7372 3044 7412
rect 7564 7372 7604 7412
rect 1228 7204 1268 7244
rect 2476 7195 2516 7235
rect 2851 7195 2891 7235
rect 4300 7204 4340 7244
rect 5548 7195 5588 7235
rect 6124 7204 6164 7244
rect 7372 7195 7412 7235
rect 8524 7204 8564 7244
rect 9772 7195 9812 7235
rect 3532 7120 3572 7160
rect 3916 7120 3956 7160
rect 8332 7120 8372 7160
rect 10348 7120 10388 7160
rect 2668 7036 2708 7076
rect 3292 7036 3332 7076
rect 9964 7036 10004 7076
rect 10588 7036 10628 7076
rect 3676 6952 3716 6992
rect 5740 6952 5780 6992
rect 8092 6952 8132 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 1372 6616 1412 6656
rect 10588 6616 10628 6656
rect 7756 6532 7796 6572
rect 1612 6448 1652 6488
rect 4588 6448 4628 6488
rect 9964 6448 10004 6488
rect 10348 6448 10388 6488
rect 1804 6364 1844 6404
rect 3052 6364 3092 6404
rect 4099 6364 4139 6404
rect 4204 6364 4244 6404
rect 4684 6364 4724 6404
rect 5164 6364 5204 6404
rect 5683 6364 5723 6404
rect 6316 6364 6356 6404
rect 7564 6364 7604 6404
rect 3244 6280 3284 6320
rect 10204 6280 10244 6320
rect 3523 6196 3563 6236
rect 3811 6196 3851 6236
rect 5836 6196 5876 6236
rect 6115 6196 6155 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 6211 5860 6251 5900
rect 8428 5860 8468 5900
rect 2860 5776 2900 5816
rect 1420 5692 1460 5732
rect 2668 5683 2708 5723
rect 3139 5692 3179 5732
rect 3244 5692 3284 5732
rect 3628 5692 3668 5732
rect 4204 5683 4244 5723
rect 4684 5683 4724 5723
rect 6691 5692 6731 5732
rect 6796 5692 6836 5732
rect 7180 5692 7220 5732
rect 7756 5683 7796 5723
rect 8236 5683 8276 5723
rect 8611 5683 8651 5723
rect 8764 5692 8804 5732
rect 3724 5608 3764 5648
rect 4915 5608 4955 5648
rect 5260 5608 5300 5648
rect 5644 5608 5684 5648
rect 5836 5608 5876 5648
rect 7276 5608 7316 5648
rect 9292 5608 9332 5648
rect 10348 5608 10388 5648
rect 6076 5524 6116 5564
rect 9052 5524 9092 5564
rect 5020 5440 5060 5480
rect 5404 5440 5444 5480
rect 10588 5440 10628 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 4012 5104 4052 5144
rect 8428 5104 8468 5144
rect 4876 4936 4916 4976
rect 6163 4936 6203 4976
rect 6508 4936 6548 4976
rect 1720 4852 1760 4892
rect 1888 4852 1928 4892
rect 2572 4852 2612 4892
rect 3820 4852 3860 4892
rect 4366 4852 4406 4892
rect 4489 4852 4529 4892
rect 4972 4852 5012 4892
rect 5452 4852 5492 4892
rect 5940 4852 5980 4892
rect 6988 4852 7028 4892
rect 8236 4852 8276 4892
rect 1555 4768 1595 4808
rect 2044 4684 2084 4724
rect 6268 4684 6308 4724
rect 6691 4684 6731 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 1219 4348 1259 4388
rect 3628 4348 3668 4388
rect 7180 4348 7220 4388
rect 7363 4348 7403 4388
rect 1852 4264 1892 4304
rect 5452 4264 5492 4304
rect 10051 4264 10091 4304
rect 1699 4171 1739 4211
rect 2188 4180 2228 4220
rect 3436 4171 3476 4211
rect 4012 4180 4052 4220
rect 5268 4180 5308 4220
rect 5740 4180 5780 4220
rect 6988 4171 7028 4211
rect 10444 4180 10484 4220
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 3100 3592 3140 3632
rect 3484 3592 3524 3632
rect 1564 3508 1604 3548
rect 1948 3508 1988 3548
rect 1804 3424 1844 3464
rect 2188 3424 2228 3464
rect 2332 3424 2372 3464
rect 2572 3424 2612 3464
rect 2956 3424 2996 3464
rect 3340 3424 3380 3464
rect 3724 3424 3764 3464
rect 3916 3424 3956 3464
rect 4492 3424 4532 3464
rect 4780 3424 4820 3464
rect 5644 3424 5684 3464
rect 5932 3424 5972 3464
rect 6508 3424 6548 3464
rect 6796 3424 6836 3464
rect 7084 3424 7124 3464
rect 10348 3424 10388 3464
rect 2716 3256 2756 3296
rect 1315 3172 1355 3212
rect 3907 3172 3947 3212
rect 4291 3172 4331 3212
rect 5155 3172 5195 3212
rect 5443 3172 5483 3212
rect 6307 3172 6347 3212
rect 6787 3172 6827 3212
rect 10588 3172 10628 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 1180 2836 1220 2876
rect 2716 2836 2756 2876
rect 3619 2836 3659 2876
rect 3907 2836 3947 2876
rect 5059 2836 5099 2876
rect 5827 2836 5867 2876
rect 2332 2752 2372 2792
rect 4396 2752 4436 2792
rect 4684 2752 4724 2792
rect 5260 2752 5300 2792
rect 5548 2752 5588 2792
rect 6124 2752 6164 2792
rect 6412 2752 6452 2792
rect 1612 2668 1652 2708
rect 1420 2584 1460 2624
rect 1948 2584 1988 2624
rect 2188 2584 2228 2624
rect 2572 2584 2612 2624
rect 2956 2584 2996 2624
rect 3340 2584 3380 2624
rect 4396 2584 4436 2624
rect 10348 2584 10388 2624
rect 3100 2416 3140 2456
rect 10588 2416 10628 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 1180 2080 1220 2120
rect 2332 2080 2372 2120
rect 2716 2080 2756 2120
rect 10051 2080 10091 2120
rect 1564 1996 1604 2036
rect 1420 1912 1460 1952
rect 1804 1912 1844 1952
rect 2188 1912 2228 1952
rect 2572 1912 2612 1952
rect 2956 1912 2996 1952
rect 3340 1912 3380 1952
rect 3724 1912 3764 1952
rect 4300 1912 4340 1952
rect 4588 1912 4628 1952
rect 5452 1912 5492 1952
rect 5164 1828 5204 1868
rect 10444 1828 10484 1868
rect 1948 1744 1988 1784
rect 3100 1744 3140 1784
rect 4012 1744 4052 1784
rect 5740 1744 5780 1784
rect 6028 1744 6068 1784
rect 3484 1660 3524 1700
rect 4867 1660 4907 1700
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
<< metal2 >>
rect 11750 46304 11840 46324
rect 10243 46264 10252 46304
rect 10292 46264 11840 46304
rect 11750 46244 11840 46264
rect 4919 45340 4928 45380
rect 4968 45340 5010 45380
rect 5050 45340 5092 45380
rect 5132 45340 5174 45380
rect 5214 45340 5256 45380
rect 5296 45340 5305 45380
rect 11750 45296 11840 45316
rect 5635 45256 5644 45296
rect 5684 45256 8468 45296
rect 11011 45256 11020 45296
rect 11060 45256 11840 45296
rect 2371 45172 2380 45212
rect 2420 45172 3484 45212
rect 3524 45172 3533 45212
rect 3907 45172 3916 45212
rect 3956 45172 3964 45212
rect 4004 45172 4087 45212
rect 4291 45172 4300 45212
rect 4340 45172 4348 45212
rect 4388 45172 4471 45212
rect 4675 45172 4684 45212
rect 4724 45172 4732 45212
rect 4772 45172 4855 45212
rect 5107 45172 5116 45212
rect 5156 45172 5356 45212
rect 5396 45172 5405 45212
rect 5539 45172 5548 45212
rect 5588 45172 5780 45212
rect 5827 45172 5836 45212
rect 5876 45172 5884 45212
rect 5924 45172 6007 45212
rect 6211 45172 6220 45212
rect 6260 45172 6268 45212
rect 6308 45172 6391 45212
rect 6595 45172 6604 45212
rect 6644 45172 6652 45212
rect 6692 45172 6775 45212
rect 6979 45172 6988 45212
rect 7028 45172 7036 45212
rect 7076 45172 7159 45212
rect 7363 45172 7372 45212
rect 7412 45172 7420 45212
rect 7460 45172 7543 45212
rect 7747 45172 7756 45212
rect 7796 45172 7804 45212
rect 7844 45172 7927 45212
rect 8131 45172 8140 45212
rect 8180 45172 8188 45212
rect 8228 45172 8311 45212
rect 5740 45128 5780 45172
rect 2083 45088 2092 45128
rect 2132 45088 2332 45128
rect 2372 45088 2381 45128
rect 3379 45088 3388 45128
rect 3428 45088 4532 45128
rect 5443 45088 5452 45128
rect 5492 45088 5500 45128
rect 5540 45088 5623 45128
rect 5740 45088 7700 45128
rect 1193 45004 1315 45044
rect 1364 45004 1373 45044
rect 1420 45004 2131 45044
rect 2171 45004 2180 45044
rect 2537 45035 2668 45044
rect 2537 45004 2659 45035
rect 2708 45004 2717 45044
rect 2803 45004 2812 45044
rect 2852 45004 3340 45044
rect 3380 45004 3389 45044
rect 0 44960 90 44980
rect 1420 44960 1460 45004
rect 2650 44995 2659 45004
rect 2699 44995 2708 45004
rect 2650 44994 2708 44995
rect 0 44920 1460 44960
rect 3017 44920 3148 44960
rect 3188 44920 3197 44960
rect 3244 44920 3724 44960
rect 3764 44920 3773 44960
rect 4195 44920 4204 44960
rect 4244 44920 4253 44960
rect 0 44900 90 44920
rect 3244 44876 3284 44920
rect 2275 44836 2284 44876
rect 2324 44836 3284 44876
rect 739 44752 748 44792
rect 788 44752 1516 44792
rect 1556 44752 1565 44792
rect 4204 44708 4244 44920
rect 4492 44792 4532 45088
rect 4588 45004 6124 45044
rect 6164 45004 6173 45044
rect 4588 44960 4628 45004
rect 7660 44960 7700 45088
rect 8428 44960 8468 45256
rect 11750 45236 11840 45256
rect 8515 45172 8524 45212
rect 8564 45172 8572 45212
rect 8612 45172 8695 45212
rect 8899 45172 8908 45212
rect 8948 45172 8956 45212
rect 8996 45172 9079 45212
rect 9283 45172 9292 45212
rect 9332 45172 9340 45212
rect 9380 45172 9463 45212
rect 9667 45172 9676 45212
rect 9716 45172 9724 45212
rect 9764 45172 9847 45212
rect 4579 44920 4588 44960
rect 4628 44920 4637 44960
rect 4841 44920 4972 44960
rect 5012 44920 5021 44960
rect 5225 44920 5356 44960
rect 5396 44920 5405 44960
rect 5609 44920 5740 44960
rect 5780 44920 5789 44960
rect 6115 44920 6124 44960
rect 6164 44920 6173 44960
rect 6377 44920 6508 44960
rect 6548 44920 6557 44960
rect 6883 44920 6892 44960
rect 6932 44920 6941 44960
rect 7145 44920 7276 44960
rect 7316 44920 7325 44960
rect 7651 44920 7660 44960
rect 7700 44920 7709 44960
rect 7913 44920 8044 44960
rect 8084 44920 8093 44960
rect 8419 44920 8428 44960
rect 8468 44920 8477 44960
rect 8803 44920 8812 44960
rect 8852 44920 8861 44960
rect 8908 44920 9196 44960
rect 9236 44920 9245 44960
rect 9449 44920 9580 44960
rect 9620 44920 9629 44960
rect 9833 44920 9964 44960
rect 10004 44920 10013 44960
rect 10217 44920 10348 44960
rect 10388 44920 10397 44960
rect 6124 44876 6164 44920
rect 5251 44836 5260 44876
rect 5300 44836 6164 44876
rect 6892 44876 6932 44920
rect 8812 44876 8852 44920
rect 6892 44836 7756 44876
rect 7796 44836 7805 44876
rect 7939 44836 7948 44876
rect 7988 44836 8852 44876
rect 8908 44792 8948 44920
rect 4492 44752 8948 44792
rect 10579 44752 10588 44792
rect 10628 44752 11692 44792
rect 11732 44752 11741 44792
rect 4204 44668 6796 44708
rect 6836 44668 6845 44708
rect 0 44624 90 44644
rect 0 44584 2668 44624
rect 2708 44584 2717 44624
rect 3679 44584 3688 44624
rect 3728 44584 3770 44624
rect 3810 44584 3852 44624
rect 3892 44584 3934 44624
rect 3974 44584 4016 44624
rect 4056 44584 4065 44624
rect 4492 44584 5492 44624
rect 0 44564 90 44584
rect 4492 44540 4532 44584
rect 3043 44500 3052 44540
rect 3092 44500 4532 44540
rect 4588 44500 5356 44540
rect 5396 44500 5405 44540
rect 4588 44456 4628 44500
rect 5452 44456 5492 44584
rect 3859 44416 3868 44456
rect 3908 44416 4628 44456
rect 5155 44416 5164 44456
rect 5204 44416 5212 44456
rect 5252 44416 5335 44456
rect 5452 44416 5596 44456
rect 5636 44416 5645 44456
rect 6115 44416 6124 44456
rect 6164 44416 6172 44456
rect 6212 44416 6295 44456
rect 6499 44416 6508 44456
rect 6548 44416 6556 44456
rect 6596 44416 6679 44456
rect 6787 44416 6796 44456
rect 6836 44416 7036 44456
rect 7076 44416 7085 44456
rect 7267 44416 7276 44456
rect 7316 44416 7420 44456
rect 7460 44416 7469 44456
rect 7747 44416 7756 44456
rect 7796 44416 7804 44456
rect 7844 44416 7927 44456
rect 9235 44416 9244 44456
rect 9284 44416 9580 44456
rect 9620 44416 9629 44456
rect 10121 44416 10204 44456
rect 10244 44416 10252 44456
rect 10292 44416 10301 44456
rect 10579 44416 10588 44456
rect 10628 44416 11020 44456
rect 11060 44416 11069 44456
rect 163 44332 172 44372
rect 212 44332 4436 44372
rect 5107 44332 5116 44372
rect 5156 44332 5260 44372
rect 5300 44332 5309 44372
rect 5836 44332 7948 44372
rect 7988 44332 7997 44372
rect 9619 44332 9628 44372
rect 9668 44332 9964 44372
rect 10004 44332 10013 44372
rect 0 44288 90 44308
rect 4396 44288 4436 44332
rect 5836 44288 5876 44332
rect 11750 44288 11840 44308
rect 0 44248 76 44288
rect 116 44248 125 44288
rect 2345 44248 2476 44288
rect 2516 44248 2525 44288
rect 2947 44248 2956 44288
rect 2996 44248 3628 44288
rect 3668 44248 3677 44288
rect 4003 44248 4012 44288
rect 4052 44248 4061 44288
rect 4387 44248 4396 44288
rect 4436 44248 4445 44288
rect 4675 44248 4684 44288
rect 4724 44248 4828 44288
rect 4868 44248 4877 44288
rect 5443 44248 5452 44288
rect 5492 44248 5501 44288
rect 5827 44248 5836 44288
rect 5876 44248 5885 44288
rect 6281 44248 6316 44288
rect 6356 44248 6412 44288
rect 6452 44248 6461 44288
rect 6665 44248 6796 44288
rect 6836 44248 6845 44288
rect 7145 44248 7276 44288
rect 7316 44248 7325 44288
rect 7529 44248 7660 44288
rect 7700 44248 7709 44288
rect 8035 44248 8044 44288
rect 8084 44248 8276 44288
rect 8873 44248 9004 44288
rect 9044 44248 9053 44288
rect 9257 44248 9388 44288
rect 9428 44248 9437 44288
rect 9955 44248 9964 44288
rect 10004 44248 10013 44288
rect 10217 44248 10252 44288
rect 10292 44248 10348 44288
rect 10388 44248 10397 44288
rect 11683 44248 11692 44288
rect 11732 44248 11840 44288
rect 0 44228 90 44248
rect 4012 44204 4052 44248
rect 5452 44204 5492 44248
rect 643 44164 652 44204
rect 692 44164 1315 44204
rect 1355 44164 1364 44204
rect 1804 44164 1939 44204
rect 1979 44164 1988 44204
rect 4012 44164 5396 44204
rect 5452 44164 6412 44204
rect 6452 44164 6461 44204
rect 547 43996 556 44036
rect 596 43996 1516 44036
rect 1556 43996 1565 44036
rect 0 43952 90 43972
rect 0 43912 76 43952
rect 116 43912 125 43952
rect 0 43892 90 43912
rect 0 43616 90 43636
rect 1804 43616 1844 44164
rect 5356 44120 5396 44164
rect 8236 44120 8276 44248
rect 2707 44080 2716 44120
rect 2756 44080 4972 44120
rect 5012 44080 5021 44120
rect 5356 44080 6220 44120
rect 6260 44080 6269 44120
rect 7171 44080 7180 44120
rect 7220 44080 8044 44120
rect 8084 44080 8093 44120
rect 8227 44080 8236 44120
rect 8276 44080 8524 44120
rect 8564 44080 8573 44120
rect 1891 43996 1900 44036
rect 1940 43996 2140 44036
rect 2180 43996 2189 44036
rect 2938 43996 2947 44036
rect 2987 43996 2996 44036
rect 3113 43996 3235 44036
rect 3284 43996 3293 44036
rect 4243 43996 4252 44036
rect 4292 43996 4492 44036
rect 4532 43996 4541 44036
rect 4627 43996 4636 44036
rect 4676 43996 5492 44036
rect 5827 43996 5836 44036
rect 5876 43996 7852 44036
rect 7892 43996 7901 44036
rect 8131 43996 8140 44036
rect 8180 43996 8227 44036
rect 8267 43996 8311 44036
rect 2956 43952 2996 43996
rect 5452 43952 5492 43996
rect 9964 43952 10004 44248
rect 11750 44228 11840 44248
rect 2956 43912 4684 43952
rect 4724 43912 4733 43952
rect 4780 43912 5356 43952
rect 5396 43912 5405 43952
rect 5452 43912 6316 43952
rect 6356 43912 6365 43952
rect 6412 43912 10004 43952
rect 4780 43868 4820 43912
rect 6412 43868 6452 43912
rect 4300 43828 4820 43868
rect 4919 43828 4928 43868
rect 4968 43828 5010 43868
rect 5050 43828 5092 43868
rect 5132 43828 5174 43868
rect 5214 43828 5256 43868
rect 5296 43828 5305 43868
rect 5635 43828 5644 43868
rect 5684 43828 6452 43868
rect 4300 43784 4340 43828
rect 4108 43744 4340 43784
rect 4387 43744 4396 43784
rect 4436 43744 5740 43784
rect 5780 43744 5789 43784
rect 6665 43744 6796 43784
rect 6836 43744 10828 43784
rect 10868 43744 10877 43784
rect 4108 43700 4148 43744
rect 6700 43700 6740 43744
rect 2345 43660 2467 43700
rect 2516 43660 2525 43700
rect 3475 43660 3484 43700
rect 3524 43660 3724 43700
rect 3764 43660 3773 43700
rect 4099 43660 4108 43700
rect 4148 43660 4157 43700
rect 6394 43660 6403 43700
rect 6443 43660 6691 43700
rect 6731 43660 6740 43700
rect 7651 43660 7660 43700
rect 7700 43660 8035 43700
rect 8075 43660 8515 43700
rect 8555 43660 8564 43700
rect 8873 43660 8995 43700
rect 9044 43660 9053 43700
rect 9257 43660 9379 43700
rect 9428 43660 9437 43700
rect 9004 43616 9044 43660
rect 0 43576 1268 43616
rect 1804 43576 1940 43616
rect 3427 43576 3436 43616
rect 3476 43576 4436 43616
rect 4675 43576 4684 43616
rect 4724 43576 4876 43616
rect 4916 43576 4925 43616
rect 5347 43576 5356 43616
rect 5396 43576 5684 43616
rect 5731 43576 5740 43616
rect 5780 43576 7084 43616
rect 7124 43576 7276 43616
rect 7316 43576 7372 43616
rect 7412 43576 7564 43616
rect 7604 43576 7660 43616
rect 7700 43576 8140 43616
rect 8180 43576 8189 43616
rect 9004 43576 9676 43616
rect 9716 43576 9725 43616
rect 0 43556 90 43576
rect 1228 43532 1268 43576
rect 1210 43523 1268 43532
rect 1210 43483 1219 43523
rect 1259 43483 1268 43523
rect 1673 43492 1795 43532
rect 1844 43492 1853 43532
rect 1210 43482 1268 43483
rect 1363 43408 1372 43448
rect 1412 43408 1708 43448
rect 1748 43408 1757 43448
rect 1900 43364 1940 43576
rect 3244 43492 4300 43532
rect 4340 43492 4349 43532
rect 3244 43448 3284 43492
rect 4396 43448 4436 43576
rect 5644 43448 5684 43576
rect 5827 43492 5836 43532
rect 5876 43492 10348 43532
rect 10388 43492 10397 43532
rect 2851 43408 2860 43448
rect 2900 43408 2909 43448
rect 3235 43408 3244 43448
rect 3284 43408 3293 43448
rect 3532 43408 3580 43448
rect 3620 43408 3629 43448
rect 3859 43408 3868 43448
rect 3908 43408 4204 43448
rect 4244 43408 4253 43448
rect 4387 43408 4396 43448
rect 4436 43408 4445 43448
rect 4579 43408 4588 43448
rect 4628 43408 5116 43448
rect 5156 43408 5165 43448
rect 5347 43408 5356 43448
rect 5396 43408 5405 43448
rect 5644 43408 6028 43448
rect 6068 43408 6316 43448
rect 6356 43408 6365 43448
rect 8105 43408 8236 43448
rect 8276 43408 8285 43448
rect 8515 43408 8524 43448
rect 8564 43408 9196 43448
rect 9236 43408 9245 43448
rect 9955 43408 9964 43448
rect 10004 43408 10013 43448
rect 10339 43408 10348 43448
rect 10388 43408 10540 43448
rect 10580 43408 10589 43448
rect 844 43324 1940 43364
rect 0 43280 90 43300
rect 844 43280 884 43324
rect 2860 43280 2900 43408
rect 3532 43364 3572 43408
rect 5356 43364 5396 43408
rect 3017 43324 3100 43364
rect 3140 43324 3148 43364
rect 3188 43324 3197 43364
rect 3427 43324 3436 43364
rect 3476 43324 3572 43364
rect 3715 43324 3724 43364
rect 3764 43324 4532 43364
rect 4627 43324 4636 43364
rect 4676 43324 4780 43364
rect 4820 43324 4829 43364
rect 5356 43324 8716 43364
rect 8756 43324 8765 43364
rect 4492 43280 4532 43324
rect 9964 43280 10004 43408
rect 10195 43324 10204 43364
rect 10244 43324 11060 43364
rect 11020 43280 11060 43324
rect 11750 43280 11840 43300
rect 0 43240 884 43280
rect 931 43240 940 43280
rect 980 43240 1996 43280
rect 2036 43240 2045 43280
rect 2860 43240 4340 43280
rect 4492 43240 7180 43280
rect 7220 43240 7229 43280
rect 7276 43240 10004 43280
rect 10579 43240 10588 43280
rect 10628 43240 10924 43280
rect 10964 43240 10973 43280
rect 11020 43240 11840 43280
rect 0 43220 90 43240
rect 4300 43196 4340 43240
rect 7276 43196 7316 43240
rect 11750 43220 11840 43240
rect 4300 43156 5836 43196
rect 5876 43156 5885 43196
rect 7075 43156 7084 43196
rect 7124 43156 7316 43196
rect 3679 43072 3688 43112
rect 3728 43072 3770 43112
rect 3810 43072 3852 43112
rect 3892 43072 3934 43112
rect 3974 43072 4016 43112
rect 4056 43072 4065 43112
rect 4483 43072 4492 43112
rect 4532 43072 9868 43112
rect 9908 43072 9917 43112
rect 1708 42988 7372 43028
rect 7412 42988 7421 43028
rect 0 42944 90 42964
rect 1708 42944 1748 42988
rect 0 42904 1324 42944
rect 1364 42904 1373 42944
rect 1699 42904 1708 42944
rect 1748 42904 1757 42944
rect 3401 42904 3484 42944
rect 3524 42904 3532 42944
rect 3572 42904 3581 42944
rect 4771 42904 4780 42944
rect 4820 42904 5204 42944
rect 5417 42904 5500 42944
rect 5540 42904 5548 42944
rect 5588 42904 5597 42944
rect 5923 42904 5932 42944
rect 5972 42904 8756 42944
rect 0 42884 90 42904
rect 5164 42860 5204 42904
rect 3532 42820 5108 42860
rect 5164 42820 7468 42860
rect 7508 42820 7517 42860
rect 3532 42776 3572 42820
rect 5068 42776 5108 42820
rect 1987 42736 1996 42776
rect 2036 42736 2764 42776
rect 2804 42736 2813 42776
rect 3523 42736 3532 42776
rect 3572 42736 3581 42776
rect 3715 42736 3724 42776
rect 3764 42736 4828 42776
rect 4868 42736 4877 42776
rect 5059 42736 5068 42776
rect 5108 42736 5117 42776
rect 5251 42736 5260 42776
rect 5300 42736 6988 42776
rect 7028 42736 7037 42776
rect 8227 42736 8236 42776
rect 8276 42736 8428 42776
rect 8468 42736 8477 42776
rect 8716 42692 8756 42904
rect 9833 42736 9964 42776
rect 10004 42736 10013 42776
rect 10217 42736 10348 42776
rect 10388 42736 10397 42776
rect 1193 42652 1315 42692
rect 1364 42652 1373 42692
rect 1507 42652 1516 42692
rect 1556 42652 2083 42692
rect 2123 42652 2132 42692
rect 2179 42652 2188 42692
rect 2228 42652 3874 42692
rect 3914 42652 3923 42692
rect 4012 42652 4354 42692
rect 4394 42652 4403 42692
rect 4579 42652 4588 42692
rect 4628 42652 5548 42692
rect 5588 42652 6796 42692
rect 6836 42652 6845 42692
rect 8707 42652 8716 42692
rect 8756 42652 9388 42692
rect 9428 42652 9437 42692
rect 0 42608 90 42628
rect 4012 42608 4052 42652
rect 0 42568 1804 42608
rect 1844 42568 1853 42608
rect 2371 42568 2380 42608
rect 2420 42568 4052 42608
rect 6211 42568 6220 42608
rect 6260 42568 6508 42608
rect 6548 42568 6700 42608
rect 6740 42568 6749 42608
rect 7075 42568 7084 42608
rect 7124 42568 7564 42608
rect 7604 42568 7613 42608
rect 7843 42568 7852 42608
rect 7892 42568 7948 42608
rect 7988 42568 8023 42608
rect 9004 42568 9196 42608
rect 9236 42568 9676 42608
rect 9716 42568 9725 42608
rect 10195 42568 10204 42608
rect 10244 42568 11692 42608
rect 11732 42568 11741 42608
rect 0 42548 90 42568
rect 9004 42524 9044 42568
rect 2275 42484 2284 42524
rect 2324 42484 2333 42524
rect 2995 42484 3004 42524
rect 3044 42484 3188 42524
rect 3322 42484 3331 42524
rect 3371 42484 3916 42524
rect 3956 42484 3965 42524
rect 4051 42484 4060 42524
rect 4100 42484 4484 42524
rect 4531 42484 4540 42524
rect 4580 42484 4588 42524
rect 4628 42484 4711 42524
rect 5722 42484 5731 42524
rect 5771 42484 5780 42524
rect 5914 42484 5923 42524
rect 5972 42484 6103 42524
rect 6298 42484 6307 42524
rect 6347 42484 6508 42524
rect 6548 42484 6557 42524
rect 6883 42484 6892 42524
rect 6932 42484 7276 42524
rect 7316 42484 7363 42524
rect 7403 42484 7447 42524
rect 7642 42484 7651 42524
rect 7691 42484 7700 42524
rect 8803 42484 8812 42524
rect 8852 42484 8995 42524
rect 9035 42484 9044 42524
rect 9466 42484 9475 42524
rect 9515 42484 9964 42524
rect 10004 42484 10013 42524
rect 10579 42484 10588 42524
rect 10628 42484 11212 42524
rect 11252 42484 11261 42524
rect 2284 42440 2324 42484
rect 3148 42440 3188 42484
rect 4444 42440 4484 42484
rect 5740 42440 5780 42484
rect 7660 42440 7700 42484
rect 2284 42400 2900 42440
rect 3148 42400 3244 42440
rect 3284 42400 3293 42440
rect 4444 42400 5588 42440
rect 5705 42400 5836 42440
rect 5876 42400 6220 42440
rect 6260 42400 7700 42440
rect 2860 42356 2900 42400
rect 5548 42356 5588 42400
rect 2860 42316 4780 42356
rect 4820 42316 4829 42356
rect 4919 42316 4928 42356
rect 4968 42316 5010 42356
rect 5050 42316 5092 42356
rect 5132 42316 5174 42356
rect 5214 42316 5256 42356
rect 5296 42316 5305 42356
rect 5548 42316 5972 42356
rect 0 42272 90 42292
rect 5932 42272 5972 42316
rect 11750 42272 11840 42292
rect 0 42232 652 42272
rect 692 42232 701 42272
rect 4675 42232 4684 42272
rect 4724 42232 5780 42272
rect 5932 42232 9388 42272
rect 9428 42232 9437 42272
rect 11683 42232 11692 42272
rect 11732 42232 11840 42272
rect 0 42212 90 42232
rect 2275 42148 2284 42188
rect 2324 42148 3148 42188
rect 3188 42148 3197 42188
rect 3436 42148 4492 42188
rect 4532 42148 4541 42188
rect 4723 42148 4732 42188
rect 4772 42148 5644 42188
rect 5684 42148 5693 42188
rect 3436 42104 3476 42148
rect 5740 42104 5780 42232
rect 11750 42212 11840 42232
rect 7939 42148 7948 42188
rect 7988 42148 7996 42188
rect 8036 42148 8119 42188
rect 8297 42148 8419 42188
rect 8468 42148 8477 42188
rect 8707 42148 8716 42188
rect 8756 42148 9628 42188
rect 9668 42148 9677 42188
rect 1027 42064 1036 42104
rect 1076 42064 1460 42104
rect 1699 42064 1708 42104
rect 1748 42064 3476 42104
rect 3523 42064 3532 42104
rect 3572 42064 3676 42104
rect 3716 42064 3725 42104
rect 4867 42064 4876 42104
rect 4916 42064 5548 42104
rect 5588 42064 5597 42104
rect 5644 42064 5932 42104
rect 5972 42064 7180 42104
rect 7220 42064 8716 42104
rect 8756 42064 8765 42104
rect 8969 42064 9004 42104
rect 9044 42064 9100 42104
rect 9140 42064 10060 42104
rect 10100 42064 10109 42104
rect 1420 42020 1460 42064
rect 5644 42020 5684 42064
rect 259 41980 268 42020
rect 308 41980 1315 42020
rect 1355 41980 1364 42020
rect 1420 41980 2083 42020
rect 2123 41980 2132 42020
rect 2842 41980 2851 42020
rect 2891 41980 2900 42020
rect 3139 41980 3148 42020
rect 3188 42011 3572 42020
rect 3188 41980 3523 42011
rect 0 41936 90 41956
rect 2860 41936 2900 41980
rect 3514 41971 3523 41980
rect 3563 41971 3572 42011
rect 3514 41970 3572 41971
rect 3994 42011 4052 42020
rect 3994 41971 4003 42011
rect 4043 41971 4052 42011
rect 4771 41980 4780 42020
rect 4820 42011 5204 42020
rect 4820 41980 5155 42011
rect 3994 41970 4052 41971
rect 5146 41971 5155 41980
rect 5195 41971 5204 42011
rect 5635 41980 5644 42020
rect 5684 41980 5693 42020
rect 6307 41980 6316 42020
rect 6356 41980 6412 42020
rect 6452 41980 6487 42020
rect 7660 42011 9292 42020
rect 5146 41970 5204 41971
rect 7700 41980 9292 42011
rect 9332 41980 9908 42020
rect 9955 41980 9964 42020
rect 10004 41980 10060 42020
rect 10100 41980 11404 42020
rect 11444 41980 11453 42020
rect 0 41896 2900 41936
rect 0 41876 90 41896
rect 4012 41852 4052 41970
rect 7660 41962 7700 41971
rect 9868 41936 9908 41980
rect 4147 41896 4156 41936
rect 4196 41896 4436 41936
rect 4483 41896 4492 41936
rect 4532 41896 4588 41936
rect 4628 41896 4663 41936
rect 5299 41896 5308 41936
rect 5348 41896 5452 41936
rect 5492 41896 5501 41936
rect 7747 41896 7756 41936
rect 7796 41896 8236 41936
rect 8276 41896 8285 41936
rect 9100 41896 9292 41936
rect 9332 41896 9341 41936
rect 9859 41896 9868 41936
rect 9908 41896 9917 41936
rect 10217 41896 10348 41936
rect 10388 41896 10397 41936
rect 10579 41896 10588 41936
rect 10628 41896 11116 41936
rect 11156 41896 11165 41936
rect 2921 41812 3052 41852
rect 3092 41812 3101 41852
rect 3148 41812 4052 41852
rect 4396 41852 4436 41896
rect 9100 41852 9140 41896
rect 4396 41812 7604 41852
rect 7721 41812 7852 41852
rect 7892 41812 7901 41852
rect 7948 41812 9044 41852
rect 9091 41812 9100 41852
rect 9140 41812 9149 41852
rect 9523 41812 9532 41852
rect 9572 41812 11692 41852
rect 11732 41812 11741 41852
rect 3148 41768 3188 41812
rect 1795 41728 1804 41768
rect 1844 41728 3188 41768
rect 7564 41768 7604 41812
rect 7948 41768 7988 41812
rect 7564 41728 7988 41768
rect 9004 41768 9044 41812
rect 9004 41728 9196 41768
rect 9236 41728 9245 41768
rect 0 41600 90 41620
rect 0 41560 2188 41600
rect 2228 41560 2237 41600
rect 3679 41560 3688 41600
rect 3728 41560 3770 41600
rect 3810 41560 3852 41600
rect 3892 41560 3934 41600
rect 3974 41560 4016 41600
rect 4056 41560 4065 41600
rect 0 41540 90 41560
rect 1036 41308 1516 41348
rect 1556 41308 1565 41348
rect 1996 41308 5836 41348
rect 5876 41308 6316 41348
rect 6356 41308 6452 41348
rect 0 41264 90 41284
rect 1036 41264 1076 41308
rect 0 41224 1076 41264
rect 1132 41224 1228 41264
rect 1268 41224 1277 41264
rect 0 41204 90 41224
rect 1132 41180 1172 41224
rect 1996 41180 2036 41308
rect 3139 41224 3148 41264
rect 3188 41224 3340 41264
rect 3380 41224 3389 41264
rect 5356 41224 6124 41264
rect 6164 41224 6173 41264
rect 451 41140 460 41180
rect 500 41140 1172 41180
rect 1411 41140 1420 41180
rect 1460 41140 1612 41180
rect 1652 41140 2036 41180
rect 2860 41180 2900 41189
rect 5072 41180 5112 41189
rect 3427 41140 3436 41180
rect 3476 41140 3820 41180
rect 3860 41140 3869 41180
rect 5068 41140 5072 41180
rect 2860 41096 2900 41140
rect 5068 41131 5112 41140
rect 5068 41096 5108 41131
rect 2860 41056 3532 41096
rect 3572 41056 5108 41096
rect 1459 40972 1468 41012
rect 1508 40972 1612 41012
rect 1652 40972 1661 41012
rect 2921 40972 3052 41012
rect 3092 40972 3101 41012
rect 3322 40972 3331 41012
rect 3371 40972 3619 41012
rect 3659 40972 3668 41012
rect 4675 40972 4684 41012
rect 4724 40972 5260 41012
rect 5300 40972 5309 41012
rect 0 40928 90 40948
rect 3628 40928 3668 40972
rect 5356 40928 5396 41224
rect 6412 41180 6452 41308
rect 11750 41264 11840 41284
rect 9833 41224 9964 41264
rect 10004 41224 10013 41264
rect 10339 41224 10348 41264
rect 10388 41224 10636 41264
rect 10676 41224 10685 41264
rect 11683 41224 11692 41264
rect 11732 41224 11840 41264
rect 11750 41204 11840 41224
rect 7660 41180 7700 41189
rect 9292 41180 9332 41189
rect 0 40888 1324 40928
rect 1364 40888 1373 40928
rect 3628 40888 5396 40928
rect 5548 41140 5602 41180
rect 5642 41140 5651 41180
rect 6403 41140 6412 41180
rect 6452 41140 6461 41180
rect 7529 41140 7660 41180
rect 7700 41140 7709 41180
rect 7756 41140 8044 41180
rect 8084 41140 8093 41180
rect 9161 41140 9292 41180
rect 9332 41140 9341 41180
rect 0 40868 90 40888
rect 4919 40804 4928 40844
rect 4968 40804 5010 40844
rect 5050 40804 5092 40844
rect 5132 40804 5174 40844
rect 5214 40804 5256 40844
rect 5296 40804 5305 40844
rect 5548 40676 5588 41140
rect 7660 41131 7700 41140
rect 5657 40972 5740 41012
rect 5780 40972 5788 41012
rect 5828 40972 5837 41012
rect 6202 40972 6211 41012
rect 6251 40972 6892 41012
rect 6932 40972 6941 41012
rect 7756 40928 7796 41140
rect 9292 41131 9332 41140
rect 10195 41056 10204 41096
rect 10244 41056 11020 41096
rect 11060 41056 11069 41096
rect 7843 40972 7852 41012
rect 7892 40972 7901 41012
rect 9353 40972 9484 41012
rect 9524 40972 9533 41012
rect 9754 40972 9763 41012
rect 9803 40972 10060 41012
rect 10100 40972 10109 41012
rect 10579 40972 10588 41012
rect 10628 40972 11500 41012
rect 11540 40972 11549 41012
rect 6115 40888 6124 40928
rect 6164 40888 7796 40928
rect 7852 40676 7892 40972
rect 5539 40636 5548 40676
rect 5588 40636 5597 40676
rect 5971 40636 5980 40676
rect 6020 40636 7084 40676
rect 7124 40636 7133 40676
rect 7852 40636 9044 40676
rect 9571 40636 9580 40676
rect 9620 40636 9629 40676
rect 0 40592 90 40612
rect 0 40552 1804 40592
rect 1844 40552 1853 40592
rect 3523 40552 3532 40592
rect 3572 40552 3860 40592
rect 0 40532 90 40552
rect 3820 40508 3860 40552
rect 4876 40552 6068 40592
rect 7555 40552 7564 40592
rect 7604 40552 7892 40592
rect 1193 40468 1315 40508
rect 1364 40468 1373 40508
rect 2083 40468 2092 40508
rect 2132 40468 2380 40508
rect 2420 40468 2429 40508
rect 2860 40499 3380 40508
rect 2860 40468 3340 40499
rect 2860 40340 2900 40468
rect 3802 40468 3811 40508
rect 3851 40468 3860 40508
rect 3907 40468 3916 40508
rect 3956 40468 4108 40508
rect 4148 40468 4157 40508
rect 4265 40468 4300 40508
rect 4340 40468 4396 40508
rect 4436 40468 4445 40508
rect 4876 40499 4916 40552
rect 3340 40450 3380 40459
rect 5225 40468 5356 40508
rect 5396 40468 5405 40508
rect 4876 40450 4916 40459
rect 5356 40450 5396 40459
rect 6028 40424 6068 40552
rect 7852 40508 7892 40552
rect 9004 40508 9044 40636
rect 9580 40508 9620 40636
rect 6115 40468 6124 40508
rect 6164 40468 6295 40508
rect 7372 40499 7412 40508
rect 7834 40468 7843 40508
rect 7883 40468 7892 40508
rect 7939 40468 7948 40508
rect 7988 40468 8119 40508
rect 8323 40468 8332 40508
rect 8372 40468 8620 40508
rect 8660 40468 8669 40508
rect 8777 40468 8908 40508
rect 8948 40468 8957 40508
rect 9004 40499 9428 40508
rect 9004 40468 9388 40499
rect 7372 40424 7412 40459
rect 8908 40450 8948 40459
rect 9580 40499 10292 40508
rect 9580 40468 10243 40499
rect 9388 40450 9428 40459
rect 10234 40459 10243 40468
rect 10283 40459 10292 40499
rect 10234 40458 10292 40459
rect 4291 40384 4300 40424
rect 4340 40384 4396 40424
rect 4436 40384 4471 40424
rect 5705 40384 5740 40424
rect 5780 40384 5836 40424
rect 5876 40384 5885 40424
rect 6028 40384 6260 40424
rect 7372 40384 7660 40424
rect 7700 40384 8372 40424
rect 8419 40384 8428 40424
rect 8468 40384 8524 40424
rect 8564 40384 8599 40424
rect 9833 40384 9964 40424
rect 10004 40384 10013 40424
rect 10339 40384 10348 40424
rect 10388 40384 10396 40424
rect 10436 40384 10519 40424
rect 6220 40340 6260 40384
rect 8332 40340 8372 40384
rect 1123 40300 1132 40340
rect 1172 40300 1516 40340
rect 1556 40300 1565 40340
rect 2563 40300 2572 40340
rect 2612 40300 2900 40340
rect 3427 40300 3436 40340
rect 3476 40300 6124 40340
rect 6164 40300 6173 40340
rect 6220 40300 8276 40340
rect 8323 40300 8332 40340
rect 8372 40300 8381 40340
rect 0 40256 90 40276
rect 8236 40256 8276 40300
rect 11750 40256 11840 40276
rect 0 40216 1036 40256
rect 1076 40216 1085 40256
rect 4291 40216 4300 40256
rect 4340 40216 7948 40256
rect 7988 40216 7997 40256
rect 8236 40216 8908 40256
rect 8948 40216 8957 40256
rect 10915 40216 10924 40256
rect 10964 40216 11840 40256
rect 0 40196 90 40216
rect 11750 40196 11840 40216
rect 3679 40048 3688 40088
rect 3728 40048 3770 40088
rect 3810 40048 3852 40088
rect 3892 40048 3934 40088
rect 3974 40048 4016 40088
rect 4056 40048 4065 40088
rect 0 39920 90 39940
rect 0 39880 268 39920
rect 308 39880 317 39920
rect 4003 39880 4012 39920
rect 4052 39880 5300 39920
rect 0 39860 90 39880
rect 1507 39796 1516 39836
rect 1556 39796 5204 39836
rect 5164 39752 5204 39796
rect 3715 39712 3724 39752
rect 3764 39712 4108 39752
rect 4148 39712 4157 39752
rect 5155 39712 5164 39752
rect 5204 39712 5213 39752
rect 2668 39668 2708 39677
rect 4300 39668 4340 39677
rect 5260 39668 5300 39880
rect 5788 39880 11692 39920
rect 11732 39880 11741 39920
rect 5788 39752 5828 39880
rect 6259 39796 6268 39836
rect 6308 39796 8044 39836
rect 8084 39796 8093 39836
rect 5683 39712 5692 39752
rect 5732 39712 5828 39752
rect 5897 39712 6028 39752
rect 6068 39712 6077 39752
rect 6595 39712 6604 39752
rect 6644 39712 6653 39752
rect 8297 39712 8428 39752
rect 8468 39712 8477 39752
rect 9737 39712 9868 39752
rect 9908 39712 9917 39752
rect 1289 39628 1420 39668
rect 1460 39628 1469 39668
rect 2537 39628 2668 39668
rect 2708 39628 2717 39668
rect 3043 39628 3052 39668
rect 3092 39628 3235 39668
rect 3275 39628 3284 39668
rect 3331 39628 3340 39668
rect 3380 39628 3389 39668
rect 3811 39628 3820 39668
rect 3860 39628 4052 39668
rect 4169 39628 4300 39668
rect 4340 39628 4349 39668
rect 4675 39628 4684 39668
rect 4724 39628 4788 39668
rect 4828 39628 4855 39668
rect 5260 39628 5536 39668
rect 5576 39628 6124 39668
rect 6164 39628 6173 39668
rect 2668 39619 2708 39628
rect 0 39584 90 39604
rect 3340 39584 3380 39628
rect 0 39544 844 39584
rect 884 39544 893 39584
rect 2947 39544 2956 39584
rect 2996 39544 3380 39584
rect 0 39524 90 39544
rect 4012 39500 4052 39628
rect 4300 39619 4340 39628
rect 4483 39544 4492 39584
rect 4532 39544 5404 39584
rect 5444 39544 5453 39584
rect 2851 39460 2860 39500
rect 2900 39460 3031 39500
rect 4012 39460 4396 39500
rect 4436 39460 4445 39500
rect 4771 39460 4780 39500
rect 4820 39460 4972 39500
rect 5012 39460 5021 39500
rect 6355 39460 6364 39500
rect 6404 39460 6508 39500
rect 6548 39460 6557 39500
rect 6604 39416 6644 39712
rect 9004 39668 9044 39677
rect 7787 39628 7852 39668
rect 7892 39628 7918 39668
rect 7958 39628 7967 39668
rect 8032 39628 8041 39668
rect 8081 39628 8140 39668
rect 8180 39628 8221 39668
rect 8489 39628 8524 39668
rect 8564 39628 8620 39668
rect 8660 39628 8669 39668
rect 8899 39628 8908 39668
rect 8948 39628 9004 39668
rect 9044 39628 9079 39668
rect 9475 39628 9484 39668
rect 9532 39628 9655 39668
rect 10186 39628 10195 39668
rect 10235 39628 10244 39668
rect 9004 39619 9044 39628
rect 10204 39584 10244 39628
rect 9676 39544 10244 39584
rect 9676 39500 9716 39544
rect 6761 39460 6883 39500
rect 6932 39460 6941 39500
rect 6988 39460 7075 39500
rect 7115 39460 7124 39500
rect 7267 39460 7276 39500
rect 7316 39460 7363 39500
rect 7403 39460 7447 39500
rect 9667 39460 9676 39500
rect 9716 39460 9725 39500
rect 10099 39460 10108 39500
rect 10148 39460 10156 39500
rect 10196 39460 10279 39500
rect 10387 39460 10396 39500
rect 10436 39460 10444 39500
rect 10484 39460 10567 39500
rect 1420 39376 3436 39416
rect 3476 39376 3485 39416
rect 4204 39376 6644 39416
rect 0 39248 90 39268
rect 0 39208 1324 39248
rect 1364 39208 1373 39248
rect 0 39188 90 39208
rect 1420 38996 1460 39376
rect 2563 39292 2572 39332
rect 2612 39292 3820 39332
rect 3860 39292 3869 39332
rect 4204 39248 4244 39376
rect 6988 39332 7028 39460
rect 4291 39292 4300 39332
rect 4340 39292 4780 39332
rect 4820 39292 4829 39332
rect 4919 39292 4928 39332
rect 4968 39292 5010 39332
rect 5050 39292 5092 39332
rect 5132 39292 5174 39332
rect 5214 39292 5256 39332
rect 5296 39292 5305 39332
rect 5347 39292 5356 39332
rect 5396 39292 5492 39332
rect 5539 39292 5548 39332
rect 5588 39292 7028 39332
rect 1516 39208 4244 39248
rect 1411 38956 1420 38996
rect 1460 38956 1469 38996
rect 0 38912 90 38932
rect 1516 38912 1556 39208
rect 5452 39164 5492 39292
rect 11750 39248 11840 39268
rect 7939 39208 7948 39248
rect 7988 39208 8372 39248
rect 11203 39208 11212 39248
rect 11252 39208 11840 39248
rect 3187 39124 3196 39164
rect 3236 39124 5396 39164
rect 5443 39124 5452 39164
rect 5492 39124 5501 39164
rect 5836 39124 6796 39164
rect 6836 39124 6845 39164
rect 5356 39080 5396 39124
rect 5836 39080 5876 39124
rect 2851 39040 2860 39080
rect 2900 39040 3148 39080
rect 3188 39040 3197 39080
rect 3811 39040 3820 39080
rect 3860 39040 5300 39080
rect 5356 39040 5876 39080
rect 5993 39040 6124 39080
rect 6164 39040 7468 39080
rect 7508 39040 7517 39080
rect 1795 38956 1804 38996
rect 1844 38956 2668 38996
rect 2708 38956 2717 38996
rect 2921 38987 3052 38996
rect 2921 38956 3043 38987
rect 3092 38956 3101 38996
rect 3401 38987 3532 38996
rect 3401 38956 3523 38987
rect 3572 38956 3581 38996
rect 3881 38956 4012 38996
rect 4052 38956 4300 38996
rect 4340 38956 4349 38996
rect 5260 38987 5300 39040
rect 6124 38996 6164 39040
rect 8332 38996 8372 39208
rect 11750 39188 11840 39208
rect 9955 39124 9964 39164
rect 10004 39124 10196 39164
rect 10156 38996 10196 39124
rect 2668 38938 2708 38947
rect 3034 38947 3043 38956
rect 3083 38947 3092 38956
rect 3034 38946 3092 38947
rect 3514 38947 3523 38956
rect 3563 38947 3572 38956
rect 3514 38946 3572 38947
rect 5260 38938 5300 38947
rect 5356 38987 5684 38996
rect 5356 38956 5635 38987
rect 0 38872 1556 38912
rect 3619 38872 3628 38912
rect 3668 38872 3676 38912
rect 3716 38872 3799 38912
rect 4195 38872 4204 38912
rect 4244 38872 5204 38912
rect 0 38852 90 38872
rect 5164 38828 5204 38872
rect 5356 38828 5396 38956
rect 5626 38947 5635 38956
rect 5675 38947 5684 38987
rect 6115 38956 6124 38996
rect 6164 38956 6173 38996
rect 7372 38987 7700 38996
rect 5626 38946 5684 38947
rect 7412 38956 7700 38987
rect 8214 38956 8223 38996
rect 8263 38956 8276 38996
rect 8323 38956 8332 38996
rect 8372 38956 8381 38996
rect 8585 38956 8716 38996
rect 8756 38956 8765 38996
rect 8899 38956 8908 38996
rect 8948 38987 9332 38996
rect 8948 38956 9292 38987
rect 7372 38938 7412 38947
rect 7660 38912 7700 38956
rect 8236 38912 8276 38956
rect 9641 38956 9772 38996
rect 9812 38956 9821 38996
rect 10138 38987 10196 38996
rect 9292 38938 9332 38947
rect 9772 38938 9812 38947
rect 10138 38947 10147 38987
rect 10187 38947 10196 38987
rect 10138 38946 10196 38947
rect 5779 38872 5788 38912
rect 5828 38872 5836 38912
rect 5876 38872 5959 38912
rect 7651 38872 7660 38912
rect 7700 38872 7756 38912
rect 7796 38872 7831 38912
rect 8236 38872 8428 38912
rect 8468 38872 8477 38912
rect 8524 38872 8812 38912
rect 8852 38872 8861 38912
rect 10291 38872 10300 38912
rect 10340 38872 10444 38912
rect 10484 38872 10493 38912
rect 8524 38828 8564 38872
rect 5164 38788 5396 38828
rect 8515 38788 8524 38828
rect 8564 38788 8573 38828
rect 7433 38704 7564 38744
rect 7604 38704 7613 38744
rect 7987 38704 7996 38744
rect 8036 38704 8620 38744
rect 8660 38704 9292 38744
rect 9332 38704 9341 38744
rect 2860 38620 6028 38660
rect 6068 38620 6077 38660
rect 0 38576 90 38596
rect 2860 38576 2900 38620
rect 0 38536 2900 38576
rect 3679 38536 3688 38576
rect 3728 38536 3770 38576
rect 3810 38536 3852 38576
rect 3892 38536 3934 38576
rect 3974 38536 4016 38576
rect 4056 38536 4065 38576
rect 5347 38536 5356 38576
rect 5396 38536 8140 38576
rect 8180 38536 8716 38576
rect 8756 38536 8765 38576
rect 0 38516 90 38536
rect 2467 38452 2476 38492
rect 2516 38452 6124 38492
rect 6164 38452 6173 38492
rect 8297 38368 8428 38408
rect 8468 38368 8477 38408
rect 9763 38368 9772 38408
rect 9812 38368 10252 38408
rect 10292 38368 10301 38408
rect 2227 38284 2236 38324
rect 2276 38284 5356 38324
rect 5396 38284 5405 38324
rect 5731 38284 5740 38324
rect 5780 38284 7028 38324
rect 0 38240 90 38260
rect 0 38200 1516 38240
rect 1556 38200 1565 38240
rect 1987 38200 1996 38240
rect 2036 38200 2045 38240
rect 3628 38200 5492 38240
rect 0 38180 90 38200
rect 1996 38156 2036 38200
rect 3628 38156 3668 38200
rect 5452 38156 5492 38200
rect 6988 38156 7028 38284
rect 11750 38240 11840 38260
rect 9283 38200 9292 38240
rect 9332 38200 10100 38240
rect 10435 38200 10444 38240
rect 10484 38200 10732 38240
rect 10772 38200 10964 38240
rect 11011 38200 11020 38240
rect 11060 38200 11840 38240
rect 8236 38156 8276 38165
rect 10060 38156 10100 38200
rect 10924 38156 10964 38200
rect 11750 38180 11840 38200
rect 835 38116 844 38156
rect 884 38116 1315 38156
rect 1355 38116 1364 38156
rect 1411 38116 1420 38156
rect 1460 38116 2036 38156
rect 2345 38116 2380 38156
rect 2420 38116 2476 38156
rect 2516 38116 2525 38156
rect 4169 38116 4204 38156
rect 4244 38116 4300 38156
rect 4340 38116 4349 38156
rect 5731 38116 5740 38156
rect 5780 38116 5875 38156
rect 5915 38116 5924 38156
rect 6019 38116 6028 38156
rect 6068 38116 6370 38156
rect 6410 38116 6419 38156
rect 6979 38116 6988 38156
rect 7028 38116 7084 38156
rect 7124 38116 7188 38156
rect 8276 38116 8620 38156
rect 8660 38116 8669 38156
rect 8803 38116 8812 38156
rect 8852 38116 9868 38156
rect 9908 38116 9917 38156
rect 10915 38116 10924 38156
rect 10964 38116 10973 38156
rect 3628 38107 3668 38116
rect 5452 38072 5492 38116
rect 8236 38107 8276 38116
rect 10060 38107 10100 38116
rect 1481 38032 1603 38072
rect 1652 38032 1661 38072
rect 3724 38032 4148 38072
rect 5452 38032 5780 38072
rect 5827 38032 5836 38072
rect 5876 38032 6556 38072
rect 6596 38032 6605 38072
rect 0 37904 90 37924
rect 3724 37904 3764 38032
rect 3811 37948 3820 37988
rect 3860 37948 3869 37988
rect 0 37864 1996 37904
rect 2036 37864 2045 37904
rect 2371 37864 2380 37904
rect 2420 37864 3764 37904
rect 0 37844 90 37864
rect 739 37696 748 37736
rect 788 37696 2900 37736
rect 2860 37652 2900 37696
rect 1219 37612 1228 37652
rect 1268 37612 2516 37652
rect 2860 37612 3571 37652
rect 3611 37612 3620 37652
rect 0 37568 90 37588
rect 0 37528 364 37568
rect 404 37528 413 37568
rect 1027 37528 1036 37568
rect 1076 37528 2036 37568
rect 0 37508 90 37528
rect 1996 37484 2036 37528
rect 2476 37484 2516 37612
rect 3820 37568 3860 37948
rect 3091 37528 3100 37568
rect 3140 37528 3284 37568
rect 3820 37528 4052 37568
rect 3244 37484 3284 37528
rect 4012 37484 4052 37528
rect 4108 37484 4148 38032
rect 5635 37948 5644 37988
rect 5684 37948 5693 37988
rect 4919 37780 4928 37820
rect 4968 37780 5010 37820
rect 5050 37780 5092 37820
rect 5132 37780 5174 37820
rect 5214 37780 5256 37820
rect 5296 37780 5305 37820
rect 5644 37484 5684 37948
rect 5740 37904 5780 38032
rect 6067 37948 6076 37988
rect 6116 37948 6316 37988
rect 6356 37948 6365 37988
rect 5740 37864 9004 37904
rect 9044 37864 9053 37904
rect 5731 37612 5740 37652
rect 5780 37612 5911 37652
rect 6019 37612 6028 37652
rect 6068 37612 6892 37652
rect 6932 37612 8227 37652
rect 8267 37612 8276 37652
rect 7372 37528 7660 37568
rect 7700 37528 7709 37568
rect 1193 37444 1315 37484
rect 1364 37444 1373 37484
rect 1978 37475 2036 37484
rect 1978 37435 1987 37475
rect 2027 37435 2036 37475
rect 2131 37444 2140 37484
rect 2180 37444 2284 37484
rect 2324 37444 2333 37484
rect 2458 37475 2516 37484
rect 1978 37434 2036 37435
rect 2458 37435 2467 37475
rect 2507 37435 2516 37475
rect 2611 37444 2620 37484
rect 2660 37444 2764 37484
rect 2804 37444 2813 37484
rect 2938 37475 2956 37484
rect 2458 37434 2516 37435
rect 2938 37435 2947 37475
rect 2996 37444 3127 37484
rect 3235 37444 3244 37484
rect 3284 37444 3293 37484
rect 3757 37444 3766 37484
rect 3806 37444 3860 37484
rect 3994 37444 4003 37484
rect 4043 37444 4052 37484
rect 4099 37444 4108 37484
rect 4148 37444 4157 37484
rect 4483 37444 4492 37484
rect 4532 37444 4541 37484
rect 4937 37444 5068 37484
rect 5108 37444 5117 37484
rect 5548 37475 5684 37484
rect 2987 37435 2996 37444
rect 2938 37434 2996 37435
rect 3820 37400 3860 37444
rect 3820 37360 4300 37400
rect 4340 37360 4349 37400
rect 4492 37316 4532 37444
rect 5068 37426 5108 37435
rect 5588 37444 5684 37475
rect 5993 37444 6124 37484
rect 6164 37444 6173 37484
rect 7372 37475 7412 37528
rect 5548 37426 5588 37435
rect 7625 37475 7756 37484
rect 7625 37444 7747 37475
rect 7796 37444 7805 37484
rect 7891 37444 7900 37484
rect 7940 37444 7948 37484
rect 7988 37444 8071 37484
rect 8995 37444 9004 37484
rect 9044 37475 9175 37484
rect 9044 37444 9096 37475
rect 7372 37426 7412 37435
rect 7738 37435 7747 37444
rect 7787 37435 7796 37444
rect 7738 37434 7796 37435
rect 9136 37444 9175 37475
rect 9859 37444 9868 37484
rect 9908 37444 10348 37484
rect 10388 37444 10397 37484
rect 9096 37426 9136 37435
rect 4579 37360 4588 37400
rect 4628 37360 4780 37400
rect 4820 37360 4829 37400
rect 8515 37360 8524 37400
rect 8564 37360 8812 37400
rect 8852 37360 8861 37400
rect 8524 37316 8564 37360
rect 172 37276 4204 37316
rect 4244 37276 4253 37316
rect 4492 37276 5644 37316
rect 5684 37276 5693 37316
rect 7075 37276 7084 37316
rect 7124 37276 8564 37316
rect 8755 37276 8764 37316
rect 8804 37276 9580 37316
rect 9620 37276 9629 37316
rect 0 37232 90 37252
rect 172 37232 212 37276
rect 11750 37232 11840 37252
rect 0 37192 212 37232
rect 1385 37192 1516 37232
rect 1556 37192 1565 37232
rect 7555 37192 7564 37232
rect 7604 37192 8716 37232
rect 8756 37192 8765 37232
rect 8899 37192 8908 37232
rect 8948 37192 8957 37232
rect 11107 37192 11116 37232
rect 11156 37192 11840 37232
rect 0 37172 90 37192
rect 8908 37148 8948 37192
rect 11750 37172 11840 37192
rect 5539 37108 5548 37148
rect 5588 37108 8948 37148
rect 3679 37024 3688 37064
rect 3728 37024 3770 37064
rect 3810 37024 3852 37064
rect 3892 37024 3934 37064
rect 3974 37024 4016 37064
rect 4056 37024 4065 37064
rect 8803 37024 8812 37064
rect 8852 37024 10060 37064
rect 10100 37024 10109 37064
rect 2275 36940 2284 36980
rect 2324 36940 8524 36980
rect 8564 36940 8573 36980
rect 0 36896 90 36916
rect 0 36856 1324 36896
rect 1364 36856 1373 36896
rect 4867 36856 4876 36896
rect 4916 36856 7508 36896
rect 0 36836 90 36856
rect 1516 36772 3532 36812
rect 3572 36772 3581 36812
rect 3628 36772 4108 36812
rect 4148 36772 4157 36812
rect 5260 36772 5548 36812
rect 5588 36772 5597 36812
rect 5731 36772 5740 36812
rect 5780 36772 5789 36812
rect 451 36604 460 36644
rect 500 36604 844 36644
rect 884 36604 1324 36644
rect 1364 36604 1373 36644
rect 0 36560 90 36580
rect 1516 36560 1556 36772
rect 3628 36728 3668 36772
rect 5260 36728 5300 36772
rect 5740 36728 5780 36772
rect 2860 36688 3532 36728
rect 3572 36688 3668 36728
rect 4204 36688 4876 36728
rect 4916 36688 4925 36728
rect 5164 36688 5300 36728
rect 5513 36688 5644 36728
rect 5684 36688 5693 36728
rect 5740 36688 7412 36728
rect 2572 36644 2612 36653
rect 2860 36644 2900 36688
rect 4108 36644 4148 36653
rect 4204 36644 4244 36688
rect 5164 36644 5204 36688
rect 6220 36644 6260 36688
rect 7372 36644 7412 36688
rect 7468 36644 7508 36856
rect 7756 36728 7796 36940
rect 7747 36688 7756 36728
rect 7796 36688 7805 36728
rect 9833 36688 9964 36728
rect 10004 36688 10013 36728
rect 10339 36688 10348 36728
rect 10388 36688 11308 36728
rect 11348 36688 11357 36728
rect 8332 36644 8372 36653
rect 2441 36604 2572 36644
rect 2612 36604 2621 36644
rect 2668 36604 2900 36644
rect 3034 36604 3043 36644
rect 3083 36604 3092 36644
rect 3139 36604 3148 36644
rect 3188 36604 3197 36644
rect 3619 36604 3628 36644
rect 3668 36604 4052 36644
rect 2572 36595 2612 36604
rect 0 36520 1556 36560
rect 0 36500 90 36520
rect 2668 36476 2708 36604
rect 3052 36560 3092 36604
rect 2755 36520 2764 36560
rect 2804 36520 3092 36560
rect 2467 36436 2476 36476
rect 2516 36436 2708 36476
rect 3148 36476 3188 36604
rect 3148 36436 3532 36476
rect 3572 36436 3581 36476
rect 4012 36392 4052 36604
rect 4148 36604 4204 36644
rect 4244 36604 4279 36644
rect 4579 36604 4588 36644
rect 4636 36604 4759 36644
rect 5146 36604 5155 36644
rect 5195 36604 5204 36644
rect 5251 36604 5260 36644
rect 5300 36604 5548 36644
rect 5588 36604 5597 36644
rect 5731 36604 5740 36644
rect 5780 36604 5911 36644
rect 6730 36604 6739 36644
rect 6779 36604 7124 36644
rect 7258 36604 7267 36644
rect 7307 36604 7316 36644
rect 7363 36604 7372 36644
rect 7412 36604 7421 36644
rect 7468 36604 7852 36644
rect 7892 36604 7901 36644
rect 8131 36604 8140 36644
rect 8180 36604 8332 36644
rect 4108 36595 4148 36604
rect 6220 36595 6260 36604
rect 7084 36560 7124 36604
rect 7276 36560 7316 36604
rect 8332 36595 8372 36604
rect 8620 36604 8820 36644
rect 8860 36604 8869 36644
rect 9004 36604 9235 36644
rect 9275 36604 9284 36644
rect 7084 36520 7180 36560
rect 7220 36520 7229 36560
rect 7276 36520 7372 36560
rect 7412 36520 7421 36560
rect 4291 36436 4300 36476
rect 4340 36436 4780 36476
rect 4820 36436 4829 36476
rect 6883 36436 6892 36476
rect 6932 36436 7756 36476
rect 7796 36436 7805 36476
rect 4012 36352 4396 36392
rect 4436 36352 4445 36392
rect 4919 36268 4928 36308
rect 4968 36268 5010 36308
rect 5050 36268 5092 36308
rect 5132 36268 5174 36308
rect 5214 36268 5256 36308
rect 5296 36268 5305 36308
rect 0 36224 90 36244
rect 0 36184 3052 36224
rect 3092 36184 3101 36224
rect 4396 36184 6220 36224
rect 6260 36184 6892 36224
rect 6932 36184 6941 36224
rect 0 36164 90 36184
rect 4396 36140 4436 36184
rect 8620 36140 8660 36604
rect 9004 36476 9044 36604
rect 10195 36520 10204 36560
rect 10244 36520 11020 36560
rect 11060 36520 11069 36560
rect 8995 36436 9004 36476
rect 9044 36436 9053 36476
rect 9427 36436 9436 36476
rect 9476 36436 9484 36476
rect 9524 36436 9607 36476
rect 10579 36436 10588 36476
rect 10628 36436 11116 36476
rect 11156 36436 11165 36476
rect 11750 36224 11840 36244
rect 11491 36184 11500 36224
rect 11540 36184 11840 36224
rect 11750 36164 11840 36184
rect 1843 36100 1852 36140
rect 1892 36100 4204 36140
rect 4244 36100 4253 36140
rect 4378 36100 4387 36140
rect 4427 36100 4436 36140
rect 4780 36100 5644 36140
rect 5684 36100 5693 36140
rect 5932 36100 6836 36140
rect 8611 36100 8620 36140
rect 8660 36100 8669 36140
rect 10051 36100 10060 36140
rect 10100 36100 10109 36140
rect 10522 36100 10531 36140
rect 10571 36100 10828 36140
rect 10868 36100 10877 36140
rect 1363 36016 1372 36056
rect 1412 36016 1996 36056
rect 2036 36016 2045 36056
rect 2563 36016 2572 36056
rect 2612 36016 3572 36056
rect 3532 35972 3572 36016
rect 4780 35972 4820 36100
rect 5164 36016 5740 36056
rect 5780 36016 5789 36056
rect 5164 35972 5204 36016
rect 5932 35972 5972 36100
rect 6796 36056 6836 36100
rect 10060 36056 10100 36100
rect 6124 36016 6740 36056
rect 6796 36016 9484 36056
rect 9524 36016 9533 36056
rect 10060 36016 10292 36056
rect 6124 35972 6164 36016
rect 6700 35972 6740 36016
rect 10252 35972 10292 36016
rect 451 35932 460 35972
rect 500 35963 1268 35972
rect 500 35932 1219 35963
rect 1210 35923 1219 35932
rect 1259 35923 1268 35963
rect 1315 35932 1324 35972
rect 1364 35963 1748 35972
rect 1364 35932 1699 35963
rect 1210 35922 1268 35923
rect 1690 35923 1699 35932
rect 1739 35923 1748 35963
rect 1690 35922 1748 35923
rect 1804 35963 2228 35972
rect 1804 35932 2179 35963
rect 0 35888 90 35908
rect 0 35848 212 35888
rect 0 35828 90 35848
rect 172 35720 212 35848
rect 1804 35804 1844 35932
rect 2170 35923 2179 35932
rect 2219 35923 2228 35963
rect 2537 35932 2668 35972
rect 2708 35932 2717 35972
rect 3523 35932 3532 35972
rect 3572 35963 3956 35972
rect 3572 35932 3916 35963
rect 2170 35922 2228 35923
rect 4666 35932 4675 35972
rect 4715 35932 4724 35972
rect 4771 35932 4780 35972
rect 4820 35932 4829 35972
rect 5155 35932 5164 35972
rect 5204 35932 5213 35972
rect 5740 35963 5972 35972
rect 3916 35914 3956 35923
rect 2323 35848 2332 35888
rect 2372 35848 3436 35888
rect 3476 35848 3485 35888
rect 1411 35764 1420 35804
rect 1460 35764 1844 35804
rect 4099 35764 4108 35804
rect 4148 35764 4588 35804
rect 4628 35764 4637 35804
rect 4684 35720 4724 35932
rect 5164 35888 5204 35932
rect 5780 35932 5972 35963
rect 6019 35932 6028 35972
rect 6068 35932 6164 35972
rect 6220 35963 6260 35972
rect 5740 35914 5780 35923
rect 6442 35932 6451 35972
rect 6491 35963 6644 35972
rect 6491 35932 6595 35963
rect 4771 35848 4780 35888
rect 4820 35848 5204 35888
rect 5251 35848 5260 35888
rect 5300 35848 5431 35888
rect 6220 35804 6260 35923
rect 6586 35923 6595 35932
rect 6635 35923 6644 35963
rect 6700 35932 7180 35972
rect 7220 35932 7229 35972
rect 8393 35963 8524 35972
rect 8393 35932 8428 35963
rect 6586 35922 6644 35923
rect 8468 35932 8524 35963
rect 8564 35932 8573 35972
rect 8995 35932 9004 35972
rect 9044 35932 10060 35972
rect 10100 35932 10109 35972
rect 10243 35932 10252 35972
rect 10292 35932 11500 35972
rect 11540 35932 11549 35972
rect 8428 35914 8468 35923
rect 9004 35914 9044 35923
rect 6691 35848 6700 35888
rect 6740 35848 6748 35888
rect 6788 35848 6871 35888
rect 5155 35764 5164 35804
rect 5204 35764 6260 35804
rect 7171 35764 7180 35804
rect 7220 35764 8812 35804
rect 8852 35764 8861 35804
rect 172 35680 2956 35720
rect 2996 35680 3005 35720
rect 3100 35680 4724 35720
rect 0 35552 90 35572
rect 3100 35552 3140 35680
rect 0 35512 1228 35552
rect 1268 35512 1277 35552
rect 2956 35512 3140 35552
rect 3679 35512 3688 35552
rect 3728 35512 3770 35552
rect 3810 35512 3852 35552
rect 3892 35512 3934 35552
rect 3974 35512 4016 35552
rect 4056 35512 4065 35552
rect 0 35492 90 35512
rect 2956 35384 2996 35512
rect 3043 35428 3052 35468
rect 3092 35428 4628 35468
rect 1459 35344 1468 35384
rect 1508 35344 2188 35384
rect 2228 35344 2237 35384
rect 2659 35344 2668 35384
rect 2708 35344 2804 35384
rect 2956 35344 3052 35384
rect 3092 35344 3101 35384
rect 3715 35344 3724 35384
rect 3764 35344 4148 35384
rect 2764 35300 2804 35344
rect 2764 35260 4052 35300
rect 0 35216 90 35236
rect 0 35176 1036 35216
rect 1076 35176 1085 35216
rect 1219 35176 1228 35216
rect 1268 35176 1804 35216
rect 1844 35176 2284 35216
rect 2324 35176 2333 35216
rect 2860 35176 3052 35216
rect 3092 35176 3724 35216
rect 3764 35176 3773 35216
rect 0 35156 90 35176
rect 2860 35132 2900 35176
rect 4012 35132 4052 35260
rect 4108 35216 4148 35344
rect 4588 35300 4628 35428
rect 7468 35428 9196 35468
rect 9236 35428 9245 35468
rect 5155 35344 5164 35384
rect 5204 35344 5452 35384
rect 5492 35344 5501 35384
rect 7468 35300 7508 35428
rect 4588 35260 5780 35300
rect 5875 35260 5884 35300
rect 5924 35260 7508 35300
rect 7564 35344 11596 35384
rect 11636 35344 11645 35384
rect 5740 35216 5780 35260
rect 7564 35216 7604 35344
rect 11750 35216 11840 35236
rect 4108 35176 5300 35216
rect 5635 35176 5644 35216
rect 5684 35176 5693 35216
rect 5740 35176 6028 35216
rect 6068 35176 6077 35216
rect 6259 35176 6268 35216
rect 6308 35176 7604 35216
rect 8131 35176 8140 35216
rect 8180 35176 8756 35216
rect 10217 35176 10348 35216
rect 10388 35176 10397 35216
rect 11011 35176 11020 35216
rect 11060 35176 11840 35216
rect 5260 35132 5300 35176
rect 5644 35132 5684 35176
rect 7660 35132 7700 35141
rect 8716 35132 8756 35176
rect 11750 35156 11840 35176
rect 9964 35132 10004 35141
rect 835 35092 844 35132
rect 884 35092 1612 35132
rect 1652 35092 2668 35132
rect 2708 35092 2717 35132
rect 2860 35083 2900 35092
rect 2956 35092 3187 35132
rect 3227 35092 3236 35132
rect 4003 35092 4012 35132
rect 4052 35092 4061 35132
rect 5300 35092 5356 35132
rect 5396 35092 5431 35132
rect 5644 35092 6412 35132
rect 6452 35092 6508 35132
rect 6548 35092 6557 35132
rect 7747 35092 7756 35132
rect 7796 35092 8536 35132
rect 8576 35092 8585 35132
rect 8707 35092 8716 35132
rect 8756 35092 8765 35132
rect 9833 35092 9964 35132
rect 10004 35092 10013 35132
rect 2956 34964 2996 35092
rect 1795 34924 1804 34964
rect 1844 34924 2996 34964
rect 3244 35008 3668 35048
rect 0 34880 90 34900
rect 3244 34880 3284 35008
rect 3379 34924 3388 34964
rect 3428 34924 3437 34964
rect 0 34840 3284 34880
rect 0 34820 90 34840
rect 3388 34796 3428 34924
rect 3628 34880 3668 35008
rect 4012 34964 4052 35092
rect 5260 35083 5300 35092
rect 5644 34964 5684 35092
rect 7660 35048 7700 35092
rect 9964 35048 10004 35092
rect 7075 35008 7084 35048
rect 7124 35008 8371 35048
rect 8411 35008 8524 35048
rect 8564 35008 10004 35048
rect 3785 34924 3811 34964
rect 3851 34924 3916 34964
rect 3956 34924 3965 34964
rect 4012 34924 5684 34964
rect 7721 34924 7852 34964
rect 7892 34924 7901 34964
rect 9859 34924 9868 34964
rect 9908 34924 10156 34964
rect 10196 34924 10205 34964
rect 10579 34924 10588 34964
rect 10628 34924 11212 34964
rect 11252 34924 11261 34964
rect 3628 34840 7756 34880
rect 7796 34840 7805 34880
rect 3388 34756 4868 34796
rect 4919 34756 4928 34796
rect 4968 34756 5010 34796
rect 5050 34756 5092 34796
rect 5132 34756 5174 34796
rect 5214 34756 5256 34796
rect 5296 34756 5305 34796
rect 4828 34712 4868 34756
rect 2275 34672 2284 34712
rect 2324 34672 2476 34712
rect 2516 34672 2525 34712
rect 4828 34672 8585 34712
rect 8545 34628 8585 34672
rect 7385 34588 7468 34628
rect 7508 34588 7516 34628
rect 7556 34588 7565 34628
rect 8545 34588 8660 34628
rect 10522 34588 10531 34628
rect 10571 34588 10924 34628
rect 10964 34588 10973 34628
rect 0 34544 90 34564
rect 0 34504 1036 34544
rect 1076 34504 1085 34544
rect 1996 34504 2860 34544
rect 2900 34504 2909 34544
rect 3427 34504 3436 34544
rect 3476 34504 3860 34544
rect 0 34484 90 34504
rect 1996 34460 2036 34504
rect 1097 34451 1228 34460
rect 1097 34420 1219 34451
rect 1268 34420 1277 34460
rect 1865 34420 1996 34460
rect 2036 34420 2045 34460
rect 3244 34451 3532 34460
rect 1210 34411 1219 34420
rect 1259 34411 1268 34420
rect 1210 34410 1268 34411
rect 3284 34420 3532 34451
rect 3572 34420 3581 34460
rect 3244 34402 3284 34411
rect 1363 34336 1372 34376
rect 1412 34336 1748 34376
rect 1795 34336 1804 34376
rect 1844 34336 2188 34376
rect 2228 34336 2237 34376
rect 3427 34336 3436 34376
rect 3476 34336 3628 34376
rect 3668 34336 3677 34376
rect 0 34208 90 34228
rect 0 34168 76 34208
rect 116 34168 125 34208
rect 0 34148 90 34168
rect 1708 34124 1748 34336
rect 3820 34292 3860 34504
rect 3916 34504 4492 34544
rect 4532 34504 5588 34544
rect 7241 34504 7372 34544
rect 7412 34504 7421 34544
rect 8131 34504 8140 34544
rect 8180 34504 8564 34544
rect 3916 34460 3956 34504
rect 5548 34460 5588 34504
rect 8524 34460 8564 34504
rect 3907 34420 3916 34460
rect 3956 34420 3965 34460
rect 5164 34451 5356 34460
rect 5204 34420 5356 34451
rect 5396 34420 5405 34460
rect 5548 34420 5932 34460
rect 5972 34420 5981 34460
rect 7075 34420 7084 34460
rect 7124 34451 7255 34460
rect 7124 34420 7180 34451
rect 5164 34402 5204 34411
rect 5548 34376 5588 34420
rect 7220 34420 7255 34451
rect 7555 34420 7564 34460
rect 7604 34420 8035 34460
rect 8075 34420 8084 34460
rect 8131 34420 8140 34460
rect 8180 34420 8189 34460
rect 8515 34420 8524 34460
rect 8564 34420 8573 34460
rect 7180 34402 7220 34411
rect 8140 34376 8180 34420
rect 8620 34376 8660 34588
rect 8707 34504 8716 34544
rect 8756 34504 9620 34544
rect 9100 34451 9388 34460
rect 9140 34420 9388 34451
rect 9428 34420 9437 34460
rect 9580 34451 9620 34504
rect 9100 34402 9140 34411
rect 9802 34420 9811 34460
rect 9851 34451 10004 34460
rect 9851 34420 9955 34451
rect 9580 34402 9620 34411
rect 9946 34411 9955 34420
rect 9995 34411 10004 34451
rect 9946 34410 10004 34411
rect 5539 34336 5548 34376
rect 5588 34336 5597 34376
rect 7625 34336 7756 34376
rect 7796 34336 7805 34376
rect 8044 34336 8180 34376
rect 8611 34336 8620 34376
rect 8660 34336 8669 34376
rect 10099 34336 10108 34376
rect 10148 34336 10924 34376
rect 10964 34336 10973 34376
rect 8044 34292 8084 34336
rect 3820 34252 7084 34292
rect 7124 34252 8084 34292
rect 8620 34292 8660 34336
rect 8620 34252 9676 34292
rect 9716 34252 9725 34292
rect 8044 34208 8084 34252
rect 11750 34208 11840 34228
rect 3427 34168 3436 34208
rect 3476 34168 4492 34208
rect 4532 34168 4541 34208
rect 5225 34168 5356 34208
rect 5396 34168 5405 34208
rect 5779 34168 5788 34208
rect 5828 34168 6892 34208
rect 6932 34168 6941 34208
rect 8044 34168 8716 34208
rect 8756 34168 8765 34208
rect 11107 34168 11116 34208
rect 11156 34168 11840 34208
rect 11750 34148 11840 34168
rect 1708 34084 8428 34124
rect 8468 34084 8477 34124
rect 3679 34000 3688 34040
rect 3728 34000 3770 34040
rect 3810 34000 3852 34040
rect 3892 34000 3934 34040
rect 3974 34000 4016 34040
rect 4056 34000 4065 34040
rect 0 33872 90 33892
rect 0 33832 1516 33872
rect 1556 33832 1565 33872
rect 3964 33832 8660 33872
rect 0 33812 90 33832
rect 3964 33704 4004 33832
rect 4867 33748 4876 33788
rect 4916 33748 7028 33788
rect 6988 33704 7028 33748
rect 3331 33664 3340 33704
rect 3380 33664 3628 33704
rect 3668 33664 3677 33704
rect 3955 33664 3964 33704
rect 4004 33664 4013 33704
rect 4435 33664 4444 33704
rect 4484 33664 5644 33704
rect 5684 33664 5693 33704
rect 6211 33664 6220 33704
rect 6260 33664 6412 33704
rect 6452 33664 6461 33704
rect 6508 33664 6748 33704
rect 6788 33664 6797 33704
rect 6979 33664 6988 33704
rect 7028 33664 7037 33704
rect 7171 33664 7180 33704
rect 7220 33664 7351 33704
rect 7692 33664 7756 33704
rect 7796 33664 7852 33704
rect 7892 33664 8236 33704
rect 8276 33664 8285 33704
rect 2956 33620 2996 33629
rect 3340 33620 3380 33664
rect 6028 33620 6068 33629
rect 6508 33620 6548 33664
rect 8620 33620 8660 33832
rect 8707 33748 8716 33788
rect 8756 33748 9332 33788
rect 8707 33664 8716 33704
rect 8756 33664 9004 33704
rect 9044 33664 9053 33704
rect 9292 33620 9332 33748
rect 739 33580 748 33620
rect 788 33580 1171 33620
rect 1211 33580 1220 33620
rect 1699 33580 1708 33620
rect 1748 33580 1996 33620
rect 2036 33580 2045 33620
rect 2860 33580 2956 33620
rect 2996 33580 3052 33620
rect 3092 33580 3101 33620
rect 3293 33580 3328 33620
rect 3368 33580 3380 33620
rect 3427 33580 3436 33620
rect 3476 33580 3778 33620
rect 3818 33580 3827 33620
rect 4169 33580 4288 33620
rect 4340 33580 4349 33620
rect 4579 33580 4588 33620
rect 4628 33580 4780 33620
rect 4820 33580 4829 33620
rect 6115 33580 6124 33620
rect 6164 33580 6548 33620
rect 6787 33580 6796 33620
rect 6836 33580 7468 33620
rect 7508 33580 7517 33620
rect 7843 33580 7852 33620
rect 7892 33580 8227 33620
rect 8267 33580 8276 33620
rect 8323 33580 8332 33620
rect 8372 33580 8524 33620
rect 8564 33580 8573 33620
rect 8620 33580 8716 33620
rect 8756 33580 8812 33620
rect 8852 33580 8887 33620
rect 9737 33580 9811 33620
rect 9851 33580 9868 33620
rect 9908 33580 9917 33620
rect 9964 33580 10099 33620
rect 10139 33580 10148 33620
rect 0 33536 90 33556
rect 2860 33536 2900 33580
rect 2956 33571 2996 33580
rect 6028 33536 6068 33580
rect 9292 33571 9332 33580
rect 0 33496 1804 33536
rect 1844 33496 1853 33536
rect 2563 33496 2572 33536
rect 2612 33496 2900 33536
rect 3523 33496 3532 33536
rect 3572 33496 6404 33536
rect 6643 33496 6652 33536
rect 6692 33496 8140 33536
rect 8180 33496 8189 33536
rect 0 33476 90 33496
rect 1363 33412 1372 33452
rect 1412 33412 2900 33452
rect 3139 33412 3148 33452
rect 3188 33412 3340 33452
rect 3380 33412 3389 33452
rect 3475 33412 3484 33452
rect 3524 33412 3533 33452
rect 6089 33412 6220 33452
rect 6260 33412 6269 33452
rect 1372 33244 1516 33284
rect 1556 33244 1565 33284
rect 0 33200 90 33220
rect 0 33140 116 33200
rect 76 33032 116 33140
rect 1372 33116 1412 33244
rect 2860 33200 2900 33412
rect 3484 33368 3524 33412
rect 6364 33368 6404 33496
rect 9964 33452 10004 33580
rect 7258 33412 7267 33452
rect 7307 33412 7468 33452
rect 7508 33412 7517 33452
rect 9955 33412 9964 33452
rect 10004 33412 10013 33452
rect 10291 33412 10300 33452
rect 10340 33412 11116 33452
rect 11156 33412 11165 33452
rect 3484 33328 5396 33368
rect 6364 33328 7852 33368
rect 7892 33328 7901 33368
rect 5356 33284 5396 33328
rect 2947 33244 2956 33284
rect 2996 33244 3628 33284
rect 3668 33244 3677 33284
rect 4919 33244 4928 33284
rect 4968 33244 5010 33284
rect 5050 33244 5092 33284
rect 5132 33244 5174 33284
rect 5214 33244 5256 33284
rect 5296 33244 5305 33284
rect 5356 33244 5972 33284
rect 5932 33200 5972 33244
rect 11750 33200 11840 33220
rect 2860 33160 5876 33200
rect 5932 33160 10252 33200
rect 10292 33160 10301 33200
rect 11203 33160 11212 33200
rect 11252 33160 11840 33200
rect 1372 33076 1516 33116
rect 1556 33076 1565 33116
rect 5443 33076 5452 33116
rect 5492 33076 5501 33116
rect 76 32992 1364 33032
rect 1411 32992 1420 33032
rect 1460 32992 2956 33032
rect 2996 32992 3005 33032
rect 3244 32992 3916 33032
rect 3956 32992 3965 33032
rect 4780 32992 5260 33032
rect 5300 32992 5309 33032
rect 1324 32948 1364 32992
rect 1306 32908 1315 32948
rect 1355 32908 1364 32948
rect 1961 32908 1996 32948
rect 2036 32908 2092 32948
rect 2132 32908 2141 32948
rect 3244 32939 3284 32992
rect 3331 32908 3340 32948
rect 3380 32908 3715 32948
rect 3755 32908 3764 32948
rect 3811 32908 3820 32948
rect 3860 32908 3869 32948
rect 4169 32908 4204 32948
rect 4244 32908 4300 32948
rect 4340 32908 4349 32948
rect 4780 32939 4820 32992
rect 5452 32948 5492 33076
rect 5836 33032 5876 33160
rect 11750 33140 11840 33160
rect 6019 33076 6028 33116
rect 6068 33076 6796 33116
rect 6836 33076 6845 33116
rect 8236 33076 8524 33116
rect 8564 33076 8573 33116
rect 9763 33076 9772 33116
rect 9812 33076 9821 33116
rect 10522 33076 10531 33116
rect 10571 33076 11404 33116
rect 11444 33076 11453 33116
rect 5635 32992 5644 33032
rect 5684 32992 5780 33032
rect 5836 32992 6452 33032
rect 7747 32992 7756 33032
rect 7796 32992 8084 33032
rect 5740 32948 5780 32992
rect 0 32864 90 32884
rect 3244 32864 3284 32899
rect 3820 32864 3860 32908
rect 5225 32939 5356 32948
rect 5225 32908 5260 32939
rect 4780 32890 4820 32899
rect 5300 32908 5356 32939
rect 5396 32908 5405 32948
rect 5452 32939 5684 32948
rect 5452 32908 5635 32939
rect 5260 32890 5300 32899
rect 5626 32899 5635 32908
rect 5675 32899 5684 32939
rect 5740 32908 6316 32948
rect 6356 32908 6365 32948
rect 5626 32898 5684 32899
rect 0 32824 1132 32864
rect 1172 32824 1181 32864
rect 2659 32824 2668 32864
rect 2708 32824 3284 32864
rect 3523 32824 3532 32864
rect 3572 32824 3860 32864
rect 4291 32824 4300 32864
rect 4340 32824 4349 32864
rect 5779 32824 5788 32864
rect 5828 32824 6124 32864
rect 6164 32824 6173 32864
rect 0 32804 90 32824
rect 4300 32780 4340 32824
rect 2851 32740 2860 32780
rect 2900 32740 4340 32780
rect 6316 32780 6356 32908
rect 6412 32864 6452 32992
rect 8044 32948 8084 32992
rect 8236 32948 8276 33076
rect 8323 32992 8332 33032
rect 8372 32992 9140 33032
rect 7564 32939 7604 32948
rect 8026 32908 8035 32948
rect 8075 32908 8084 32948
rect 8131 32908 8140 32948
rect 8180 32908 8372 32948
rect 7564 32864 7604 32899
rect 6412 32824 6508 32864
rect 6548 32824 6557 32864
rect 7564 32824 8236 32864
rect 8276 32824 8285 32864
rect 6316 32740 6796 32780
rect 6836 32740 6845 32780
rect 1481 32656 1516 32696
rect 1556 32656 1612 32696
rect 1652 32656 1661 32696
rect 3427 32656 3436 32696
rect 3476 32656 3485 32696
rect 3619 32656 3628 32696
rect 3668 32656 4204 32696
rect 4244 32656 4253 32696
rect 2947 32572 2956 32612
rect 2996 32572 3244 32612
rect 3284 32572 3293 32612
rect 0 32528 90 32548
rect 0 32488 1324 32528
rect 1364 32488 1373 32528
rect 0 32468 90 32488
rect 3436 32276 3476 32656
rect 4300 32612 4340 32740
rect 8332 32696 8372 32908
rect 8428 32908 8528 32948
rect 8568 32908 9004 32948
rect 9044 32908 9053 32948
rect 9100 32939 9140 32992
rect 9772 32948 9812 33076
rect 8428 32780 8468 32908
rect 9100 32864 9140 32899
rect 9580 32939 9620 32948
rect 9772 32939 10004 32948
rect 9772 32908 9955 32939
rect 8585 32824 8620 32864
rect 8660 32824 8716 32864
rect 8756 32824 8765 32864
rect 9091 32824 9100 32864
rect 9140 32824 9216 32864
rect 8716 32780 8756 32824
rect 8428 32740 8524 32780
rect 8564 32740 8573 32780
rect 8716 32740 9292 32780
rect 9332 32740 9341 32780
rect 8332 32656 8756 32696
rect 8716 32612 8756 32656
rect 4300 32572 8524 32612
rect 8564 32572 8573 32612
rect 8707 32572 8716 32612
rect 8756 32572 8765 32612
rect 3679 32488 3688 32528
rect 3728 32488 3770 32528
rect 3810 32488 3852 32528
rect 3892 32488 3934 32528
rect 3974 32488 4016 32528
rect 4056 32488 4065 32528
rect 4300 32360 4340 32572
rect 9580 32360 9620 32899
rect 9946 32899 9955 32908
rect 9995 32899 10004 32939
rect 9946 32898 10004 32899
rect 10051 32824 10060 32864
rect 10100 32824 10108 32864
rect 10148 32824 10231 32864
rect 4003 32320 4012 32360
rect 4052 32320 4340 32360
rect 7843 32320 7852 32360
rect 7892 32320 9620 32360
rect 9676 32320 10732 32360
rect 10772 32320 10781 32360
rect 9676 32276 9716 32320
rect 3436 32236 4148 32276
rect 0 32192 90 32212
rect 0 32152 460 32192
rect 500 32152 509 32192
rect 3139 32152 3148 32192
rect 3188 32152 3436 32192
rect 3476 32152 3532 32192
rect 3572 32152 3636 32192
rect 0 32132 90 32152
rect 2476 32108 2516 32117
rect 4012 32108 4052 32117
rect 4108 32108 4148 32236
rect 9292 32236 9716 32276
rect 9811 32236 9820 32276
rect 9860 32236 10868 32276
rect 9292 32192 9332 32236
rect 10828 32192 10868 32236
rect 11750 32192 11840 32212
rect 4195 32152 4204 32192
rect 4244 32152 6452 32192
rect 6412 32108 6452 32152
rect 7660 32152 8179 32192
rect 8219 32152 8236 32192
rect 8276 32152 8285 32192
rect 8611 32152 8620 32192
rect 8660 32152 9004 32192
rect 9044 32152 9053 32192
rect 9283 32152 9292 32192
rect 9332 32152 9341 32192
rect 9449 32152 9580 32192
rect 9620 32152 9629 32192
rect 9955 32152 9964 32192
rect 10004 32152 10156 32192
rect 10196 32152 10205 32192
rect 10339 32152 10348 32192
rect 10388 32152 10397 32192
rect 10828 32152 11840 32192
rect 7660 32108 7700 32152
rect 9292 32108 9332 32152
rect 10348 32108 10388 32152
rect 11750 32132 11840 32152
rect 1219 32068 1228 32108
rect 1268 32068 1420 32108
rect 1460 32068 1469 32108
rect 2516 32068 2668 32108
rect 2708 32068 2717 32108
rect 2860 32068 2947 32108
rect 2987 32068 2996 32108
rect 3043 32068 3052 32108
rect 3092 32068 3101 32108
rect 3523 32068 3532 32108
rect 3572 32068 3581 32108
rect 3881 32068 4012 32108
rect 4052 32068 4061 32108
rect 4108 32068 4500 32108
rect 4540 32068 4549 32108
rect 4684 32068 4819 32108
rect 4859 32068 4868 32108
rect 5164 32068 5314 32108
rect 5354 32068 5363 32108
rect 5827 32068 5836 32108
rect 5876 32068 6028 32108
rect 6068 32068 6077 32108
rect 6403 32068 6412 32108
rect 6452 32068 6461 32108
rect 8222 32068 8332 32108
rect 8384 32068 8402 32108
rect 8515 32068 8524 32108
rect 8564 32068 9332 32108
rect 10243 32068 10252 32108
rect 10292 32068 10388 32108
rect 2476 32059 2516 32068
rect 2860 32024 2900 32068
rect 2659 31984 2668 32024
rect 2708 31984 2900 32024
rect 3052 31940 3092 32068
rect 1507 31900 1516 31940
rect 1556 31900 3092 31940
rect 3532 31940 3572 32068
rect 4012 32059 4052 32068
rect 4684 31940 4724 32068
rect 3532 31900 4300 31940
rect 4340 31900 4349 31940
rect 4675 31900 4684 31940
rect 4724 31900 4733 31940
rect 4867 31900 4876 31940
rect 4916 31900 5020 31940
rect 5060 31900 5069 31940
rect 0 31856 90 31876
rect 5164 31856 5204 32068
rect 6028 32024 6068 32068
rect 7660 32059 7700 32068
rect 6028 31984 6892 32024
rect 6932 31984 6941 32024
rect 10195 31984 10204 32024
rect 10244 31984 11020 32024
rect 11060 31984 11069 32024
rect 5491 31900 5500 31940
rect 5540 31900 5644 31940
rect 5684 31900 5693 31940
rect 5993 31900 6115 31940
rect 6164 31900 6173 31940
rect 8969 31900 9091 31940
rect 9140 31900 9149 31940
rect 10579 31900 10588 31940
rect 10628 31900 11212 31940
rect 11252 31900 11261 31940
rect 0 31816 5204 31856
rect 0 31796 90 31816
rect 6124 31772 6164 31900
rect 835 31732 844 31772
rect 884 31732 1420 31772
rect 1460 31732 1469 31772
rect 2659 31732 2668 31772
rect 2708 31732 2956 31772
rect 2996 31732 3005 31772
rect 4919 31732 4928 31772
rect 4968 31732 5010 31772
rect 5050 31732 5092 31772
rect 5132 31732 5174 31772
rect 5214 31732 5256 31772
rect 5296 31732 5305 31772
rect 6124 31732 6932 31772
rect 355 31648 364 31688
rect 404 31648 2612 31688
rect 2572 31604 2612 31648
rect 1900 31564 2324 31604
rect 2572 31564 2620 31604
rect 2660 31564 2669 31604
rect 3187 31564 3196 31604
rect 3236 31564 4780 31604
rect 4820 31564 4829 31604
rect 5155 31564 5164 31604
rect 5204 31564 5396 31604
rect 0 31520 90 31540
rect 1900 31520 1940 31564
rect 0 31480 1940 31520
rect 2284 31520 2324 31564
rect 2284 31480 3436 31520
rect 3476 31480 3485 31520
rect 4003 31480 4012 31520
rect 4052 31480 4061 31520
rect 0 31460 90 31480
rect 4012 31436 4052 31480
rect 5356 31436 5396 31564
rect 6892 31520 6932 31732
rect 7267 31648 7276 31688
rect 7316 31648 10828 31688
rect 10868 31648 10877 31688
rect 7066 31564 7075 31604
rect 7115 31564 7756 31604
rect 7796 31564 7805 31604
rect 8105 31564 8179 31604
rect 8219 31564 8236 31604
rect 8276 31564 8285 31604
rect 1193 31396 1315 31436
rect 1364 31396 1373 31436
rect 1420 31427 2036 31436
rect 1420 31396 1987 31427
rect 1420 31352 1460 31396
rect 1978 31387 1987 31396
rect 2027 31387 2036 31427
rect 1978 31386 2036 31387
rect 2458 31427 2516 31436
rect 2458 31387 2467 31427
rect 2507 31387 2516 31427
rect 2659 31396 2668 31436
rect 2708 31396 3427 31436
rect 3467 31396 3476 31436
rect 3523 31396 3532 31436
rect 3572 31396 3703 31436
rect 3907 31396 3916 31436
rect 3956 31396 3965 31436
rect 4012 31427 4532 31436
rect 4012 31396 4492 31427
rect 2458 31386 2516 31387
rect 1027 31312 1036 31352
rect 1076 31312 1460 31352
rect 2131 31312 2140 31352
rect 2180 31312 2228 31352
rect 0 31184 90 31204
rect 2188 31184 2228 31312
rect 0 31144 1228 31184
rect 1268 31144 1277 31184
rect 1385 31144 1516 31184
rect 1556 31144 1565 31184
rect 2179 31144 2188 31184
rect 2228 31144 2237 31184
rect 0 31124 90 31144
rect 2476 31100 2516 31386
rect 3916 31352 3956 31396
rect 4675 31396 4684 31436
rect 4724 31427 5012 31436
rect 4724 31396 4972 31427
rect 4492 31378 4532 31387
rect 4972 31378 5012 31387
rect 5338 31427 5396 31436
rect 5338 31387 5347 31427
rect 5387 31387 5396 31427
rect 5338 31386 5396 31387
rect 5740 31480 6220 31520
rect 6260 31480 6269 31520
rect 6892 31480 7124 31520
rect 7267 31480 7276 31520
rect 7316 31480 7447 31520
rect 7699 31480 7708 31520
rect 7748 31480 8620 31520
rect 8660 31480 8669 31520
rect 2851 31312 2860 31352
rect 2900 31312 2956 31352
rect 2996 31312 3031 31352
rect 3139 31312 3148 31352
rect 3188 31312 3956 31352
rect 4003 31312 4012 31352
rect 4052 31312 4061 31352
rect 5491 31312 5500 31352
rect 5540 31312 5548 31352
rect 5588 31312 5671 31352
rect 4012 31268 4052 31312
rect 4012 31228 4300 31268
rect 4340 31228 4780 31268
rect 4820 31228 4829 31268
rect 5740 31184 5780 31480
rect 5827 31312 5836 31352
rect 5876 31312 5885 31352
rect 3619 31144 3628 31184
rect 3668 31144 5780 31184
rect 451 31060 460 31100
rect 500 31060 2516 31100
rect 3679 30976 3688 31016
rect 3728 30976 3770 31016
rect 3810 30976 3852 31016
rect 3892 30976 3934 31016
rect 3974 30976 4016 31016
rect 4056 30976 4065 31016
rect 5836 30932 5876 31312
rect 6028 31268 6068 31480
rect 7084 31436 7124 31480
rect 6115 31396 6124 31436
rect 6164 31396 6508 31436
rect 6548 31396 6557 31436
rect 7075 31396 7084 31436
rect 7124 31396 7133 31436
rect 7546 31427 7604 31436
rect 7546 31387 7555 31427
rect 7595 31387 7604 31427
rect 8602 31396 8611 31436
rect 8651 31396 8660 31436
rect 8707 31396 8716 31436
rect 8756 31396 8887 31436
rect 8995 31396 9004 31436
rect 9044 31396 9100 31436
rect 9140 31396 9175 31436
rect 9571 31396 9580 31436
rect 9620 31427 9751 31436
rect 9620 31396 9676 31427
rect 7546 31386 7604 31387
rect 7564 31268 7604 31386
rect 8249 31354 8332 31394
rect 8411 31354 8429 31394
rect 6019 31228 6028 31268
rect 6068 31228 6077 31268
rect 7555 31228 7564 31268
rect 7604 31228 7613 31268
rect 6067 31144 6076 31184
rect 6116 31144 6604 31184
rect 6644 31144 6653 31184
rect 1411 30892 1420 30932
rect 1460 30892 5876 30932
rect 0 30848 90 30868
rect 8620 30848 8660 31396
rect 9716 31396 9751 31427
rect 10025 31396 10156 31436
rect 10196 31396 10205 31436
rect 9676 31378 9716 31387
rect 10156 31378 10196 31387
rect 9161 31312 9196 31352
rect 9236 31312 9292 31352
rect 9332 31312 9341 31352
rect 11750 31184 11840 31204
rect 10156 31144 10387 31184
rect 10427 31144 10436 31184
rect 11011 31144 11020 31184
rect 11060 31144 11840 31184
rect 0 30808 1324 30848
rect 1364 30808 1373 30848
rect 8620 30808 9292 30848
rect 9332 30808 9341 30848
rect 0 30788 90 30808
rect 10156 30764 10196 31144
rect 11750 31124 11840 31144
rect 10339 30808 10348 30848
rect 10388 30808 10396 30848
rect 10436 30808 10519 30848
rect 1507 30724 1516 30764
rect 1556 30724 2860 30764
rect 2900 30724 2909 30764
rect 3235 30724 3244 30764
rect 3284 30724 4628 30764
rect 7171 30724 7180 30764
rect 7220 30724 7892 30764
rect 1891 30640 1900 30680
rect 1940 30640 2708 30680
rect 2668 30596 2708 30640
rect 3586 30640 3628 30680
rect 3668 30640 3677 30680
rect 3859 30640 3868 30680
rect 3908 30640 4012 30680
rect 4052 30640 4061 30680
rect 3586 30596 3626 30640
rect 4588 30596 4628 30724
rect 6019 30640 6028 30680
rect 6068 30640 7220 30680
rect 5836 30596 5876 30605
rect 7180 30596 7220 30640
rect 7468 30596 7508 30605
rect 7852 30596 7892 30724
rect 10060 30724 10196 30764
rect 10060 30638 10100 30724
rect 10147 30640 10156 30680
rect 10196 30640 10205 30680
rect 9100 30596 9140 30605
rect 9994 30598 10003 30638
rect 10043 30598 10100 30638
rect 1411 30556 1420 30596
rect 1460 30556 1996 30596
rect 2036 30556 2045 30596
rect 2668 30547 2708 30556
rect 2956 30556 3340 30596
rect 3380 30556 3389 30596
rect 3450 30556 3459 30596
rect 3499 30556 3524 30596
rect 3568 30556 3577 30596
rect 3617 30556 3626 30596
rect 3703 30556 3712 30596
rect 3752 30556 3764 30596
rect 3811 30556 3820 30596
rect 3860 30556 4204 30596
rect 4244 30556 4253 30596
rect 4387 30556 4396 30596
rect 4436 30556 4445 30596
rect 4579 30556 4588 30596
rect 4628 30556 4637 30596
rect 6211 30556 6220 30596
rect 6260 30556 6796 30596
rect 6836 30556 6845 30596
rect 7171 30556 7180 30596
rect 7220 30556 7229 30596
rect 7433 30556 7468 30596
rect 7508 30556 7564 30596
rect 7604 30556 7613 30596
rect 7843 30556 7852 30596
rect 7892 30556 8044 30596
rect 8084 30556 8093 30596
rect 8803 30556 8812 30596
rect 8852 30556 9100 30596
rect 9140 30556 9868 30596
rect 9908 30556 9917 30596
rect 0 30512 90 30532
rect 0 30472 748 30512
rect 788 30472 797 30512
rect 0 30452 90 30472
rect 2956 30428 2996 30556
rect 3484 30428 3524 30556
rect 2851 30388 2860 30428
rect 2900 30388 2956 30428
rect 2996 30388 3031 30428
rect 3235 30388 3244 30428
rect 3284 30388 3415 30428
rect 3484 30388 3628 30428
rect 3668 30388 3677 30428
rect 3724 30344 3764 30556
rect 4396 30512 4436 30556
rect 4195 30472 4204 30512
rect 4244 30472 4436 30512
rect 5836 30512 5876 30556
rect 7468 30512 7508 30556
rect 9100 30547 9140 30556
rect 5836 30472 7372 30512
rect 7412 30472 7508 30512
rect 10156 30428 10196 30640
rect 4169 30388 4300 30428
rect 4340 30388 4349 30428
rect 5897 30388 6028 30428
rect 6068 30388 6077 30428
rect 7529 30388 7660 30428
rect 7700 30388 7709 30428
rect 9802 30388 9811 30428
rect 9851 30388 9868 30428
rect 9908 30388 9991 30428
rect 10060 30388 10196 30428
rect 10060 30344 10100 30388
rect 3331 30304 3340 30344
rect 3380 30304 3764 30344
rect 9475 30304 9484 30344
rect 9524 30304 10100 30344
rect 4919 30220 4928 30260
rect 4968 30220 5010 30260
rect 5050 30220 5092 30260
rect 5132 30220 5174 30260
rect 5214 30220 5256 30260
rect 5296 30220 5305 30260
rect 0 30176 90 30196
rect 11750 30176 11840 30196
rect 0 30136 1420 30176
rect 1460 30136 1469 30176
rect 2668 30136 4012 30176
rect 4052 30136 4061 30176
rect 4108 30136 4436 30176
rect 11203 30136 11212 30176
rect 11252 30136 11840 30176
rect 0 30116 90 30136
rect 2668 30092 2708 30136
rect 4108 30092 4148 30136
rect 2659 30052 2668 30092
rect 2708 30052 2717 30092
rect 3100 30052 4148 30092
rect 3100 29924 3140 30052
rect 4396 30050 4436 30136
rect 11750 30116 11840 30136
rect 4867 30052 4876 30092
rect 4916 30052 5212 30092
rect 5252 30052 5261 30092
rect 7843 30052 7852 30092
rect 7892 30052 7901 30092
rect 10147 30052 10156 30092
rect 10196 30052 10540 30092
rect 10580 30052 10589 30092
rect 4378 30010 4387 30050
rect 4427 30010 4436 30050
rect 3203 29968 3244 30008
rect 3284 29968 3293 30008
rect 3811 29968 3820 30008
rect 3860 29968 4292 30008
rect 3203 29924 3243 29968
rect 4252 29924 4292 29968
rect 4611 29968 4972 30008
rect 5012 29968 5021 30008
rect 4611 29924 4651 29968
rect 7852 29924 7892 30052
rect 8707 29968 8716 30008
rect 8756 29968 9004 30008
rect 9044 29968 9053 30008
rect 835 29884 844 29924
rect 884 29884 1228 29924
rect 1268 29884 1277 29924
rect 1891 29884 1900 29924
rect 1940 29915 2516 29924
rect 1940 29884 2476 29915
rect 2476 29866 2516 29875
rect 2978 29866 2987 29906
rect 3027 29866 3039 29906
rect 3095 29884 3104 29924
rect 3144 29884 3153 29924
rect 3203 29884 3226 29924
rect 3266 29884 3275 29924
rect 3427 29884 3436 29924
rect 3476 29884 3485 29924
rect 3628 29884 3724 29924
rect 3764 29884 3773 29924
rect 4003 29884 4012 29924
rect 4052 29884 4156 29924
rect 4196 29884 4205 29924
rect 4252 29884 4457 29924
rect 4497 29884 4506 29924
rect 4602 29884 4611 29924
rect 4651 29884 4660 29924
rect 4762 29915 4780 29924
rect 0 29840 90 29860
rect 2999 29840 3039 29866
rect 0 29800 1324 29840
rect 1364 29800 1373 29840
rect 2999 29800 3052 29840
rect 3092 29800 3101 29840
rect 0 29780 90 29800
rect 3436 29756 3476 29884
rect 3052 29716 3476 29756
rect 3052 29588 3092 29716
rect 3139 29632 3148 29672
rect 3188 29632 3499 29672
rect 3459 29588 3499 29632
rect 3628 29588 3668 29884
rect 4762 29875 4771 29915
rect 4820 29884 4951 29924
rect 5993 29884 6028 29924
rect 6068 29884 6115 29924
rect 6155 29884 6173 29924
rect 6216 29884 6225 29924
rect 6265 29884 6274 29924
rect 6473 29884 6604 29924
rect 6644 29884 6653 29924
rect 7180 29915 7372 29924
rect 4811 29875 4820 29884
rect 4762 29874 4820 29875
rect 6220 29840 6260 29884
rect 7220 29884 7372 29915
rect 7412 29884 7421 29924
rect 7529 29884 7660 29924
rect 7700 29884 7709 29924
rect 7852 29915 8084 29924
rect 7852 29884 8035 29915
rect 7180 29866 7220 29875
rect 7660 29866 7700 29875
rect 8026 29875 8035 29884
rect 8075 29875 8084 29915
rect 9091 29884 9100 29924
rect 9140 29884 9484 29924
rect 9524 29884 9533 29924
rect 10051 29884 10060 29924
rect 10100 29915 10388 29924
rect 10100 29884 10348 29915
rect 8026 29874 8084 29875
rect 10348 29866 10388 29875
rect 4291 29800 4300 29840
rect 4340 29800 4349 29840
rect 4867 29800 4876 29840
rect 4916 29800 4924 29840
rect 4964 29800 5047 29840
rect 5155 29800 5164 29840
rect 5204 29800 5452 29840
rect 5492 29800 5501 29840
rect 5827 29800 5836 29840
rect 5876 29800 5932 29840
rect 5972 29800 6007 29840
rect 6124 29800 6260 29840
rect 6403 29800 6412 29840
rect 6452 29800 6700 29840
rect 6740 29800 6749 29840
rect 8179 29800 8188 29840
rect 8228 29800 8236 29840
rect 8276 29800 8359 29840
rect 8585 29800 8716 29840
rect 8756 29800 8765 29840
rect 3785 29632 3820 29672
rect 3860 29632 3916 29672
rect 3956 29632 3965 29672
rect 3052 29548 3188 29588
rect 3459 29548 3668 29588
rect 0 29504 90 29524
rect 0 29464 2900 29504
rect 0 29444 90 29464
rect 2860 29252 2900 29464
rect 3148 29336 3188 29548
rect 3679 29464 3688 29504
rect 3728 29464 3770 29504
rect 3810 29464 3852 29504
rect 3892 29464 3934 29504
rect 3974 29464 4016 29504
rect 4056 29464 4065 29504
rect 4300 29336 4340 29800
rect 6124 29756 6164 29800
rect 4387 29716 4396 29756
rect 4436 29716 5492 29756
rect 5539 29716 5548 29756
rect 5588 29716 6164 29756
rect 5452 29672 5492 29716
rect 5452 29632 5596 29672
rect 5636 29632 5645 29672
rect 8947 29632 8956 29672
rect 8996 29632 10828 29672
rect 10868 29632 10877 29672
rect 3130 29296 3139 29336
rect 3179 29296 3188 29336
rect 4195 29296 4204 29336
rect 4244 29296 4340 29336
rect 259 29212 268 29252
rect 308 29212 2804 29252
rect 2860 29212 5164 29252
rect 5204 29212 5213 29252
rect 5644 29212 6604 29252
rect 6644 29212 6653 29252
rect 8524 29212 8716 29252
rect 8756 29212 9004 29252
rect 9044 29212 9053 29252
rect 0 29168 90 29188
rect 2764 29168 2804 29212
rect 0 29128 1516 29168
rect 1556 29128 1565 29168
rect 2371 29128 2380 29168
rect 2459 29128 2551 29168
rect 2755 29128 2764 29168
rect 2804 29128 2813 29168
rect 3398 29128 4300 29168
rect 4340 29128 4349 29168
rect 4771 29128 4780 29168
rect 4820 29128 5164 29168
rect 5204 29128 5548 29168
rect 5588 29128 5597 29168
rect 0 29108 90 29128
rect 3398 29084 3438 29128
rect 5644 29084 5684 29212
rect 739 29044 748 29084
rect 788 29044 1171 29084
rect 1211 29044 1220 29084
rect 1315 29044 1324 29084
rect 1364 29044 1666 29084
rect 1706 29044 1715 29084
rect 2467 29044 2476 29084
rect 2516 29044 2584 29084
rect 2624 29044 2647 29084
rect 3017 29044 3139 29084
rect 3188 29044 3197 29084
rect 3248 29044 3257 29084
rect 3297 29044 3306 29084
rect 3380 29044 3389 29084
rect 3429 29044 3438 29084
rect 3514 29044 3523 29084
rect 3563 29044 3619 29084
rect 3691 29044 3700 29084
rect 3740 29044 3749 29084
rect 3898 29044 3907 29084
rect 3947 29044 3956 29084
rect 4099 29044 4108 29084
rect 4148 29044 4204 29084
rect 4244 29044 4279 29084
rect 4483 29044 4492 29084
rect 4532 29044 4675 29084
rect 4715 29044 4724 29084
rect 4771 29044 4780 29084
rect 4820 29044 4829 29084
rect 5225 29044 5260 29084
rect 5300 29044 5356 29084
rect 5396 29044 5684 29084
rect 5740 29128 5932 29168
rect 5972 29128 6412 29168
rect 6452 29128 6461 29168
rect 7075 29128 7084 29168
rect 7124 29128 7468 29168
rect 7508 29128 7517 29168
rect 5740 29084 5780 29128
rect 8524 29084 8564 29212
rect 11750 29168 11840 29188
rect 9161 29128 9196 29168
rect 9236 29128 9292 29168
rect 9332 29128 9341 29168
rect 10217 29128 10348 29168
rect 10388 29128 10397 29168
rect 10819 29128 10828 29168
rect 10868 29128 11840 29168
rect 11750 29108 11840 29128
rect 8812 29084 8852 29093
rect 6106 29044 6220 29084
rect 6268 29044 6286 29084
rect 6442 29044 6451 29084
rect 6491 29044 6547 29084
rect 6587 29044 6631 29084
rect 7555 29044 7564 29084
rect 7604 29044 8564 29084
rect 8681 29044 8812 29084
rect 8852 29044 8861 29084
rect 9997 29044 10006 29084
rect 10046 29044 10252 29084
rect 10292 29044 10301 29084
rect 3266 29000 3306 29044
rect 3532 29000 3572 29044
rect 3709 29000 3749 29044
rect 3916 29000 3956 29044
rect 4780 29000 4820 29044
rect 5740 29035 5780 29044
rect 8812 29035 8852 29044
rect 1843 28960 1852 29000
rect 1892 28960 2572 29000
rect 2612 28960 2621 29000
rect 2851 28960 2860 29000
rect 2900 28960 3004 29000
rect 3044 28960 3053 29000
rect 3219 28960 3244 29000
rect 3284 28960 3306 29000
rect 3523 28960 3532 29000
rect 3572 28960 3581 29000
rect 3709 28960 3724 29000
rect 3764 28960 3796 29000
rect 3916 28960 4204 29000
rect 4244 28960 4253 29000
rect 4387 28960 4396 29000
rect 4436 28960 4820 29000
rect 6316 28960 7468 29000
rect 7508 28960 7517 29000
rect 6316 28916 6356 28960
rect 1363 28876 1372 28916
rect 1412 28876 2180 28916
rect 0 28832 90 28852
rect 2140 28832 2180 28876
rect 5356 28876 6356 28916
rect 6739 28876 6748 28916
rect 6788 28876 6796 28916
rect 6836 28876 6919 28916
rect 7066 28876 7075 28916
rect 7115 28876 7124 28916
rect 8995 28876 9004 28916
rect 9044 28876 9053 28916
rect 9523 28876 9532 28916
rect 9572 28876 9620 28916
rect 9667 28876 9676 28916
rect 9716 28876 9811 28916
rect 9851 28876 9860 28916
rect 10579 28876 10588 28916
rect 10628 28876 11500 28916
rect 11540 28876 11549 28916
rect 0 28792 1708 28832
rect 1748 28792 1757 28832
rect 2140 28792 3572 28832
rect 0 28772 90 28792
rect 3532 28664 3572 28792
rect 4919 28708 4928 28748
rect 4968 28708 5010 28748
rect 5050 28708 5092 28748
rect 5132 28708 5174 28748
rect 5214 28708 5256 28748
rect 5296 28708 5305 28748
rect 5356 28664 5396 28876
rect 7084 28832 7124 28876
rect 6019 28792 6028 28832
rect 6068 28792 7124 28832
rect 8428 28792 8524 28832
rect 8564 28792 8573 28832
rect 7267 28708 7276 28748
rect 7316 28708 7325 28748
rect 76 28624 3340 28664
rect 3380 28624 3389 28664
rect 3532 28624 5396 28664
rect 7276 28664 7316 28708
rect 7276 28624 7604 28664
rect 76 28516 116 28624
rect 7564 28580 7604 28624
rect 8428 28580 8468 28792
rect 2659 28540 2668 28580
rect 2708 28540 2860 28580
rect 2900 28540 2909 28580
rect 3593 28540 3724 28580
rect 3764 28540 3773 28580
rect 4195 28540 4204 28580
rect 4244 28540 4628 28580
rect 6211 28540 6220 28580
rect 6260 28540 6269 28580
rect 6761 28540 6883 28580
rect 6932 28540 6941 28580
rect 7075 28540 7084 28580
rect 7124 28540 7171 28580
rect 7211 28540 7276 28580
rect 7316 28540 7380 28580
rect 7546 28540 7555 28580
rect 7595 28540 7660 28580
rect 7700 28540 7764 28580
rect 7930 28540 7939 28580
rect 7979 28540 8468 28580
rect 0 28456 116 28516
rect 2467 28456 2476 28496
rect 2516 28456 3187 28496
rect 3227 28456 3236 28496
rect 3427 28456 3436 28496
rect 3476 28456 3628 28496
rect 3668 28456 3677 28496
rect 3825 28456 3834 28496
rect 3874 28456 4108 28496
rect 4148 28456 4157 28496
rect 0 28436 90 28456
rect 4588 28412 4628 28540
rect 6220 28412 6260 28540
rect 9004 28496 9044 28876
rect 9580 28664 9620 28876
rect 9580 28624 10924 28664
rect 10964 28624 10973 28664
rect 10121 28540 10252 28580
rect 10292 28540 10301 28580
rect 10522 28540 10531 28580
rect 10571 28540 11404 28580
rect 11444 28540 11453 28580
rect 7843 28456 7852 28496
rect 7892 28456 7901 28496
rect 8524 28456 9044 28496
rect 9667 28456 9676 28496
rect 9716 28456 10444 28496
rect 10484 28456 10493 28496
rect 7852 28412 7892 28456
rect 8524 28412 8564 28456
rect 1219 28372 1228 28412
rect 1268 28372 1420 28412
rect 1460 28372 1708 28412
rect 1748 28372 1757 28412
rect 2668 28403 2708 28412
rect 3230 28372 3340 28412
rect 3392 28372 3410 28412
rect 3514 28372 3523 28412
rect 3563 28372 3572 28412
rect 3881 28372 4012 28412
rect 4052 28372 4061 28412
rect 4186 28372 4195 28412
rect 4235 28372 4244 28412
rect 4474 28372 4483 28412
rect 4523 28372 4532 28412
rect 4579 28372 4588 28412
rect 4628 28372 4637 28412
rect 4771 28372 4780 28412
rect 4820 28372 4972 28412
rect 5012 28372 5021 28412
rect 5548 28403 5932 28412
rect 2668 28244 2708 28363
rect 3532 28328 3572 28372
rect 4204 28328 4244 28372
rect 3532 28288 4108 28328
rect 4148 28288 4244 28328
rect 2668 28204 4300 28244
rect 4340 28204 4349 28244
rect 0 28160 90 28180
rect 0 28120 460 28160
rect 500 28120 509 28160
rect 0 28100 90 28120
rect 3679 27952 3688 27992
rect 3728 27952 3770 27992
rect 3810 27952 3852 27992
rect 3892 27952 3934 27992
rect 3974 27952 4016 27992
rect 4056 27952 4065 27992
rect 0 27824 90 27844
rect 4492 27824 4532 28372
rect 5588 28372 5932 28403
rect 5972 28372 5981 28412
rect 6028 28403 6068 28412
rect 5548 28354 5588 28363
rect 6220 28403 6452 28412
rect 6220 28372 6403 28403
rect 5059 28288 5068 28328
rect 5108 28288 5356 28328
rect 5396 28288 5405 28328
rect 6028 27824 6068 28363
rect 6394 28363 6403 28372
rect 6443 28363 6452 28403
rect 6394 28362 6452 28363
rect 7276 28372 7892 28412
rect 8506 28372 8515 28412
rect 8555 28372 8564 28412
rect 8611 28372 8620 28412
rect 8660 28372 8669 28412
rect 8716 28372 9004 28412
rect 9044 28372 9053 28412
rect 9283 28372 9292 28412
rect 9332 28403 9620 28412
rect 9332 28372 9580 28403
rect 7276 28328 7316 28372
rect 8620 28328 8660 28372
rect 6547 28288 6556 28328
rect 6596 28288 6604 28328
rect 6644 28288 6727 28328
rect 7171 28288 7180 28328
rect 7220 28288 7316 28328
rect 7721 28288 7852 28328
rect 7892 28288 7901 28328
rect 8105 28288 8140 28328
rect 8180 28288 8236 28328
rect 8276 28288 8285 28328
rect 8524 28288 8660 28328
rect 8524 28244 8564 28288
rect 6403 28204 6412 28244
rect 6452 28204 8564 28244
rect 8716 28160 8756 28372
rect 9580 28354 9620 28363
rect 10060 28403 10100 28412
rect 10060 28328 10100 28363
rect 9091 28288 9100 28328
rect 9140 28288 9187 28328
rect 9859 28288 9868 28328
rect 9908 28288 10004 28328
rect 10060 28288 10388 28328
rect 9100 28244 9140 28288
rect 9091 28204 9100 28244
rect 9140 28204 9149 28244
rect 8131 28120 8140 28160
rect 8180 28120 8524 28160
rect 8564 28120 8756 28160
rect 9964 28076 10004 28288
rect 9955 28036 9964 28076
rect 10004 28036 10013 28076
rect 10348 27824 10388 28288
rect 11750 28160 11840 28180
rect 10915 28120 10924 28160
rect 10964 28120 11840 28160
rect 11750 28100 11840 28120
rect 0 27784 1036 27824
rect 1076 27784 1085 27824
rect 3907 27784 3916 27824
rect 3956 27784 4532 27824
rect 5923 27784 5932 27824
rect 5972 27784 6068 27824
rect 10339 27784 10348 27824
rect 10388 27784 10397 27824
rect 0 27764 90 27784
rect 1507 27700 1516 27740
rect 1556 27700 4148 27740
rect 4339 27700 4348 27740
rect 4388 27700 5740 27740
rect 5780 27700 5789 27740
rect 7372 27700 7604 27740
rect 7939 27700 7948 27740
rect 7988 27700 11404 27740
rect 11444 27700 11453 27740
rect 4108 27656 4148 27700
rect 7372 27656 7412 27700
rect 1891 27616 1900 27656
rect 1940 27616 2131 27656
rect 2171 27616 2180 27656
rect 2371 27616 2380 27656
rect 2420 27616 2429 27656
rect 4099 27616 4108 27656
rect 4148 27616 4157 27656
rect 5740 27616 7412 27656
rect 2380 27572 2420 27616
rect 3724 27572 3764 27581
rect 5740 27572 5780 27616
rect 7468 27572 7508 27581
rect 355 27532 364 27572
rect 404 27532 1171 27572
rect 1211 27532 1220 27572
rect 2317 27532 2326 27572
rect 2366 27532 2420 27572
rect 2467 27532 2476 27572
rect 2516 27532 2525 27572
rect 2851 27532 2860 27572
rect 2900 27532 3724 27572
rect 4457 27532 4492 27572
rect 4532 27532 4588 27572
rect 4628 27532 4637 27572
rect 6211 27532 6220 27572
rect 6260 27532 6269 27572
rect 7171 27532 7180 27572
rect 7220 27532 7468 27572
rect 7564 27572 7604 27700
rect 7747 27616 7756 27656
rect 7796 27616 8140 27656
rect 8180 27616 8189 27656
rect 8908 27572 8948 27700
rect 10156 27572 10196 27581
rect 7564 27532 8371 27572
rect 8411 27532 8420 27572
rect 8899 27532 8908 27572
rect 8948 27532 8957 27572
rect 10051 27532 10060 27572
rect 10100 27532 10156 27572
rect 10196 27532 10231 27572
rect 0 27488 90 27508
rect 2476 27488 2516 27532
rect 3724 27488 3764 27532
rect 5740 27488 5780 27532
rect 0 27448 1036 27488
rect 1076 27448 1085 27488
rect 1987 27448 1996 27488
rect 2036 27448 2900 27488
rect 3724 27448 5780 27488
rect 0 27428 90 27448
rect 2860 27404 2900 27448
rect 6220 27404 6260 27532
rect 7468 27523 7508 27532
rect 10156 27523 10196 27532
rect 7651 27448 7660 27488
rect 7700 27448 8140 27488
rect 8180 27448 8189 27488
rect 8332 27448 9676 27488
rect 9716 27448 9725 27488
rect 1363 27364 1372 27404
rect 1412 27364 1420 27404
rect 1460 27364 1543 27404
rect 1786 27364 1795 27404
rect 1835 27364 2284 27404
rect 2324 27364 2333 27404
rect 2860 27364 6028 27404
rect 6068 27364 6260 27404
rect 7930 27364 7939 27404
rect 7979 27364 7988 27404
rect 8105 27364 8227 27404
rect 8276 27364 8285 27404
rect 7948 27320 7988 27364
rect 8332 27320 8372 27448
rect 8563 27364 8572 27404
rect 8612 27364 10348 27404
rect 10388 27364 10397 27404
rect 1708 27280 2860 27320
rect 2900 27280 2909 27320
rect 5635 27280 5644 27320
rect 5684 27280 7084 27320
rect 7124 27280 7133 27320
rect 7948 27280 8372 27320
rect 0 27152 90 27172
rect 0 27112 1324 27152
rect 1364 27112 1373 27152
rect 0 27092 90 27112
rect 1708 27068 1748 27280
rect 4291 27196 4300 27236
rect 4340 27196 4436 27236
rect 4919 27196 4928 27236
rect 4968 27196 5010 27236
rect 5050 27196 5092 27236
rect 5132 27196 5174 27236
rect 5214 27196 5256 27236
rect 5296 27196 5305 27236
rect 4396 27152 4436 27196
rect 11750 27152 11840 27172
rect 1795 27112 1804 27152
rect 1844 27112 3039 27152
rect 4396 27112 7180 27152
rect 7220 27112 7229 27152
rect 11491 27112 11500 27152
rect 11540 27112 11840 27152
rect 1699 27028 1708 27068
rect 1748 27028 1757 27068
rect 2131 27028 2140 27068
rect 2180 27028 2668 27068
rect 2708 27028 2717 27068
rect 2999 26984 3039 27112
rect 3091 27028 3100 27068
rect 3140 27028 3532 27068
rect 3572 27028 3581 27068
rect 4553 27028 4684 27068
rect 4724 27028 4733 27068
rect 2611 26944 2620 26984
rect 2660 26944 2860 26984
rect 2900 26944 2909 26984
rect 2999 26944 4492 26984
rect 4532 26944 4541 26984
rect 3244 26900 3284 26944
rect 1097 26891 1228 26900
rect 1097 26860 1219 26891
rect 1268 26860 1277 26900
rect 1865 26891 1996 26900
rect 1865 26860 1987 26891
rect 2036 26860 2045 26900
rect 2441 26891 2572 26900
rect 2441 26860 2467 26891
rect 1210 26851 1219 26860
rect 1259 26851 1268 26860
rect 1210 26850 1268 26851
rect 1978 26851 1987 26860
rect 2027 26851 2036 26860
rect 1978 26850 2036 26851
rect 2458 26851 2467 26860
rect 2507 26860 2572 26891
rect 2612 26860 2900 26900
rect 2947 26860 2956 26900
rect 2996 26860 3127 26900
rect 3235 26860 3244 26900
rect 3284 26860 3293 26900
rect 4492 26891 4532 26900
rect 2507 26851 2516 26860
rect 2458 26850 2516 26851
rect 0 26816 90 26836
rect 0 26776 268 26816
rect 308 26776 317 26816
rect 1363 26776 1372 26816
rect 1412 26776 1748 26816
rect 0 26756 90 26776
rect 1708 26648 1748 26776
rect 2476 26732 2516 26850
rect 1795 26692 1804 26732
rect 1844 26692 2516 26732
rect 2860 26732 2900 26860
rect 4579 26860 4588 26900
rect 4628 26860 4876 26900
rect 4916 26860 4972 26900
rect 5012 26860 5021 26900
rect 6124 26891 6164 27112
rect 11750 27092 11840 27112
rect 6499 27028 6508 27068
rect 6548 27028 6740 27068
rect 8323 27028 8332 27068
rect 8372 27028 8381 27068
rect 6307 26944 6316 26984
rect 6356 26944 6644 26984
rect 6604 26900 6644 26944
rect 6700 26900 6740 27028
rect 8332 26900 8372 27028
rect 4492 26816 4532 26851
rect 6586 26860 6595 26900
rect 6635 26860 6644 26900
rect 6691 26860 6700 26900
rect 6740 26860 6749 26900
rect 6953 26860 7084 26900
rect 7124 26860 7133 26900
rect 7363 26860 7372 26900
rect 7412 26891 7700 26900
rect 7412 26860 7660 26891
rect 6124 26816 6164 26851
rect 8009 26860 8140 26900
rect 8180 26860 8189 26900
rect 8332 26891 8564 26900
rect 8332 26860 8515 26891
rect 7660 26842 7700 26851
rect 8140 26842 8180 26851
rect 8506 26851 8515 26860
rect 8555 26851 8564 26891
rect 8803 26860 8812 26900
rect 8852 26860 9100 26900
rect 9140 26860 9149 26900
rect 10217 26860 10348 26900
rect 10388 26860 10397 26900
rect 8506 26850 8564 26851
rect 10348 26842 10388 26851
rect 4492 26776 6164 26816
rect 7171 26776 7180 26816
rect 7220 26776 7229 26816
rect 8611 26776 8620 26816
rect 8660 26776 8668 26816
rect 8708 26776 8791 26816
rect 7180 26732 7220 26776
rect 2860 26692 4588 26732
rect 4628 26692 4637 26732
rect 7049 26692 7180 26732
rect 7220 26692 8428 26732
rect 8468 26692 8477 26732
rect 1708 26608 4684 26648
rect 4724 26608 4733 26648
rect 10409 26608 10540 26648
rect 10580 26608 10589 26648
rect 1027 26524 1036 26564
rect 1076 26524 5068 26564
rect 5108 26524 5117 26564
rect 0 26480 90 26500
rect 0 26440 1516 26480
rect 1556 26440 1565 26480
rect 3679 26440 3688 26480
rect 3728 26440 3770 26480
rect 3810 26440 3852 26480
rect 3892 26440 3934 26480
rect 3974 26440 4016 26480
rect 4056 26440 4065 26480
rect 0 26420 90 26440
rect 4684 26356 7660 26396
rect 7700 26356 7709 26396
rect 4684 26312 4724 26356
rect 2467 26272 2476 26312
rect 2516 26272 3340 26312
rect 3380 26272 3389 26312
rect 3436 26272 4300 26312
rect 4340 26272 4349 26312
rect 4627 26272 4636 26312
rect 4676 26272 4724 26312
rect 4771 26272 4780 26312
rect 4820 26272 5020 26312
rect 5060 26272 5069 26312
rect 9619 26272 9628 26312
rect 9668 26272 10636 26312
rect 10676 26272 10685 26312
rect 3436 26228 3476 26272
rect 1372 26188 3476 26228
rect 4300 26188 4724 26228
rect 5251 26188 5260 26228
rect 5300 26188 6796 26228
rect 6836 26188 6932 26228
rect 6979 26188 6988 26228
rect 7028 26188 10004 26228
rect 10195 26188 10204 26228
rect 10244 26188 11060 26228
rect 0 26144 90 26164
rect 1372 26144 1412 26188
rect 4300 26144 4340 26188
rect 0 26104 748 26144
rect 788 26104 797 26144
rect 1363 26104 1372 26144
rect 1412 26104 1421 26144
rect 1891 26104 1900 26144
rect 1940 26104 2572 26144
rect 2612 26104 2900 26144
rect 3667 26104 3676 26144
rect 3716 26104 4340 26144
rect 4387 26104 4396 26144
rect 4436 26104 4445 26144
rect 0 26084 90 26104
rect 2860 26060 2900 26104
rect 3052 26060 3092 26069
rect 643 26020 652 26060
rect 692 26020 1171 26060
rect 1211 26020 1220 26060
rect 1795 26020 1804 26060
rect 1844 26020 1996 26060
rect 2036 26020 2045 26060
rect 2860 26020 3052 26060
rect 3331 26020 3340 26060
rect 3380 26020 3475 26060
rect 3515 26020 3524 26060
rect 3881 26020 3916 26060
rect 3956 26020 4012 26060
rect 4052 26020 4061 26060
rect 4169 26020 4195 26060
rect 4235 26020 4300 26060
rect 4340 26020 4349 26060
rect 3052 26011 3092 26020
rect 4396 25976 4436 26104
rect 3148 25936 4436 25976
rect 4684 25976 4724 26188
rect 6892 26144 6932 26188
rect 9964 26144 10004 26188
rect 11020 26144 11060 26188
rect 11750 26144 11840 26164
rect 4771 26104 4780 26144
rect 4820 26104 5068 26144
rect 5108 26104 5117 26144
rect 5443 26104 5452 26144
rect 5492 26104 5932 26144
rect 5972 26104 5981 26144
rect 6307 26104 6316 26144
rect 6356 26104 6700 26144
rect 6740 26104 6749 26144
rect 6883 26104 6892 26144
rect 6932 26104 6941 26144
rect 7555 26104 7564 26144
rect 7604 26104 9044 26144
rect 9091 26104 9100 26144
rect 9140 26104 9388 26144
rect 9428 26104 9437 26144
rect 9955 26104 9964 26144
rect 10004 26104 10013 26144
rect 10339 26104 10348 26144
rect 10388 26104 10397 26144
rect 11020 26104 11840 26144
rect 9004 26060 9044 26104
rect 4963 26020 4972 26060
rect 5012 26020 7756 26060
rect 7796 26020 7805 26060
rect 10348 26060 10388 26104
rect 11750 26084 11840 26104
rect 10348 26020 11636 26060
rect 9004 26011 9044 26020
rect 11596 25976 11636 26020
rect 4684 25936 6508 25976
rect 6548 25936 6557 25976
rect 6700 25936 7276 25976
rect 7316 25936 7468 25976
rect 7508 25936 7517 25976
rect 10579 25936 10588 25976
rect 10628 25936 11404 25976
rect 11444 25936 11453 25976
rect 11596 25936 11692 25976
rect 11732 25936 11741 25976
rect 3148 25892 3188 25936
rect 6700 25892 6740 25936
rect 1516 25852 3188 25892
rect 3235 25852 3244 25892
rect 3284 25852 3820 25892
rect 3860 25852 3869 25892
rect 3977 25852 4108 25892
rect 4148 25852 4157 25892
rect 5129 25852 5251 25892
rect 5300 25852 5309 25892
rect 5644 25852 5731 25892
rect 5771 25852 5780 25892
rect 6106 25852 6115 25892
rect 6155 25852 6164 25892
rect 6682 25852 6691 25892
rect 6731 25852 6740 25892
rect 7258 25852 7267 25892
rect 7307 25852 7316 25892
rect 7546 25852 7555 25892
rect 7595 25852 7948 25892
rect 7988 25852 7997 25892
rect 9187 25852 9196 25892
rect 9236 25852 9484 25892
rect 9524 25852 9533 25892
rect 0 25808 90 25828
rect 1516 25808 1556 25852
rect 5644 25808 5684 25852
rect 6124 25808 6164 25852
rect 7276 25808 7316 25852
rect 0 25768 1556 25808
rect 2275 25768 2284 25808
rect 2324 25768 5684 25808
rect 5731 25768 5740 25808
rect 5780 25768 6892 25808
rect 6932 25768 6941 25808
rect 7276 25768 7756 25808
rect 7796 25768 9580 25808
rect 9620 25768 9629 25808
rect 0 25748 90 25768
rect 5644 25724 5684 25768
rect 4919 25684 4928 25724
rect 4968 25684 5010 25724
rect 5050 25684 5092 25724
rect 5132 25684 5174 25724
rect 5214 25684 5256 25724
rect 5296 25684 5305 25724
rect 5644 25684 7276 25724
rect 7316 25684 7325 25724
rect 4716 25516 4732 25556
rect 4772 25516 4838 25556
rect 4878 25516 4896 25556
rect 6691 25516 6700 25556
rect 6740 25516 6892 25556
rect 6932 25516 6941 25556
rect 9667 25516 9676 25556
rect 9716 25516 9908 25556
rect 0 25472 90 25492
rect 0 25432 364 25472
rect 404 25432 413 25472
rect 3139 25432 3148 25472
rect 3188 25432 3476 25472
rect 0 25412 90 25432
rect 3436 25388 3476 25432
rect 3628 25432 4108 25472
rect 4148 25432 4157 25472
rect 4265 25432 4300 25472
rect 4340 25432 4396 25472
rect 4436 25432 4445 25472
rect 7459 25432 7468 25472
rect 7508 25432 7517 25472
rect 3628 25388 3668 25432
rect 7468 25388 7508 25432
rect 9868 25388 9908 25516
rect 1219 25348 1228 25388
rect 1268 25348 1804 25388
rect 1844 25348 1853 25388
rect 2441 25379 2572 25388
rect 2441 25348 2476 25379
rect 2516 25348 2572 25379
rect 2612 25348 2621 25388
rect 2825 25348 2947 25388
rect 2996 25348 3005 25388
rect 3139 25348 3148 25388
rect 3188 25348 3244 25388
rect 3284 25348 3319 25388
rect 3427 25348 3436 25388
rect 3476 25348 3485 25388
rect 3552 25348 3561 25388
rect 3601 25348 3668 25388
rect 3715 25348 3724 25388
rect 3764 25348 3820 25388
rect 3860 25348 3895 25388
rect 4003 25348 4012 25388
rect 4052 25348 4061 25388
rect 4265 25348 4291 25388
rect 4331 25348 4396 25388
rect 4436 25348 4445 25388
rect 4954 25348 4963 25388
rect 5003 25348 5012 25388
rect 2476 25330 2516 25339
rect 4012 25304 4052 25348
rect 4972 25304 5012 25348
rect 5068 25379 5500 25388
rect 5108 25348 5500 25379
rect 5540 25348 5549 25388
rect 5635 25348 5644 25388
rect 5684 25348 5693 25388
rect 5897 25348 6028 25388
rect 6068 25348 6077 25388
rect 7276 25379 7316 25388
rect 5068 25330 5108 25339
rect 5644 25304 5684 25348
rect 3907 25264 3916 25304
rect 3956 25264 4052 25304
rect 4099 25264 4108 25304
rect 4148 25264 5012 25304
rect 5347 25264 5356 25304
rect 5396 25264 5684 25304
rect 7468 25348 7939 25388
rect 7979 25348 7988 25388
rect 8035 25348 8044 25388
rect 8084 25348 8093 25388
rect 8323 25348 8332 25388
rect 8372 25348 8428 25388
rect 8468 25348 8503 25388
rect 9004 25379 9044 25388
rect 7276 25304 7316 25339
rect 8044 25304 8084 25348
rect 9353 25348 9484 25388
rect 9524 25348 9533 25388
rect 9850 25379 9908 25388
rect 7276 25264 7564 25304
rect 7604 25264 7613 25304
rect 7939 25264 7948 25304
rect 7988 25264 8084 25304
rect 8393 25264 8524 25304
rect 8564 25264 8573 25304
rect 5356 25220 5396 25264
rect 9004 25220 9044 25339
rect 9484 25330 9524 25339
rect 9850 25339 9859 25379
rect 9899 25339 9908 25379
rect 10003 25348 10012 25388
rect 10052 25348 10348 25388
rect 10388 25348 10397 25388
rect 9850 25338 9908 25339
rect 10339 25264 10348 25304
rect 10388 25264 11596 25304
rect 11636 25264 11645 25304
rect 2275 25180 2284 25220
rect 2324 25180 2668 25220
rect 2708 25180 5396 25220
rect 7363 25180 7372 25220
rect 7412 25180 8716 25220
rect 8756 25180 9044 25220
rect 0 25136 90 25156
rect 11750 25136 11840 25156
rect 0 25096 1228 25136
rect 1268 25096 1277 25136
rect 3427 25096 3436 25136
rect 3476 25096 3485 25136
rect 5347 25096 5356 25136
rect 5396 25096 5405 25136
rect 10579 25096 10588 25136
rect 10628 25096 11840 25136
rect 0 25076 90 25096
rect 0 24800 90 24820
rect 0 24760 652 24800
rect 692 24760 701 24800
rect 2659 24760 2668 24800
rect 2708 24760 2956 24800
rect 2996 24760 3005 24800
rect 0 24740 90 24760
rect 2476 24548 2516 24557
rect 3436 24548 3476 25096
rect 3679 24928 3688 24968
rect 3728 24928 3770 24968
rect 3810 24928 3852 24968
rect 3892 24928 3934 24968
rect 3974 24928 4016 24968
rect 4056 24928 4065 24968
rect 5356 24716 5396 25096
rect 11750 25076 11840 25096
rect 7171 24844 7180 24884
rect 7220 24844 8140 24884
rect 8180 24844 8189 24884
rect 3628 24676 5396 24716
rect 5452 24760 7508 24800
rect 3628 24632 3668 24676
rect 5452 24632 5492 24760
rect 6019 24676 6028 24716
rect 6068 24676 6077 24716
rect 3610 24592 3619 24632
rect 3659 24592 3668 24632
rect 3811 24592 3820 24632
rect 3860 24592 4323 24632
rect 4363 24592 4372 24632
rect 4579 24592 4588 24632
rect 4628 24592 5492 24632
rect 5836 24548 5876 24557
rect 6028 24548 6068 24676
rect 7468 24632 7508 24760
rect 10531 24676 10540 24716
rect 10580 24676 11692 24716
rect 11732 24676 11741 24716
rect 6787 24592 6796 24632
rect 6836 24592 7084 24632
rect 7124 24592 7133 24632
rect 7468 24592 8380 24632
rect 8420 24592 8429 24632
rect 7372 24548 7412 24557
rect 10348 24548 10388 24557
rect 835 24508 844 24548
rect 884 24508 1228 24548
rect 1268 24508 1996 24548
rect 2036 24508 2045 24548
rect 2371 24508 2380 24548
rect 2420 24508 2476 24548
rect 2516 24508 2551 24548
rect 2921 24508 3052 24548
rect 3092 24508 3101 24548
rect 3185 24508 3194 24548
rect 3234 24508 3244 24548
rect 3284 24508 3374 24548
rect 3436 24508 3496 24548
rect 3536 24508 3545 24548
rect 3595 24508 3724 24548
rect 3764 24508 3773 24548
rect 3820 24508 4204 24548
rect 4244 24508 4253 24548
rect 4387 24508 4396 24548
rect 4461 24508 4567 24548
rect 4611 24508 4628 24548
rect 4668 24508 4677 24548
rect 5801 24508 5836 24548
rect 5876 24508 5932 24548
rect 5972 24508 5981 24548
rect 6028 24508 6307 24548
rect 6347 24508 6356 24548
rect 6403 24508 6412 24548
rect 6452 24508 6836 24548
rect 6883 24508 6892 24548
rect 6932 24508 7172 24548
rect 7241 24508 7372 24548
rect 7412 24508 7421 24548
rect 7738 24508 7852 24548
rect 7900 24508 7918 24548
rect 8074 24508 8083 24548
rect 8123 24508 8179 24548
rect 8219 24508 8263 24548
rect 9091 24508 9100 24548
rect 9140 24508 9388 24548
rect 9428 24508 10060 24548
rect 10100 24508 10109 24548
rect 10243 24508 10252 24548
rect 10292 24508 10348 24548
rect 10388 24508 10828 24548
rect 10868 24508 10877 24548
rect 2476 24499 2516 24508
rect 0 24464 90 24484
rect 3052 24464 3092 24508
rect 3595 24464 3635 24508
rect 0 24424 652 24464
rect 692 24424 701 24464
rect 3052 24424 3635 24464
rect 0 24404 90 24424
rect 3820 24380 3860 24508
rect 4611 24464 4651 24508
rect 5836 24499 5876 24508
rect 4483 24424 4492 24464
rect 4532 24424 4651 24464
rect 6796 24464 6836 24508
rect 7132 24464 7172 24508
rect 7372 24499 7412 24508
rect 10348 24499 10388 24508
rect 6796 24424 6988 24464
rect 7028 24424 7037 24464
rect 7132 24424 7180 24464
rect 7220 24424 7229 24464
rect 8227 24424 8236 24464
rect 8276 24424 8716 24464
rect 8756 24424 8765 24464
rect 2537 24340 2572 24380
rect 2612 24340 2668 24380
rect 2708 24340 2717 24380
rect 3331 24340 3340 24380
rect 3380 24340 3860 24380
rect 3907 24340 3916 24380
rect 3956 24340 4108 24380
rect 4148 24340 4157 24380
rect 4919 24172 4928 24212
rect 4968 24172 5010 24212
rect 5050 24172 5092 24212
rect 5132 24172 5174 24212
rect 5214 24172 5256 24212
rect 5296 24172 5305 24212
rect 0 24128 90 24148
rect 11750 24128 11840 24148
rect 0 24088 748 24128
rect 788 24088 797 24128
rect 5164 24088 6028 24128
rect 6068 24088 6796 24128
rect 6836 24088 6845 24128
rect 11395 24088 11404 24128
rect 11444 24088 11840 24128
rect 0 24068 90 24088
rect 5164 24044 5204 24088
rect 11750 24068 11840 24088
rect 1420 24004 2572 24044
rect 2612 24004 2621 24044
rect 3235 24004 3244 24044
rect 3284 24004 4012 24044
rect 4052 24004 4061 24044
rect 4387 24004 4396 24044
rect 4436 24004 4780 24044
rect 4820 24004 4829 24044
rect 5146 24004 5155 24044
rect 5195 24004 5204 24044
rect 5609 24004 5731 24044
rect 5780 24004 6700 24044
rect 6740 24004 6749 24044
rect 7363 24004 7372 24044
rect 7412 24004 7852 24044
rect 7892 24004 7901 24044
rect 8410 24004 8419 24044
rect 8459 24004 9004 24044
rect 9044 24004 9053 24044
rect 1420 23876 1460 24004
rect 1577 23920 1708 23960
rect 1748 23920 1757 23960
rect 2237 23920 2284 23960
rect 2324 23920 2333 23960
rect 2380 23920 3052 23960
rect 3092 23920 3101 23960
rect 3244 23920 4244 23960
rect 4339 23920 4348 23960
rect 4388 23920 4972 23960
rect 5012 23920 5021 23960
rect 5923 23920 5932 23960
rect 5972 23920 7220 23960
rect 7459 23920 7468 23960
rect 7508 23920 7564 23960
rect 7604 23920 7639 23960
rect 7747 23920 7756 23960
rect 7796 23920 7852 23960
rect 7892 23920 7927 23960
rect 8611 23920 8620 23960
rect 8660 23920 9676 23960
rect 9716 23920 9964 23960
rect 10004 23920 10013 23960
rect 2284 23876 2324 23920
rect 2380 23876 2420 23920
rect 1315 23836 1324 23876
rect 1364 23836 1460 23876
rect 1507 23836 1516 23876
rect 1556 23836 1603 23876
rect 1643 23836 2092 23876
rect 2132 23836 2141 23876
rect 2266 23836 2275 23876
rect 2315 23836 2324 23876
rect 2371 23836 2380 23876
rect 2420 23836 2429 23876
rect 2476 23836 2764 23876
rect 2804 23836 2813 23876
rect 0 23792 90 23812
rect 2476 23792 2516 23836
rect 0 23752 460 23792
rect 500 23752 509 23792
rect 1996 23752 2516 23792
rect 2851 23752 2860 23792
rect 2900 23752 2956 23792
rect 2996 23752 3031 23792
rect 0 23732 90 23752
rect 1996 23708 2036 23752
rect 3244 23708 3284 23920
rect 4204 23876 4244 23920
rect 3339 23867 3476 23876
rect 3379 23836 3476 23867
rect 3339 23818 3379 23827
rect 1987 23668 1996 23708
rect 2036 23668 2045 23708
rect 2860 23668 3284 23708
rect 1699 23584 1708 23624
rect 1748 23584 2284 23624
rect 2324 23584 2333 23624
rect 0 23456 90 23476
rect 2860 23456 2900 23668
rect 0 23416 2900 23456
rect 0 23396 90 23416
rect 3436 23288 3476 23836
rect 3820 23867 3860 23876
rect 3820 23792 3860 23827
rect 4186 23867 4244 23876
rect 4186 23827 4195 23867
rect 4235 23827 4244 23867
rect 4637 23836 4684 23876
rect 4724 23836 4733 23876
rect 4867 23836 4876 23876
rect 4916 23836 5356 23876
rect 5396 23836 5405 23876
rect 5923 23836 5932 23876
rect 5972 23836 6124 23876
rect 6164 23836 6173 23876
rect 7180 23867 7220 23920
rect 4186 23826 4244 23827
rect 4684 23792 4724 23836
rect 8611 23836 8620 23876
rect 8660 23867 9580 23876
rect 8660 23836 9100 23867
rect 7180 23818 7220 23827
rect 9140 23836 9580 23867
rect 9620 23836 9629 23876
rect 10051 23836 10060 23876
rect 10100 23836 10348 23876
rect 10388 23836 10397 23876
rect 9100 23818 9140 23827
rect 3820 23752 4108 23792
rect 4148 23752 4157 23792
rect 4675 23752 4684 23792
rect 4724 23752 4733 23792
rect 5251 23752 5260 23792
rect 5300 23752 5356 23792
rect 5396 23752 5431 23792
rect 8323 23752 8332 23792
rect 8372 23752 8381 23792
rect 8332 23708 8372 23752
rect 5059 23668 5068 23708
rect 5108 23668 7468 23708
rect 7508 23668 7517 23708
rect 8332 23668 8620 23708
rect 8660 23668 8669 23708
rect 7747 23584 7756 23624
rect 7796 23584 8044 23624
rect 8084 23584 8093 23624
rect 8899 23584 8908 23624
rect 8948 23584 8957 23624
rect 3679 23416 3688 23456
rect 3728 23416 3770 23456
rect 3810 23416 3852 23456
rect 3892 23416 3934 23456
rect 3974 23416 4016 23456
rect 4056 23416 4065 23456
rect 7747 23416 7756 23456
rect 7796 23416 8428 23456
rect 8468 23416 8477 23456
rect 8908 23288 8948 23584
rect 3427 23248 3436 23288
rect 3476 23248 3485 23288
rect 4195 23248 4204 23288
rect 4244 23248 4253 23288
rect 5779 23248 5788 23288
rect 5828 23248 6028 23288
rect 6068 23248 6077 23288
rect 8092 23248 8948 23288
rect 4204 23204 4244 23248
rect 652 23164 1460 23204
rect 0 23120 90 23140
rect 652 23120 692 23164
rect 1420 23120 1460 23164
rect 3709 23164 4244 23204
rect 5059 23164 5068 23204
rect 5108 23164 5356 23204
rect 5396 23164 5405 23204
rect 0 23080 692 23120
rect 739 23080 748 23120
rect 788 23080 1364 23120
rect 1420 23080 3380 23120
rect 0 23060 90 23080
rect 1324 23036 1364 23080
rect 3340 23036 3380 23080
rect 643 22996 652 23036
rect 692 22996 1171 23036
rect 1211 22996 1220 23036
rect 1324 22996 1666 23036
rect 1706 22996 1715 23036
rect 1987 22996 1996 23036
rect 2036 22996 2146 23036
rect 2186 22996 2195 23036
rect 2563 22996 2572 23036
rect 2612 22996 2764 23036
rect 2804 22996 2813 23036
rect 3034 22996 3043 23036
rect 3083 22996 3244 23036
rect 3284 22996 3293 23036
rect 3340 22996 3586 23036
rect 3626 22996 3635 23036
rect 1996 22952 2036 22996
rect 3709 22952 3749 23164
rect 8092 23120 8132 23248
rect 8611 23164 8620 23204
rect 8660 23164 10100 23204
rect 4003 23080 4012 23120
rect 4052 23080 4876 23120
rect 4916 23080 5300 23120
rect 6115 23080 6124 23120
rect 6164 23080 6295 23120
rect 6403 23080 6412 23120
rect 6452 23080 6604 23120
rect 6644 23080 6653 23120
rect 8044 23080 8132 23120
rect 8419 23080 8428 23120
rect 8468 23080 8524 23120
rect 8564 23080 8599 23120
rect 5260 23036 5300 23080
rect 8044 23036 8084 23080
rect 9100 23036 9140 23045
rect 10060 23036 10100 23164
rect 11750 23120 11840 23140
rect 10627 23080 10636 23120
rect 10676 23080 11840 23120
rect 11750 23060 11840 23080
rect 4012 22996 4066 23036
rect 4106 22996 4115 23036
rect 4387 22996 4396 23036
rect 4436 22996 4588 23036
rect 4628 22996 4637 23036
rect 4867 22996 4876 23036
rect 4916 22996 5068 23036
rect 5108 22996 5117 23036
rect 5251 22996 5260 23036
rect 5300 22996 5309 23036
rect 5513 22996 5644 23036
rect 5684 22996 5693 23036
rect 6967 22996 6976 23036
rect 7016 22996 7028 23036
rect 7123 22996 7132 23036
rect 7172 22996 7468 23036
rect 7508 22996 7517 23036
rect 8026 22996 8035 23036
rect 8075 22996 8084 23036
rect 8131 22996 8140 23036
rect 8180 22996 8189 23036
rect 8323 22996 8332 23036
rect 8372 22996 8620 23036
rect 8660 22996 8669 23036
rect 8995 22996 9004 23036
rect 9044 22996 9100 23036
rect 9140 22996 9196 23036
rect 9236 22996 9300 23036
rect 9610 22996 9619 23036
rect 9659 22996 9716 23036
rect 4012 22952 4052 22996
rect 5068 22952 5108 22996
rect 6988 22952 7028 22996
rect 1123 22912 1132 22952
rect 1172 22912 2036 22952
rect 2083 22912 2092 22952
rect 2132 22912 2332 22952
rect 2372 22912 2381 22952
rect 3139 22912 3148 22952
rect 3188 22912 3340 22952
rect 3380 22912 3749 22952
rect 4003 22912 4012 22952
rect 4052 22912 4061 22952
rect 5068 22912 5452 22952
rect 5492 22912 5501 22952
rect 6988 22912 7180 22952
rect 7220 22912 7229 22952
rect 1363 22828 1372 22868
rect 1412 22828 1708 22868
rect 1748 22828 1757 22868
rect 1843 22828 1852 22868
rect 1892 22828 3052 22868
rect 3092 22828 3101 22868
rect 3715 22828 3724 22868
rect 3764 22828 3772 22868
rect 3812 22828 3895 22868
rect 4243 22828 4252 22868
rect 4292 22828 4436 22868
rect 4666 22828 4675 22868
rect 4715 22828 4780 22868
rect 4820 22828 4855 22868
rect 4963 22828 4972 22868
rect 5012 22828 5492 22868
rect 5731 22828 5740 22868
rect 5780 22828 5884 22868
rect 5924 22828 5933 22868
rect 6211 22828 6220 22868
rect 6260 22828 6403 22868
rect 6443 22828 6452 22868
rect 6691 22828 6700 22868
rect 6740 22828 7555 22868
rect 7595 22828 7852 22868
rect 7892 22828 7901 22868
rect 0 22784 90 22804
rect 0 22744 1228 22784
rect 1268 22744 1277 22784
rect 0 22724 90 22744
rect 4396 22700 4436 22828
rect 5452 22700 5492 22828
rect 6412 22784 6452 22828
rect 6412 22744 6508 22784
rect 6548 22744 6557 22784
rect 8140 22700 8180 22996
rect 9100 22987 9140 22996
rect 4387 22660 4396 22700
rect 4436 22660 4445 22700
rect 4919 22660 4928 22700
rect 4968 22660 5010 22700
rect 5050 22660 5092 22700
rect 5132 22660 5174 22700
rect 5214 22660 5256 22700
rect 5296 22660 5305 22700
rect 5443 22660 5452 22700
rect 5492 22660 8180 22700
rect 9676 22532 9716 22996
rect 9868 22996 9907 23036
rect 9947 22996 9956 23036
rect 10060 22996 10444 23036
rect 10484 22996 10493 23036
rect 9868 22868 9908 22996
rect 9763 22828 9772 22868
rect 9812 22828 9908 22868
rect 10099 22828 10108 22868
rect 10148 22828 11596 22868
rect 11636 22828 11645 22868
rect 2083 22492 2092 22532
rect 2132 22492 2860 22532
rect 2900 22492 2909 22532
rect 5731 22492 5740 22532
rect 5780 22492 6124 22532
rect 6164 22492 6173 22532
rect 7555 22492 7564 22532
rect 7604 22492 7747 22532
rect 7787 22492 7796 22532
rect 7913 22492 8035 22532
rect 8084 22492 8093 22532
rect 9676 22492 9868 22532
rect 9908 22492 9917 22532
rect 10505 22492 10588 22532
rect 10628 22492 10636 22532
rect 10676 22492 10685 22532
rect 0 22448 90 22468
rect 0 22408 76 22448
rect 116 22408 125 22448
rect 2659 22408 2668 22448
rect 2708 22408 4052 22448
rect 5251 22408 5260 22448
rect 5300 22408 10732 22448
rect 10772 22408 10781 22448
rect 0 22388 90 22408
rect 4012 22364 4052 22408
rect 1219 22324 1228 22364
rect 1268 22324 1804 22364
rect 1844 22324 1996 22364
rect 2036 22324 2045 22364
rect 2476 22355 2516 22364
rect 2563 22324 2572 22364
rect 2612 22324 3148 22364
rect 3188 22324 3197 22364
rect 3244 22324 3257 22364
rect 3297 22324 3306 22364
rect 3401 22324 3532 22364
rect 3572 22324 3581 22364
rect 3994 22324 4003 22364
rect 4043 22324 4052 22364
rect 4099 22324 4108 22364
rect 4148 22324 4157 22364
rect 4483 22324 4492 22364
rect 4532 22324 5012 22364
rect 5059 22324 5068 22364
rect 5108 22324 5239 22364
rect 5548 22355 6164 22364
rect 2476 22280 2516 22315
rect 3244 22280 3284 22324
rect 4108 22280 4148 22324
rect 2476 22240 2668 22280
rect 2708 22240 2717 22280
rect 2851 22240 2860 22280
rect 2900 22240 3284 22280
rect 3595 22240 4148 22280
rect 4291 22240 4300 22280
rect 4340 22240 4588 22280
rect 4628 22240 4637 22280
rect 2851 22156 2860 22196
rect 2900 22156 2956 22196
rect 2996 22156 3031 22196
rect 0 22112 90 22132
rect 0 22072 556 22112
rect 596 22072 605 22112
rect 0 22052 90 22072
rect 0 21776 90 21796
rect 0 21736 364 21776
rect 404 21736 413 21776
rect 2659 21736 2668 21776
rect 2708 21736 2764 21776
rect 2804 21736 2839 21776
rect 0 21716 90 21736
rect 2999 21652 3436 21692
rect 3476 21652 3485 21692
rect 2999 21608 3039 21652
rect 3595 21608 3635 22240
rect 4972 22196 5012 22324
rect 5068 22306 5108 22315
rect 5588 22324 6164 22355
rect 5548 22306 5588 22315
rect 6124 22280 6164 22324
rect 6106 22240 6115 22280
rect 6155 22240 6164 22280
rect 6220 22355 6356 22364
rect 6220 22324 6316 22355
rect 6220 22196 6260 22324
rect 6595 22324 6604 22364
rect 6644 22324 7084 22364
rect 7124 22324 7564 22364
rect 7604 22324 7613 22364
rect 8035 22324 8044 22364
rect 8084 22324 8428 22364
rect 8468 22324 8477 22364
rect 9571 22324 9580 22364
rect 9620 22355 9751 22364
rect 9620 22324 9676 22355
rect 6316 22306 6356 22315
rect 9716 22324 9751 22355
rect 9676 22306 9716 22315
rect 10051 22240 10060 22280
rect 10100 22240 10109 22280
rect 10339 22240 10348 22280
rect 10388 22240 11404 22280
rect 11444 22240 11453 22280
rect 10060 22196 10100 22240
rect 4841 22156 4972 22196
rect 5012 22156 5452 22196
rect 5492 22156 5501 22196
rect 6115 22156 6124 22196
rect 6164 22156 6260 22196
rect 7555 22156 7564 22196
rect 7604 22156 10100 22196
rect 11750 22112 11840 22132
rect 3715 22072 3724 22112
rect 3764 22072 4300 22112
rect 4340 22072 4349 22112
rect 10588 22072 11840 22112
rect 3679 21904 3688 21944
rect 3728 21904 3770 21944
rect 3810 21904 3852 21944
rect 3892 21904 3934 21944
rect 3974 21904 4016 21944
rect 4056 21904 4065 21944
rect 5635 21820 5644 21860
rect 5684 21820 8756 21860
rect 8716 21776 8756 21820
rect 10588 21776 10628 22072
rect 11750 22052 11840 22072
rect 8707 21736 8716 21776
rect 8756 21736 8765 21776
rect 10579 21736 10588 21776
rect 10628 21736 10637 21776
rect 5059 21652 5068 21692
rect 5108 21652 5117 21692
rect 5932 21652 6356 21692
rect 1363 21568 1372 21608
rect 1412 21568 1900 21608
rect 1940 21568 1949 21608
rect 1996 21568 3039 21608
rect 3427 21568 3436 21608
rect 3476 21568 3628 21608
rect 3668 21568 3677 21608
rect 3881 21568 4012 21608
rect 4052 21568 4972 21608
rect 5012 21568 5021 21608
rect 1996 21524 2036 21568
rect 2956 21524 2996 21568
rect 4012 21524 4052 21568
rect 5068 21524 5108 21652
rect 5155 21568 5164 21608
rect 5204 21568 5396 21608
rect 5356 21524 5396 21568
rect 5932 21524 5972 21652
rect 6316 21608 6356 21652
rect 6316 21568 6691 21608
rect 6731 21568 6740 21608
rect 8201 21568 8332 21608
rect 8372 21568 8381 21608
rect 10217 21568 10348 21608
rect 10388 21568 10397 21608
rect 6019 21526 6028 21566
rect 6068 21526 6199 21566
rect 451 21484 460 21524
rect 500 21484 1171 21524
rect 1211 21484 1220 21524
rect 1987 21484 1996 21524
rect 2036 21484 2045 21524
rect 2153 21484 2275 21524
rect 2324 21484 2333 21524
rect 2938 21484 2947 21524
rect 2987 21484 2996 21524
rect 3043 21484 3052 21524
rect 3092 21484 3476 21524
rect 3523 21484 3532 21524
rect 3572 21484 3581 21524
rect 4099 21484 4108 21524
rect 4148 21484 4500 21524
rect 4540 21484 4549 21524
rect 4963 21484 4972 21524
rect 5012 21484 5021 21524
rect 5068 21484 5227 21524
rect 5267 21484 5276 21524
rect 5338 21484 5347 21524
rect 5387 21484 5396 21524
rect 5443 21484 5452 21524
rect 5492 21484 5923 21524
rect 5963 21484 5972 21524
rect 6892 21524 6932 21533
rect 8908 21524 8948 21533
rect 6028 21508 6068 21517
rect 6595 21484 6604 21524
rect 6644 21484 6892 21524
rect 8035 21484 8044 21524
rect 8084 21484 8140 21524
rect 8180 21484 8215 21524
rect 10025 21484 10060 21524
rect 10100 21484 10156 21524
rect 10196 21484 10205 21524
rect 0 21440 90 21460
rect 0 21400 652 21440
rect 692 21400 701 21440
rect 2371 21400 2380 21440
rect 2420 21400 2668 21440
rect 2708 21400 2717 21440
rect 0 21380 90 21400
rect 3436 21272 3476 21484
rect 3532 21356 3572 21484
rect 4012 21475 4052 21484
rect 4972 21440 5012 21484
rect 6892 21440 6932 21484
rect 8908 21440 8948 21484
rect 4972 21400 5644 21440
rect 5684 21400 5693 21440
rect 5827 21400 5836 21440
rect 5876 21400 6355 21440
rect 6395 21400 6404 21440
rect 6892 21400 8908 21440
rect 8948 21400 8957 21440
rect 3532 21316 4300 21356
rect 4340 21316 4349 21356
rect 4553 21316 4684 21356
rect 4724 21316 4733 21356
rect 3436 21232 3916 21272
rect 3956 21232 3965 21272
rect 4919 21148 4928 21188
rect 4968 21148 5010 21188
rect 5050 21148 5092 21188
rect 5132 21148 5174 21188
rect 5214 21148 5256 21188
rect 5296 21148 5305 21188
rect 0 21104 90 21124
rect 0 21064 268 21104
rect 308 21064 317 21104
rect 1372 21064 3628 21104
rect 3668 21064 3677 21104
rect 0 21044 90 21064
rect 1372 21020 1412 21064
rect 1363 20980 1372 21020
rect 1412 20980 1421 21020
rect 1699 20980 1708 21020
rect 1748 20980 2092 21020
rect 2132 20980 2324 21020
rect 2284 20936 2324 20980
rect 5356 20936 5396 21400
rect 5683 21316 5692 21356
rect 5732 21347 5876 21356
rect 5732 21316 5827 21347
rect 5818 21307 5827 21316
rect 5867 21307 5876 21347
rect 8563 21316 8572 21356
rect 8612 21316 8660 21356
rect 5818 21306 5876 21307
rect 8620 21104 8660 21316
rect 11750 21104 11840 21124
rect 8620 21064 11840 21104
rect 11750 21044 11840 21064
rect 5539 20980 5548 21020
rect 5588 20980 5932 21020
rect 5972 20980 5981 21020
rect 6490 20980 6499 21020
rect 6539 20980 6700 21020
rect 6740 20980 6749 21020
rect 7066 20980 7075 21020
rect 7115 20980 7852 21020
rect 7892 20980 7901 21020
rect 1507 20896 1516 20936
rect 1556 20896 1900 20936
rect 1940 20896 2228 20936
rect 2275 20896 2284 20936
rect 2324 20896 2333 20936
rect 3209 20896 3244 20936
rect 3284 20896 3340 20936
rect 3380 20896 3389 20936
rect 3820 20896 5396 20936
rect 5731 20896 5740 20936
rect 5780 20896 7276 20936
rect 7316 20896 7325 20936
rect 8716 20896 9100 20936
rect 9140 20896 9149 20936
rect 2188 20852 2228 20896
rect 3820 20852 3860 20896
rect 5932 20852 5972 20896
rect 8716 20852 8756 20896
rect 1097 20843 1228 20852
rect 1097 20812 1219 20843
rect 1268 20812 1277 20852
rect 1891 20812 1900 20852
rect 1940 20812 1949 20852
rect 2170 20812 2179 20852
rect 2219 20812 2228 20852
rect 2851 20812 2860 20852
rect 2900 20812 2909 20852
rect 3017 20812 3139 20852
rect 3188 20812 3197 20852
rect 3802 20812 3811 20852
rect 3851 20812 3860 20852
rect 3907 20812 3916 20852
rect 3956 20812 4087 20852
rect 4156 20812 4300 20852
rect 4340 20812 4349 20852
rect 4876 20843 4916 20852
rect 1210 20803 1219 20812
rect 1259 20803 1268 20812
rect 1210 20802 1268 20803
rect 0 20768 90 20788
rect 1900 20768 1940 20812
rect 2860 20768 2900 20812
rect 3820 20768 3860 20812
rect 4156 20768 4196 20812
rect 5196 20812 5260 20852
rect 5300 20843 5452 20852
rect 5300 20812 5356 20843
rect 0 20728 460 20768
rect 500 20728 509 20768
rect 1900 20728 2092 20768
rect 2132 20728 3860 20768
rect 3916 20728 4196 20768
rect 4291 20728 4300 20768
rect 4340 20728 4396 20768
rect 4436 20728 4471 20768
rect 0 20708 90 20728
rect 3916 20684 3956 20728
rect 4876 20684 4916 20803
rect 5396 20812 5452 20843
rect 5492 20812 5501 20852
rect 5635 20812 5644 20852
rect 5684 20812 5687 20852
rect 5727 20812 5815 20852
rect 5923 20812 5932 20852
rect 5972 20812 5981 20852
rect 6115 20812 6124 20852
rect 6164 20812 6167 20852
rect 6207 20812 6295 20852
rect 6403 20812 6412 20852
rect 6452 20812 6461 20852
rect 6595 20812 6604 20852
rect 6644 20843 7508 20852
rect 6644 20812 7468 20843
rect 5356 20794 5396 20803
rect 5705 20728 5827 20768
rect 5876 20728 5885 20768
rect 6019 20728 6028 20768
rect 6068 20728 6307 20768
rect 6347 20728 6356 20768
rect 6412 20684 6452 20812
rect 8707 20812 8716 20852
rect 8756 20812 8765 20852
rect 8899 20812 8908 20852
rect 8948 20843 9140 20852
rect 8948 20812 9100 20843
rect 7468 20794 7508 20803
rect 10339 20812 10348 20852
rect 10388 20812 10636 20852
rect 10676 20812 11308 20852
rect 11348 20812 11357 20852
rect 9100 20794 9140 20803
rect 6691 20728 6700 20768
rect 6740 20728 6749 20768
rect 6700 20684 6740 20728
rect 3436 20644 3628 20684
rect 3668 20644 3956 20684
rect 4003 20644 4012 20684
rect 4052 20644 4916 20684
rect 5443 20644 5452 20684
rect 5492 20644 6452 20684
rect 6499 20644 6508 20684
rect 6548 20644 6740 20684
rect 8777 20644 8908 20684
rect 8948 20644 8957 20684
rect 2563 20560 2572 20600
rect 2612 20560 3148 20600
rect 3188 20560 3197 20600
rect 3436 20516 3476 20644
rect 4876 20600 4916 20644
rect 3523 20560 3532 20600
rect 3572 20560 4108 20600
rect 4148 20560 4157 20600
rect 4876 20560 5836 20600
rect 5876 20560 5885 20600
rect 3436 20476 3626 20516
rect 0 20432 90 20452
rect 0 20392 1228 20432
rect 1268 20392 1277 20432
rect 0 20372 90 20392
rect 3586 20348 3626 20476
rect 3679 20392 3688 20432
rect 3728 20392 3770 20432
rect 3810 20392 3852 20432
rect 3892 20392 3934 20432
rect 3974 20392 4016 20432
rect 4056 20392 4065 20432
rect 3586 20308 3956 20348
rect 3916 20264 3956 20308
rect 2668 20224 2860 20264
rect 2900 20224 2909 20264
rect 3907 20224 3916 20264
rect 3956 20224 3965 20264
rect 5923 20224 5932 20264
rect 5972 20224 6124 20264
rect 6164 20224 6173 20264
rect 2668 20180 2708 20224
rect 1795 20140 1804 20180
rect 1844 20140 2708 20180
rect 2755 20140 2764 20180
rect 2804 20140 2813 20180
rect 3139 20140 3148 20180
rect 3188 20140 3572 20180
rect 5155 20140 5164 20180
rect 5204 20140 5644 20180
rect 5684 20140 5693 20180
rect 8755 20140 8764 20180
rect 8804 20140 10292 20180
rect 0 20096 90 20116
rect 2764 20096 2804 20140
rect 3532 20096 3572 20140
rect 10252 20096 10292 20140
rect 11750 20096 11840 20116
rect 0 20056 1516 20096
rect 1556 20056 1565 20096
rect 2764 20056 3401 20096
rect 3523 20056 3532 20096
rect 3572 20056 3581 20096
rect 4684 20056 5068 20096
rect 5108 20056 5117 20096
rect 5164 20056 5356 20096
rect 5396 20056 5405 20096
rect 5731 20056 5740 20096
rect 5780 20056 5789 20096
rect 8393 20056 8524 20096
rect 8564 20056 8573 20096
rect 8620 20056 9868 20096
rect 9908 20056 9917 20096
rect 10252 20056 11840 20096
rect 0 20036 90 20056
rect 3361 20012 3401 20056
rect 4108 20012 4148 20021
rect 4684 20012 4724 20056
rect 5164 20012 5204 20056
rect 5740 20012 5780 20056
rect 7852 20012 7892 20021
rect 8620 20012 8660 20056
rect 11750 20036 11840 20056
rect 10156 20012 10196 20021
rect 547 19972 556 20012
rect 596 19972 1171 20012
rect 1211 19972 1220 20012
rect 1673 19972 1804 20012
rect 1844 19972 1853 20012
rect 1961 19972 2092 20012
rect 2132 19972 2141 20012
rect 2275 19972 2284 20012
rect 2324 19972 2371 20012
rect 2411 19972 2455 20012
rect 3034 19971 3043 20011
rect 3083 19971 3092 20011
rect 3139 19972 3148 20012
rect 3188 19972 3319 20012
rect 3361 19972 3628 20012
rect 3668 19972 3677 20012
rect 3977 19972 4108 20012
rect 4148 19972 4157 20012
rect 4618 19972 4627 20012
rect 4667 19972 4724 20012
rect 4771 19972 4780 20012
rect 4820 19972 4972 20012
rect 5012 19972 5021 20012
rect 5088 19972 5097 20012
rect 5137 19972 5204 20012
rect 5251 19972 5260 20012
rect 5300 19972 5431 20012
rect 5548 19972 5596 20012
rect 5636 19972 5645 20012
rect 5731 19972 5740 20012
rect 5780 19972 5827 20012
rect 5923 19972 5932 20012
rect 5972 19972 5981 20012
rect 6115 19972 6124 20012
rect 6164 19972 6173 20012
rect 6595 19972 6604 20012
rect 6644 19972 7084 20012
rect 7124 19972 7133 20012
rect 7892 19972 8660 20012
rect 8899 19972 8908 20012
rect 8948 19972 9100 20012
rect 9140 19972 9149 20012
rect 9571 19972 9580 20012
rect 9620 19972 10156 20012
rect 1123 19888 1132 19928
rect 1172 19888 2476 19928
rect 2516 19888 2668 19928
rect 2708 19888 2717 19928
rect 1363 19804 1372 19844
rect 1412 19804 1804 19844
rect 1844 19804 1853 19844
rect 0 19760 90 19780
rect 3052 19760 3092 19971
rect 4108 19963 4148 19972
rect 5548 19928 5588 19972
rect 5932 19928 5972 19972
rect 4780 19888 5588 19928
rect 5923 19888 5932 19928
rect 5972 19888 6019 19928
rect 4780 19844 4820 19888
rect 6124 19844 6164 19972
rect 4771 19804 4780 19844
rect 4820 19804 4829 19844
rect 5321 19804 5443 19844
rect 5492 19804 5501 19844
rect 6028 19804 6164 19844
rect 6377 19804 6403 19844
rect 6443 19804 6508 19844
rect 6548 19804 6557 19844
rect 6028 19760 6068 19804
rect 0 19720 556 19760
rect 596 19720 605 19760
rect 3052 19720 5932 19760
rect 5972 19720 6068 19760
rect 0 19700 90 19720
rect 1411 19636 1420 19676
rect 1460 19636 3052 19676
rect 3092 19636 3101 19676
rect 4919 19636 4928 19676
rect 4968 19636 5010 19676
rect 5050 19636 5092 19676
rect 5132 19636 5174 19676
rect 5214 19636 5256 19676
rect 5296 19636 5305 19676
rect 1891 19552 1900 19592
rect 1940 19552 3044 19592
rect 3004 19508 3044 19552
rect 259 19468 268 19508
rect 308 19468 2900 19508
rect 3004 19468 3196 19508
rect 3236 19468 3245 19508
rect 3516 19468 3532 19508
rect 3572 19468 3676 19508
rect 3716 19468 7028 19508
rect 0 19424 90 19444
rect 2860 19424 2900 19468
rect 0 19384 940 19424
rect 980 19384 989 19424
rect 2563 19384 2572 19424
rect 2612 19384 2743 19424
rect 2860 19384 3092 19424
rect 3619 19384 3628 19424
rect 3668 19384 4532 19424
rect 4627 19384 4636 19424
rect 4676 19384 6356 19424
rect 6595 19384 6604 19424
rect 6644 19384 6653 19424
rect 0 19364 90 19384
rect 3052 19340 3092 19384
rect 4492 19340 4532 19384
rect 355 19300 364 19340
rect 404 19331 1268 19340
rect 404 19300 1219 19331
rect 1210 19291 1219 19300
rect 1259 19291 1268 19331
rect 1363 19300 1372 19340
rect 1412 19300 1420 19340
rect 1460 19300 1543 19340
rect 2092 19300 2140 19340
rect 2180 19300 2189 19340
rect 2458 19300 2467 19340
rect 2507 19300 2516 19340
rect 1210 19290 1268 19291
rect 1699 19216 1708 19256
rect 1748 19216 1996 19256
rect 2036 19216 2045 19256
rect 2092 19172 2132 19300
rect 2476 19256 2516 19300
rect 3034 19331 3092 19340
rect 3034 19291 3043 19331
rect 3083 19291 3092 19331
rect 3034 19290 3092 19291
rect 3514 19331 3724 19340
rect 3514 19291 3523 19331
rect 3563 19300 3724 19331
rect 3764 19300 3773 19340
rect 3881 19331 4012 19340
rect 3881 19300 4003 19331
rect 4052 19300 4061 19340
rect 4474 19331 4532 19340
rect 3563 19291 3572 19300
rect 3514 19290 3572 19291
rect 3994 19291 4003 19300
rect 4043 19291 4052 19300
rect 3994 19290 4052 19291
rect 4474 19291 4483 19331
rect 4523 19291 4532 19331
rect 5033 19300 5164 19340
rect 5204 19300 5213 19340
rect 4474 19290 4532 19291
rect 2476 19216 2572 19256
rect 2612 19216 2764 19256
rect 2804 19216 2813 19256
rect 4108 19216 4156 19256
rect 4196 19216 4205 19256
rect 2083 19132 2092 19172
rect 2132 19132 2141 19172
rect 2851 19132 2860 19172
rect 2900 19132 3148 19172
rect 3188 19132 3197 19172
rect 0 19088 90 19108
rect 4108 19088 4148 19216
rect 6316 19172 6356 19384
rect 6604 19340 6644 19384
rect 6988 19340 7028 19468
rect 7852 19424 7892 19972
rect 10156 19963 10196 19972
rect 7939 19888 7948 19928
rect 7988 19888 8236 19928
rect 8276 19888 8620 19928
rect 8660 19888 8669 19928
rect 8035 19804 8044 19844
rect 8084 19804 8093 19844
rect 9667 19804 9676 19844
rect 9716 19804 10348 19844
rect 10388 19804 10397 19844
rect 7084 19384 7892 19424
rect 6412 19331 6452 19340
rect 6604 19300 6883 19340
rect 6923 19300 6932 19340
rect 6979 19300 6988 19340
rect 7028 19300 7037 19340
rect 6412 19256 6452 19291
rect 7084 19256 7124 19384
rect 8044 19340 8084 19804
rect 8611 19468 8620 19508
rect 8660 19468 9868 19508
rect 9908 19468 9917 19508
rect 7363 19300 7372 19340
rect 7412 19300 7660 19340
rect 7700 19300 7709 19340
rect 7948 19331 7988 19340
rect 8044 19331 8468 19340
rect 8044 19300 8428 19331
rect 7948 19256 7988 19291
rect 8428 19282 8468 19291
rect 9292 19331 9580 19340
rect 9332 19300 9580 19331
rect 9620 19300 9629 19340
rect 10243 19300 10252 19340
rect 10292 19300 10540 19340
rect 10580 19300 10636 19340
rect 10676 19300 10685 19340
rect 9292 19282 9332 19291
rect 6412 19216 7124 19256
rect 7337 19216 7468 19256
rect 7508 19216 7517 19256
rect 7948 19216 8140 19256
rect 8180 19216 8189 19256
rect 8803 19216 8812 19256
rect 8852 19216 9100 19256
rect 9140 19216 9149 19256
rect 9100 19172 9140 19216
rect 6316 19132 7276 19172
rect 7316 19132 7325 19172
rect 9100 19132 9484 19172
rect 9524 19132 9533 19172
rect 11750 19088 11840 19108
rect 0 19048 1420 19088
rect 1460 19048 1469 19088
rect 1939 19048 1948 19088
rect 1988 19048 2036 19088
rect 2659 19048 2668 19088
rect 2708 19048 4148 19088
rect 9091 19048 9100 19088
rect 9140 19048 9149 19088
rect 10627 19048 10636 19088
rect 10676 19048 11840 19088
rect 0 19028 90 19048
rect 1996 18836 2036 19048
rect 9100 19004 9140 19048
rect 11750 19028 11840 19048
rect 7459 18964 7468 19004
rect 7508 18964 9140 19004
rect 3679 18880 3688 18920
rect 3728 18880 3770 18920
rect 3810 18880 3852 18920
rect 3892 18880 3934 18920
rect 3974 18880 4016 18920
rect 4056 18880 4065 18920
rect 1996 18796 5644 18836
rect 5684 18796 5693 18836
rect 8131 18796 8140 18836
rect 8180 18796 8660 18836
rect 0 18752 90 18772
rect 0 18712 748 18752
rect 788 18712 797 18752
rect 2275 18712 2284 18752
rect 2324 18712 3532 18752
rect 3572 18712 3581 18752
rect 4204 18712 4820 18752
rect 7315 18712 7324 18752
rect 7364 18712 8524 18752
rect 8564 18712 8573 18752
rect 0 18692 90 18712
rect 1411 18628 1420 18668
rect 1460 18628 3956 18668
rect 1363 18544 1372 18584
rect 1412 18544 1708 18584
rect 1748 18544 1757 18584
rect 1891 18544 1900 18584
rect 1940 18544 2476 18584
rect 2516 18544 2525 18584
rect 3916 18542 3956 18628
rect 4204 18584 4244 18712
rect 4780 18668 4820 18712
rect 4339 18628 4348 18668
rect 4388 18628 4684 18668
rect 4724 18628 4733 18668
rect 4780 18628 6700 18668
rect 6740 18628 7412 18668
rect 4051 18544 4060 18584
rect 4100 18544 4244 18584
rect 4579 18544 4588 18584
rect 4628 18544 4637 18584
rect 4963 18544 4972 18584
rect 5012 18544 5021 18584
rect 6953 18544 7084 18584
rect 7124 18544 7133 18584
rect 3898 18533 3956 18542
rect 3052 18500 3092 18509
rect 643 18460 652 18500
rect 692 18460 1171 18500
rect 1211 18460 1220 18500
rect 1507 18460 1516 18500
rect 1556 18460 1987 18500
rect 2027 18460 2036 18500
rect 2083 18460 2092 18500
rect 2132 18460 2141 18500
rect 2275 18460 2284 18500
rect 2324 18460 2572 18500
rect 2612 18460 2621 18500
rect 2921 18460 3052 18500
rect 3092 18460 3101 18500
rect 3235 18460 3244 18500
rect 3284 18460 3540 18500
rect 3580 18460 3589 18500
rect 3898 18493 3907 18533
rect 3947 18493 3956 18533
rect 3898 18492 3956 18493
rect 0 18416 90 18436
rect 2092 18416 2132 18460
rect 3052 18451 3092 18460
rect 4588 18416 4628 18544
rect 0 18376 940 18416
rect 980 18376 989 18416
rect 1987 18376 1996 18416
rect 2036 18376 2572 18416
rect 2612 18376 2621 18416
rect 2947 18376 2956 18416
rect 2996 18376 3005 18416
rect 3724 18376 4628 18416
rect 0 18356 90 18376
rect 2956 18332 2996 18376
rect 3724 18332 3764 18376
rect 2956 18292 3532 18332
rect 3572 18292 3581 18332
rect 3715 18292 3724 18332
rect 3764 18292 3773 18332
rect 4492 18292 4732 18332
rect 4772 18292 4781 18332
rect 4492 18248 4532 18292
rect 4972 18248 5012 18544
rect 6700 18500 6740 18509
rect 5155 18460 5164 18500
rect 5204 18460 5452 18500
rect 5492 18460 5501 18500
rect 5923 18460 5932 18500
rect 5972 18460 6604 18500
rect 6644 18460 6700 18500
rect 6700 18451 6740 18460
rect 7372 18416 7412 18628
rect 7468 18628 8332 18668
rect 8372 18628 8381 18668
rect 7468 18584 7508 18628
rect 8620 18584 8660 18796
rect 7459 18544 7468 18584
rect 7508 18544 7517 18584
rect 7651 18544 7660 18584
rect 7700 18544 8236 18584
rect 8276 18544 8524 18584
rect 8564 18544 8573 18584
rect 8620 18544 9140 18584
rect 9100 18500 9140 18544
rect 7459 18460 7468 18500
rect 7508 18460 8035 18500
rect 8075 18460 8084 18500
rect 8131 18460 8140 18500
rect 8180 18460 8189 18500
rect 8585 18460 8620 18500
rect 8660 18460 8716 18500
rect 8756 18460 8765 18500
rect 9545 18460 9619 18500
rect 9659 18460 9676 18500
rect 9716 18460 9725 18500
rect 9859 18460 9868 18500
rect 9947 18460 10039 18500
rect 8140 18416 8180 18460
rect 9100 18451 9140 18460
rect 7372 18376 7852 18416
rect 7892 18376 7901 18416
rect 8092 18376 8180 18416
rect 5129 18292 5251 18332
rect 5300 18292 5309 18332
rect 6595 18292 6604 18332
rect 6644 18292 6892 18332
rect 6932 18292 6941 18332
rect 7337 18292 7459 18332
rect 7508 18292 7517 18332
rect 8092 18248 8132 18376
rect 9763 18292 9772 18332
rect 9812 18292 9821 18332
rect 10099 18292 10108 18332
rect 10148 18292 10540 18332
rect 10580 18292 10589 18332
rect 2947 18208 2956 18248
rect 2996 18208 4532 18248
rect 4780 18208 5012 18248
rect 5347 18208 5356 18248
rect 5396 18208 8132 18248
rect 4780 18164 4820 18208
rect 3628 18124 4820 18164
rect 4919 18124 4928 18164
rect 4968 18124 5010 18164
rect 5050 18124 5092 18164
rect 5132 18124 5174 18164
rect 5214 18124 5256 18164
rect 5296 18124 5305 18164
rect 0 18080 90 18100
rect 0 18040 364 18080
rect 404 18040 413 18080
rect 0 18020 90 18040
rect 3628 17996 3668 18124
rect 3619 17956 3628 17996
rect 3668 17956 3677 17996
rect 4483 17956 4492 17996
rect 4532 17956 5588 17996
rect 5635 17956 5644 17996
rect 5684 17956 5693 17996
rect 6089 17956 6220 17996
rect 6260 17956 6269 17996
rect 9353 17956 9484 17996
rect 9524 17956 9533 17996
rect 1123 17872 1132 17912
rect 1172 17872 1372 17912
rect 1412 17872 1421 17912
rect 1891 17872 1900 17912
rect 1940 17872 2420 17912
rect 2380 17828 2420 17872
rect 3148 17872 3532 17912
rect 3572 17872 3581 17912
rect 4387 17872 4396 17912
rect 4436 17872 5356 17912
rect 5396 17872 5405 17912
rect 451 17788 460 17828
rect 500 17819 1268 17828
rect 500 17788 1219 17819
rect 1210 17779 1219 17788
rect 1259 17779 1268 17819
rect 1882 17788 1891 17828
rect 1931 17788 1940 17828
rect 1987 17788 1996 17828
rect 2036 17788 2167 17828
rect 2371 17788 2380 17828
rect 2420 17788 2429 17828
rect 2921 17819 3052 17828
rect 2921 17788 2956 17819
rect 1210 17778 1268 17779
rect 0 17744 90 17764
rect 1900 17744 1940 17788
rect 2996 17788 3052 17819
rect 3092 17788 3101 17828
rect 2956 17770 2996 17779
rect 0 17704 76 17744
rect 116 17704 125 17744
rect 1891 17704 1900 17744
rect 1940 17704 1987 17744
rect 2275 17704 2284 17744
rect 2324 17704 2476 17744
rect 2516 17704 2525 17744
rect 0 17684 90 17704
rect 3148 17660 3188 17872
rect 3532 17828 3572 17872
rect 4972 17828 5012 17872
rect 3305 17788 3436 17828
rect 3476 17788 3485 17828
rect 3532 17788 3916 17828
rect 3956 17788 3965 17828
rect 4012 17788 4099 17828
rect 4139 17788 4148 17828
rect 4195 17788 4204 17828
rect 4244 17788 4253 17828
rect 4474 17788 4483 17828
rect 4523 17788 4532 17828
rect 4579 17788 4588 17828
rect 4628 17788 4780 17828
rect 4820 17788 4829 17828
rect 4963 17788 4972 17828
rect 5012 17788 5021 17828
rect 5548 17819 5588 17956
rect 5644 17912 5684 17956
rect 5644 17872 6548 17912
rect 6595 17872 6604 17912
rect 6644 17872 6653 17912
rect 7267 17872 7276 17912
rect 7316 17872 7660 17912
rect 7700 17872 7892 17912
rect 3436 17770 3476 17779
rect 4012 17744 4052 17788
rect 4204 17744 4244 17788
rect 4492 17744 4532 17788
rect 5635 17788 5644 17828
rect 5684 17819 6068 17828
rect 5684 17788 6028 17819
rect 5548 17770 5588 17779
rect 6028 17770 6068 17779
rect 3523 17704 3532 17744
rect 3572 17704 4052 17744
rect 4099 17704 4108 17744
rect 4148 17704 4244 17744
rect 4483 17704 4492 17744
rect 4532 17704 4579 17744
rect 4937 17704 5068 17744
rect 5108 17704 5117 17744
rect 6403 17704 6412 17744
rect 6452 17704 6461 17744
rect 3043 17620 3052 17660
rect 3092 17620 3188 17660
rect 4195 17536 4204 17576
rect 4244 17536 4300 17576
rect 4340 17536 4375 17576
rect 6412 17492 6452 17704
rect 6508 17660 6548 17872
rect 6604 17828 6644 17872
rect 7852 17828 7892 17872
rect 6604 17788 7747 17828
rect 7787 17788 7796 17828
rect 7843 17788 7852 17828
rect 7892 17788 7901 17828
rect 8105 17788 8236 17828
rect 8276 17788 8285 17828
rect 8681 17788 8812 17828
rect 8852 17788 8861 17828
rect 9161 17788 9292 17828
rect 9332 17788 9341 17828
rect 8812 17744 8852 17779
rect 9292 17770 9332 17779
rect 9772 17744 9812 18292
rect 11750 18080 11840 18100
rect 10723 18040 10732 18080
rect 10772 18040 11840 18080
rect 11750 18020 11840 18040
rect 10505 17956 10588 17996
rect 10628 17956 10636 17996
rect 10676 17956 10685 17996
rect 6595 17704 6604 17744
rect 6644 17704 7468 17744
rect 7508 17704 7517 17744
rect 8131 17704 8140 17744
rect 8180 17704 8332 17744
rect 8372 17704 8381 17744
rect 8812 17704 9196 17744
rect 9236 17704 9245 17744
rect 9772 17704 9868 17744
rect 9908 17704 9917 17744
rect 10339 17704 10348 17744
rect 10388 17704 10397 17744
rect 10348 17660 10388 17704
rect 6508 17620 10388 17660
rect 7267 17536 7276 17576
rect 7316 17536 9628 17576
rect 9668 17536 9677 17576
rect 6412 17452 8140 17492
rect 8180 17452 8189 17492
rect 0 17408 90 17428
rect 0 17368 460 17408
rect 500 17368 509 17408
rect 3679 17368 3688 17408
rect 3728 17368 3770 17408
rect 3810 17368 3852 17408
rect 3892 17368 3934 17408
rect 3974 17368 4016 17408
rect 4056 17368 4065 17408
rect 4108 17368 4876 17408
rect 4916 17368 4925 17408
rect 0 17348 90 17368
rect 3139 17116 3148 17156
rect 3188 17116 3532 17156
rect 3572 17116 4052 17156
rect 0 17072 90 17092
rect 0 17032 1420 17072
rect 1460 17032 1469 17072
rect 3532 17032 3628 17072
rect 3668 17032 3677 17072
rect 3785 17032 3907 17072
rect 3956 17032 3965 17072
rect 0 17012 90 17032
rect 2956 16988 2996 16997
rect 3532 16988 3572 17032
rect 4012 16988 4052 17116
rect 4108 17072 4148 17368
rect 4492 17284 5836 17324
rect 5876 17284 5885 17324
rect 10531 17284 10540 17324
rect 10580 17284 10924 17324
rect 10964 17284 10973 17324
rect 4099 17032 4108 17072
rect 4148 17032 4157 17072
rect 4492 16988 4532 17284
rect 4771 17200 4780 17240
rect 4820 17200 5251 17240
rect 5291 17200 5300 17240
rect 6787 17200 6796 17240
rect 6836 17200 7948 17240
rect 7988 17200 7997 17240
rect 9161 17200 9292 17240
rect 9332 17200 9341 17240
rect 10579 17200 10588 17240
rect 10628 17200 10732 17240
rect 10772 17200 10781 17240
rect 4579 17116 4588 17156
rect 4628 17116 5069 17156
rect 6307 17116 6316 17156
rect 6356 17116 10388 17156
rect 5029 17072 5069 17116
rect 10348 17072 10388 17116
rect 11750 17072 11840 17092
rect 4867 17032 4876 17072
rect 4916 17032 4925 17072
rect 5029 17032 5396 17072
rect 5731 17032 5740 17072
rect 5780 17032 5828 17072
rect 6211 17032 6220 17072
rect 6260 17032 6508 17072
rect 6548 17032 6557 17072
rect 7075 17032 7084 17072
rect 7124 17032 7892 17072
rect 9475 17032 9484 17072
rect 9524 17032 10156 17072
rect 10196 17032 10205 17072
rect 10339 17032 10348 17072
rect 10388 17032 10397 17072
rect 11203 17032 11212 17072
rect 11252 17032 11840 17072
rect 4876 16988 4916 17032
rect 5356 16988 5396 17032
rect 5548 16988 5588 16997
rect 5788 16988 5828 17032
rect 7852 16988 7892 17032
rect 11750 17012 11840 17032
rect 9100 16988 9140 16997
rect 547 16948 556 16988
rect 596 16948 1171 16988
rect 1211 16948 1220 16988
rect 1699 16948 1708 16988
rect 1748 16948 1757 16988
rect 2825 16948 2956 16988
rect 2996 16948 3005 16988
rect 3244 16948 3287 16988
rect 3327 16948 3336 16988
rect 3418 16948 3427 16988
rect 3467 16948 3476 16988
rect 3523 16948 3532 16988
rect 3572 16948 3581 16988
rect 3715 16948 3724 16988
rect 3764 16948 3767 16988
rect 3807 16948 3895 16988
rect 4003 16948 4012 16988
rect 4052 16948 4061 16988
rect 4282 16948 4291 16988
rect 4331 16948 4532 16988
rect 4579 16948 4588 16988
rect 4628 16948 4637 16988
rect 4771 16948 4780 16988
rect 4820 16948 4829 16988
rect 4876 16948 4902 16988
rect 4942 16948 4963 16988
rect 5020 16948 5029 16988
rect 5069 16948 5164 16988
rect 5204 16948 5246 16988
rect 5286 16948 5295 16988
rect 5356 16948 5548 16988
rect 5770 16948 5779 16988
rect 5819 16948 5828 16988
rect 5873 16948 5882 16988
rect 5922 16948 5932 16988
rect 5972 16948 6062 16988
rect 7171 16948 7180 16988
rect 7232 16948 7330 16988
rect 7370 16948 7401 16988
rect 7843 16948 7852 16988
rect 7892 16948 7901 16988
rect 8803 16948 8812 16988
rect 8852 16948 9100 16988
rect 9140 16948 9144 16988
rect 9283 16948 9292 16988
rect 9332 16948 9427 16988
rect 9467 16948 9476 16988
rect 9667 16948 9676 16988
rect 9716 16948 9868 16988
rect 9908 16948 9917 16988
rect 1708 16904 1748 16948
rect 2956 16939 2996 16948
rect 163 16864 172 16904
rect 212 16864 1748 16904
rect 3244 16904 3284 16948
rect 3436 16904 3476 16948
rect 4012 16904 4052 16948
rect 4588 16904 4628 16948
rect 3244 16864 3340 16904
rect 3380 16864 3389 16904
rect 3436 16864 3628 16904
rect 3668 16864 3677 16904
rect 4012 16864 4628 16904
rect 4396 16820 4436 16864
rect 1363 16780 1372 16820
rect 1412 16780 1804 16820
rect 1844 16780 1996 16820
rect 2036 16780 2045 16820
rect 3610 16780 3619 16820
rect 3659 16780 4012 16820
rect 4052 16780 4061 16820
rect 4387 16780 4396 16820
rect 4436 16780 4512 16820
rect 0 16736 90 16756
rect 4780 16736 4820 16948
rect 5548 16939 5588 16948
rect 9100 16939 9144 16948
rect 9104 16904 9144 16939
rect 5827 16864 5836 16904
rect 5876 16864 6268 16904
rect 6308 16864 6317 16904
rect 9104 16864 9628 16904
rect 9668 16864 9677 16904
rect 5059 16780 5068 16820
rect 5108 16780 5117 16820
rect 5251 16780 5260 16820
rect 5300 16780 5452 16820
rect 5492 16780 5501 16820
rect 6019 16780 6028 16820
rect 6068 16780 6077 16820
rect 6211 16780 6220 16820
rect 6260 16780 7027 16820
rect 7067 16780 7076 16820
rect 7180 16780 7516 16820
rect 7556 16780 7565 16820
rect 9785 16780 9868 16820
rect 9908 16780 9916 16820
rect 9956 16780 9965 16820
rect 0 16696 652 16736
rect 692 16696 701 16736
rect 4300 16696 4820 16736
rect 5068 16736 5108 16780
rect 5068 16696 5356 16736
rect 5396 16696 5405 16736
rect 0 16676 90 16696
rect 1027 16528 1036 16568
rect 1076 16528 1085 16568
rect 1036 16484 1076 16528
rect 4300 16484 4340 16696
rect 4919 16612 4928 16652
rect 4968 16612 5010 16652
rect 5050 16612 5092 16652
rect 5132 16612 5174 16652
rect 5214 16612 5256 16652
rect 5296 16612 5305 16652
rect 4387 16528 4396 16568
rect 4436 16528 5932 16568
rect 5972 16528 5981 16568
rect 1036 16444 1612 16484
rect 1652 16444 1844 16484
rect 4090 16444 4099 16484
rect 4139 16444 4340 16484
rect 0 16400 90 16420
rect 0 16360 1036 16400
rect 1076 16360 1085 16400
rect 0 16340 90 16360
rect 1804 16316 1844 16444
rect 3235 16360 3244 16400
rect 3284 16360 3293 16400
rect 4003 16360 4012 16400
rect 4052 16360 4532 16400
rect 3244 16316 3284 16360
rect 4492 16316 4532 16360
rect 4828 16316 4868 16528
rect 4937 16444 4972 16484
rect 5012 16444 5059 16484
rect 5099 16444 5117 16484
rect 5443 16444 5452 16484
rect 5492 16444 5644 16484
rect 5684 16444 5693 16484
rect 6028 16400 6068 16780
rect 7180 16400 7220 16780
rect 7459 16696 7468 16736
rect 7508 16696 7948 16736
rect 7988 16696 9292 16736
rect 9332 16696 9341 16736
rect 9484 16528 9676 16568
rect 9716 16528 9725 16568
rect 4972 16360 6068 16400
rect 6124 16360 7220 16400
rect 7468 16444 7564 16484
rect 7604 16444 7613 16484
rect 4972 16316 5012 16360
rect 6124 16316 6164 16360
rect 7468 16316 7508 16444
rect 9484 16400 9524 16528
rect 9571 16444 9580 16484
rect 9620 16444 10156 16484
rect 10196 16444 10205 16484
rect 7747 16360 7756 16400
rect 7796 16360 8372 16400
rect 8611 16360 8620 16400
rect 8660 16360 9859 16400
rect 9899 16360 9908 16400
rect 8332 16316 8372 16360
rect 739 16276 748 16316
rect 788 16307 1268 16316
rect 788 16276 1219 16307
rect 1210 16267 1219 16276
rect 1259 16267 1268 16307
rect 1795 16276 1804 16316
rect 1844 16276 1853 16316
rect 2921 16276 2956 16316
rect 2996 16307 3092 16316
rect 2996 16276 3052 16307
rect 1210 16266 1268 16267
rect 3209 16276 3340 16316
rect 3380 16276 3916 16316
rect 3956 16276 3965 16316
rect 4060 16276 4107 16316
rect 4147 16276 4156 16316
rect 4258 16295 4267 16316
rect 4204 16276 4267 16295
rect 4307 16276 4316 16316
rect 4483 16276 4492 16316
rect 4532 16276 4541 16316
rect 4723 16276 4732 16316
rect 4772 16276 4781 16316
rect 4828 16276 4867 16316
rect 4907 16276 4916 16316
rect 4963 16276 4972 16316
rect 5012 16276 5021 16316
rect 5347 16276 5356 16316
rect 5396 16307 6164 16316
rect 5396 16276 5644 16307
rect 3052 16258 3092 16267
rect 4060 16232 4100 16276
rect 4204 16255 4316 16276
rect 67 16192 76 16232
rect 116 16192 212 16232
rect 1363 16192 1372 16232
rect 1412 16192 2860 16232
rect 2900 16192 2909 16232
rect 3497 16192 3532 16232
rect 3572 16192 3628 16232
rect 3668 16192 3677 16232
rect 4060 16192 4108 16232
rect 4148 16192 4157 16232
rect 172 16148 212 16192
rect 4204 16148 4244 16255
rect 4732 16232 4772 16276
rect 5684 16276 6164 16307
rect 6883 16276 6892 16316
rect 6932 16276 6941 16316
rect 7075 16276 7084 16316
rect 7124 16276 7508 16316
rect 7555 16276 7564 16316
rect 7604 16276 7843 16316
rect 7883 16276 7892 16316
rect 7939 16276 7948 16316
rect 7988 16276 7997 16316
rect 8201 16276 8332 16316
rect 8372 16276 8381 16316
rect 8803 16276 8812 16316
rect 8852 16307 9004 16316
rect 8852 16276 8908 16307
rect 5644 16258 5684 16267
rect 6892 16232 6932 16276
rect 7948 16232 7988 16276
rect 8948 16276 9004 16307
rect 9044 16276 9108 16316
rect 9257 16276 9388 16316
rect 9428 16276 9437 16316
rect 9667 16276 9676 16316
rect 9716 16276 10252 16316
rect 10292 16276 10301 16316
rect 8908 16258 8948 16267
rect 9388 16258 9428 16267
rect 4378 16192 4387 16232
rect 4427 16192 4484 16232
rect 4579 16192 4588 16232
rect 4628 16192 4637 16232
rect 4732 16192 4876 16232
rect 4916 16192 4925 16232
rect 5731 16192 5740 16232
rect 5780 16192 7468 16232
rect 7508 16192 7517 16232
rect 7747 16192 7756 16232
rect 7796 16192 7988 16232
rect 8297 16192 8428 16232
rect 8468 16192 8477 16232
rect 4444 16148 4484 16192
rect 172 16108 3388 16148
rect 3428 16108 3437 16148
rect 4204 16108 4340 16148
rect 4387 16108 4396 16148
rect 4436 16108 4484 16148
rect 0 16064 90 16084
rect 4300 16064 4340 16108
rect 0 16024 212 16064
rect 4291 16024 4300 16064
rect 4340 16024 4349 16064
rect 0 16004 90 16024
rect 172 15896 212 16024
rect 4588 15896 4628 16192
rect 11750 16064 11840 16084
rect 10723 16024 10732 16064
rect 10772 16024 11840 16064
rect 11750 16004 11840 16024
rect 172 15856 2900 15896
rect 3679 15856 3688 15896
rect 3728 15856 3770 15896
rect 3810 15856 3852 15896
rect 3892 15856 3934 15896
rect 3974 15856 4016 15896
rect 4056 15856 4065 15896
rect 4588 15856 5644 15896
rect 5684 15856 5693 15896
rect 0 15728 90 15748
rect 2860 15728 2900 15856
rect 3724 15772 9868 15812
rect 9908 15772 9917 15812
rect 0 15688 1324 15728
rect 1364 15688 1373 15728
rect 1891 15688 1900 15728
rect 1940 15688 2668 15728
rect 2708 15688 2717 15728
rect 2860 15688 3196 15728
rect 3236 15688 3245 15728
rect 0 15668 90 15688
rect 1411 15604 1420 15644
rect 1460 15604 2812 15644
rect 2852 15604 2861 15644
rect 3043 15604 3052 15644
rect 3092 15604 3628 15644
rect 3668 15604 3677 15644
rect 3724 15560 3764 15772
rect 4003 15688 4012 15728
rect 4052 15688 5356 15728
rect 5396 15688 5405 15728
rect 7433 15688 7564 15728
rect 7604 15688 7613 15728
rect 9379 15688 9388 15728
rect 9428 15688 9772 15728
rect 9812 15688 9821 15728
rect 10579 15688 10588 15728
rect 10628 15688 11212 15728
rect 11252 15688 11261 15728
rect 4108 15604 4732 15644
rect 4772 15604 4781 15644
rect 7171 15604 7180 15644
rect 7220 15604 10388 15644
rect 2921 15520 2956 15560
rect 2996 15520 3052 15560
rect 3092 15520 3101 15560
rect 3427 15520 3436 15560
rect 3476 15520 3764 15560
rect 3811 15520 3820 15560
rect 3860 15520 3991 15560
rect 2476 15476 2516 15485
rect 163 15436 172 15476
rect 212 15436 1228 15476
rect 1268 15436 1940 15476
rect 1987 15436 1996 15476
rect 2036 15436 2476 15476
rect 2516 15436 4012 15476
rect 4052 15436 4061 15476
rect 0 15392 90 15412
rect 1900 15392 1940 15436
rect 2476 15427 2516 15436
rect 0 15352 788 15392
rect 1891 15352 1900 15392
rect 1940 15352 1949 15392
rect 2572 15352 3580 15392
rect 3620 15352 3629 15392
rect 0 15332 90 15352
rect 748 15308 788 15352
rect 2572 15308 2612 15352
rect 748 15268 2612 15308
rect 3436 15268 3964 15308
rect 4004 15268 4013 15308
rect 3436 15224 3476 15268
rect 67 15184 76 15224
rect 116 15184 3476 15224
rect 4108 15140 4148 15604
rect 10348 15560 10388 15604
rect 4195 15520 4204 15560
rect 4244 15520 4300 15560
rect 4340 15520 4375 15560
rect 4492 15520 4588 15560
rect 4628 15520 4637 15560
rect 4963 15520 4972 15560
rect 5012 15520 5740 15560
rect 5780 15520 5789 15560
rect 7372 15520 8620 15560
rect 8660 15520 9620 15560
rect 10025 15520 10156 15560
rect 10196 15520 10205 15560
rect 10339 15520 10348 15560
rect 10388 15520 10397 15560
rect 4217 15268 4300 15308
rect 4340 15268 4348 15308
rect 4388 15268 4397 15308
rect 4492 15224 4532 15520
rect 7372 15476 7412 15520
rect 9580 15476 9620 15520
rect 5129 15436 5260 15476
rect 5300 15436 5309 15476
rect 6019 15436 6028 15476
rect 6068 15436 6124 15476
rect 6164 15436 6199 15476
rect 7459 15436 7468 15476
rect 7508 15436 8332 15476
rect 8372 15436 8381 15476
rect 7372 15427 7412 15436
rect 9580 15427 9620 15436
rect 172 15100 4148 15140
rect 4204 15184 4532 15224
rect 4588 15268 5116 15308
rect 5156 15268 5165 15308
rect 8995 15268 9004 15308
rect 9044 15268 9916 15308
rect 9956 15268 9965 15308
rect 0 15056 90 15076
rect 0 15016 76 15056
rect 116 15016 125 15056
rect 0 14996 90 15016
rect 0 14720 90 14740
rect 172 14720 212 15100
rect 4204 14972 4244 15184
rect 355 14932 364 14972
rect 404 14932 1564 14972
rect 1604 14932 1613 14972
rect 1699 14932 1708 14972
rect 1748 14932 2852 14972
rect 4195 14932 4204 14972
rect 4244 14932 4253 14972
rect 4361 14932 4492 14972
rect 4532 14932 4541 14972
rect 451 14848 460 14888
rect 500 14848 1948 14888
rect 1988 14848 1997 14888
rect 2812 14804 2852 14932
rect 4588 14888 4628 15268
rect 4919 15100 4928 15140
rect 4968 15100 5010 15140
rect 5050 15100 5092 15140
rect 5132 15100 5174 15140
rect 5214 15100 5256 15140
rect 5296 15100 5305 15140
rect 11750 15056 11840 15076
rect 10627 15016 10636 15056
rect 10676 15016 11840 15056
rect 11750 14996 11840 15016
rect 3619 14848 3628 14888
rect 3668 14848 4628 14888
rect 7468 14932 7948 14972
rect 7988 14932 8428 14972
rect 8468 14932 8477 14972
rect 10579 14932 10588 14972
rect 10628 14932 10732 14972
rect 10772 14932 10781 14972
rect 7468 14804 7508 14932
rect 7555 14848 7564 14888
rect 7604 14848 7892 14888
rect 7852 14804 7892 14848
rect 2458 14764 2467 14804
rect 2507 14764 2516 14804
rect 2563 14764 2572 14804
rect 2612 14764 2743 14804
rect 2812 14764 2860 14804
rect 2900 14764 2956 14804
rect 2996 14764 3031 14804
rect 3532 14795 3724 14804
rect 2476 14720 2516 14764
rect 3572 14764 3724 14795
rect 3764 14764 3773 14804
rect 4012 14795 4052 14804
rect 3532 14746 3572 14755
rect 0 14680 212 14720
rect 931 14680 940 14720
rect 980 14680 1228 14720
rect 1268 14680 1277 14720
rect 1795 14680 1804 14720
rect 1844 14680 1853 14720
rect 2179 14680 2188 14720
rect 2228 14680 2284 14720
rect 2324 14680 2359 14720
rect 2476 14680 2668 14720
rect 2708 14680 2717 14720
rect 3043 14680 3052 14720
rect 3092 14680 3223 14720
rect 0 14660 90 14680
rect 1804 14636 1844 14680
rect 4012 14636 4052 14755
rect 4684 14795 5356 14804
rect 4724 14764 5356 14795
rect 5396 14764 5405 14804
rect 5731 14764 5740 14804
rect 5780 14764 5932 14804
rect 5972 14764 6028 14804
rect 6068 14764 6124 14804
rect 6164 14764 6228 14804
rect 7372 14795 7564 14804
rect 4684 14746 4724 14755
rect 7412 14764 7564 14795
rect 7604 14764 7668 14804
rect 7834 14764 7843 14804
rect 7883 14764 7892 14804
rect 7939 14764 7948 14804
rect 7988 14764 8119 14804
rect 8201 14764 8332 14804
rect 8372 14764 8381 14804
rect 8777 14764 8908 14804
rect 8948 14764 8957 14804
rect 9257 14764 9388 14804
rect 9428 14764 9437 14804
rect 7372 14746 7412 14755
rect 8908 14746 8948 14755
rect 9388 14746 9428 14755
rect 8419 14680 8428 14720
rect 8468 14680 8812 14720
rect 8852 14680 8861 14720
rect 9610 14680 9619 14720
rect 9659 14680 9964 14720
rect 10004 14680 10013 14720
rect 10339 14680 10348 14720
rect 10388 14680 11020 14720
rect 11060 14680 11069 14720
rect 1804 14596 2900 14636
rect 3331 14596 3340 14636
rect 3380 14596 4052 14636
rect 2860 14552 2900 14596
rect 1459 14512 1468 14552
rect 1508 14512 2228 14552
rect 2860 14512 5548 14552
rect 5588 14512 5597 14552
rect 8611 14512 8620 14552
rect 8660 14512 9724 14552
rect 9764 14512 9773 14552
rect 2188 14468 2228 14512
rect 2188 14428 6220 14468
rect 6260 14428 6269 14468
rect 0 14384 90 14404
rect 0 14344 212 14384
rect 3679 14344 3688 14384
rect 3728 14344 3770 14384
rect 3810 14344 3852 14384
rect 3892 14344 3934 14384
rect 3974 14344 4016 14384
rect 4056 14344 4065 14384
rect 0 14324 90 14344
rect 172 14216 212 14344
rect 5068 14260 10540 14300
rect 10580 14260 10589 14300
rect 172 14176 4828 14216
rect 4868 14176 4877 14216
rect 643 14092 652 14132
rect 692 14092 1180 14132
rect 1220 14092 1229 14132
rect 1315 14092 1324 14132
rect 1364 14092 1556 14132
rect 0 14048 90 14068
rect 0 14008 556 14048
rect 596 14008 605 14048
rect 1289 14008 1420 14048
rect 1460 14008 1469 14048
rect 0 13988 90 14008
rect 1516 13880 1556 14092
rect 1804 14092 2572 14132
rect 2612 14092 2621 14132
rect 3715 14092 3724 14132
rect 3764 14092 4876 14132
rect 4916 14092 4925 14132
rect 1804 14048 1844 14092
rect 5068 14048 5108 14260
rect 5779 14176 5788 14216
rect 5828 14176 7180 14216
rect 7220 14176 7229 14216
rect 9187 14176 9196 14216
rect 9236 14176 9388 14216
rect 9428 14176 9437 14216
rect 10505 14176 10588 14216
rect 10628 14176 10636 14216
rect 10676 14176 10685 14216
rect 6185 14092 6268 14132
rect 6308 14092 6316 14132
rect 6356 14092 6365 14132
rect 10195 14092 10204 14132
rect 10244 14092 11060 14132
rect 11020 14048 11060 14092
rect 11750 14048 11840 14068
rect 1795 14008 1804 14048
rect 1844 14008 1853 14048
rect 2179 14008 2188 14048
rect 2228 14008 2237 14048
rect 2851 14008 2860 14048
rect 2900 14008 3052 14048
rect 3092 14008 3101 14048
rect 4330 14008 4339 14048
rect 4379 14008 4684 14048
rect 4724 14008 4733 14048
rect 5059 14008 5068 14048
rect 5108 14008 5117 14048
rect 5539 14008 5548 14048
rect 5588 14008 5740 14048
rect 5780 14008 5789 14048
rect 6019 14008 6028 14048
rect 6068 14008 7468 14048
rect 7508 14008 7517 14048
rect 9449 14008 9532 14048
rect 9572 14008 9580 14048
rect 9620 14008 9629 14048
rect 9955 14008 9964 14048
rect 10004 14008 10060 14048
rect 10100 14008 10135 14048
rect 10339 14008 10348 14048
rect 10388 14008 10540 14048
rect 10580 14008 10589 14048
rect 11020 14008 11840 14048
rect 1516 13840 1948 13880
rect 1988 13840 1997 13880
rect 2188 13796 2228 14008
rect 3628 13964 3668 13973
rect 7468 13964 7508 14008
rect 11750 13988 11840 14008
rect 9004 13964 9044 13973
rect 2275 13924 2284 13964
rect 2324 13924 2563 13964
rect 2603 13924 2612 13964
rect 2659 13924 2668 13964
rect 2708 13924 2764 13964
rect 2804 13924 2839 13964
rect 3043 13924 3052 13964
rect 3092 13924 3148 13964
rect 3188 13924 3223 13964
rect 3497 13924 3628 13964
rect 3668 13924 3677 13964
rect 4138 13924 4147 13964
rect 4187 13924 4204 13964
rect 4244 13924 4327 13964
rect 7171 13924 7180 13964
rect 7259 13924 7351 13964
rect 7468 13924 7756 13964
rect 7796 13924 7805 13964
rect 8419 13924 8428 13964
rect 8468 13924 9004 13964
rect 9367 13924 9376 13964
rect 9416 13924 10252 13964
rect 10292 13924 10301 13964
rect 3628 13915 3668 13924
rect 9004 13915 9044 13924
rect 4300 13840 8620 13880
rect 8660 13840 8669 13880
rect 4300 13796 4340 13840
rect 1027 13756 1036 13796
rect 1076 13756 1564 13796
rect 1604 13756 1613 13796
rect 2188 13756 4340 13796
rect 4435 13756 4444 13796
rect 4484 13756 4492 13796
rect 4532 13756 4615 13796
rect 7411 13756 7420 13796
rect 7460 13756 10348 13796
rect 10388 13756 10397 13796
rect 0 13712 90 13732
rect 0 13672 1324 13712
rect 1364 13672 1373 13712
rect 0 13652 90 13672
rect 4919 13588 4928 13628
rect 4968 13588 5010 13628
rect 5050 13588 5092 13628
rect 5132 13588 5174 13628
rect 5214 13588 5256 13628
rect 5296 13588 5305 13628
rect 7084 13588 8948 13628
rect 1411 13504 1420 13544
rect 1460 13504 6028 13544
rect 6068 13504 6077 13544
rect 7084 13460 7124 13588
rect 2851 13420 2860 13460
rect 2900 13420 3340 13460
rect 3380 13420 3389 13460
rect 4483 13420 4492 13460
rect 4532 13420 4780 13460
rect 4820 13420 4829 13460
rect 5932 13420 7124 13460
rect 7276 13504 7660 13544
rect 7700 13504 7709 13544
rect 0 13376 90 13396
rect 0 13336 652 13376
rect 692 13336 701 13376
rect 2860 13336 3724 13376
rect 3764 13336 3773 13376
rect 4300 13336 5876 13376
rect 0 13316 90 13336
rect 2860 13292 2900 13336
rect 1411 13252 1420 13292
rect 1460 13252 1612 13292
rect 1652 13252 1661 13292
rect 2668 13283 2900 13292
rect 2708 13252 2900 13283
rect 3043 13252 3052 13292
rect 3092 13252 3101 13292
rect 4300 13283 4340 13336
rect 2668 13234 2708 13243
rect 3052 13124 3092 13252
rect 4675 13252 4684 13292
rect 4724 13252 4733 13292
rect 4300 13234 4340 13243
rect 4684 13124 4724 13252
rect 2851 13084 2860 13124
rect 2900 13084 2909 13124
rect 3052 13084 3340 13124
rect 3380 13084 4724 13124
rect 5836 13124 5876 13336
rect 5932 13283 5972 13420
rect 6115 13336 6124 13376
rect 6164 13336 7028 13376
rect 6988 13292 7028 13336
rect 7276 13292 7316 13504
rect 7363 13336 7372 13376
rect 7412 13336 8812 13376
rect 8852 13336 8861 13376
rect 8908 13292 8948 13588
rect 10243 13336 10252 13376
rect 10292 13336 10348 13376
rect 10388 13336 10423 13376
rect 6979 13252 6988 13292
rect 7028 13252 7037 13292
rect 7258 13252 7267 13292
rect 7307 13252 7316 13292
rect 7372 13252 8044 13292
rect 8084 13252 8812 13292
rect 8852 13252 8861 13292
rect 8908 13252 9292 13292
rect 9332 13283 10100 13292
rect 9332 13252 10060 13283
rect 5932 13234 5972 13243
rect 7372 13208 7412 13252
rect 10060 13234 10100 13243
rect 7171 13168 7180 13208
rect 7220 13168 7412 13208
rect 8035 13168 8044 13208
rect 8084 13168 8093 13208
rect 8419 13168 8428 13208
rect 8468 13168 9100 13208
rect 9140 13168 9149 13208
rect 5836 13084 7564 13124
rect 7604 13084 7613 13124
rect 7673 13084 7756 13124
rect 7796 13084 7804 13124
rect 7844 13084 7853 13124
rect 0 13040 90 13060
rect 2860 13040 2900 13084
rect 0 13000 748 13040
rect 788 13000 797 13040
rect 2275 13000 2284 13040
rect 2324 13000 2900 13040
rect 0 12980 90 13000
rect 3052 12956 3092 13084
rect 8044 13040 8084 13168
rect 8659 13084 8668 13124
rect 8708 13084 10388 13124
rect 3715 13000 3724 13040
rect 3764 13000 3773 13040
rect 3907 13000 3916 13040
rect 3956 13000 4684 13040
rect 4724 13000 4733 13040
rect 7651 13000 7660 13040
rect 7700 13000 8084 13040
rect 10348 13040 10388 13084
rect 11750 13040 11840 13060
rect 10348 13000 11840 13040
rect 3724 12956 3764 13000
rect 11750 12980 11840 13000
rect 1603 12916 1612 12956
rect 1652 12916 3092 12956
rect 3331 12916 3340 12956
rect 3380 12916 3764 12956
rect 3679 12832 3688 12872
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 4056 12832 4065 12872
rect 4108 12832 11788 12872
rect 11828 12832 11837 12872
rect 1420 12748 3532 12788
rect 3572 12748 3581 12788
rect 0 12704 90 12724
rect 1420 12704 1460 12748
rect 4108 12704 4148 12832
rect 5059 12748 5068 12788
rect 5108 12748 11116 12788
rect 11156 12748 11165 12788
rect 0 12664 1460 12704
rect 2851 12664 2860 12704
rect 2900 12664 3031 12704
rect 3715 12664 3724 12704
rect 3764 12664 4148 12704
rect 4204 12664 6076 12704
rect 6116 12664 6125 12704
rect 8969 12664 9100 12704
rect 9140 12664 9149 12704
rect 0 12644 90 12664
rect 4204 12620 4244 12664
rect 2537 12580 2668 12620
rect 2708 12580 2717 12620
rect 3907 12580 3916 12620
rect 3956 12580 4244 12620
rect 4300 12580 6124 12620
rect 6164 12580 6173 12620
rect 8777 12580 8908 12620
rect 8948 12580 8957 12620
rect 9196 12580 9964 12620
rect 10004 12580 10013 12620
rect 2476 12452 2516 12461
rect 3052 12452 3092 12461
rect 4300 12452 4340 12580
rect 9196 12536 9236 12580
rect 4675 12496 4684 12536
rect 4724 12496 4780 12536
rect 4820 12496 4855 12536
rect 5059 12496 5068 12536
rect 5108 12496 5239 12536
rect 5443 12496 5452 12536
rect 5492 12496 5836 12536
rect 5876 12496 5885 12536
rect 5932 12496 6316 12536
rect 6356 12496 6365 12536
rect 7468 12496 9236 12536
rect 1097 12412 1228 12452
rect 1268 12412 1277 12452
rect 2516 12412 2764 12452
rect 2804 12412 3052 12452
rect 3092 12412 3340 12452
rect 3380 12412 3389 12452
rect 3619 12412 3628 12452
rect 3668 12412 4300 12452
rect 4340 12412 4396 12452
rect 4436 12412 4500 12452
rect 2476 12403 2516 12412
rect 3052 12403 3092 12412
rect 0 12368 90 12388
rect 0 12328 212 12368
rect 0 12308 90 12328
rect 172 12200 212 12328
rect 3148 12328 5212 12368
rect 5252 12328 5261 12368
rect 3148 12284 3188 12328
rect 451 12244 460 12284
rect 500 12244 3188 12284
rect 3340 12244 4444 12284
rect 4484 12244 4493 12284
rect 4819 12244 4828 12284
rect 4868 12244 4877 12284
rect 3340 12200 3380 12244
rect 172 12160 3380 12200
rect 4828 12116 4868 12244
rect 844 12076 4868 12116
rect 4919 12076 4928 12116
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 5296 12076 5305 12116
rect 5635 12076 5644 12116
rect 5684 12076 5693 12116
rect 0 12032 90 12052
rect 844 12032 884 12076
rect 5644 12032 5684 12076
rect 0 11992 884 12032
rect 1795 11992 1804 12032
rect 1844 11992 4340 12032
rect 0 11972 90 11992
rect 2921 11908 2956 11948
rect 2996 11908 3052 11948
rect 3092 11908 3101 11948
rect 3449 11908 3532 11948
rect 3572 11908 3580 11948
rect 3620 11908 3629 11948
rect 2851 11824 2860 11864
rect 2900 11824 3956 11864
rect 1481 11740 1516 11780
rect 1556 11740 1612 11780
rect 1652 11740 1661 11780
rect 1987 11740 1996 11780
rect 2036 11740 2668 11780
rect 2708 11771 2804 11780
rect 2708 11740 2764 11771
rect 3469 11740 3478 11780
rect 3518 11740 3628 11780
rect 3668 11740 3677 11780
rect 2764 11722 2804 11731
rect 0 11696 90 11716
rect 3916 11696 3956 11824
rect 4300 11780 4340 11992
rect 4876 11992 5684 12032
rect 4876 11780 4916 11992
rect 5932 11948 5972 12496
rect 7468 12452 7508 12496
rect 9292 12452 9332 12461
rect 7213 12412 7222 12452
rect 7262 12412 7508 12452
rect 7555 12412 7564 12452
rect 7604 12412 8083 12452
rect 8123 12412 8132 12452
rect 9161 12412 9292 12452
rect 9332 12412 9341 12452
rect 10243 12412 10252 12452
rect 10292 12412 10540 12452
rect 10580 12412 10589 12452
rect 9292 12403 9332 12412
rect 6403 12244 6412 12284
rect 6452 12244 7027 12284
rect 7067 12244 7076 12284
rect 7555 12244 7564 12284
rect 7604 12244 8284 12284
rect 8324 12244 8333 12284
rect 11750 12032 11840 12052
rect 10627 11992 10636 12032
rect 10676 11992 11840 12032
rect 11750 11972 11840 11992
rect 5923 11908 5932 11948
rect 5972 11908 5981 11948
rect 7721 11908 7804 11948
rect 7844 11908 7852 11948
rect 7892 11908 7901 11948
rect 8419 11908 8428 11948
rect 8468 11908 10060 11948
rect 10100 11908 10540 11948
rect 10580 11908 10589 11948
rect 5260 11824 5932 11864
rect 5972 11824 6700 11864
rect 6740 11824 6749 11864
rect 8044 11824 8660 11864
rect 4043 11740 4108 11780
rect 4148 11740 4174 11780
rect 4214 11740 4223 11780
rect 4291 11740 4300 11780
rect 4340 11740 4349 11780
rect 4675 11740 4684 11780
rect 4724 11740 4876 11780
rect 4916 11740 4925 11780
rect 5260 11771 5300 11824
rect 5609 11740 5740 11780
rect 5780 11740 5789 11780
rect 6115 11740 6124 11780
rect 6164 11740 6220 11780
rect 6260 11740 6295 11780
rect 7433 11771 7564 11780
rect 7433 11740 7468 11771
rect 5260 11722 5300 11731
rect 5740 11722 5780 11731
rect 7508 11740 7564 11771
rect 7604 11740 7613 11780
rect 7468 11722 7508 11731
rect 8044 11696 8084 11824
rect 8620 11780 8660 11824
rect 8602 11740 8611 11780
rect 8660 11740 8791 11780
rect 0 11656 172 11696
rect 212 11656 221 11696
rect 3274 11656 3283 11696
rect 3323 11656 3532 11696
rect 3572 11656 3581 11696
rect 3689 11656 3820 11696
rect 3860 11656 3869 11696
rect 3916 11656 4492 11696
rect 4532 11656 4780 11696
rect 4820 11656 4829 11696
rect 8035 11656 8044 11696
rect 8084 11656 8093 11696
rect 8227 11656 8236 11696
rect 8276 11656 8372 11696
rect 8899 11656 8908 11696
rect 8948 11656 8957 11696
rect 0 11636 90 11656
rect 8044 11612 8084 11656
rect 1987 11572 1996 11612
rect 2036 11572 8084 11612
rect 8332 11528 8372 11656
rect 8524 11572 8812 11612
rect 8852 11572 8861 11612
rect 8524 11528 8564 11572
rect 3907 11488 3916 11528
rect 3956 11488 3965 11528
rect 7529 11488 7660 11528
rect 7700 11488 7709 11528
rect 8332 11488 8564 11528
rect 3916 11444 3956 11488
rect 3523 11404 3532 11444
rect 3572 11404 3956 11444
rect 4963 11404 4972 11444
rect 5012 11404 11404 11444
rect 11444 11404 11453 11444
rect 0 11360 90 11380
rect 0 11320 1228 11360
rect 1268 11320 1277 11360
rect 3679 11320 3688 11360
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 4056 11320 4065 11360
rect 6691 11320 6700 11360
rect 6740 11320 11500 11360
rect 11540 11320 11549 11360
rect 0 11300 90 11320
rect 2467 11236 2476 11276
rect 2516 11236 6740 11276
rect 6700 11192 6740 11236
rect 547 11152 556 11192
rect 596 11152 1180 11192
rect 1220 11152 1229 11192
rect 1315 11152 1324 11192
rect 1364 11152 1564 11192
rect 1604 11152 1613 11192
rect 3619 11152 3628 11192
rect 3668 11152 4300 11192
rect 4340 11152 4349 11192
rect 5705 11152 5740 11192
rect 5780 11152 5836 11192
rect 5876 11152 5885 11192
rect 6115 11152 6124 11192
rect 6164 11152 6508 11192
rect 6548 11152 6557 11192
rect 6700 11152 6836 11192
rect 1420 11068 2860 11108
rect 2900 11068 2909 11108
rect 4483 11068 4492 11108
rect 4532 11068 6740 11108
rect 0 11024 90 11044
rect 1420 11024 1460 11068
rect 6700 11024 6740 11068
rect 0 10984 1132 11024
rect 1172 10984 1181 11024
rect 1411 10984 1420 11024
rect 1460 10984 1469 11024
rect 1795 10984 1804 11024
rect 1844 10984 2956 11024
rect 2996 10984 3005 11024
rect 3689 10984 3820 11024
rect 3860 10984 3869 11024
rect 4051 10984 4060 11024
rect 4100 10984 4972 11024
rect 5012 10984 5021 11024
rect 6211 10984 6220 11024
rect 6260 10984 6356 11024
rect 6691 10984 6700 11024
rect 6740 10984 6749 11024
rect 0 10964 90 10984
rect 3436 10940 3476 10949
rect 5644 10940 5684 10949
rect 6316 10940 6356 10984
rect 6796 10940 6836 11152
rect 7276 11152 9580 11192
rect 9620 11152 10540 11192
rect 10580 11152 10589 11192
rect 7276 10940 7316 11152
rect 11750 11024 11840 11044
rect 9283 10984 9292 11024
rect 9332 10984 9341 11024
rect 10243 10984 10252 11024
rect 10292 10984 11840 11024
rect 11750 10964 11840 10984
rect 2153 10900 2188 10940
rect 2228 10900 2284 10940
rect 2324 10900 2333 10940
rect 2851 10900 2860 10940
rect 2900 10900 3436 10940
rect 4265 10900 4396 10940
rect 4436 10900 4445 10940
rect 5731 10900 5740 10940
rect 5780 10900 6211 10940
rect 6251 10900 6260 10940
rect 6307 10900 6316 10940
rect 6356 10900 6508 10940
rect 6548 10900 6557 10940
rect 6787 10900 6796 10940
rect 6836 10900 6845 10940
rect 7316 10900 7468 10940
rect 7508 10900 7517 10940
rect 7651 10900 7660 10940
rect 7700 10900 7764 10940
rect 7804 10900 7831 10940
rect 8602 10900 8611 10940
rect 8660 10900 8791 10940
rect 3436 10891 3476 10900
rect 5644 10856 5684 10900
rect 7276 10891 7316 10900
rect 5356 10816 6412 10856
rect 6452 10816 6461 10856
rect 7756 10816 8084 10856
rect 8218 10816 8227 10856
rect 8267 10816 8716 10856
rect 8756 10816 9196 10856
rect 9236 10816 9245 10856
rect 2275 10732 2284 10772
rect 2324 10732 3820 10772
rect 3860 10732 3869 10772
rect 4780 10732 4876 10772
rect 4916 10732 4925 10772
rect 0 10688 90 10708
rect 0 10648 1036 10688
rect 1076 10648 1085 10688
rect 0 10628 90 10648
rect 643 10396 652 10436
rect 692 10396 1180 10436
rect 1220 10396 1229 10436
rect 3715 10396 3724 10436
rect 3764 10396 4108 10436
rect 4148 10396 4157 10436
rect 0 10352 90 10372
rect 0 10312 460 10352
rect 500 10312 509 10352
rect 739 10312 748 10352
rect 788 10312 1564 10352
rect 1604 10312 1613 10352
rect 0 10292 90 10312
rect 4780 10268 4820 10732
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 5356 10436 5396 10816
rect 7756 10772 7796 10816
rect 5539 10732 5548 10772
rect 5588 10732 7796 10772
rect 7939 10732 7948 10772
rect 7988 10732 7997 10772
rect 5251 10396 5260 10436
rect 5300 10396 5396 10436
rect 5356 10312 5932 10352
rect 5972 10312 6988 10352
rect 7028 10312 7037 10352
rect 2153 10228 2284 10268
rect 2324 10228 2333 10268
rect 3532 10259 3572 10268
rect 4282 10228 4291 10268
rect 4331 10228 4340 10268
rect 4387 10228 4396 10268
rect 4436 10228 4588 10268
rect 4628 10228 4637 10268
rect 4745 10228 4780 10268
rect 4820 10228 4876 10268
rect 4916 10228 4925 10268
rect 5356 10259 5396 10312
rect 1289 10144 1420 10184
rect 1460 10144 1469 10184
rect 1673 10144 1804 10184
rect 1844 10144 1853 10184
rect 3532 10100 3572 10219
rect 4300 10184 4340 10228
rect 5705 10228 5836 10268
rect 5876 10228 5885 10268
rect 6019 10228 6028 10268
rect 6068 10228 7028 10268
rect 5356 10210 5396 10219
rect 5836 10210 5876 10219
rect 4291 10144 4300 10184
rect 4340 10144 4387 10184
rect 4483 10144 4492 10184
rect 4532 10144 4876 10184
rect 4916 10144 4925 10184
rect 6058 10144 6067 10184
rect 6107 10144 6412 10184
rect 6452 10144 6461 10184
rect 6665 10144 6700 10184
rect 6740 10144 6796 10184
rect 6836 10144 6845 10184
rect 6988 10100 7028 10228
rect 7948 10184 7988 10732
rect 8044 10436 8084 10816
rect 8044 10396 8380 10436
rect 8420 10396 8429 10436
rect 10121 10396 10204 10436
rect 10244 10396 10252 10436
rect 10292 10396 10301 10436
rect 10505 10396 10588 10436
rect 10628 10396 10636 10436
rect 10676 10396 10685 10436
rect 9964 10228 11692 10268
rect 11732 10228 11741 10268
rect 9964 10184 10004 10228
rect 7948 10144 8236 10184
rect 8276 10144 8285 10184
rect 8489 10144 8620 10184
rect 8660 10144 8669 10184
rect 8777 10144 8908 10184
rect 8948 10144 8957 10184
rect 9139 10144 9148 10184
rect 9188 10144 9908 10184
rect 9955 10144 9964 10184
rect 10004 10144 10013 10184
rect 10217 10144 10348 10184
rect 10388 10144 10397 10184
rect 9868 10100 9908 10144
rect 3401 10060 3532 10100
rect 3572 10060 5260 10100
rect 5300 10060 5309 10100
rect 6041 10060 6124 10100
rect 6164 10060 6172 10100
rect 6212 10060 6221 10100
rect 6988 10060 7996 10100
rect 8036 10060 8045 10100
rect 9161 10060 9292 10100
rect 9332 10060 9341 10100
rect 9868 10060 10772 10100
rect 0 10016 90 10036
rect 10732 10016 10772 10060
rect 11750 10016 11840 10036
rect 0 9976 1076 10016
rect 2947 9976 2956 10016
rect 2996 9976 4396 10016
rect 4436 9976 4445 10016
rect 6316 9976 6556 10016
rect 6596 9976 6605 10016
rect 10732 9976 11840 10016
rect 0 9956 90 9976
rect 1036 9932 1076 9976
rect 6316 9932 6356 9976
rect 11750 9956 11840 9976
rect 1036 9892 6356 9932
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 4867 9808 4876 9848
rect 4916 9808 6932 9848
rect 3436 9724 5740 9764
rect 5780 9724 5789 9764
rect 0 9680 90 9700
rect 3436 9680 3476 9724
rect 0 9640 3052 9680
rect 3092 9640 3101 9680
rect 3427 9640 3436 9680
rect 3476 9640 3485 9680
rect 5443 9640 5452 9680
rect 5492 9640 5836 9680
rect 5876 9640 5885 9680
rect 0 9620 90 9640
rect 163 9556 172 9596
rect 212 9556 1180 9596
rect 1220 9556 1229 9596
rect 1315 9556 1324 9596
rect 1364 9556 1564 9596
rect 1604 9556 1613 9596
rect 1708 9556 3580 9596
rect 3620 9556 3629 9596
rect 1289 9472 1420 9512
rect 1460 9472 1469 9512
rect 1708 9428 1748 9556
rect 6892 9512 6932 9808
rect 8170 9640 8179 9680
rect 8219 9640 8620 9680
rect 8660 9640 8669 9680
rect 7084 9556 8332 9596
rect 8372 9556 8381 9596
rect 1795 9472 1804 9512
rect 1844 9472 2956 9512
rect 2996 9472 3005 9512
rect 3811 9472 3820 9512
rect 3860 9472 4780 9512
rect 4820 9472 4829 9512
rect 6115 9472 6124 9512
rect 6164 9472 6173 9512
rect 6883 9472 6892 9512
rect 6932 9472 6941 9512
rect 3244 9428 3284 9437
rect 5260 9428 5300 9437
rect 1123 9388 1132 9428
rect 1172 9388 1748 9428
rect 1987 9388 1996 9428
rect 2036 9388 2284 9428
rect 2324 9388 2333 9428
rect 3284 9388 3820 9428
rect 3860 9388 3869 9428
rect 4003 9388 4012 9428
rect 4052 9388 4061 9428
rect 5129 9388 5260 9428
rect 5300 9388 5740 9428
rect 5780 9388 5789 9428
rect 3244 9379 3284 9388
rect 0 9344 90 9364
rect 0 9304 2956 9344
rect 2996 9304 3005 9344
rect 0 9284 90 9304
rect 4012 9176 4052 9388
rect 5260 9379 5300 9388
rect 4387 9220 4396 9260
rect 4436 9220 5884 9260
rect 5924 9220 5933 9260
rect 2467 9136 2476 9176
rect 2516 9136 4052 9176
rect 0 9008 90 9028
rect 0 8968 748 9008
rect 788 8968 797 9008
rect 1324 8968 1804 9008
rect 1844 8968 2284 9008
rect 2324 8968 2333 9008
rect 0 8948 90 8968
rect 1324 8756 1364 8968
rect 1459 8884 1468 8924
rect 1508 8884 2860 8924
rect 2900 8884 2909 8924
rect 3628 8756 3668 9136
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 6124 8924 6164 9472
rect 6394 9388 6403 9428
rect 6443 9388 6452 9428
rect 6499 9388 6508 9428
rect 6548 9388 6679 9428
rect 6857 9388 6988 9428
rect 7028 9388 7037 9428
rect 6412 9344 6452 9388
rect 7084 9344 7124 9556
rect 9379 9472 9388 9512
rect 9428 9472 10099 9512
rect 10139 9472 10148 9512
rect 7468 9428 7508 9437
rect 8524 9428 8564 9437
rect 7337 9388 7468 9428
rect 7508 9388 7517 9428
rect 7978 9388 7987 9428
rect 8027 9388 8276 9428
rect 8323 9388 8332 9428
rect 8372 9388 8524 9428
rect 9641 9388 9772 9428
rect 9812 9388 9821 9428
rect 10217 9388 10294 9428
rect 10334 9388 10348 9428
rect 10388 9388 10828 9428
rect 10868 9388 10877 9428
rect 7468 9379 7508 9388
rect 6412 9304 7124 9344
rect 8236 8924 8276 9388
rect 8524 9379 8564 9388
rect 11750 9008 11840 9028
rect 10627 8968 10636 9008
rect 10676 8968 11840 9008
rect 11750 8948 11840 8968
rect 3715 8884 3724 8924
rect 3764 8884 4300 8924
rect 4340 8884 4349 8924
rect 6124 8884 6652 8924
rect 6692 8884 6701 8924
rect 6892 8884 7468 8924
rect 7508 8884 7517 8924
rect 8236 8884 8428 8924
rect 8468 8884 8477 8924
rect 6892 8840 6932 8884
rect 5443 8800 5452 8840
rect 5492 8800 5972 8840
rect 6307 8800 6316 8840
rect 6356 8800 6932 8840
rect 6988 8800 10444 8840
rect 10484 8800 10493 8840
rect 5932 8756 5972 8800
rect 6988 8756 7028 8800
rect 1306 8747 1364 8756
rect 1306 8707 1315 8747
rect 1355 8707 1364 8747
rect 1673 8747 1804 8756
rect 1673 8716 1795 8747
rect 1844 8716 2284 8756
rect 2324 8716 2764 8756
rect 2804 8716 2813 8756
rect 3401 8716 3532 8756
rect 3572 8716 3581 8756
rect 3628 8716 4012 8756
rect 4052 8716 4061 8756
rect 5260 8747 5300 8756
rect 1306 8706 1364 8707
rect 1786 8707 1795 8716
rect 1835 8707 1844 8716
rect 1786 8706 1844 8707
rect 3532 8698 3572 8707
rect 5923 8716 5932 8756
rect 5972 8716 5981 8756
rect 6202 8716 6211 8756
rect 6251 8716 6508 8756
rect 6548 8716 6557 8756
rect 6979 8716 6988 8756
rect 7028 8716 7037 8756
rect 8201 8747 8332 8756
rect 8201 8716 8236 8747
rect 0 8672 90 8692
rect 0 8632 556 8672
rect 596 8632 605 8672
rect 1939 8632 1948 8672
rect 1988 8632 2860 8672
rect 2900 8632 2909 8672
rect 0 8612 90 8632
rect 5260 8588 5300 8707
rect 8276 8716 8332 8747
rect 8372 8716 8381 8756
rect 9091 8716 9100 8756
rect 9140 8716 9772 8756
rect 9812 8716 9821 8756
rect 10217 8716 10348 8756
rect 10388 8716 10397 8756
rect 8236 8698 8276 8707
rect 10348 8698 10388 8707
rect 8585 8632 8716 8672
rect 8756 8632 8765 8672
rect 8947 8632 8956 8672
rect 8996 8632 10252 8672
rect 10292 8632 10301 8672
rect 4483 8548 4492 8588
rect 4532 8548 7180 8588
rect 7220 8548 7229 8588
rect 10409 8464 10540 8504
rect 10580 8464 10589 8504
rect 0 8336 90 8356
rect 0 8296 2900 8336
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 0 8276 90 8296
rect 2860 8252 2900 8296
rect 2860 8212 4532 8252
rect 4492 8168 4532 8212
rect 172 8128 2900 8168
rect 2947 8128 2956 8168
rect 2996 8128 3244 8168
rect 3284 8128 3293 8168
rect 4492 8128 6172 8168
rect 6212 8128 6221 8168
rect 8899 8128 8908 8168
rect 8948 8128 9004 8168
rect 9044 8128 9079 8168
rect 0 8000 90 8020
rect 172 8000 212 8128
rect 2860 8084 2900 8128
rect 2860 8044 4724 8084
rect 5635 8044 5644 8084
rect 5684 8044 6068 8084
rect 8297 8044 8332 8084
rect 8372 8044 8428 8084
rect 8468 8044 8477 8084
rect 4684 8000 4724 8044
rect 6028 8000 6068 8044
rect 11750 8000 11840 8020
rect 0 7960 212 8000
rect 931 7960 940 8000
rect 980 7960 1132 8000
rect 1172 7960 1228 8000
rect 1268 7960 1277 8000
rect 4684 7960 5396 8000
rect 6019 7960 6028 8000
rect 6068 7960 6077 8000
rect 6281 7960 6412 8000
rect 6452 7960 6461 8000
rect 6508 7960 6556 8000
rect 6596 7960 6605 8000
rect 6787 7960 6796 8000
rect 6836 7960 7276 8000
rect 7316 7960 7325 8000
rect 7651 7960 7660 8000
rect 7700 7960 8428 8000
rect 8468 7960 8477 8000
rect 10243 7960 10252 8000
rect 10292 7960 11840 8000
rect 0 7940 90 7960
rect 2764 7916 2804 7925
rect 4396 7916 4436 7925
rect 5356 7916 5396 7960
rect 6508 7916 6548 7960
rect 1481 7876 1516 7916
rect 1556 7876 1612 7916
rect 1652 7876 1661 7916
rect 2633 7876 2668 7916
rect 2708 7876 2764 7916
rect 2851 7876 2860 7916
rect 2900 7876 3148 7916
rect 3188 7876 3197 7916
rect 4361 7876 4396 7916
rect 4436 7876 4492 7916
rect 4532 7876 4541 7916
rect 4963 7876 4972 7916
rect 5012 7876 5021 7916
rect 5129 7876 5251 7916
rect 5300 7876 5309 7916
rect 5356 7876 6548 7916
rect 7625 7876 7756 7916
rect 7796 7876 7805 7916
rect 7913 7876 7948 7916
rect 7988 7876 8035 7916
rect 8075 7876 8093 7916
rect 2764 7867 2804 7876
rect 4396 7867 4436 7876
rect 4972 7832 5012 7876
rect 8140 7832 8180 7960
rect 11750 7940 11840 7960
rect 9196 7916 9236 7925
rect 9236 7876 10388 7916
rect 10435 7876 10444 7916
rect 10484 7876 10615 7916
rect 9196 7867 9236 7876
rect 10348 7832 10388 7876
rect 4579 7792 4588 7832
rect 4628 7792 5012 7832
rect 5347 7792 5356 7832
rect 5396 7792 8084 7832
rect 8131 7792 8140 7832
rect 8180 7792 8189 7832
rect 10339 7792 10348 7832
rect 10388 7792 10397 7832
rect 8044 7748 8084 7792
rect 4483 7708 4492 7748
rect 4532 7708 5788 7748
rect 5828 7708 5837 7748
rect 8044 7708 8620 7748
rect 8660 7708 10060 7748
rect 10100 7708 10109 7748
rect 0 7664 90 7684
rect 0 7624 3436 7664
rect 3476 7624 3485 7664
rect 0 7604 90 7624
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 2275 7372 2284 7412
rect 2324 7372 2900 7412
rect 2995 7372 3004 7412
rect 3044 7372 3628 7412
rect 3668 7372 3677 7412
rect 5635 7372 5644 7412
rect 5684 7372 7508 7412
rect 7555 7372 7564 7412
rect 7604 7372 7756 7412
rect 7796 7372 7805 7412
rect 0 7328 90 7348
rect 2860 7328 2900 7372
rect 0 7288 1420 7328
rect 1460 7288 1469 7328
rect 2380 7288 2804 7328
rect 2860 7288 6164 7328
rect 0 7268 90 7288
rect 1193 7204 1228 7244
rect 1268 7204 1324 7244
rect 1364 7204 1373 7244
rect 2380 7160 2420 7288
rect 2764 7244 2804 7288
rect 4300 7244 4340 7288
rect 6124 7244 6164 7288
rect 7468 7244 7508 7372
rect 2476 7235 2668 7244
rect 2516 7204 2668 7235
rect 2708 7204 2717 7244
rect 2764 7235 2964 7244
rect 2764 7204 2851 7235
rect 2476 7186 2516 7195
rect 2842 7195 2851 7204
rect 2891 7204 2964 7235
rect 4291 7204 4300 7244
rect 4340 7204 4349 7244
rect 5548 7235 5740 7244
rect 2891 7195 2900 7204
rect 2842 7194 2900 7195
rect 5588 7204 5740 7235
rect 5780 7204 5789 7244
rect 6115 7204 6124 7244
rect 6164 7204 6173 7244
rect 7171 7204 7180 7244
rect 7220 7235 7412 7244
rect 7220 7204 7372 7235
rect 5548 7186 5588 7195
rect 7468 7204 8524 7244
rect 8564 7204 8620 7244
rect 8660 7204 8724 7244
rect 8812 7204 9388 7244
rect 9428 7235 9812 7244
rect 9428 7204 9772 7235
rect 1699 7120 1708 7160
rect 1748 7120 2420 7160
rect 3523 7120 3532 7160
rect 3572 7120 3724 7160
rect 3764 7120 3773 7160
rect 3907 7120 3916 7160
rect 3956 7120 4148 7160
rect 1507 7036 1516 7076
rect 1556 7036 2668 7076
rect 2708 7036 2717 7076
rect 3043 7036 3052 7076
rect 3092 7036 3292 7076
rect 3332 7036 3341 7076
rect 0 6992 90 7012
rect 0 6952 1804 6992
rect 1844 6952 1853 6992
rect 2947 6952 2956 6992
rect 2996 6952 3676 6992
rect 3716 6952 3725 6992
rect 0 6932 90 6952
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 4108 6740 4148 7120
rect 7372 7076 7412 7195
rect 8812 7160 8852 7204
rect 9772 7186 9812 7195
rect 8201 7120 8332 7160
rect 8372 7120 8381 7160
rect 8428 7120 8852 7160
rect 10339 7120 10348 7160
rect 10388 7120 10540 7160
rect 10580 7120 10589 7160
rect 8428 7076 8468 7120
rect 7372 7036 7564 7076
rect 7604 7036 8468 7076
rect 8707 7036 8716 7076
rect 8756 7036 9964 7076
rect 10004 7036 10013 7076
rect 10505 7036 10588 7076
rect 10628 7036 10636 7076
rect 10676 7036 10685 7076
rect 11750 6992 11840 7012
rect 5609 6952 5740 6992
rect 5780 6952 5789 6992
rect 6019 6952 6028 6992
rect 6068 6952 8092 6992
rect 8132 6952 8141 6992
rect 10588 6952 11840 6992
rect 4012 6700 4148 6740
rect 0 6656 90 6676
rect 4012 6656 4052 6700
rect 10588 6656 10628 6952
rect 11750 6932 11840 6952
rect 0 6616 172 6656
rect 212 6616 221 6656
rect 739 6616 748 6656
rect 788 6616 1372 6656
rect 1412 6616 1421 6656
rect 4003 6616 4012 6656
rect 4052 6616 4061 6656
rect 10579 6616 10588 6656
rect 10628 6616 10637 6656
rect 0 6596 90 6616
rect 3052 6532 3532 6572
rect 3572 6532 3581 6572
rect 7747 6532 7756 6572
rect 7796 6532 10388 6572
rect 1481 6448 1612 6488
rect 1652 6448 1661 6488
rect 3052 6404 3092 6532
rect 10348 6488 10388 6532
rect 3331 6448 3340 6488
rect 3380 6448 4244 6488
rect 4457 6448 4588 6488
rect 4628 6448 4637 6488
rect 9833 6448 9964 6488
rect 10004 6448 10013 6488
rect 10339 6448 10348 6488
rect 10388 6448 10397 6488
rect 4204 6404 4244 6448
rect 5164 6404 5204 6413
rect 7564 6404 7604 6413
rect 1699 6364 1708 6404
rect 1748 6364 1804 6404
rect 1844 6364 1879 6404
rect 2892 6364 2956 6404
rect 2996 6364 3052 6404
rect 3052 6355 3092 6364
rect 3244 6364 4099 6404
rect 4139 6364 4148 6404
rect 4195 6364 4204 6404
rect 4244 6364 4253 6404
rect 4675 6364 4684 6404
rect 4724 6364 4780 6404
rect 4820 6364 4855 6404
rect 5609 6364 5683 6404
rect 5723 6364 5740 6404
rect 5780 6364 5789 6404
rect 6211 6364 6220 6404
rect 6260 6364 6316 6404
rect 6356 6364 6391 6404
rect 7433 6364 7564 6404
rect 7604 6364 7613 6404
rect 0 6320 90 6340
rect 3244 6320 3284 6364
rect 5164 6320 5204 6364
rect 7564 6355 7604 6364
rect 0 6280 2476 6320
rect 2516 6280 2525 6320
rect 3235 6280 3244 6320
rect 3284 6280 3293 6320
rect 4099 6280 4108 6320
rect 4148 6280 7276 6320
rect 7316 6280 7325 6320
rect 10195 6280 10204 6320
rect 10244 6280 11692 6320
rect 11732 6280 11741 6320
rect 0 6260 90 6280
rect 3514 6196 3523 6236
rect 3563 6196 3811 6236
rect 3851 6196 3860 6236
rect 5705 6196 5836 6236
rect 5876 6196 5885 6236
rect 6106 6196 6115 6236
rect 6155 6196 10732 6236
rect 10772 6196 10781 6236
rect 3820 6152 3860 6196
rect 6220 6152 6260 6196
rect 3820 6112 4012 6152
rect 4052 6112 6260 6152
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 0 5984 90 6004
rect 0 5944 1228 5984
rect 1268 5944 1277 5984
rect 0 5924 90 5944
rect 6220 5900 6260 6112
rect 11750 5984 11840 6004
rect 11683 5944 11692 5984
rect 11732 5944 11840 5984
rect 11750 5924 11840 5944
rect 2083 5860 2092 5900
rect 2132 5860 4588 5900
rect 4628 5860 4637 5900
rect 6202 5860 6211 5900
rect 6251 5860 6260 5900
rect 6691 5860 6700 5900
rect 6740 5860 6836 5900
rect 8419 5860 8428 5900
rect 8468 5860 8477 5900
rect 2851 5776 2860 5816
rect 2900 5776 3188 5816
rect 3148 5732 3188 5776
rect 3628 5732 3668 5860
rect 4108 5776 4780 5816
rect 4820 5776 4829 5816
rect 1385 5692 1420 5732
rect 1460 5692 1516 5732
rect 1556 5692 1565 5732
rect 2633 5723 2764 5732
rect 2633 5692 2668 5723
rect 2708 5692 2764 5723
rect 2804 5692 2813 5732
rect 3130 5692 3139 5732
rect 3179 5692 3188 5732
rect 3235 5692 3244 5732
rect 3284 5692 3293 5732
rect 3619 5692 3628 5732
rect 3668 5692 3677 5732
rect 2668 5674 2708 5683
rect 0 5648 90 5668
rect 3244 5648 3284 5692
rect 4108 5648 4148 5776
rect 6796 5732 6836 5860
rect 8428 5816 8468 5860
rect 8428 5776 9044 5816
rect 4204 5723 4300 5732
rect 4244 5692 4300 5723
rect 4340 5692 4375 5732
rect 4553 5692 4588 5732
rect 4628 5723 4724 5732
rect 4628 5692 4684 5723
rect 4204 5674 4244 5683
rect 6682 5692 6691 5732
rect 6731 5692 6740 5732
rect 6787 5692 6796 5732
rect 6836 5692 6845 5732
rect 7049 5692 7180 5732
rect 7220 5692 7229 5732
rect 7625 5692 7756 5732
rect 7796 5692 7805 5732
rect 8201 5723 8332 5732
rect 8201 5692 8236 5723
rect 4684 5674 4724 5683
rect 0 5608 940 5648
rect 980 5608 989 5648
rect 1891 5608 1900 5648
rect 1940 5608 2572 5648
rect 2612 5608 2621 5648
rect 2764 5608 3284 5648
rect 3715 5608 3724 5648
rect 3764 5608 4148 5648
rect 4906 5608 4915 5648
rect 4955 5608 5260 5648
rect 5300 5608 5309 5648
rect 5513 5608 5644 5648
rect 5684 5608 5693 5648
rect 5827 5608 5836 5648
rect 5876 5608 6007 5648
rect 0 5588 90 5608
rect 2764 5564 2804 5608
rect 2179 5524 2188 5564
rect 2228 5524 2804 5564
rect 3724 5480 3764 5608
rect 6700 5564 6740 5692
rect 7756 5674 7796 5683
rect 8276 5692 8332 5723
rect 8372 5692 8381 5732
rect 8489 5723 8620 5732
rect 8489 5692 8611 5723
rect 8660 5692 8669 5732
rect 8755 5692 8764 5732
rect 8804 5692 8812 5732
rect 8852 5692 8935 5732
rect 8236 5674 8276 5683
rect 8602 5683 8611 5692
rect 8651 5683 8660 5692
rect 8602 5682 8660 5683
rect 9004 5648 9044 5776
rect 7145 5608 7276 5648
rect 7316 5608 7325 5648
rect 9004 5608 9292 5648
rect 9332 5608 9341 5648
rect 10339 5608 10348 5648
rect 10388 5608 10397 5648
rect 6067 5524 6076 5564
rect 6116 5524 6412 5564
rect 6452 5524 6461 5564
rect 6691 5524 6700 5564
rect 6740 5524 6749 5564
rect 7075 5524 7084 5564
rect 7124 5524 9052 5564
rect 9092 5524 9101 5564
rect 835 5440 844 5480
rect 884 5440 3764 5480
rect 4771 5440 4780 5480
rect 4820 5440 5020 5480
rect 5060 5440 5069 5480
rect 5164 5440 5404 5480
rect 5444 5440 5453 5480
rect 5164 5396 5204 5440
rect 4780 5356 5204 5396
rect 0 5312 90 5332
rect 0 5272 1324 5312
rect 1364 5272 1373 5312
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 4579 5272 4588 5312
rect 4628 5272 4637 5312
rect 0 5252 90 5272
rect 4588 5228 4628 5272
rect 4012 5188 4628 5228
rect 4012 5144 4052 5188
rect 4003 5104 4012 5144
rect 4052 5104 4061 5144
rect 4780 5060 4820 5356
rect 5635 5272 5644 5312
rect 5684 5272 9004 5312
rect 9044 5272 9053 5312
rect 10348 5228 10388 5608
rect 10579 5440 10588 5480
rect 10628 5440 11692 5480
rect 11732 5440 11741 5480
rect 4963 5188 4972 5228
rect 5012 5188 10388 5228
rect 8297 5104 8332 5144
rect 8372 5104 8428 5144
rect 8468 5104 8477 5144
rect 2860 5020 4820 5060
rect 7468 5020 8620 5060
rect 8660 5020 8669 5060
rect 0 4976 90 4996
rect 2860 4976 2900 5020
rect 0 4936 2900 4976
rect 4745 4936 4876 4976
rect 4916 4936 4925 4976
rect 6154 4936 6163 4976
rect 6203 4936 6508 4976
rect 6548 4936 6557 4976
rect 0 4916 90 4936
rect 3820 4892 3860 4901
rect 5452 4892 5492 4901
rect 7468 4892 7508 5020
rect 11750 4976 11840 4996
rect 11683 4936 11692 4976
rect 11732 4936 11840 4976
rect 11750 4916 11840 4936
rect 8236 4892 8276 4901
rect 1507 4852 1516 4892
rect 1556 4852 1720 4892
rect 1760 4852 1769 4892
rect 1879 4852 1888 4892
rect 1928 4852 2036 4892
rect 2537 4852 2572 4892
rect 2612 4852 2668 4892
rect 2708 4852 2717 4892
rect 2851 4852 2860 4892
rect 2900 4852 3820 4892
rect 3907 4852 3916 4892
rect 3956 4852 4366 4892
rect 4406 4852 4415 4892
rect 4480 4852 4489 4892
rect 4529 4852 4588 4892
rect 4628 4852 4669 4892
rect 4841 4852 4972 4892
rect 5012 4852 5021 4892
rect 5923 4852 5932 4892
rect 5980 4852 6103 4892
rect 6979 4852 6988 4892
rect 7028 4852 7508 4892
rect 8105 4852 8236 4892
rect 8276 4852 8285 4892
rect 1996 4808 2036 4852
rect 3820 4843 3860 4852
rect 5452 4808 5492 4852
rect 8236 4843 8276 4852
rect 1546 4768 1555 4808
rect 1595 4768 1900 4808
rect 1940 4768 1949 4808
rect 1996 4768 2228 4808
rect 5452 4768 7756 4808
rect 7796 4768 7805 4808
rect 1961 4684 2044 4724
rect 2084 4684 2092 4724
rect 2132 4684 2141 4724
rect 0 4640 90 4660
rect 2188 4640 2228 4768
rect 2563 4684 2572 4724
rect 2612 4684 3956 4724
rect 3916 4640 3956 4684
rect 4108 4684 6268 4724
rect 6308 4684 6317 4724
rect 6682 4684 6691 4724
rect 6731 4684 6740 4724
rect 4108 4640 4148 4684
rect 6700 4640 6740 4684
rect 0 4600 460 4640
rect 500 4600 509 4640
rect 2188 4600 2900 4640
rect 3916 4600 4148 4640
rect 4579 4600 4588 4640
rect 4628 4600 6740 4640
rect 0 4580 90 4600
rect 2860 4556 2900 4600
rect 2860 4516 4724 4556
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 4684 4472 4724 4516
rect 6700 4472 6740 4600
rect 1228 4432 1612 4472
rect 1652 4432 4588 4472
rect 4628 4432 4637 4472
rect 4684 4432 6220 4472
rect 6260 4432 6269 4472
rect 6700 4432 7412 4472
rect 1228 4388 1268 4432
rect 7372 4388 7412 4432
rect 1123 4348 1132 4388
rect 1172 4348 1219 4388
rect 1259 4348 1303 4388
rect 1507 4348 1516 4388
rect 1556 4348 2228 4388
rect 3619 4348 3628 4388
rect 3668 4348 3916 4388
rect 3956 4348 3965 4388
rect 6691 4348 6700 4388
rect 6740 4348 7180 4388
rect 7220 4348 7229 4388
rect 7354 4348 7363 4388
rect 7403 4348 7412 4388
rect 0 4304 90 4324
rect 0 4264 844 4304
rect 884 4264 893 4304
rect 1769 4264 1852 4304
rect 1892 4264 1900 4304
rect 1940 4264 1949 4304
rect 0 4244 90 4264
rect 2188 4220 2228 4348
rect 2860 4264 3572 4304
rect 5443 4264 5452 4304
rect 5492 4264 5932 4304
rect 5972 4264 5981 4304
rect 9929 4264 10051 4304
rect 10100 4264 10109 4304
rect 1690 4211 1748 4220
rect 1690 4171 1699 4211
rect 1739 4171 1748 4211
rect 2179 4180 2188 4220
rect 2228 4180 2237 4220
rect 1690 4170 1748 4171
rect 1708 4136 1748 4170
rect 2860 4136 2900 4264
rect 3532 4220 3572 4264
rect 1708 4096 2188 4136
rect 2228 4096 2668 4136
rect 2708 4096 2900 4136
rect 3436 4211 3476 4220
rect 3532 4180 4012 4220
rect 4052 4180 4061 4220
rect 5259 4180 5268 4220
rect 5308 4180 5396 4220
rect 5731 4180 5740 4220
rect 5780 4180 6220 4220
rect 6260 4180 6269 4220
rect 6988 4211 8236 4220
rect 3436 4052 3476 4171
rect 5356 4052 5396 4180
rect 7028 4180 8236 4211
rect 8276 4180 8285 4220
rect 10435 4180 10444 4220
rect 10484 4180 11252 4220
rect 6988 4052 7028 4171
rect 3436 4012 7028 4052
rect 0 3968 90 3988
rect 11212 3968 11252 4180
rect 11750 3968 11840 3988
rect 0 3928 1132 3968
rect 1172 3928 1181 3968
rect 11212 3928 11840 3968
rect 0 3908 90 3928
rect 11750 3908 11840 3928
rect 172 3760 2900 3800
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 0 3632 90 3652
rect 172 3632 212 3760
rect 1027 3676 1036 3716
rect 1076 3676 1988 3716
rect 0 3592 212 3632
rect 0 3572 90 3592
rect 1948 3548 1988 3676
rect 2860 3632 2900 3760
rect 2860 3592 3100 3632
rect 3140 3592 3149 3632
rect 3427 3592 3436 3632
rect 3476 3592 3484 3632
rect 3524 3592 3607 3632
rect 3724 3592 11596 3632
rect 11636 3592 11645 3632
rect 1411 3508 1420 3548
rect 1460 3508 1564 3548
rect 1604 3508 1613 3548
rect 1939 3508 1948 3548
rect 1988 3508 1997 3548
rect 2860 3508 3244 3548
rect 3284 3508 3293 3548
rect 2860 3464 2900 3508
rect 3724 3464 3764 3592
rect 5731 3508 5740 3548
rect 5780 3508 10388 3548
rect 10348 3464 10388 3508
rect 1603 3424 1612 3464
rect 1652 3424 1804 3464
rect 1844 3424 1853 3464
rect 2057 3424 2188 3464
rect 2228 3424 2237 3464
rect 2323 3424 2332 3464
rect 2372 3424 2381 3464
rect 2563 3424 2572 3464
rect 2612 3424 2900 3464
rect 2947 3424 2956 3464
rect 2996 3424 3005 3464
rect 3209 3424 3340 3464
rect 3380 3424 3389 3464
rect 3715 3424 3724 3464
rect 3764 3424 3773 3464
rect 3907 3424 3916 3464
rect 3956 3424 4108 3464
rect 4148 3424 4157 3464
rect 4457 3424 4492 3464
rect 4532 3424 4588 3464
rect 4628 3424 4780 3464
rect 4820 3424 5548 3464
rect 5588 3424 5644 3464
rect 5684 3424 5932 3464
rect 5972 3424 6508 3464
rect 6548 3424 6557 3464
rect 6787 3424 6796 3464
rect 6836 3424 6988 3464
rect 7028 3424 7084 3464
rect 7124 3424 7159 3464
rect 10339 3424 10348 3464
rect 10388 3424 10397 3464
rect 2332 3380 2372 3424
rect 1219 3340 1228 3380
rect 1268 3340 2372 3380
rect 2956 3380 2996 3424
rect 2956 3340 10924 3380
rect 10964 3340 10973 3380
rect 0 3296 90 3316
rect 0 3256 1036 3296
rect 1076 3256 1085 3296
rect 1315 3256 1324 3296
rect 1364 3256 2716 3296
rect 2756 3256 2765 3296
rect 0 3236 90 3256
rect 1306 3172 1315 3212
rect 1355 3172 1420 3212
rect 1460 3172 1495 3212
rect 3427 3172 3436 3212
rect 3476 3172 3907 3212
rect 3947 3172 3956 3212
rect 4282 3172 4291 3212
rect 4331 3172 5155 3212
rect 5195 3172 5443 3212
rect 5483 3172 6307 3212
rect 6347 3172 6787 3212
rect 6827 3172 6836 3212
rect 10579 3172 10588 3212
rect 10628 3172 11692 3212
rect 11732 3172 11741 3212
rect 1420 3128 1460 3172
rect 4300 3128 4340 3172
rect 1420 3088 4340 3128
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 0 2960 90 2980
rect 0 2920 1364 2960
rect 0 2900 90 2920
rect 1324 2876 1364 2920
rect 5356 2876 5396 3172
rect 11750 2960 11840 2980
rect 11683 2920 11692 2960
rect 11732 2920 11840 2960
rect 11750 2900 11840 2920
rect 163 2836 172 2876
rect 212 2836 1180 2876
rect 1220 2836 1229 2876
rect 1324 2836 2716 2876
rect 2756 2836 2765 2876
rect 3427 2836 3436 2876
rect 3476 2836 3619 2876
rect 3659 2836 3907 2876
rect 3947 2836 3956 2876
rect 5050 2836 5059 2876
rect 5099 2836 5740 2876
rect 5780 2836 5827 2876
rect 5867 2836 5876 2876
rect 1123 2752 1132 2792
rect 1172 2752 2332 2792
rect 2372 2752 2381 2792
rect 2860 2752 4396 2792
rect 4436 2752 4684 2792
rect 4724 2752 5260 2792
rect 5300 2752 5548 2792
rect 5588 2752 6124 2792
rect 6164 2752 6412 2792
rect 6452 2752 6508 2792
rect 6548 2752 6612 2792
rect 2860 2708 2900 2752
rect 1481 2668 1612 2708
rect 1652 2668 2900 2708
rect 2956 2668 4492 2708
rect 4532 2668 4541 2708
rect 0 2624 90 2644
rect 2956 2624 2996 2668
rect 0 2584 1172 2624
rect 1385 2584 1420 2624
rect 1460 2584 1516 2624
rect 1556 2584 1565 2624
rect 1795 2584 1804 2624
rect 1844 2584 1948 2624
rect 1988 2584 1997 2624
rect 2179 2584 2188 2624
rect 2228 2584 2359 2624
rect 2441 2584 2572 2624
rect 2612 2584 2621 2624
rect 2947 2584 2956 2624
rect 2996 2584 3005 2624
rect 3331 2584 3340 2624
rect 3380 2584 3389 2624
rect 4265 2584 4396 2624
rect 4436 2584 4445 2624
rect 10217 2584 10252 2624
rect 10292 2584 10348 2624
rect 10388 2584 10397 2624
rect 0 2564 90 2584
rect 1132 2540 1172 2584
rect 3340 2540 3380 2584
rect 1132 2500 1900 2540
rect 1940 2500 1949 2540
rect 3340 2500 7756 2540
rect 7796 2500 7805 2540
rect 1516 2416 3100 2456
rect 3140 2416 3149 2456
rect 10579 2416 10588 2456
rect 10628 2416 11692 2456
rect 11732 2416 11741 2456
rect 0 2288 90 2308
rect 1516 2288 1556 2416
rect 0 2248 1556 2288
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 0 2228 90 2248
rect 1804 2164 6124 2204
rect 6164 2164 6173 2204
rect 451 2080 460 2120
rect 500 2080 1180 2120
rect 1220 2080 1229 2120
rect 547 1996 556 2036
rect 596 1996 1564 2036
rect 1604 1996 1613 2036
rect 1804 1952 1844 2164
rect 1891 2080 1900 2120
rect 1940 2080 2332 2120
rect 2372 2080 2381 2120
rect 2467 2080 2476 2120
rect 2516 2080 2716 2120
rect 2756 2080 2765 2120
rect 3244 2080 6028 2120
rect 6068 2080 6077 2120
rect 8707 2080 8716 2120
rect 8756 2080 10051 2120
rect 10091 2080 10100 2120
rect 3244 2036 3284 2080
rect 2572 1996 3284 2036
rect 3340 1996 4588 2036
rect 4628 1996 4637 2036
rect 2572 1952 2612 1996
rect 3340 1952 3380 1996
rect 11750 1952 11840 1972
rect 1289 1912 1420 1952
rect 1460 1912 1469 1952
rect 1795 1912 1804 1952
rect 1844 1912 1853 1952
rect 2179 1912 2188 1952
rect 2228 1912 2237 1952
rect 2563 1912 2572 1952
rect 2612 1912 2621 1952
rect 2825 1912 2956 1952
rect 2996 1912 3005 1952
rect 3331 1912 3340 1952
rect 3380 1912 3389 1952
rect 3593 1912 3724 1952
rect 3764 1912 3773 1952
rect 4265 1912 4300 1952
rect 4340 1912 4396 1952
rect 4436 1912 4588 1952
rect 4628 1912 5452 1952
rect 5492 1912 5501 1952
rect 11683 1912 11692 1952
rect 11732 1912 11840 1952
rect 2188 1868 2228 1912
rect 11750 1892 11840 1912
rect 1027 1828 1036 1868
rect 1076 1828 2132 1868
rect 2188 1828 4780 1868
rect 4820 1828 4829 1868
rect 5155 1828 5164 1868
rect 5204 1828 5548 1868
rect 5588 1828 5597 1868
rect 10313 1828 10444 1868
rect 10484 1828 10493 1868
rect 2092 1784 2132 1828
rect 931 1744 940 1784
rect 980 1744 1948 1784
rect 1988 1744 1997 1784
rect 2092 1744 3100 1784
rect 3140 1744 3149 1784
rect 3427 1744 3436 1784
rect 3476 1744 4012 1784
rect 4052 1744 5740 1784
rect 5780 1744 6028 1784
rect 6068 1744 6077 1784
rect 2860 1660 3484 1700
rect 3524 1660 3533 1700
rect 4858 1660 4867 1700
rect 4907 1660 4916 1700
rect 2860 1616 2900 1660
rect 835 1576 844 1616
rect 884 1576 2900 1616
rect 4876 1616 4916 1660
rect 4876 1576 5740 1616
rect 5780 1576 5789 1616
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 7939 1408 7948 1448
rect 7988 1408 8908 1448
rect 8948 1408 8957 1448
rect 11750 944 11840 964
rect 10435 904 10444 944
rect 10484 904 11840 944
rect 11750 884 11840 904
<< via2 >>
rect 10252 46264 10292 46304
rect 4928 45340 4968 45380
rect 5010 45340 5050 45380
rect 5092 45340 5132 45380
rect 5174 45340 5214 45380
rect 5256 45340 5296 45380
rect 5644 45256 5684 45296
rect 11020 45256 11060 45296
rect 2380 45172 2420 45212
rect 3916 45172 3956 45212
rect 4300 45172 4340 45212
rect 4684 45172 4724 45212
rect 5356 45172 5396 45212
rect 5548 45172 5588 45212
rect 5836 45172 5876 45212
rect 6220 45172 6260 45212
rect 6604 45172 6644 45212
rect 6988 45172 7028 45212
rect 7372 45172 7412 45212
rect 7756 45172 7796 45212
rect 8140 45172 8180 45212
rect 2092 45088 2132 45128
rect 5452 45088 5492 45128
rect 1324 45004 1355 45044
rect 1355 45004 1364 45044
rect 2668 45035 2708 45044
rect 2668 45004 2699 45035
rect 2699 45004 2708 45035
rect 3340 45004 3380 45044
rect 3148 44920 3188 44960
rect 2284 44836 2324 44876
rect 748 44752 788 44792
rect 6124 45004 6164 45044
rect 8524 45172 8564 45212
rect 8908 45172 8948 45212
rect 9292 45172 9332 45212
rect 9676 45172 9716 45212
rect 4972 44920 5012 44960
rect 5356 44920 5396 44960
rect 5740 44920 5780 44960
rect 6508 44920 6548 44960
rect 7276 44920 7316 44960
rect 8044 44920 8084 44960
rect 9580 44920 9620 44960
rect 9964 44920 10004 44960
rect 10348 44920 10388 44960
rect 5260 44836 5300 44876
rect 7756 44836 7796 44876
rect 7948 44836 7988 44876
rect 11692 44752 11732 44792
rect 6796 44668 6836 44708
rect 2668 44584 2708 44624
rect 3688 44584 3728 44624
rect 3770 44584 3810 44624
rect 3852 44584 3892 44624
rect 3934 44584 3974 44624
rect 4016 44584 4056 44624
rect 3052 44500 3092 44540
rect 5356 44500 5396 44540
rect 5164 44416 5204 44456
rect 6124 44416 6164 44456
rect 6508 44416 6548 44456
rect 6796 44416 6836 44456
rect 7276 44416 7316 44456
rect 7756 44416 7796 44456
rect 9580 44416 9620 44456
rect 10252 44416 10292 44456
rect 11020 44416 11060 44456
rect 172 44332 212 44372
rect 5260 44332 5300 44372
rect 7948 44332 7988 44372
rect 9964 44332 10004 44372
rect 76 44248 116 44288
rect 2476 44248 2516 44288
rect 2956 44248 2996 44288
rect 4684 44248 4724 44288
rect 6316 44248 6356 44288
rect 6796 44248 6836 44288
rect 7276 44248 7316 44288
rect 7660 44248 7700 44288
rect 9004 44248 9044 44288
rect 9388 44248 9428 44288
rect 10252 44248 10292 44288
rect 11692 44248 11732 44288
rect 652 44164 692 44204
rect 6412 44164 6452 44204
rect 556 43996 596 44036
rect 76 43912 116 43952
rect 4972 44080 5012 44120
rect 6220 44080 6260 44120
rect 7180 44080 7220 44120
rect 8044 44080 8084 44120
rect 8236 44080 8276 44120
rect 1900 43996 1940 44036
rect 3244 43996 3275 44036
rect 3275 43996 3284 44036
rect 4492 43996 4532 44036
rect 5836 43996 5876 44036
rect 7852 43996 7892 44036
rect 8140 43996 8180 44036
rect 4684 43912 4724 43952
rect 5356 43912 5396 43952
rect 6316 43912 6356 43952
rect 4928 43828 4968 43868
rect 5010 43828 5050 43868
rect 5092 43828 5132 43868
rect 5174 43828 5214 43868
rect 5256 43828 5296 43868
rect 5644 43828 5684 43868
rect 4396 43744 4436 43784
rect 5740 43744 5780 43784
rect 6796 43744 6836 43784
rect 10828 43744 10868 43784
rect 2476 43660 2507 43700
rect 2507 43660 2516 43700
rect 3724 43660 3764 43700
rect 7660 43660 7700 43700
rect 9004 43660 9035 43700
rect 9035 43660 9044 43700
rect 9388 43660 9419 43700
rect 9419 43660 9428 43700
rect 3436 43576 3476 43616
rect 4684 43576 4724 43616
rect 5356 43576 5396 43616
rect 7276 43576 7316 43616
rect 7564 43576 7604 43616
rect 8140 43576 8180 43616
rect 1804 43492 1835 43532
rect 1835 43492 1844 43532
rect 1708 43408 1748 43448
rect 4300 43492 4340 43532
rect 5836 43492 5876 43532
rect 10348 43492 10388 43532
rect 4204 43408 4244 43448
rect 4588 43408 4628 43448
rect 8236 43408 8276 43448
rect 9196 43408 9236 43448
rect 10540 43408 10580 43448
rect 3148 43324 3188 43364
rect 3436 43324 3476 43364
rect 3724 43324 3764 43364
rect 4780 43324 4820 43364
rect 8716 43324 8756 43364
rect 940 43240 980 43280
rect 7180 43240 7220 43280
rect 10924 43240 10964 43280
rect 5836 43156 5876 43196
rect 7084 43156 7124 43196
rect 3688 43072 3728 43112
rect 3770 43072 3810 43112
rect 3852 43072 3892 43112
rect 3934 43072 3974 43112
rect 4016 43072 4056 43112
rect 4492 43072 4532 43112
rect 9868 43072 9908 43112
rect 7372 42988 7412 43028
rect 1324 42904 1364 42944
rect 3532 42904 3572 42944
rect 4780 42904 4820 42944
rect 5548 42904 5588 42944
rect 5932 42904 5972 42944
rect 7468 42820 7508 42860
rect 1996 42736 2036 42776
rect 3532 42736 3572 42776
rect 6988 42736 7028 42776
rect 8236 42736 8276 42776
rect 9964 42736 10004 42776
rect 10348 42736 10388 42776
rect 1324 42652 1355 42692
rect 1355 42652 1364 42692
rect 1516 42652 1556 42692
rect 2188 42652 2228 42692
rect 4588 42652 4628 42692
rect 5548 42652 5588 42692
rect 9388 42652 9428 42692
rect 1804 42568 1844 42608
rect 2380 42568 2420 42608
rect 6220 42568 6260 42608
rect 6700 42568 6740 42608
rect 7564 42568 7604 42608
rect 7852 42568 7892 42608
rect 9196 42568 9236 42608
rect 11692 42568 11732 42608
rect 3916 42484 3956 42524
rect 4588 42484 4628 42524
rect 5932 42484 5963 42524
rect 5963 42484 5972 42524
rect 6508 42484 6548 42524
rect 6892 42484 6932 42524
rect 7276 42484 7316 42524
rect 8812 42484 8852 42524
rect 9964 42484 10004 42524
rect 11212 42484 11252 42524
rect 3244 42400 3284 42440
rect 5836 42400 5876 42440
rect 6220 42400 6260 42440
rect 4780 42316 4820 42356
rect 4928 42316 4968 42356
rect 5010 42316 5050 42356
rect 5092 42316 5132 42356
rect 5174 42316 5214 42356
rect 5256 42316 5296 42356
rect 652 42232 692 42272
rect 4684 42232 4724 42272
rect 9388 42232 9428 42272
rect 11692 42232 11732 42272
rect 3148 42148 3188 42188
rect 4492 42148 4532 42188
rect 5644 42148 5684 42188
rect 7948 42148 7988 42188
rect 8428 42148 8459 42188
rect 8459 42148 8468 42188
rect 8716 42148 8756 42188
rect 1036 42064 1076 42104
rect 3532 42064 3572 42104
rect 5548 42064 5588 42104
rect 7180 42064 7220 42104
rect 9100 42064 9140 42104
rect 10060 42064 10100 42104
rect 268 41980 308 42020
rect 3148 41980 3188 42020
rect 4780 41980 4820 42020
rect 6316 41980 6356 42020
rect 9292 41980 9332 42020
rect 9964 41980 10004 42020
rect 11404 41980 11444 42020
rect 4588 41896 4628 41936
rect 5452 41896 5492 41936
rect 7756 41896 7796 41936
rect 10348 41896 10388 41936
rect 11116 41896 11156 41936
rect 3052 41812 3092 41852
rect 7852 41812 7892 41852
rect 9100 41812 9140 41852
rect 11692 41812 11732 41852
rect 1804 41728 1844 41768
rect 9196 41728 9236 41768
rect 2188 41560 2228 41600
rect 3688 41560 3728 41600
rect 3770 41560 3810 41600
rect 3852 41560 3892 41600
rect 3934 41560 3974 41600
rect 4016 41560 4056 41600
rect 1516 41308 1556 41348
rect 5836 41308 5876 41348
rect 6316 41308 6356 41348
rect 3148 41224 3188 41264
rect 460 41140 500 41180
rect 1420 41140 1460 41180
rect 3436 41140 3476 41180
rect 3532 41056 3572 41096
rect 1612 40972 1652 41012
rect 3052 40972 3092 41012
rect 4684 40972 4724 41012
rect 9964 41224 10004 41264
rect 10636 41224 10676 41264
rect 11692 41224 11732 41264
rect 1324 40888 1364 40928
rect 7660 41140 7700 41180
rect 9292 41140 9332 41180
rect 4928 40804 4968 40844
rect 5010 40804 5050 40844
rect 5092 40804 5132 40844
rect 5174 40804 5214 40844
rect 5256 40804 5296 40844
rect 5740 40972 5780 41012
rect 6892 40972 6932 41012
rect 11020 41056 11060 41096
rect 9484 40972 9524 41012
rect 10060 40972 10100 41012
rect 11500 40972 11540 41012
rect 6124 40888 6164 40928
rect 7084 40636 7124 40676
rect 1804 40552 1844 40592
rect 1324 40468 1355 40508
rect 1355 40468 1364 40508
rect 2380 40468 2420 40508
rect 4108 40468 4148 40508
rect 4396 40468 4436 40508
rect 5356 40499 5396 40508
rect 5356 40468 5396 40499
rect 6124 40468 6164 40508
rect 7948 40468 7988 40508
rect 8620 40468 8660 40508
rect 8908 40499 8948 40508
rect 8908 40468 8948 40499
rect 4300 40384 4340 40424
rect 5836 40384 5876 40424
rect 7660 40384 7700 40424
rect 8524 40384 8564 40424
rect 9964 40384 10004 40424
rect 10348 40384 10388 40424
rect 1132 40300 1172 40340
rect 2572 40300 2612 40340
rect 3436 40300 3476 40340
rect 6124 40300 6164 40340
rect 8332 40300 8372 40340
rect 1036 40216 1076 40256
rect 4300 40216 4340 40256
rect 7948 40216 7988 40256
rect 8908 40216 8948 40256
rect 10924 40216 10964 40256
rect 3688 40048 3728 40088
rect 3770 40048 3810 40088
rect 3852 40048 3892 40088
rect 3934 40048 3974 40088
rect 4016 40048 4056 40088
rect 268 39880 308 39920
rect 4012 39880 4052 39920
rect 1516 39796 1556 39836
rect 4108 39712 4148 39752
rect 11692 39880 11732 39920
rect 8044 39796 8084 39836
rect 6028 39712 6068 39752
rect 8428 39712 8468 39752
rect 9868 39712 9908 39752
rect 1420 39628 1460 39668
rect 2668 39628 2708 39668
rect 3052 39628 3092 39668
rect 4300 39628 4340 39668
rect 4684 39628 4724 39668
rect 6124 39628 6164 39668
rect 844 39544 884 39584
rect 2956 39544 2996 39584
rect 4492 39544 4532 39584
rect 2860 39460 2900 39500
rect 4396 39460 4436 39500
rect 4780 39460 4820 39500
rect 6508 39460 6548 39500
rect 7852 39628 7892 39668
rect 8140 39628 8180 39668
rect 8620 39628 8660 39668
rect 8908 39628 8948 39668
rect 9484 39628 9492 39668
rect 9492 39628 9524 39668
rect 6892 39460 6923 39500
rect 6923 39460 6932 39500
rect 7276 39460 7316 39500
rect 10156 39460 10196 39500
rect 10444 39460 10484 39500
rect 3436 39376 3476 39416
rect 1324 39208 1364 39248
rect 2572 39292 2612 39332
rect 3820 39292 3860 39332
rect 4300 39292 4340 39332
rect 4780 39292 4820 39332
rect 4928 39292 4968 39332
rect 5010 39292 5050 39332
rect 5092 39292 5132 39332
rect 5174 39292 5214 39332
rect 5256 39292 5296 39332
rect 5356 39292 5396 39332
rect 5548 39292 5588 39332
rect 7948 39208 7988 39248
rect 11212 39208 11252 39248
rect 6796 39124 6836 39164
rect 3148 39040 3188 39080
rect 3820 39040 3860 39080
rect 6124 39040 6164 39080
rect 7468 39040 7508 39080
rect 1804 38956 1844 38996
rect 2668 38987 2708 38996
rect 2668 38956 2708 38987
rect 3052 38987 3092 38996
rect 3052 38956 3083 38987
rect 3083 38956 3092 38987
rect 3532 38987 3572 38996
rect 3532 38956 3563 38987
rect 3563 38956 3572 38987
rect 4012 38956 4052 38996
rect 4300 38956 4340 38996
rect 3628 38872 3668 38912
rect 4204 38872 4244 38912
rect 8716 38956 8756 38996
rect 8908 38956 8948 38996
rect 9772 38987 9812 38996
rect 9772 38956 9812 38987
rect 5836 38872 5876 38912
rect 7660 38872 7700 38912
rect 8428 38872 8468 38912
rect 10444 38872 10484 38912
rect 8524 38788 8564 38828
rect 7564 38704 7604 38744
rect 8620 38704 8660 38744
rect 9292 38704 9332 38744
rect 6028 38620 6068 38660
rect 3688 38536 3728 38576
rect 3770 38536 3810 38576
rect 3852 38536 3892 38576
rect 3934 38536 3974 38576
rect 4016 38536 4056 38576
rect 5356 38536 5396 38576
rect 8140 38536 8180 38576
rect 8716 38536 8756 38576
rect 2476 38452 2516 38492
rect 6124 38452 6164 38492
rect 8428 38368 8468 38408
rect 9772 38368 9812 38408
rect 5356 38284 5396 38324
rect 5740 38284 5780 38324
rect 1516 38200 1556 38240
rect 9292 38200 9332 38240
rect 10732 38200 10772 38240
rect 11020 38200 11060 38240
rect 844 38116 884 38156
rect 1420 38116 1460 38156
rect 2476 38116 2516 38156
rect 4300 38116 4340 38156
rect 5740 38116 5780 38156
rect 6028 38116 6068 38156
rect 7084 38116 7124 38156
rect 8620 38116 8660 38156
rect 9868 38116 9908 38156
rect 10924 38116 10964 38156
rect 1612 38032 1643 38072
rect 1643 38032 1652 38072
rect 5836 38032 5876 38072
rect 1996 37864 2036 37904
rect 2380 37864 2420 37904
rect 748 37696 788 37736
rect 1228 37612 1268 37652
rect 364 37528 404 37568
rect 1036 37528 1076 37568
rect 4928 37780 4968 37820
rect 5010 37780 5050 37820
rect 5092 37780 5132 37820
rect 5174 37780 5214 37820
rect 5256 37780 5296 37820
rect 6316 37948 6356 37988
rect 9004 37864 9044 37904
rect 5740 37612 5780 37652
rect 6028 37612 6068 37652
rect 6892 37612 6932 37652
rect 7660 37528 7700 37568
rect 1324 37444 1355 37484
rect 1355 37444 1364 37484
rect 2284 37444 2324 37484
rect 2764 37444 2804 37484
rect 2956 37475 2996 37484
rect 2956 37444 2987 37475
rect 2987 37444 2996 37475
rect 3244 37444 3284 37484
rect 5068 37475 5108 37484
rect 5068 37444 5108 37475
rect 4300 37360 4340 37400
rect 6124 37444 6164 37484
rect 7756 37475 7796 37484
rect 7756 37444 7787 37475
rect 7787 37444 7796 37475
rect 7948 37444 7988 37484
rect 9004 37444 9044 37484
rect 9868 37444 9908 37484
rect 4780 37360 4820 37400
rect 8812 37360 8852 37400
rect 4204 37276 4244 37316
rect 5644 37276 5684 37316
rect 7084 37276 7124 37316
rect 9580 37276 9620 37316
rect 1516 37192 1556 37232
rect 8716 37192 8756 37232
rect 11116 37192 11156 37232
rect 5548 37108 5588 37148
rect 3688 37024 3728 37064
rect 3770 37024 3810 37064
rect 3852 37024 3892 37064
rect 3934 37024 3974 37064
rect 4016 37024 4056 37064
rect 8812 37024 8852 37064
rect 10060 37024 10100 37064
rect 2284 36940 2324 36980
rect 8524 36940 8564 36980
rect 1324 36856 1364 36896
rect 4876 36856 4916 36896
rect 3532 36772 3572 36812
rect 4108 36772 4148 36812
rect 5548 36772 5588 36812
rect 5740 36772 5780 36812
rect 460 36604 500 36644
rect 844 36604 884 36644
rect 4876 36688 4916 36728
rect 5644 36688 5684 36728
rect 9964 36688 10004 36728
rect 11308 36688 11348 36728
rect 2572 36604 2612 36644
rect 2476 36436 2516 36476
rect 3532 36436 3572 36476
rect 4204 36604 4244 36644
rect 4588 36604 4596 36644
rect 4596 36604 4628 36644
rect 5548 36604 5588 36644
rect 5740 36604 5780 36644
rect 8140 36604 8180 36644
rect 7180 36520 7220 36560
rect 7372 36520 7412 36560
rect 4300 36436 4340 36476
rect 7756 36436 7796 36476
rect 4396 36352 4436 36392
rect 4928 36268 4968 36308
rect 5010 36268 5050 36308
rect 5092 36268 5132 36308
rect 5174 36268 5214 36308
rect 5256 36268 5296 36308
rect 3052 36184 3092 36224
rect 6220 36184 6260 36224
rect 6892 36184 6932 36224
rect 11020 36520 11060 36560
rect 9484 36436 9524 36476
rect 11116 36436 11156 36476
rect 11500 36184 11540 36224
rect 4204 36100 4244 36140
rect 5644 36100 5684 36140
rect 10060 36100 10100 36140
rect 10828 36100 10868 36140
rect 1996 36016 2036 36056
rect 2572 36016 2612 36056
rect 5740 36016 5780 36056
rect 9484 36016 9524 36056
rect 460 35932 500 35972
rect 1324 35932 1364 35972
rect 2668 35932 2708 35972
rect 3532 35932 3572 35972
rect 3436 35848 3476 35888
rect 1420 35764 1460 35804
rect 4588 35764 4628 35804
rect 6028 35932 6068 35972
rect 4780 35848 4820 35888
rect 5260 35848 5300 35888
rect 8524 35932 8564 35972
rect 9004 35963 9044 35972
rect 9004 35932 9044 35963
rect 10060 35932 10100 35972
rect 11500 35932 11540 35972
rect 6700 35848 6740 35888
rect 5164 35764 5204 35804
rect 7180 35764 7220 35804
rect 2956 35680 2996 35720
rect 1228 35512 1268 35552
rect 3688 35512 3728 35552
rect 3770 35512 3810 35552
rect 3852 35512 3892 35552
rect 3934 35512 3974 35552
rect 4016 35512 4056 35552
rect 3052 35428 3092 35468
rect 2188 35344 2228 35384
rect 2668 35344 2708 35384
rect 3724 35344 3764 35384
rect 1036 35176 1076 35216
rect 1804 35176 1844 35216
rect 2284 35176 2324 35216
rect 3052 35176 3092 35216
rect 3724 35176 3764 35216
rect 9196 35428 9236 35468
rect 5164 35344 5204 35384
rect 11596 35344 11636 35384
rect 6028 35176 6068 35216
rect 8140 35176 8180 35216
rect 10348 35176 10388 35216
rect 11020 35176 11060 35216
rect 844 35092 884 35132
rect 2668 35092 2708 35132
rect 5356 35092 5396 35132
rect 6508 35092 6548 35132
rect 7756 35092 7796 35132
rect 9964 35092 10004 35132
rect 1804 34924 1844 34964
rect 7084 35008 7124 35048
rect 8524 35008 8564 35048
rect 3916 34924 3956 34964
rect 7852 34924 7892 34964
rect 9868 34924 9908 34964
rect 11212 34924 11252 34964
rect 7756 34840 7796 34880
rect 4928 34756 4968 34796
rect 5010 34756 5050 34796
rect 5092 34756 5132 34796
rect 5174 34756 5214 34796
rect 5256 34756 5296 34796
rect 2284 34672 2324 34712
rect 2476 34672 2516 34712
rect 7468 34588 7508 34628
rect 10924 34588 10964 34628
rect 1036 34504 1076 34544
rect 2860 34504 2900 34544
rect 3436 34504 3476 34544
rect 1228 34451 1268 34460
rect 1228 34420 1259 34451
rect 1259 34420 1268 34451
rect 1996 34420 2036 34460
rect 3532 34420 3572 34460
rect 2188 34336 2228 34376
rect 3436 34336 3476 34376
rect 3628 34336 3668 34376
rect 76 34168 116 34208
rect 4492 34504 4532 34544
rect 7372 34504 7412 34544
rect 8140 34504 8180 34544
rect 5356 34420 5396 34460
rect 7084 34420 7124 34460
rect 7564 34420 7604 34460
rect 8716 34504 8756 34544
rect 9388 34420 9428 34460
rect 7756 34336 7796 34376
rect 10924 34336 10964 34376
rect 7084 34252 7124 34292
rect 9676 34252 9716 34292
rect 4492 34168 4532 34208
rect 5356 34168 5396 34208
rect 6892 34168 6932 34208
rect 8716 34168 8756 34208
rect 11116 34168 11156 34208
rect 8428 34084 8468 34124
rect 3688 34000 3728 34040
rect 3770 34000 3810 34040
rect 3852 34000 3892 34040
rect 3934 34000 3974 34040
rect 4016 34000 4056 34040
rect 1516 33832 1556 33872
rect 4876 33748 4916 33788
rect 3340 33664 3380 33704
rect 3628 33664 3668 33704
rect 5644 33664 5684 33704
rect 6220 33664 6260 33704
rect 7180 33664 7220 33704
rect 7756 33664 7796 33704
rect 8236 33664 8276 33704
rect 8716 33748 8756 33788
rect 9004 33664 9044 33704
rect 748 33580 788 33620
rect 1996 33580 2036 33620
rect 3052 33580 3092 33620
rect 3436 33580 3476 33620
rect 4300 33580 4328 33620
rect 4328 33580 4340 33620
rect 4588 33580 4628 33620
rect 6124 33580 6164 33620
rect 6796 33580 6836 33620
rect 7852 33580 7892 33620
rect 8524 33580 8564 33620
rect 8716 33580 8756 33620
rect 9868 33580 9908 33620
rect 1804 33496 1844 33536
rect 2572 33496 2612 33536
rect 3532 33496 3572 33536
rect 8140 33496 8180 33536
rect 3340 33412 3380 33452
rect 6220 33412 6260 33452
rect 1516 33244 1556 33284
rect 7468 33412 7508 33452
rect 11116 33412 11156 33452
rect 7852 33328 7892 33368
rect 2956 33244 2996 33284
rect 3628 33244 3668 33284
rect 4928 33244 4968 33284
rect 5010 33244 5050 33284
rect 5092 33244 5132 33284
rect 5174 33244 5214 33284
rect 5256 33244 5296 33284
rect 10252 33160 10292 33200
rect 11212 33160 11252 33200
rect 1420 32992 1460 33032
rect 2956 32992 2996 33032
rect 3916 32992 3956 33032
rect 5260 32992 5300 33032
rect 2092 32908 2132 32948
rect 3340 32908 3380 32948
rect 4300 32908 4340 32948
rect 6028 33076 6068 33116
rect 6796 33076 6836 33116
rect 8524 33076 8564 33116
rect 11404 33076 11444 33116
rect 5644 32992 5684 33032
rect 5356 32908 5396 32948
rect 1132 32824 1172 32864
rect 2668 32824 2708 32864
rect 3532 32824 3572 32864
rect 6124 32824 6164 32864
rect 2860 32740 2900 32780
rect 8332 32992 8372 33032
rect 6508 32824 6548 32864
rect 8236 32824 8276 32864
rect 6796 32740 6836 32780
rect 1612 32656 1652 32696
rect 3628 32656 3668 32696
rect 4204 32656 4244 32696
rect 2956 32572 2996 32612
rect 3244 32572 3284 32612
rect 1324 32488 1364 32528
rect 9004 32908 9044 32948
rect 8716 32824 8756 32864
rect 9100 32824 9140 32864
rect 8524 32740 8564 32780
rect 9292 32740 9332 32780
rect 8524 32572 8564 32612
rect 8716 32572 8756 32612
rect 3688 32488 3728 32528
rect 3770 32488 3810 32528
rect 3852 32488 3892 32528
rect 3934 32488 3974 32528
rect 4016 32488 4056 32528
rect 10060 32824 10100 32864
rect 4012 32320 4052 32360
rect 10732 32320 10772 32360
rect 460 32152 500 32192
rect 3148 32152 3188 32192
rect 3532 32152 3572 32192
rect 4204 32152 4244 32192
rect 8236 32152 8276 32192
rect 8620 32152 8660 32192
rect 9580 32152 9620 32192
rect 10156 32152 10196 32192
rect 1420 32068 1460 32108
rect 2668 32068 2708 32108
rect 4012 32068 4052 32108
rect 6028 32068 6068 32108
rect 8332 32068 8344 32108
rect 8344 32068 8372 32108
rect 8524 32068 8564 32108
rect 10252 32068 10292 32108
rect 1516 31900 1556 31940
rect 4300 31900 4340 31940
rect 4876 31900 4916 31940
rect 6892 31984 6932 32024
rect 11020 31984 11060 32024
rect 5644 31900 5684 31940
rect 6124 31900 6155 31940
rect 6155 31900 6164 31940
rect 9100 31900 9131 31940
rect 9131 31900 9140 31940
rect 11212 31900 11252 31940
rect 844 31732 884 31772
rect 1420 31732 1460 31772
rect 2668 31732 2708 31772
rect 2956 31732 2996 31772
rect 4928 31732 4968 31772
rect 5010 31732 5050 31772
rect 5092 31732 5132 31772
rect 5174 31732 5214 31772
rect 5256 31732 5296 31772
rect 364 31648 404 31688
rect 4780 31564 4820 31604
rect 3436 31480 3476 31520
rect 4012 31480 4052 31520
rect 7276 31648 7316 31688
rect 10828 31648 10868 31688
rect 7756 31564 7796 31604
rect 8236 31564 8276 31604
rect 1324 31396 1355 31436
rect 1355 31396 1364 31436
rect 2668 31396 2708 31436
rect 3532 31396 3572 31436
rect 1036 31312 1076 31352
rect 1228 31144 1268 31184
rect 1516 31144 1556 31184
rect 2188 31144 2228 31184
rect 4684 31396 4724 31436
rect 7276 31480 7316 31520
rect 8620 31480 8660 31520
rect 2860 31312 2900 31352
rect 3148 31312 3188 31352
rect 5548 31312 5588 31352
rect 4300 31228 4340 31268
rect 4780 31228 4820 31268
rect 3628 31144 3668 31184
rect 460 31060 500 31100
rect 3688 30976 3728 31016
rect 3770 30976 3810 31016
rect 3852 30976 3892 31016
rect 3934 30976 3974 31016
rect 4016 30976 4056 31016
rect 6124 31396 6164 31436
rect 7084 31396 7124 31436
rect 8716 31396 8756 31436
rect 9004 31396 9044 31436
rect 9580 31396 9620 31436
rect 8332 31354 8371 31394
rect 8371 31354 8372 31394
rect 6028 31228 6068 31268
rect 7564 31228 7604 31268
rect 6604 31144 6644 31184
rect 1420 30892 1460 30932
rect 10156 31427 10196 31436
rect 10156 31396 10196 31427
rect 9292 31312 9332 31352
rect 11020 31144 11060 31184
rect 1324 30808 1364 30848
rect 10348 30808 10388 30848
rect 1516 30724 1556 30764
rect 2860 30724 2900 30764
rect 3244 30724 3284 30764
rect 7180 30724 7220 30764
rect 1900 30640 1940 30680
rect 3628 30640 3668 30680
rect 4012 30640 4052 30680
rect 6028 30640 6068 30680
rect 1996 30556 2036 30596
rect 3820 30556 3860 30596
rect 6796 30556 6836 30596
rect 7180 30556 7220 30596
rect 7564 30556 7604 30596
rect 8044 30556 8084 30596
rect 8812 30556 8852 30596
rect 9868 30556 9908 30596
rect 748 30472 788 30512
rect 2956 30388 2996 30428
rect 3244 30388 3284 30428
rect 3628 30388 3668 30428
rect 4204 30472 4244 30512
rect 7372 30472 7412 30512
rect 4300 30388 4340 30428
rect 6028 30388 6068 30428
rect 7660 30388 7700 30428
rect 9868 30388 9908 30428
rect 3340 30304 3380 30344
rect 9484 30304 9524 30344
rect 4928 30220 4968 30260
rect 5010 30220 5050 30260
rect 5092 30220 5132 30260
rect 5174 30220 5214 30260
rect 5256 30220 5296 30260
rect 1420 30136 1460 30176
rect 4012 30136 4052 30176
rect 11212 30136 11252 30176
rect 4876 30052 4916 30092
rect 10156 30052 10196 30092
rect 3244 29968 3284 30008
rect 3820 29968 3860 30008
rect 4972 29968 5012 30008
rect 8716 29968 8756 30008
rect 9004 29968 9044 30008
rect 844 29884 884 29924
rect 1900 29884 1940 29924
rect 4012 29884 4052 29924
rect 4780 29915 4820 29924
rect 1324 29800 1364 29840
rect 3052 29800 3092 29840
rect 4780 29884 4811 29915
rect 4811 29884 4820 29915
rect 6028 29884 6068 29924
rect 6604 29884 6644 29924
rect 7372 29884 7412 29924
rect 7660 29915 7700 29924
rect 7660 29884 7700 29915
rect 9484 29884 9524 29924
rect 10060 29884 10100 29924
rect 4876 29800 4916 29840
rect 5164 29800 5204 29840
rect 5932 29800 5972 29840
rect 6412 29800 6452 29840
rect 8236 29800 8276 29840
rect 8716 29800 8756 29840
rect 3820 29632 3860 29672
rect 3688 29464 3728 29504
rect 3770 29464 3810 29504
rect 3852 29464 3892 29504
rect 3934 29464 3974 29504
rect 4016 29464 4056 29504
rect 4396 29716 4436 29756
rect 5548 29716 5588 29756
rect 10828 29632 10868 29672
rect 268 29212 308 29252
rect 5164 29212 5204 29252
rect 6604 29212 6644 29252
rect 8716 29212 8756 29252
rect 9004 29212 9044 29252
rect 1516 29128 1556 29168
rect 2380 29128 2419 29168
rect 2419 29128 2420 29168
rect 4300 29128 4340 29168
rect 4780 29128 4820 29168
rect 5548 29128 5588 29168
rect 748 29044 788 29084
rect 1324 29044 1364 29084
rect 2476 29044 2516 29084
rect 3148 29044 3179 29084
rect 3179 29044 3188 29084
rect 4108 29044 4148 29084
rect 4492 29044 4532 29084
rect 5356 29044 5396 29084
rect 5932 29128 5972 29168
rect 6412 29128 6452 29168
rect 7468 29128 7508 29168
rect 9196 29128 9236 29168
rect 10348 29128 10388 29168
rect 10828 29128 10868 29168
rect 6220 29044 6228 29084
rect 6228 29044 6260 29084
rect 8812 29044 8852 29084
rect 10252 29044 10292 29084
rect 2572 28960 2612 29000
rect 2860 28960 2900 29000
rect 3244 28960 3284 29000
rect 3532 28960 3572 29000
rect 3724 28960 3764 29000
rect 4204 28960 4244 29000
rect 4396 28960 4436 29000
rect 7468 28960 7508 29000
rect 6796 28876 6836 28916
rect 9676 28876 9716 28916
rect 11500 28876 11540 28916
rect 1708 28792 1748 28832
rect 4928 28708 4968 28748
rect 5010 28708 5050 28748
rect 5092 28708 5132 28748
rect 5174 28708 5214 28748
rect 5256 28708 5296 28748
rect 6028 28792 6068 28832
rect 8524 28792 8564 28832
rect 7276 28708 7316 28748
rect 3340 28624 3380 28664
rect 2668 28540 2708 28580
rect 3724 28540 3764 28580
rect 4204 28540 4244 28580
rect 6892 28540 6923 28580
rect 6923 28540 6932 28580
rect 7084 28540 7124 28580
rect 7276 28540 7316 28580
rect 7660 28540 7700 28580
rect 2476 28456 2516 28496
rect 3436 28456 3476 28496
rect 10924 28624 10964 28664
rect 10252 28540 10292 28580
rect 11404 28540 11444 28580
rect 7852 28456 7892 28496
rect 9676 28456 9716 28496
rect 1228 28372 1268 28412
rect 1708 28372 1748 28412
rect 3340 28372 3352 28412
rect 3352 28372 3380 28412
rect 4012 28372 4052 28412
rect 4780 28372 4820 28412
rect 4108 28288 4148 28328
rect 4300 28204 4340 28244
rect 460 28120 500 28160
rect 3688 27952 3728 27992
rect 3770 27952 3810 27992
rect 3852 27952 3892 27992
rect 3934 27952 3974 27992
rect 4016 27952 4056 27992
rect 5932 28372 5972 28412
rect 5356 28288 5396 28328
rect 9292 28372 9332 28412
rect 6604 28288 6644 28328
rect 7180 28288 7220 28328
rect 7852 28288 7892 28328
rect 8236 28288 8276 28328
rect 6412 28204 6452 28244
rect 9868 28288 9908 28328
rect 9100 28204 9140 28244
rect 8140 28120 8180 28160
rect 8524 28120 8564 28160
rect 9964 28036 10004 28076
rect 10924 28120 10964 28160
rect 1036 27784 1076 27824
rect 1516 27700 1556 27740
rect 5740 27700 5780 27740
rect 7948 27700 7988 27740
rect 11404 27700 11444 27740
rect 1900 27616 1940 27656
rect 2380 27616 2420 27656
rect 364 27532 404 27572
rect 2860 27532 2900 27572
rect 4588 27532 4628 27572
rect 7180 27532 7220 27572
rect 7756 27616 7796 27656
rect 10060 27532 10100 27572
rect 1036 27448 1076 27488
rect 1996 27448 2036 27488
rect 8140 27448 8180 27488
rect 9676 27448 9716 27488
rect 1420 27364 1460 27404
rect 2284 27364 2324 27404
rect 6028 27364 6068 27404
rect 8236 27364 8267 27404
rect 8267 27364 8276 27404
rect 10348 27364 10388 27404
rect 2860 27280 2900 27320
rect 5644 27280 5684 27320
rect 7084 27280 7124 27320
rect 1324 27112 1364 27152
rect 4300 27196 4340 27236
rect 4928 27196 4968 27236
rect 5010 27196 5050 27236
rect 5092 27196 5132 27236
rect 5174 27196 5214 27236
rect 5256 27196 5296 27236
rect 1804 27112 1844 27152
rect 7180 27112 7220 27152
rect 11500 27112 11540 27152
rect 2668 27028 2708 27068
rect 3532 27028 3572 27068
rect 4684 27028 4724 27068
rect 2860 26944 2900 26984
rect 4492 26944 4532 26984
rect 1228 26891 1268 26900
rect 1228 26860 1259 26891
rect 1259 26860 1268 26891
rect 1996 26891 2036 26900
rect 1996 26860 2027 26891
rect 2027 26860 2036 26891
rect 2572 26860 2612 26900
rect 2956 26860 2996 26900
rect 268 26776 308 26816
rect 1804 26692 1844 26732
rect 4588 26860 4628 26900
rect 4972 26860 5012 26900
rect 6508 27028 6548 27068
rect 7084 26860 7124 26900
rect 7372 26860 7412 26900
rect 8140 26891 8180 26900
rect 8140 26860 8180 26891
rect 8812 26860 8852 26900
rect 9100 26860 9140 26900
rect 10348 26891 10388 26900
rect 10348 26860 10388 26891
rect 8620 26776 8660 26816
rect 4588 26692 4628 26732
rect 7180 26692 7220 26732
rect 8428 26692 8468 26732
rect 4684 26608 4724 26648
rect 10540 26608 10580 26648
rect 1036 26524 1076 26564
rect 5068 26524 5108 26564
rect 1516 26440 1556 26480
rect 3688 26440 3728 26480
rect 3770 26440 3810 26480
rect 3852 26440 3892 26480
rect 3934 26440 3974 26480
rect 4016 26440 4056 26480
rect 7660 26356 7700 26396
rect 2476 26272 2516 26312
rect 3340 26272 3380 26312
rect 4300 26272 4340 26312
rect 4780 26272 4820 26312
rect 10636 26272 10676 26312
rect 5260 26188 5300 26228
rect 6796 26188 6836 26228
rect 6988 26188 7028 26228
rect 748 26104 788 26144
rect 1900 26104 1940 26144
rect 2572 26104 2612 26144
rect 652 26020 692 26060
rect 1996 26020 2036 26060
rect 3340 26020 3380 26060
rect 3916 26020 3956 26060
rect 4300 26020 4340 26060
rect 5068 26104 5108 26144
rect 5932 26104 5972 26144
rect 6700 26104 6740 26144
rect 7564 26104 7604 26144
rect 9100 26104 9140 26144
rect 4972 26020 5012 26060
rect 6508 25936 6548 25976
rect 7276 25936 7316 25976
rect 7468 25936 7508 25976
rect 11404 25936 11444 25976
rect 11692 25936 11732 25976
rect 3820 25852 3860 25892
rect 4108 25852 4148 25892
rect 5260 25852 5291 25892
rect 5291 25852 5300 25892
rect 7948 25852 7988 25892
rect 9484 25852 9524 25892
rect 2284 25768 2324 25808
rect 5740 25768 5780 25808
rect 6892 25768 6932 25808
rect 7756 25768 7796 25808
rect 9580 25768 9620 25808
rect 4928 25684 4968 25724
rect 5010 25684 5050 25724
rect 5092 25684 5132 25724
rect 5174 25684 5214 25724
rect 5256 25684 5296 25724
rect 7276 25684 7316 25724
rect 6700 25516 6740 25556
rect 6892 25516 6932 25556
rect 364 25432 404 25472
rect 4108 25432 4148 25472
rect 4300 25432 4340 25472
rect 1804 25348 1844 25388
rect 2572 25348 2612 25388
rect 2956 25348 2987 25388
rect 2987 25348 2996 25388
rect 3148 25348 3188 25388
rect 3820 25348 3860 25388
rect 4396 25348 4436 25388
rect 6028 25348 6068 25388
rect 3916 25264 3956 25304
rect 4108 25264 4148 25304
rect 5356 25264 5396 25304
rect 8332 25348 8372 25388
rect 9484 25379 9524 25388
rect 9484 25348 9524 25379
rect 7564 25264 7604 25304
rect 7948 25264 7988 25304
rect 8524 25264 8564 25304
rect 10348 25348 10388 25388
rect 11596 25264 11636 25304
rect 2284 25180 2324 25220
rect 7372 25180 7412 25220
rect 8716 25180 8756 25220
rect 1228 25096 1268 25136
rect 652 24760 692 24800
rect 2956 24760 2996 24800
rect 3688 24928 3728 24968
rect 3770 24928 3810 24968
rect 3852 24928 3892 24968
rect 3934 24928 3974 24968
rect 4016 24928 4056 24968
rect 7180 24844 7220 24884
rect 8140 24844 8180 24884
rect 4588 24592 4628 24632
rect 11692 24676 11732 24716
rect 7084 24592 7124 24632
rect 844 24508 884 24548
rect 1996 24508 2036 24548
rect 2380 24508 2420 24548
rect 3052 24508 3092 24548
rect 3244 24508 3284 24548
rect 4396 24508 4421 24548
rect 4421 24508 4436 24548
rect 5932 24508 5972 24548
rect 6412 24508 6452 24548
rect 7372 24508 7412 24548
rect 7852 24508 7860 24548
rect 7860 24508 7892 24548
rect 9388 24508 9428 24548
rect 10060 24508 10100 24548
rect 10252 24508 10292 24548
rect 10828 24508 10868 24548
rect 652 24424 692 24464
rect 4492 24424 4532 24464
rect 6988 24424 7028 24464
rect 7180 24424 7220 24464
rect 8236 24424 8276 24464
rect 2572 24340 2612 24380
rect 3916 24340 3956 24380
rect 4928 24172 4968 24212
rect 5010 24172 5050 24212
rect 5092 24172 5132 24212
rect 5174 24172 5214 24212
rect 5256 24172 5296 24212
rect 748 24088 788 24128
rect 6028 24088 6068 24128
rect 6796 24088 6836 24128
rect 11404 24088 11444 24128
rect 2572 24004 2612 24044
rect 3244 24004 3284 24044
rect 4396 24004 4436 24044
rect 5740 24004 5771 24044
rect 5771 24004 5780 24044
rect 6700 24004 6740 24044
rect 7852 24004 7892 24044
rect 9004 24004 9044 24044
rect 1708 23920 1748 23960
rect 2284 23920 2324 23960
rect 3052 23920 3092 23960
rect 4972 23920 5012 23960
rect 5932 23920 5972 23960
rect 7468 23920 7508 23960
rect 7756 23920 7796 23960
rect 9676 23920 9716 23960
rect 9964 23920 10004 23960
rect 1516 23836 1556 23876
rect 2092 23836 2132 23876
rect 460 23752 500 23792
rect 2956 23752 2996 23792
rect 1708 23584 1748 23624
rect 2284 23584 2324 23624
rect 5356 23836 5396 23876
rect 6124 23836 6164 23876
rect 8620 23836 8660 23876
rect 9580 23836 9620 23876
rect 10060 23836 10100 23876
rect 4108 23752 4148 23792
rect 4684 23752 4724 23792
rect 5260 23752 5300 23792
rect 5068 23668 5108 23708
rect 7468 23668 7508 23708
rect 8620 23668 8660 23708
rect 7756 23584 7796 23624
rect 8044 23584 8084 23624
rect 3688 23416 3728 23456
rect 3770 23416 3810 23456
rect 3852 23416 3892 23456
rect 3934 23416 3974 23456
rect 4016 23416 4056 23456
rect 7756 23416 7796 23456
rect 8428 23416 8468 23456
rect 4204 23248 4244 23288
rect 6028 23248 6068 23288
rect 5356 23164 5396 23204
rect 748 23080 788 23120
rect 652 22996 692 23036
rect 1996 22996 2036 23036
rect 2572 22996 2612 23036
rect 3244 22996 3284 23036
rect 8620 23164 8660 23204
rect 4012 23080 4052 23120
rect 4876 23080 4916 23120
rect 6124 23080 6164 23120
rect 6412 23080 6452 23120
rect 8428 23080 8468 23120
rect 10636 23080 10676 23120
rect 4396 22996 4436 23036
rect 5644 22996 5684 23036
rect 7468 22996 7508 23036
rect 8332 22996 8372 23036
rect 9004 22996 9044 23036
rect 9196 22996 9236 23036
rect 1132 22912 1172 22952
rect 2092 22912 2132 22952
rect 3340 22912 3380 22952
rect 4012 22912 4052 22952
rect 5452 22912 5492 22952
rect 7180 22912 7220 22952
rect 1708 22828 1748 22868
rect 3052 22828 3092 22868
rect 3724 22828 3764 22868
rect 4780 22828 4820 22868
rect 4972 22828 5012 22868
rect 5740 22828 5780 22868
rect 6220 22828 6260 22868
rect 6700 22828 6740 22868
rect 7852 22828 7892 22868
rect 1228 22744 1268 22784
rect 6508 22744 6548 22784
rect 4396 22660 4436 22700
rect 4928 22660 4968 22700
rect 5010 22660 5050 22700
rect 5092 22660 5132 22700
rect 5174 22660 5214 22700
rect 5256 22660 5296 22700
rect 5452 22660 5492 22700
rect 11596 22828 11636 22868
rect 2092 22492 2132 22532
rect 2860 22492 2900 22532
rect 6124 22492 6164 22532
rect 7564 22492 7604 22532
rect 8044 22492 8075 22532
rect 8075 22492 8084 22532
rect 10636 22492 10676 22532
rect 76 22408 116 22448
rect 5260 22408 5300 22448
rect 10732 22408 10772 22448
rect 1804 22324 1844 22364
rect 1996 22324 2036 22364
rect 2572 22324 2612 22364
rect 3532 22324 3572 22364
rect 5068 22355 5108 22364
rect 5068 22324 5108 22355
rect 2668 22240 2708 22280
rect 2860 22240 2900 22280
rect 4300 22240 4340 22280
rect 2956 22156 2996 22196
rect 556 22072 596 22112
rect 364 21736 404 21776
rect 2764 21736 2804 21776
rect 3436 21652 3476 21692
rect 6604 22324 6644 22364
rect 7084 22324 7124 22364
rect 8044 22324 8084 22364
rect 9580 22324 9620 22364
rect 11404 22240 11444 22280
rect 4972 22156 5012 22196
rect 5452 22156 5492 22196
rect 6124 22156 6164 22196
rect 7564 22156 7604 22196
rect 3724 22072 3764 22112
rect 4300 22072 4340 22112
rect 3688 21904 3728 21944
rect 3770 21904 3810 21944
rect 3852 21904 3892 21944
rect 3934 21904 3974 21944
rect 4016 21904 4056 21944
rect 5644 21820 5684 21860
rect 5068 21652 5108 21692
rect 1900 21568 1940 21608
rect 3628 21568 3668 21608
rect 4012 21568 4052 21608
rect 4972 21568 5012 21608
rect 5164 21568 5204 21608
rect 8332 21568 8372 21608
rect 10348 21568 10388 21608
rect 6028 21557 6068 21566
rect 6028 21526 6068 21557
rect 460 21484 500 21524
rect 2284 21484 2315 21524
rect 2315 21484 2324 21524
rect 4108 21484 4148 21524
rect 5452 21484 5492 21524
rect 6604 21484 6644 21524
rect 8044 21484 8084 21524
rect 10060 21484 10100 21524
rect 652 21400 692 21440
rect 2668 21400 2708 21440
rect 5644 21400 5684 21440
rect 5836 21400 5876 21440
rect 8908 21400 8948 21440
rect 4300 21316 4340 21356
rect 4684 21316 4724 21356
rect 3916 21232 3956 21272
rect 4928 21148 4968 21188
rect 5010 21148 5050 21188
rect 5092 21148 5132 21188
rect 5174 21148 5214 21188
rect 5256 21148 5296 21188
rect 268 21064 308 21104
rect 3628 21064 3668 21104
rect 1708 20980 1748 21020
rect 2092 20980 2132 21020
rect 5932 20980 5972 21020
rect 6700 20980 6740 21020
rect 7852 20980 7892 21020
rect 1516 20896 1556 20936
rect 1900 20896 1940 20936
rect 3340 20896 3380 20936
rect 5740 20896 5780 20936
rect 9100 20896 9140 20936
rect 1228 20843 1268 20852
rect 1228 20812 1259 20843
rect 1259 20812 1268 20843
rect 3148 20812 3179 20852
rect 3179 20812 3188 20852
rect 3916 20812 3956 20852
rect 5260 20812 5300 20852
rect 460 20728 500 20768
rect 2092 20728 2132 20768
rect 4300 20728 4340 20768
rect 5452 20812 5492 20852
rect 5644 20812 5684 20852
rect 6124 20812 6164 20852
rect 6604 20812 6644 20852
rect 5836 20728 5867 20768
rect 5867 20728 5876 20768
rect 8908 20812 8948 20852
rect 10636 20812 10676 20852
rect 11308 20812 11348 20852
rect 3628 20644 3668 20684
rect 4012 20644 4052 20684
rect 5452 20644 5492 20684
rect 6508 20644 6548 20684
rect 8908 20644 8948 20684
rect 3148 20560 3188 20600
rect 4108 20560 4148 20600
rect 5836 20560 5876 20600
rect 1228 20392 1268 20432
rect 3688 20392 3728 20432
rect 3770 20392 3810 20432
rect 3852 20392 3892 20432
rect 3934 20392 3974 20432
rect 4016 20392 4056 20432
rect 2860 20224 2900 20264
rect 3916 20224 3956 20264
rect 6124 20224 6164 20264
rect 1804 20140 1844 20180
rect 3148 20140 3188 20180
rect 5644 20140 5684 20180
rect 1516 20056 1556 20096
rect 5068 20056 5108 20096
rect 5356 20056 5396 20096
rect 5740 20056 5780 20096
rect 8524 20056 8564 20096
rect 9868 20056 9908 20096
rect 556 19972 596 20012
rect 1804 19972 1844 20012
rect 2092 19972 2132 20012
rect 2284 19972 2324 20012
rect 3148 19972 3188 20012
rect 4108 19972 4148 20012
rect 4780 19972 4820 20012
rect 5260 19972 5300 20012
rect 7084 19972 7124 20012
rect 9100 19972 9140 20012
rect 9580 19972 9620 20012
rect 1132 19888 1172 19928
rect 2668 19888 2708 19928
rect 1804 19804 1844 19844
rect 5932 19888 5972 19928
rect 5452 19804 5483 19844
rect 5483 19804 5492 19844
rect 6508 19804 6548 19844
rect 556 19720 596 19760
rect 5932 19720 5972 19760
rect 1420 19636 1460 19676
rect 3052 19636 3092 19676
rect 4928 19636 4968 19676
rect 5010 19636 5050 19676
rect 5092 19636 5132 19676
rect 5174 19636 5214 19676
rect 5256 19636 5296 19676
rect 1900 19552 1940 19592
rect 268 19468 308 19508
rect 3532 19468 3572 19508
rect 940 19384 980 19424
rect 2572 19384 2612 19424
rect 3628 19384 3668 19424
rect 364 19300 404 19340
rect 1420 19300 1460 19340
rect 1996 19216 2036 19256
rect 3724 19300 3764 19340
rect 4012 19331 4052 19340
rect 4012 19300 4043 19331
rect 4043 19300 4052 19331
rect 5164 19300 5204 19340
rect 2572 19216 2612 19256
rect 2764 19216 2804 19256
rect 2092 19132 2132 19172
rect 3148 19132 3188 19172
rect 7948 19888 7988 19928
rect 8620 19888 8660 19928
rect 9676 19804 9716 19844
rect 9868 19468 9908 19508
rect 7660 19300 7700 19340
rect 9580 19300 9620 19340
rect 10252 19300 10292 19340
rect 10636 19300 10676 19340
rect 7468 19216 7508 19256
rect 8140 19216 8180 19256
rect 9100 19216 9140 19256
rect 7276 19132 7316 19172
rect 9484 19132 9524 19172
rect 1420 19048 1460 19088
rect 2668 19048 2708 19088
rect 10636 19048 10676 19088
rect 7468 18964 7508 19004
rect 3688 18880 3728 18920
rect 3770 18880 3810 18920
rect 3852 18880 3892 18920
rect 3934 18880 3974 18920
rect 4016 18880 4056 18920
rect 5644 18796 5684 18836
rect 8140 18796 8180 18836
rect 748 18712 788 18752
rect 2284 18712 2324 18752
rect 3532 18712 3572 18752
rect 8524 18712 8564 18752
rect 1420 18628 1460 18668
rect 1708 18544 1748 18584
rect 1900 18544 1940 18584
rect 4684 18628 4724 18668
rect 6700 18628 6740 18668
rect 7084 18544 7124 18584
rect 652 18460 692 18500
rect 1516 18460 1556 18500
rect 2284 18460 2324 18500
rect 3052 18460 3092 18500
rect 3244 18460 3284 18500
rect 940 18376 980 18416
rect 1996 18376 2036 18416
rect 2572 18376 2612 18416
rect 2956 18376 2996 18416
rect 3532 18292 3572 18332
rect 5164 18460 5204 18500
rect 5932 18460 5972 18500
rect 6604 18460 6644 18500
rect 8332 18628 8372 18668
rect 7660 18544 7700 18584
rect 8236 18544 8276 18584
rect 7468 18460 7508 18500
rect 8716 18460 8756 18500
rect 9676 18460 9716 18500
rect 9868 18460 9907 18500
rect 9907 18460 9908 18500
rect 7852 18376 7892 18416
rect 5260 18292 5291 18332
rect 5291 18292 5300 18332
rect 6604 18292 6644 18332
rect 7468 18292 7499 18332
rect 7499 18292 7508 18332
rect 10540 18292 10580 18332
rect 2956 18208 2996 18248
rect 5356 18208 5396 18248
rect 4928 18124 4968 18164
rect 5010 18124 5050 18164
rect 5092 18124 5132 18164
rect 5174 18124 5214 18164
rect 5256 18124 5296 18164
rect 364 18040 404 18080
rect 4492 17956 4532 17996
rect 5644 17956 5684 17996
rect 6220 17956 6260 17996
rect 9484 17956 9524 17996
rect 1132 17872 1172 17912
rect 1900 17872 1940 17912
rect 3532 17872 3572 17912
rect 4396 17872 4436 17912
rect 5356 17872 5396 17912
rect 460 17788 500 17828
rect 1996 17788 2036 17828
rect 3052 17788 3092 17828
rect 76 17704 116 17744
rect 1900 17704 1940 17744
rect 2284 17704 2324 17744
rect 3436 17819 3476 17828
rect 3436 17788 3476 17819
rect 4780 17788 4820 17828
rect 6604 17872 6644 17912
rect 7276 17872 7316 17912
rect 7660 17872 7700 17912
rect 5644 17788 5684 17828
rect 3532 17704 3572 17744
rect 4108 17704 4148 17744
rect 4492 17704 4532 17744
rect 5068 17704 5108 17744
rect 3052 17620 3092 17660
rect 4300 17536 4340 17576
rect 8236 17788 8276 17828
rect 8812 17819 8852 17828
rect 8812 17788 8852 17819
rect 9292 17819 9332 17828
rect 9292 17788 9332 17819
rect 10732 18040 10772 18080
rect 10636 17956 10676 17996
rect 6604 17704 6644 17744
rect 7468 17704 7508 17744
rect 8140 17704 8180 17744
rect 9196 17704 9236 17744
rect 7276 17536 7316 17576
rect 8140 17452 8180 17492
rect 460 17368 500 17408
rect 3688 17368 3728 17408
rect 3770 17368 3810 17408
rect 3852 17368 3892 17408
rect 3934 17368 3974 17408
rect 4016 17368 4056 17408
rect 4876 17368 4916 17408
rect 3532 17116 3572 17156
rect 1420 17032 1460 17072
rect 3628 17032 3668 17072
rect 3916 17032 3947 17072
rect 3947 17032 3956 17072
rect 5836 17284 5876 17324
rect 10540 17284 10580 17324
rect 10924 17284 10964 17324
rect 4780 17200 4820 17240
rect 6796 17200 6836 17240
rect 7948 17200 7988 17240
rect 9292 17200 9332 17240
rect 10732 17200 10772 17240
rect 6316 17116 6356 17156
rect 4876 17032 4916 17072
rect 5740 17032 5780 17072
rect 6220 17032 6260 17072
rect 7084 17032 7124 17072
rect 9484 17032 9524 17072
rect 11212 17032 11252 17072
rect 556 16948 596 16988
rect 2956 16948 2996 16988
rect 3724 16948 3764 16988
rect 5164 16948 5204 16988
rect 5932 16948 5972 16988
rect 7180 16948 7192 16988
rect 7192 16948 7220 16988
rect 8812 16948 8852 16988
rect 9292 16948 9332 16988
rect 9676 16948 9716 16988
rect 9868 16948 9908 16988
rect 172 16864 212 16904
rect 3340 16864 3380 16904
rect 3628 16864 3668 16904
rect 1804 16780 1844 16820
rect 1996 16780 2036 16820
rect 4012 16780 4052 16820
rect 4396 16780 4436 16820
rect 5836 16864 5876 16904
rect 5260 16780 5300 16820
rect 6220 16780 6260 16820
rect 9868 16780 9908 16820
rect 652 16696 692 16736
rect 5356 16696 5396 16736
rect 1036 16528 1076 16568
rect 4928 16612 4968 16652
rect 5010 16612 5050 16652
rect 5092 16612 5132 16652
rect 5174 16612 5214 16652
rect 5256 16612 5296 16652
rect 4396 16528 4436 16568
rect 5932 16528 5972 16568
rect 1612 16444 1652 16484
rect 1036 16360 1076 16400
rect 4012 16360 4052 16400
rect 4972 16444 5012 16484
rect 5644 16444 5684 16484
rect 7468 16696 7508 16736
rect 7948 16696 7988 16736
rect 9292 16696 9332 16736
rect 9676 16528 9716 16568
rect 7564 16444 7604 16484
rect 10156 16444 10196 16484
rect 7756 16360 7796 16400
rect 8620 16360 8660 16400
rect 748 16276 788 16316
rect 2956 16276 2996 16316
rect 3340 16276 3380 16316
rect 3916 16276 3956 16316
rect 5356 16276 5396 16316
rect 76 16192 116 16232
rect 2860 16192 2900 16232
rect 3532 16192 3572 16232
rect 4108 16192 4148 16232
rect 7084 16276 7124 16316
rect 7564 16276 7604 16316
rect 8332 16276 8372 16316
rect 8812 16276 8852 16316
rect 9004 16276 9044 16316
rect 9388 16307 9428 16316
rect 9388 16276 9428 16307
rect 9676 16276 9716 16316
rect 4876 16192 4916 16232
rect 5740 16192 5780 16232
rect 7468 16192 7508 16232
rect 7756 16192 7796 16232
rect 8428 16192 8468 16232
rect 4396 16108 4436 16148
rect 4300 16024 4340 16064
rect 10732 16024 10772 16064
rect 3688 15856 3728 15896
rect 3770 15856 3810 15896
rect 3852 15856 3892 15896
rect 3934 15856 3974 15896
rect 4016 15856 4056 15896
rect 5644 15856 5684 15896
rect 9868 15772 9908 15812
rect 1324 15688 1364 15728
rect 1900 15688 1940 15728
rect 1420 15604 1460 15644
rect 3052 15604 3092 15644
rect 3628 15604 3668 15644
rect 4012 15688 4052 15728
rect 5356 15688 5396 15728
rect 7564 15688 7604 15728
rect 9388 15688 9428 15728
rect 11212 15688 11252 15728
rect 7180 15604 7220 15644
rect 2956 15520 2996 15560
rect 3820 15520 3860 15560
rect 172 15436 212 15476
rect 1996 15436 2036 15476
rect 4012 15436 4052 15476
rect 1900 15352 1940 15392
rect 76 15184 116 15224
rect 4300 15520 4340 15560
rect 5740 15520 5780 15560
rect 8620 15520 8660 15560
rect 10156 15520 10196 15560
rect 4300 15268 4340 15308
rect 5260 15436 5300 15476
rect 6028 15436 6068 15476
rect 7468 15436 7508 15476
rect 9004 15268 9044 15308
rect 76 15016 116 15056
rect 364 14932 404 14972
rect 1708 14932 1748 14972
rect 4492 14932 4532 14972
rect 460 14848 500 14888
rect 4928 15100 4968 15140
rect 5010 15100 5050 15140
rect 5092 15100 5132 15140
rect 5174 15100 5214 15140
rect 5256 15100 5296 15140
rect 10636 15016 10676 15056
rect 3628 14848 3668 14888
rect 7948 14932 7988 14972
rect 8428 14932 8468 14972
rect 10732 14932 10772 14972
rect 2572 14764 2612 14804
rect 2860 14764 2900 14804
rect 3724 14764 3764 14804
rect 940 14680 980 14720
rect 2284 14680 2324 14720
rect 2668 14680 2708 14720
rect 3052 14680 3092 14720
rect 5356 14764 5396 14804
rect 5740 14764 5780 14804
rect 6028 14764 6068 14804
rect 7564 14764 7604 14804
rect 7948 14764 7988 14804
rect 8332 14764 8372 14804
rect 8908 14795 8948 14804
rect 8908 14764 8948 14795
rect 9388 14795 9428 14804
rect 9388 14764 9428 14795
rect 8812 14680 8852 14720
rect 11020 14680 11060 14720
rect 3340 14596 3380 14636
rect 5548 14512 5588 14552
rect 8620 14512 8660 14552
rect 6220 14428 6260 14468
rect 3688 14344 3728 14384
rect 3770 14344 3810 14384
rect 3852 14344 3892 14384
rect 3934 14344 3974 14384
rect 4016 14344 4056 14384
rect 10540 14260 10580 14300
rect 652 14092 692 14132
rect 1324 14092 1364 14132
rect 556 14008 596 14048
rect 1420 14008 1460 14048
rect 2572 14092 2612 14132
rect 3724 14092 3764 14132
rect 4876 14092 4916 14132
rect 7180 14176 7220 14216
rect 9388 14176 9428 14216
rect 10636 14176 10676 14216
rect 6316 14092 6356 14132
rect 2860 14008 2900 14048
rect 5740 14008 5780 14048
rect 7468 14008 7508 14048
rect 9580 14008 9620 14048
rect 10060 14008 10100 14048
rect 10540 14008 10580 14048
rect 2284 13924 2324 13964
rect 2764 13924 2804 13964
rect 3052 13924 3092 13964
rect 3628 13924 3668 13964
rect 4204 13924 4244 13964
rect 7180 13924 7219 13964
rect 7219 13924 7220 13964
rect 8428 13924 8468 13964
rect 10252 13924 10292 13964
rect 8620 13840 8660 13880
rect 1036 13756 1076 13796
rect 4492 13756 4532 13796
rect 10348 13756 10388 13796
rect 1324 13672 1364 13712
rect 4928 13588 4968 13628
rect 5010 13588 5050 13628
rect 5092 13588 5132 13628
rect 5174 13588 5214 13628
rect 5256 13588 5296 13628
rect 1420 13504 1460 13544
rect 6028 13504 6068 13544
rect 3340 13420 3380 13460
rect 4780 13420 4820 13460
rect 7660 13504 7700 13544
rect 652 13336 692 13376
rect 3724 13336 3764 13376
rect 1612 13252 1652 13292
rect 2860 13084 2900 13124
rect 3340 13084 3380 13124
rect 8812 13336 8852 13376
rect 10348 13336 10388 13376
rect 8044 13252 8084 13292
rect 9292 13252 9332 13292
rect 7180 13168 7220 13208
rect 9100 13168 9140 13208
rect 7564 13084 7604 13124
rect 7756 13084 7796 13124
rect 748 13000 788 13040
rect 2284 13000 2324 13040
rect 3724 13000 3764 13040
rect 3916 13000 3956 13040
rect 4684 13000 4724 13040
rect 1612 12916 1652 12956
rect 3340 12916 3380 12956
rect 3688 12832 3728 12872
rect 3770 12832 3810 12872
rect 3852 12832 3892 12872
rect 3934 12832 3974 12872
rect 4016 12832 4056 12872
rect 11788 12832 11828 12872
rect 3532 12748 3572 12788
rect 5068 12748 5108 12788
rect 11116 12748 11156 12788
rect 2860 12664 2900 12704
rect 3724 12664 3764 12704
rect 9100 12664 9140 12704
rect 2668 12580 2708 12620
rect 3916 12580 3956 12620
rect 6124 12580 6164 12620
rect 8908 12580 8948 12620
rect 9964 12580 10004 12620
rect 4780 12496 4820 12536
rect 5068 12496 5108 12536
rect 5836 12496 5876 12536
rect 1228 12412 1268 12452
rect 2764 12412 2804 12452
rect 3340 12412 3380 12452
rect 3628 12412 3668 12452
rect 4396 12412 4436 12452
rect 460 12244 500 12284
rect 4928 12076 4968 12116
rect 5010 12076 5050 12116
rect 5092 12076 5132 12116
rect 5174 12076 5214 12116
rect 5256 12076 5296 12116
rect 5644 12076 5684 12116
rect 1804 11992 1844 12032
rect 3052 11908 3092 11948
rect 3532 11908 3572 11948
rect 2860 11824 2900 11864
rect 1612 11740 1652 11780
rect 1996 11740 2036 11780
rect 2668 11740 2708 11780
rect 3628 11740 3668 11780
rect 7564 12412 7604 12452
rect 9292 12412 9332 12452
rect 10252 12412 10292 12452
rect 6412 12244 6452 12284
rect 7564 12244 7604 12284
rect 10636 11992 10676 12032
rect 7852 11908 7892 11948
rect 8428 11908 8468 11948
rect 10060 11908 10100 11948
rect 5932 11824 5972 11864
rect 6700 11824 6740 11864
rect 4108 11740 4148 11780
rect 4876 11740 4916 11780
rect 5740 11771 5780 11780
rect 5740 11740 5780 11771
rect 6124 11740 6164 11780
rect 7564 11740 7604 11780
rect 8620 11740 8651 11780
rect 8651 11740 8660 11780
rect 172 11656 212 11696
rect 3532 11656 3572 11696
rect 3820 11656 3860 11696
rect 4492 11656 4532 11696
rect 8908 11656 8948 11696
rect 1996 11572 2036 11612
rect 8812 11572 8852 11612
rect 3916 11488 3956 11528
rect 7660 11488 7700 11528
rect 3532 11404 3572 11444
rect 4972 11404 5012 11444
rect 11404 11404 11444 11444
rect 1228 11320 1268 11360
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 6700 11320 6740 11360
rect 11500 11320 11540 11360
rect 2476 11236 2516 11276
rect 556 11152 596 11192
rect 1324 11152 1364 11192
rect 4300 11152 4340 11192
rect 5740 11152 5780 11192
rect 6124 11152 6164 11192
rect 6508 11152 6548 11192
rect 2860 11068 2900 11108
rect 4492 11068 4532 11108
rect 1132 10984 1172 11024
rect 2956 10984 2996 11024
rect 3820 10984 3860 11024
rect 4972 10984 5012 11024
rect 6220 10984 6260 11024
rect 9580 11152 9620 11192
rect 9292 10984 9332 11024
rect 10252 10984 10292 11024
rect 2284 10900 2324 10940
rect 2860 10900 2900 10940
rect 4396 10900 4436 10940
rect 5740 10900 5780 10940
rect 6508 10900 6548 10940
rect 7468 10900 7508 10940
rect 7660 10900 7700 10940
rect 8620 10900 8651 10940
rect 8651 10900 8660 10940
rect 6412 10816 6452 10856
rect 8716 10816 8756 10856
rect 9196 10816 9236 10856
rect 2284 10732 2324 10772
rect 3820 10732 3860 10772
rect 4876 10732 4916 10772
rect 1036 10648 1076 10688
rect 652 10396 692 10436
rect 4108 10396 4148 10436
rect 460 10312 500 10352
rect 748 10312 788 10352
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 5548 10732 5588 10772
rect 5260 10396 5300 10436
rect 5932 10312 5972 10352
rect 6988 10312 7028 10352
rect 2284 10228 2324 10268
rect 4588 10228 4628 10268
rect 4876 10228 4916 10268
rect 1420 10144 1460 10184
rect 1804 10144 1844 10184
rect 5836 10259 5876 10268
rect 5836 10228 5876 10259
rect 6028 10228 6068 10268
rect 4300 10144 4340 10184
rect 4492 10144 4532 10184
rect 6700 10144 6740 10184
rect 10252 10396 10292 10436
rect 10636 10396 10676 10436
rect 11692 10228 11732 10268
rect 8620 10144 8660 10184
rect 8908 10144 8948 10184
rect 10348 10144 10388 10184
rect 3532 10060 3572 10100
rect 5260 10060 5300 10100
rect 6124 10060 6164 10100
rect 9292 10060 9332 10100
rect 2956 9976 2996 10016
rect 4396 9976 4436 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 4876 9808 4916 9848
rect 5740 9724 5780 9764
rect 3052 9640 3092 9680
rect 5836 9640 5876 9680
rect 172 9556 212 9596
rect 1324 9556 1364 9596
rect 1420 9472 1460 9512
rect 8620 9640 8660 9680
rect 2956 9472 2996 9512
rect 4780 9472 4820 9512
rect 1132 9388 1172 9428
rect 2284 9388 2324 9428
rect 3820 9388 3860 9428
rect 5260 9388 5300 9428
rect 5740 9388 5780 9428
rect 2956 9304 2996 9344
rect 4396 9220 4436 9260
rect 2476 9136 2516 9176
rect 748 8968 788 9008
rect 1804 8968 1844 9008
rect 2284 8968 2324 9008
rect 2860 8884 2900 8924
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 6508 9388 6548 9428
rect 6988 9388 7028 9428
rect 9388 9472 9428 9512
rect 7468 9388 7508 9428
rect 8332 9388 8372 9428
rect 9772 9388 9812 9428
rect 10348 9388 10388 9428
rect 10828 9388 10868 9428
rect 10636 8968 10676 9008
rect 4300 8884 4340 8924
rect 7468 8884 7508 8924
rect 10444 8800 10484 8840
rect 1804 8747 1844 8756
rect 1804 8716 1835 8747
rect 1835 8716 1844 8747
rect 2764 8716 2804 8756
rect 3532 8747 3572 8756
rect 3532 8716 3572 8747
rect 6508 8716 6548 8756
rect 556 8632 596 8672
rect 2860 8632 2900 8672
rect 8332 8716 8372 8756
rect 9772 8716 9812 8756
rect 10348 8747 10388 8756
rect 10348 8716 10388 8747
rect 8716 8632 8756 8672
rect 10252 8632 10292 8672
rect 4492 8548 4532 8588
rect 7180 8548 7220 8588
rect 10540 8464 10580 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 3244 8128 3284 8168
rect 8908 8128 8948 8168
rect 8332 8044 8372 8084
rect 940 7960 980 8000
rect 1132 7960 1172 8000
rect 6412 7960 6452 8000
rect 7276 7960 7316 8000
rect 7660 7960 7700 8000
rect 8428 7960 8468 8000
rect 10252 7960 10292 8000
rect 1612 7876 1652 7916
rect 2668 7876 2708 7916
rect 2860 7876 2900 7916
rect 4492 7876 4532 7916
rect 5260 7876 5291 7916
rect 5291 7876 5300 7916
rect 7756 7876 7796 7916
rect 7948 7876 7988 7916
rect 10444 7876 10484 7916
rect 10348 7792 10388 7832
rect 4492 7708 4532 7748
rect 8620 7708 8660 7748
rect 10060 7708 10100 7748
rect 3436 7624 3476 7664
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 2284 7372 2324 7412
rect 3628 7372 3668 7412
rect 5644 7372 5684 7412
rect 7756 7372 7796 7412
rect 1420 7288 1460 7328
rect 1324 7204 1364 7244
rect 2668 7204 2708 7244
rect 5740 7204 5780 7244
rect 7180 7204 7220 7244
rect 8620 7204 8660 7244
rect 9388 7204 9428 7244
rect 1708 7120 1748 7160
rect 3724 7120 3764 7160
rect 1516 7036 1556 7076
rect 3052 7036 3092 7076
rect 1804 6952 1844 6992
rect 2956 6952 2996 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 8332 7120 8372 7160
rect 10540 7120 10580 7160
rect 7564 7036 7604 7076
rect 8716 7036 8756 7076
rect 10636 7036 10676 7076
rect 5740 6952 5780 6992
rect 6028 6952 6068 6992
rect 172 6616 212 6656
rect 748 6616 788 6656
rect 4012 6616 4052 6656
rect 3532 6532 3572 6572
rect 1612 6448 1652 6488
rect 3340 6448 3380 6488
rect 4588 6448 4628 6488
rect 9964 6448 10004 6488
rect 1708 6364 1748 6404
rect 2956 6364 2996 6404
rect 4780 6364 4820 6404
rect 5740 6364 5780 6404
rect 6220 6364 6260 6404
rect 7564 6364 7604 6404
rect 2476 6280 2516 6320
rect 4108 6280 4148 6320
rect 7276 6280 7316 6320
rect 11692 6280 11732 6320
rect 5836 6196 5876 6236
rect 10732 6196 10772 6236
rect 4012 6112 4052 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 1228 5944 1268 5984
rect 11692 5944 11732 5984
rect 2092 5860 2132 5900
rect 4588 5860 4628 5900
rect 6700 5860 6740 5900
rect 4780 5776 4820 5816
rect 1516 5692 1556 5732
rect 2764 5692 2804 5732
rect 4300 5692 4340 5732
rect 4588 5692 4628 5732
rect 7180 5692 7220 5732
rect 7756 5723 7796 5732
rect 7756 5692 7796 5723
rect 940 5608 980 5648
rect 1900 5608 1940 5648
rect 2572 5608 2612 5648
rect 5644 5608 5684 5648
rect 5836 5608 5876 5648
rect 2188 5524 2228 5564
rect 8332 5692 8372 5732
rect 8620 5723 8660 5732
rect 8620 5692 8651 5723
rect 8651 5692 8660 5723
rect 8812 5692 8852 5732
rect 7276 5608 7316 5648
rect 6412 5524 6452 5564
rect 6700 5524 6740 5564
rect 7084 5524 7124 5564
rect 844 5440 884 5480
rect 4780 5440 4820 5480
rect 1324 5272 1364 5312
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 4588 5272 4628 5312
rect 5644 5272 5684 5312
rect 9004 5272 9044 5312
rect 11692 5440 11732 5480
rect 4972 5188 5012 5228
rect 8332 5104 8372 5144
rect 8620 5020 8660 5060
rect 4876 4936 4916 4976
rect 11692 4936 11732 4976
rect 1516 4852 1556 4892
rect 2668 4852 2708 4892
rect 2860 4852 2900 4892
rect 3916 4852 3956 4892
rect 4588 4852 4628 4892
rect 4972 4852 5012 4892
rect 5932 4852 5940 4892
rect 5940 4852 5972 4892
rect 8236 4852 8276 4892
rect 1900 4768 1940 4808
rect 7756 4768 7796 4808
rect 2092 4684 2132 4724
rect 2572 4684 2612 4724
rect 460 4600 500 4640
rect 4588 4600 4628 4640
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 1612 4432 1652 4472
rect 4588 4432 4628 4472
rect 6220 4432 6260 4472
rect 1132 4348 1172 4388
rect 1516 4348 1556 4388
rect 3916 4348 3956 4388
rect 6700 4348 6740 4388
rect 844 4264 884 4304
rect 1900 4264 1940 4304
rect 5932 4264 5972 4304
rect 10060 4264 10091 4304
rect 10091 4264 10100 4304
rect 2188 4096 2228 4136
rect 2668 4096 2708 4136
rect 6220 4180 6260 4220
rect 8236 4180 8276 4220
rect 1132 3928 1172 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 1036 3676 1076 3716
rect 3436 3592 3476 3632
rect 11596 3592 11636 3632
rect 1420 3508 1460 3548
rect 3244 3508 3284 3548
rect 5740 3508 5780 3548
rect 1612 3424 1652 3464
rect 2188 3424 2228 3464
rect 3340 3424 3380 3464
rect 4108 3424 4148 3464
rect 4588 3424 4628 3464
rect 5548 3424 5588 3464
rect 6988 3424 7028 3464
rect 1228 3340 1268 3380
rect 10924 3340 10964 3380
rect 1036 3256 1076 3296
rect 1324 3256 1364 3296
rect 1420 3172 1460 3212
rect 3436 3172 3476 3212
rect 11692 3172 11732 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 11692 2920 11732 2960
rect 172 2836 212 2876
rect 3436 2836 3476 2876
rect 5740 2836 5780 2876
rect 1132 2752 1172 2792
rect 6508 2752 6548 2792
rect 1612 2668 1652 2708
rect 4492 2668 4532 2708
rect 1516 2584 1556 2624
rect 1804 2584 1844 2624
rect 2188 2584 2228 2624
rect 2572 2584 2612 2624
rect 4396 2584 4436 2624
rect 10252 2584 10292 2624
rect 1900 2500 1940 2540
rect 7756 2500 7796 2540
rect 11692 2416 11732 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 6124 2164 6164 2204
rect 460 2080 500 2120
rect 556 1996 596 2036
rect 1900 2080 1940 2120
rect 2476 2080 2516 2120
rect 6028 2080 6068 2120
rect 8716 2080 8756 2120
rect 4588 1996 4628 2036
rect 1420 1912 1460 1952
rect 2956 1912 2996 1952
rect 3724 1912 3764 1952
rect 4396 1912 4436 1952
rect 11692 1912 11732 1952
rect 1036 1828 1076 1868
rect 4780 1828 4820 1868
rect 5548 1828 5588 1868
rect 10444 1828 10484 1868
rect 940 1744 980 1784
rect 3436 1744 3476 1784
rect 844 1576 884 1616
rect 5740 1576 5780 1616
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 7948 1408 7988 1448
rect 8908 1408 8948 1448
rect 10444 904 10484 944
<< metal3 >>
rect 1976 47280 2056 47360
rect 2360 47280 2440 47360
rect 2744 47280 2824 47360
rect 3128 47280 3208 47360
rect 3512 47280 3592 47360
rect 3896 47280 3976 47360
rect 4280 47280 4360 47360
rect 4664 47280 4744 47360
rect 5048 47280 5128 47360
rect 5432 47280 5512 47360
rect 5816 47280 5896 47360
rect 6200 47280 6280 47360
rect 6584 47280 6664 47360
rect 6968 47280 7048 47360
rect 7352 47280 7432 47360
rect 7736 47280 7816 47360
rect 8120 47280 8200 47360
rect 8504 47280 8584 47360
rect 8888 47280 8968 47360
rect 9272 47280 9352 47360
rect 9656 47280 9736 47360
rect 1996 45212 2036 47280
rect 1996 45163 2036 45172
rect 2380 45212 2420 47280
rect 2380 45163 2420 45172
rect 2092 45128 2132 45137
rect 1324 45044 1364 45053
rect 748 44792 788 44801
rect 172 44372 212 44381
rect 76 44288 116 44297
rect 76 44153 116 44248
rect 76 43952 116 43961
rect 172 43952 212 44332
rect 652 44204 692 44213
rect 116 43912 212 43952
rect 556 44036 596 44045
rect 76 43903 116 43912
rect 268 42020 308 42029
rect 268 39920 308 41980
rect 268 39871 308 39880
rect 460 41180 500 41189
rect 364 38156 404 38165
rect 364 37568 404 38116
rect 364 37519 404 37528
rect 460 36644 500 41140
rect 460 36595 500 36604
rect 460 35972 500 35981
rect 76 34208 116 34217
rect 76 34073 116 34168
rect 460 32192 500 35932
rect 460 32143 500 32152
rect 364 31688 404 31697
rect 268 29252 308 29261
rect 268 26816 308 29212
rect 364 27740 404 31648
rect 460 31100 500 31109
rect 460 28160 500 31060
rect 460 28111 500 28120
rect 364 27700 500 27740
rect 268 26767 308 26776
rect 364 27572 404 27581
rect 364 25472 404 27532
rect 364 25423 404 25432
rect 460 24380 500 27700
rect 460 24331 500 24340
rect 460 23792 500 23801
rect 76 22448 116 22457
rect 76 22313 116 22408
rect 172 22280 212 22289
rect 76 17744 116 17753
rect 76 16232 116 17704
rect 76 16183 116 16192
rect 172 16904 212 22240
rect 364 21776 404 21785
rect 268 21104 308 21113
rect 268 19508 308 21064
rect 268 19459 308 19468
rect 364 19340 404 21736
rect 460 21524 500 23752
rect 556 22280 596 43996
rect 652 42272 692 44164
rect 652 42223 692 42232
rect 748 38156 788 44752
rect 940 43280 980 43289
rect 652 38116 788 38156
rect 844 39584 884 39593
rect 844 38156 884 39544
rect 652 29252 692 38116
rect 844 38107 884 38116
rect 748 37736 788 37745
rect 748 34964 788 37696
rect 844 36644 884 36653
rect 844 35132 884 36604
rect 844 35083 884 35092
rect 748 34924 884 34964
rect 748 33620 788 33629
rect 748 30512 788 33580
rect 844 32024 884 34924
rect 844 31975 884 31984
rect 748 30463 788 30472
rect 844 31772 884 31781
rect 844 29924 884 31732
rect 844 29875 884 29884
rect 652 29212 884 29252
rect 748 29084 788 29093
rect 748 26144 788 29044
rect 748 26095 788 26104
rect 652 26060 692 26069
rect 652 24800 692 26020
rect 652 24751 692 24760
rect 844 24548 884 29212
rect 844 24499 884 24508
rect 652 24464 692 24473
rect 652 23036 692 24424
rect 844 24380 884 24389
rect 748 24128 788 24137
rect 748 23120 788 24088
rect 748 23071 788 23080
rect 652 22987 692 22996
rect 556 22231 596 22240
rect 460 21475 500 21484
rect 556 22112 596 22121
rect 364 19291 404 19300
rect 460 20768 500 20777
rect 172 15476 212 16864
rect 172 15427 212 15436
rect 364 18080 404 18089
rect 76 15224 116 15233
rect 76 15056 116 15184
rect 76 15007 116 15016
rect 364 14972 404 18040
rect 460 17828 500 20728
rect 556 20012 596 22072
rect 556 19963 596 19972
rect 652 21440 692 21449
rect 460 17779 500 17788
rect 556 19760 596 19769
rect 364 14923 404 14932
rect 460 17408 500 17417
rect 460 14888 500 17368
rect 556 16988 596 19720
rect 652 18500 692 21400
rect 652 18451 692 18460
rect 748 18752 788 18761
rect 556 16939 596 16948
rect 460 14839 500 14848
rect 652 16736 692 16745
rect 652 14132 692 16696
rect 748 16316 788 18712
rect 748 16267 788 16276
rect 652 14083 692 14092
rect 556 14048 596 14057
rect 460 12284 500 12293
rect 172 11696 212 11705
rect 172 9596 212 11656
rect 460 10352 500 12244
rect 556 11192 596 14008
rect 556 11143 596 11152
rect 652 13376 692 13385
rect 652 10436 692 13336
rect 652 10387 692 10396
rect 748 13040 788 13049
rect 460 10303 500 10312
rect 748 10352 788 13000
rect 748 10303 788 10312
rect 172 9547 212 9556
rect 748 9008 788 9017
rect 556 8672 596 8681
rect 172 6656 212 6665
rect 172 2876 212 6616
rect 172 2827 212 2836
rect 460 4640 500 4649
rect 460 2120 500 4600
rect 460 2071 500 2080
rect 556 2036 596 8632
rect 748 6656 788 8968
rect 748 6607 788 6616
rect 844 5480 884 24340
rect 940 23060 980 43240
rect 1324 42944 1364 45004
rect 1900 44036 1940 44045
rect 1804 43532 1844 43541
rect 1324 42895 1364 42904
rect 1708 43448 1748 43457
rect 1324 42692 1364 42701
rect 1036 42104 1076 42113
rect 1036 40256 1076 42064
rect 1324 40928 1364 42652
rect 1516 42692 1556 42701
rect 1516 41348 1556 42652
rect 1516 41299 1556 41308
rect 1324 40879 1364 40888
rect 1420 41180 1460 41189
rect 1324 40508 1364 40517
rect 1036 40207 1076 40216
rect 1132 40340 1172 40349
rect 1036 37568 1076 37577
rect 1036 35216 1076 37528
rect 1036 35167 1076 35176
rect 1036 34544 1076 34553
rect 1036 34409 1076 34504
rect 1132 33704 1172 40300
rect 1324 39248 1364 40468
rect 1420 39668 1460 41140
rect 1612 41012 1652 41021
rect 1612 40877 1652 40972
rect 1420 39619 1460 39628
rect 1516 39836 1556 39845
rect 1324 39199 1364 39208
rect 1516 38240 1556 39796
rect 1516 38191 1556 38200
rect 1420 38156 1460 38165
rect 1228 37652 1268 37661
rect 1228 35552 1268 37612
rect 1324 37484 1364 37493
rect 1324 36896 1364 37444
rect 1324 36847 1364 36856
rect 1228 35503 1268 35512
rect 1324 35972 1364 35981
rect 1420 35972 1460 38116
rect 1612 38072 1652 38081
rect 1516 37232 1556 37241
rect 1516 37097 1556 37192
rect 1420 35932 1556 35972
rect 1036 33664 1172 33704
rect 1228 34460 1268 34469
rect 1036 31520 1076 33664
rect 1132 33536 1172 33545
rect 1132 32864 1172 33496
rect 1132 32815 1172 32824
rect 1036 31471 1076 31480
rect 1132 32024 1172 32033
rect 1036 31352 1076 31361
rect 1036 27824 1076 31312
rect 1036 27775 1076 27784
rect 1036 27488 1076 27497
rect 1036 26564 1076 27448
rect 1036 26515 1076 26524
rect 1132 24968 1172 31984
rect 1228 31184 1268 34420
rect 1324 32528 1364 35932
rect 1420 35804 1460 35813
rect 1420 33536 1460 35764
rect 1516 33872 1556 35932
rect 1516 33823 1556 33832
rect 1420 33487 1460 33496
rect 1516 33704 1556 33713
rect 1516 33284 1556 33664
rect 1516 33235 1556 33244
rect 1324 32479 1364 32488
rect 1420 33032 1460 33041
rect 1420 32108 1460 32992
rect 1612 32864 1652 38032
rect 1708 33116 1748 43408
rect 1804 42608 1844 43492
rect 1804 42559 1844 42568
rect 1804 41768 1844 41777
rect 1804 40592 1844 41728
rect 1804 40543 1844 40552
rect 1804 38996 1844 39005
rect 1804 35216 1844 38956
rect 1804 35167 1844 35176
rect 1804 34964 1844 34973
rect 1804 33536 1844 34924
rect 1804 33487 1844 33496
rect 1900 33140 1940 43996
rect 1996 42776 2036 42785
rect 1996 37904 2036 42736
rect 1996 37855 2036 37864
rect 1996 36056 2036 36065
rect 1996 34628 2036 36016
rect 1996 34579 2036 34588
rect 1996 34460 2036 34469
rect 1996 33620 2036 34420
rect 1996 33571 2036 33580
rect 2092 33956 2132 45088
rect 2668 45044 2708 45053
rect 2284 44876 2324 44885
rect 2188 42692 2228 42701
rect 2188 41600 2228 42652
rect 2188 41551 2228 41560
rect 2284 37652 2324 44836
rect 2668 44624 2708 45004
rect 2764 44960 2804 47280
rect 3148 45128 3188 47280
rect 2764 44911 2804 44920
rect 3052 45088 3188 45128
rect 2668 44575 2708 44584
rect 3052 44540 3092 45088
rect 3340 45044 3380 45053
rect 3148 44960 3188 44969
rect 3188 44920 3284 44960
rect 3148 44911 3188 44920
rect 3052 44491 3092 44500
rect 2476 44288 2516 44297
rect 2476 43700 2516 44248
rect 2476 42692 2516 43660
rect 2476 42643 2516 42652
rect 2956 44288 2996 44297
rect 2380 42608 2420 42617
rect 2380 40508 2420 42568
rect 2380 40340 2420 40468
rect 2956 42608 2996 44248
rect 3244 44036 3284 44920
rect 3148 43364 3188 43373
rect 3148 43229 3188 43324
rect 3244 43028 3284 43996
rect 3244 42979 3284 42988
rect 2572 40340 2612 40349
rect 2380 40300 2516 40340
rect 2476 38492 2516 40300
rect 2476 38156 2516 38452
rect 2476 38107 2516 38116
rect 2572 39332 2612 40300
rect 2956 39752 2996 42568
rect 3244 42440 3284 42449
rect 3148 42188 3188 42283
rect 3148 42139 3188 42148
rect 3148 42020 3188 42029
rect 3052 41852 3092 41861
rect 3052 41717 3092 41812
rect 3148 41264 3188 41980
rect 3148 41215 3188 41224
rect 2956 39703 2996 39712
rect 3052 41012 3092 41021
rect 2572 37988 2612 39292
rect 2668 39668 2708 39677
rect 2668 38996 2708 39628
rect 3052 39668 3092 40972
rect 3052 39619 3092 39628
rect 2956 39584 2996 39593
rect 2860 39500 2900 39509
rect 2860 39365 2900 39460
rect 2668 38947 2708 38956
rect 2956 38576 2996 39544
rect 3148 39080 3188 39089
rect 2476 37948 2612 37988
rect 2764 38536 2996 38576
rect 3052 38996 3092 39005
rect 2188 37612 2324 37652
rect 2380 37904 2420 37913
rect 2188 35384 2228 37612
rect 2284 37484 2324 37493
rect 2284 37349 2324 37444
rect 2284 36980 2324 36989
rect 2284 35468 2324 36940
rect 2284 35419 2324 35428
rect 2188 35335 2228 35344
rect 1708 33067 1748 33076
rect 1804 33100 1940 33140
rect 1804 32948 1844 33100
rect 1612 32815 1652 32824
rect 1708 32908 1844 32948
rect 1900 33032 1940 33041
rect 1420 31772 1460 32068
rect 1612 32696 1652 32705
rect 1420 31723 1460 31732
rect 1516 31940 1556 31949
rect 1228 31135 1268 31144
rect 1324 31436 1364 31445
rect 1516 31436 1556 31900
rect 1228 31016 1268 31025
rect 1228 28412 1268 30976
rect 1324 30848 1364 31396
rect 1420 31396 1556 31436
rect 1420 31268 1460 31396
rect 1420 31219 1460 31228
rect 1516 31184 1556 31193
rect 1324 30799 1364 30808
rect 1420 30932 1460 30941
rect 1420 30176 1460 30892
rect 1516 30932 1556 31144
rect 1516 30883 1556 30892
rect 1420 30127 1460 30136
rect 1516 30764 1556 30773
rect 1420 30008 1460 30017
rect 1324 29840 1364 29849
rect 1324 29705 1364 29800
rect 1228 28363 1268 28372
rect 1324 29084 1364 29093
rect 1324 27152 1364 29044
rect 1420 27572 1460 29968
rect 1516 29168 1556 30724
rect 1516 29119 1556 29128
rect 1420 27523 1460 27532
rect 1516 27740 1556 27749
rect 1324 27103 1364 27112
rect 1420 27404 1460 27413
rect 1228 26900 1268 26909
rect 1228 25136 1268 26860
rect 1228 25087 1268 25096
rect 1132 24928 1268 24968
rect 1228 23060 1268 24928
rect 940 23020 1076 23060
rect 1228 23020 1364 23060
rect 940 19424 980 19433
rect 940 19289 980 19384
rect 940 18416 980 18425
rect 940 14720 980 18376
rect 1036 16568 1076 23020
rect 1132 22952 1172 22961
rect 1132 20180 1172 22912
rect 1228 22784 1268 22793
rect 1228 20852 1268 22744
rect 1228 20803 1268 20812
rect 1132 20131 1172 20140
rect 1228 20432 1268 20441
rect 1036 16519 1076 16528
rect 1132 19928 1172 19937
rect 1132 17912 1172 19888
rect 1228 19340 1268 20392
rect 1228 19291 1268 19300
rect 1324 17996 1364 23020
rect 1420 19844 1460 27364
rect 1516 26480 1556 27700
rect 1516 26431 1556 26440
rect 1516 23876 1556 23885
rect 1516 20936 1556 23836
rect 1516 20887 1556 20896
rect 1516 20096 1556 20105
rect 1516 19961 1556 20056
rect 1420 19804 1556 19844
rect 1420 19676 1460 19685
rect 1420 19340 1460 19636
rect 1420 19291 1460 19300
rect 1420 19088 1460 19097
rect 1420 18668 1460 19048
rect 1420 18619 1460 18628
rect 1516 18668 1556 19804
rect 1516 18619 1556 18628
rect 940 14671 980 14680
rect 1036 16400 1076 16409
rect 940 14552 980 14561
rect 940 8000 980 14512
rect 1036 13796 1076 16360
rect 1132 15056 1172 17872
rect 1132 15007 1172 15016
rect 1228 17956 1364 17996
rect 1516 18500 1556 18509
rect 1228 14552 1268 17956
rect 1420 17072 1460 17081
rect 1228 14503 1268 14512
rect 1324 15728 1364 15737
rect 1324 14132 1364 15688
rect 1420 15644 1460 17032
rect 1420 15595 1460 15604
rect 1324 14083 1364 14092
rect 1036 13747 1076 13756
rect 1420 14048 1460 14057
rect 1324 13712 1364 13721
rect 1228 12452 1268 12461
rect 1228 12317 1268 12412
rect 1228 11360 1268 11369
rect 1132 11024 1172 11033
rect 940 7951 980 7960
rect 1036 10688 1076 10697
rect 844 5431 884 5440
rect 940 5648 980 5657
rect 556 1987 596 1996
rect 844 4304 884 4313
rect 844 1616 884 4264
rect 940 1784 980 5608
rect 1036 3716 1076 10648
rect 1132 9428 1172 10984
rect 1228 9596 1268 11320
rect 1324 11192 1364 13672
rect 1420 13544 1460 14008
rect 1420 13495 1460 13504
rect 1324 11143 1364 11152
rect 1420 11276 1460 11285
rect 1420 10184 1460 11236
rect 1420 10135 1460 10144
rect 1324 9596 1364 9605
rect 1228 9556 1324 9596
rect 1324 9547 1364 9556
rect 1132 9379 1172 9388
rect 1420 9512 1460 9521
rect 1420 9377 1460 9472
rect 1132 8000 1172 8009
rect 1132 4388 1172 7960
rect 1420 7328 1460 7337
rect 1324 7244 1364 7253
rect 1324 7109 1364 7204
rect 1132 4339 1172 4348
rect 1228 5984 1268 5993
rect 1036 3667 1076 3676
rect 1132 3968 1172 3977
rect 1036 3296 1076 3305
rect 1036 1868 1076 3256
rect 1132 2792 1172 3928
rect 1228 3380 1268 5944
rect 1228 3331 1268 3340
rect 1324 5312 1364 5321
rect 1324 3296 1364 5272
rect 1420 3548 1460 7288
rect 1516 7076 1556 18460
rect 1612 16652 1652 32656
rect 1708 30260 1748 32908
rect 1708 30211 1748 30220
rect 1804 32780 1844 32789
rect 1708 29924 1748 29933
rect 1708 28832 1748 29884
rect 1708 28783 1748 28792
rect 1708 28412 1748 28421
rect 1708 27488 1748 28372
rect 1708 27439 1748 27448
rect 1708 27320 1748 27329
rect 1708 23960 1748 27280
rect 1804 27152 1844 32740
rect 1804 27103 1844 27112
rect 1900 30680 1940 32992
rect 2092 32948 2132 33916
rect 1900 29924 1940 30640
rect 1996 32908 2092 32948
rect 1996 30596 2036 32908
rect 2092 32899 2132 32908
rect 2188 35216 2228 35225
rect 2188 34376 2228 35176
rect 2284 35216 2324 35225
rect 2284 34712 2324 35176
rect 2284 34663 2324 34672
rect 1996 30547 2036 30556
rect 2092 31604 2132 31613
rect 1900 27656 1940 29884
rect 1804 26732 1844 26741
rect 1804 25388 1844 26692
rect 1900 26144 1940 27616
rect 1900 26095 1940 26104
rect 1996 30260 2036 30269
rect 1996 27488 2036 30220
rect 1996 26900 2036 27448
rect 1996 26060 2036 26860
rect 1996 26011 2036 26020
rect 1804 25339 1844 25348
rect 1708 23624 1748 23920
rect 1708 23575 1748 23584
rect 1804 24716 1844 24725
rect 1708 22868 1748 22879
rect 1708 22784 1748 22828
rect 1708 22735 1748 22744
rect 1804 22364 1844 24676
rect 1996 24548 2036 24557
rect 1804 22315 1844 22324
rect 1900 23120 1940 23129
rect 1900 21608 1940 23080
rect 1996 23036 2036 24508
rect 2092 23876 2132 31564
rect 2188 31436 2228 34336
rect 2380 34124 2420 37864
rect 2476 36644 2516 37948
rect 2764 37652 2804 38536
rect 2668 37612 2804 37652
rect 2668 36812 2708 37612
rect 2668 36763 2708 36772
rect 2764 37484 2804 37493
rect 2476 36595 2516 36604
rect 2572 36644 2612 36653
rect 2476 36476 2516 36485
rect 2476 34964 2516 36436
rect 2572 36056 2612 36604
rect 2572 36007 2612 36016
rect 2668 35972 2708 35981
rect 2476 34915 2516 34924
rect 2572 35468 2612 35477
rect 2284 34084 2420 34124
rect 2476 34712 2516 34721
rect 2284 31604 2324 34084
rect 2284 31555 2324 31564
rect 2380 33200 2420 33209
rect 2188 31396 2324 31436
rect 2092 23827 2132 23836
rect 2188 31184 2228 31193
rect 1996 22987 2036 22996
rect 2092 22952 2132 22961
rect 2092 22532 2132 22912
rect 2092 22483 2132 22492
rect 1900 21559 1940 21568
rect 1996 22364 2036 22373
rect 1612 16603 1652 16612
rect 1708 21020 1748 21029
rect 1708 18584 1748 20980
rect 1900 20936 1940 20945
rect 1804 20180 1844 20189
rect 1804 20012 1844 20140
rect 1804 19963 1844 19972
rect 1804 19844 1844 19853
rect 1804 19709 1844 19804
rect 1612 16484 1652 16493
rect 1612 13292 1652 16444
rect 1708 14972 1748 18544
rect 1900 19592 1940 20896
rect 1900 18584 1940 19552
rect 1996 19508 2036 22324
rect 2092 21692 2132 21701
rect 2092 21020 2132 21652
rect 2092 20971 2132 20980
rect 1996 19256 2036 19468
rect 1996 19207 2036 19216
rect 2092 20768 2132 20777
rect 2092 20012 2132 20728
rect 2092 19172 2132 19972
rect 2092 19123 2132 19132
rect 1900 17912 1940 18544
rect 2092 18668 2132 18677
rect 1900 17863 1940 17872
rect 1996 18416 2036 18425
rect 1996 17828 2036 18376
rect 1900 17744 1940 17753
rect 1708 14923 1748 14932
rect 1804 16820 1844 16829
rect 1652 13252 1748 13292
rect 1612 13243 1652 13252
rect 1612 12956 1652 12965
rect 1612 11780 1652 12916
rect 1612 8756 1652 11740
rect 1708 8840 1748 13252
rect 1804 12032 1844 16780
rect 1900 15728 1940 17704
rect 1996 16820 2036 17788
rect 1996 16771 2036 16780
rect 1900 15679 1940 15688
rect 1996 15476 2036 15485
rect 1900 15392 1940 15401
rect 1900 12704 1940 15352
rect 1900 12655 1940 12664
rect 1804 11983 1844 11992
rect 1900 12536 1940 12545
rect 1804 11528 1844 11537
rect 1804 10184 1844 11488
rect 1804 10135 1844 10144
rect 1804 10016 1844 10025
rect 1804 9008 1844 9976
rect 1804 8959 1844 8968
rect 1708 8800 1844 8840
rect 1804 8756 1844 8800
rect 1612 8716 1748 8756
rect 1516 7027 1556 7036
rect 1612 8588 1652 8597
rect 1612 7916 1652 8548
rect 1612 6656 1652 7876
rect 1516 6616 1652 6656
rect 1708 7160 1748 8716
rect 1804 8707 1844 8716
rect 1516 5732 1556 6616
rect 1612 6488 1652 6497
rect 1612 6353 1652 6448
rect 1708 6404 1748 7120
rect 1708 6355 1748 6364
rect 1804 6992 1844 7001
rect 1516 4892 1556 5692
rect 1516 4388 1556 4852
rect 1516 4339 1556 4348
rect 1612 4472 1652 4481
rect 1612 3632 1652 4432
rect 1420 3499 1460 3508
rect 1516 3592 1652 3632
rect 1324 3247 1364 3256
rect 1132 2743 1172 2752
rect 1420 3212 1460 3221
rect 1420 1952 1460 3172
rect 1516 2624 1556 3592
rect 1612 3464 1652 3473
rect 1612 2708 1652 3424
rect 1612 2659 1652 2668
rect 1516 2575 1556 2584
rect 1804 2624 1844 6952
rect 1900 5648 1940 12496
rect 1996 11780 2036 15436
rect 1996 11731 2036 11740
rect 1900 5599 1940 5608
rect 1996 11612 2036 11621
rect 1900 4808 1940 4817
rect 1900 4673 1940 4768
rect 1900 4304 1940 4313
rect 1900 4169 1940 4264
rect 1804 2575 1844 2584
rect 1900 2540 1940 2549
rect 1900 2120 1940 2500
rect 1900 2071 1940 2080
rect 1420 1903 1460 1912
rect 1036 1819 1076 1828
rect 940 1735 980 1744
rect 844 1567 884 1576
rect 1996 80 2036 11572
rect 2092 5900 2132 18628
rect 2188 11948 2228 31144
rect 2284 27404 2324 31396
rect 2284 25808 2324 27364
rect 2284 25759 2324 25768
rect 2380 29168 2420 33160
rect 2380 27656 2420 29128
rect 2476 29084 2516 34672
rect 2572 33704 2612 35428
rect 2668 35384 2708 35932
rect 2668 35335 2708 35344
rect 2668 35132 2708 35227
rect 2668 35083 2708 35092
rect 2572 33655 2612 33664
rect 2668 34964 2708 34973
rect 2572 33536 2612 33545
rect 2572 33140 2612 33496
rect 2572 33091 2612 33100
rect 2668 33032 2708 34924
rect 2476 28496 2516 29044
rect 2572 32992 2708 33032
rect 2572 29000 2612 32992
rect 2668 32864 2708 32873
rect 2668 32108 2708 32824
rect 2668 31772 2708 32068
rect 2668 31723 2708 31732
rect 2572 28951 2612 28960
rect 2668 31436 2708 31445
rect 2476 28447 2516 28456
rect 2572 28832 2612 28841
rect 2284 25220 2324 25229
rect 2284 23960 2324 25180
rect 2380 24548 2420 27616
rect 2572 26900 2612 28792
rect 2668 28580 2708 31396
rect 2668 28531 2708 28540
rect 2668 28412 2708 28421
rect 2668 27068 2708 28372
rect 2668 27019 2708 27028
rect 2572 26851 2612 26860
rect 2380 24499 2420 24508
rect 2476 26312 2516 26321
rect 2284 23911 2324 23920
rect 2284 23624 2324 23633
rect 2284 21692 2324 23584
rect 2476 23060 2516 26272
rect 2572 26144 2612 26153
rect 2572 25388 2612 26104
rect 2572 25339 2612 25348
rect 2284 21643 2324 21652
rect 2380 23020 2516 23060
rect 2572 24380 2612 24389
rect 2572 24044 2612 24340
rect 2572 23036 2612 24004
rect 2284 21524 2324 21533
rect 2284 20012 2324 21484
rect 2284 18752 2324 19972
rect 2284 18500 2324 18712
rect 2284 17744 2324 18460
rect 2284 17695 2324 17704
rect 2284 14720 2324 14729
rect 2284 14585 2324 14680
rect 2284 13964 2324 13973
rect 2284 13040 2324 13924
rect 2284 12991 2324 13000
rect 2188 11899 2228 11908
rect 2284 12872 2324 12881
rect 2284 11780 2324 12832
rect 2092 5851 2132 5860
rect 2188 11740 2324 11780
rect 2188 5564 2228 11740
rect 2284 10940 2324 10949
rect 2284 10772 2324 10900
rect 2284 10268 2324 10732
rect 2284 9428 2324 10228
rect 2284 9379 2324 9388
rect 2284 9008 2324 9017
rect 2284 7412 2324 8968
rect 2284 7363 2324 7372
rect 2188 5515 2228 5524
rect 2284 7244 2324 7253
rect 2284 5060 2324 7204
rect 2188 5020 2324 5060
rect 2092 4892 2132 4901
rect 2092 4724 2132 4852
rect 2092 4675 2132 4684
rect 2188 4136 2228 5020
rect 2188 4087 2228 4096
rect 2188 3464 2228 3473
rect 2188 3329 2228 3424
rect 2188 2876 2228 2885
rect 2188 2624 2228 2836
rect 2188 2575 2228 2584
rect 2380 80 2420 23020
rect 2572 22987 2612 22996
rect 2764 22952 2804 37444
rect 2956 37484 2996 37493
rect 2860 37316 2900 37325
rect 2860 35216 2900 37276
rect 2956 35720 2996 37444
rect 3052 36224 3092 38956
rect 3052 36175 3092 36184
rect 2956 35671 2996 35680
rect 3052 36056 3092 36065
rect 3052 35468 3092 36016
rect 3052 35384 3092 35428
rect 2860 35167 2900 35176
rect 2956 35344 3092 35384
rect 2956 34964 2996 35344
rect 2860 34924 2996 34964
rect 3052 35216 3092 35225
rect 2860 34544 2900 34924
rect 2860 34495 2900 34504
rect 2956 34628 2996 34637
rect 2956 33452 2996 34588
rect 3052 33620 3092 35176
rect 3052 33571 3092 33580
rect 3148 33452 3188 39040
rect 3244 37652 3284 42400
rect 3244 37603 3284 37612
rect 2860 33412 2996 33452
rect 3052 33412 3188 33452
rect 3244 37484 3284 37493
rect 2860 32780 2900 33412
rect 2860 32731 2900 32740
rect 2956 33284 2996 33293
rect 2956 33032 2996 33244
rect 2956 32612 2996 32992
rect 2956 32563 2996 32572
rect 2956 31772 2996 31781
rect 2860 31352 2900 31361
rect 2860 30764 2900 31312
rect 2860 30715 2900 30724
rect 2956 30596 2996 31732
rect 2956 30547 2996 30556
rect 2956 30428 2996 30437
rect 2956 30092 2996 30388
rect 2860 30052 2996 30092
rect 2860 29756 2900 30052
rect 3052 29840 3092 33412
rect 3148 33284 3188 33293
rect 3148 32360 3188 33244
rect 3244 32780 3284 37444
rect 3340 33704 3380 45004
rect 3436 44288 3476 44297
rect 3436 43616 3476 44248
rect 3436 43567 3476 43576
rect 3436 43364 3476 43404
rect 3436 43280 3476 43324
rect 3436 41180 3476 43240
rect 3532 42944 3572 47280
rect 3916 45212 3956 47280
rect 3916 45163 3956 45172
rect 4300 45212 4340 47280
rect 4300 45163 4340 45172
rect 4684 45212 4724 47280
rect 5068 46136 5108 47280
rect 5068 46096 5396 46136
rect 4928 45380 5296 45389
rect 4968 45340 5010 45380
rect 5050 45340 5092 45380
rect 5132 45340 5174 45380
rect 5214 45340 5256 45380
rect 4928 45331 5296 45340
rect 4684 45163 4724 45172
rect 5164 45212 5204 45221
rect 4588 44960 4628 44969
rect 3688 44624 4056 44633
rect 3728 44584 3770 44624
rect 3810 44584 3852 44624
rect 3892 44584 3934 44624
rect 3974 44584 4016 44624
rect 3688 44575 4056 44584
rect 4492 44120 4532 44129
rect 4492 44036 4532 44080
rect 4492 43985 4532 43996
rect 4396 43784 4436 43793
rect 3724 43700 3764 43709
rect 3724 43364 3764 43660
rect 4300 43532 4340 43541
rect 3724 43315 3764 43324
rect 4204 43448 4244 43457
rect 4204 43313 4244 43408
rect 4300 43220 4340 43492
rect 4396 43364 4436 43744
rect 4588 43448 4628 44920
rect 4972 44960 5012 44969
rect 4588 43399 4628 43408
rect 4684 44288 4724 44297
rect 4684 43952 4724 44248
rect 4972 44120 5012 44920
rect 5164 44456 5204 45172
rect 5356 45212 5396 46096
rect 5356 45163 5396 45172
rect 5452 45128 5492 47280
rect 5644 45296 5684 45305
rect 5452 45079 5492 45088
rect 5548 45212 5588 45221
rect 5356 44960 5396 44969
rect 5164 44407 5204 44416
rect 5260 44876 5300 44885
rect 5260 44372 5300 44836
rect 5356 44540 5396 44920
rect 5356 44491 5396 44500
rect 5260 44323 5300 44332
rect 4972 44071 5012 44080
rect 4684 43616 4724 43912
rect 5356 43952 5396 43961
rect 4928 43868 5296 43877
rect 4968 43828 5010 43868
rect 5050 43828 5092 43868
rect 5132 43828 5174 43868
rect 5214 43828 5256 43868
rect 4928 43819 5296 43828
rect 4396 43315 4436 43324
rect 4300 43180 4628 43220
rect 3688 43112 4056 43121
rect 3728 43072 3770 43112
rect 3810 43072 3852 43112
rect 3892 43072 3934 43112
rect 3974 43072 4016 43112
rect 3688 43063 4056 43072
rect 4492 43112 4532 43121
rect 3532 42895 3572 42904
rect 3916 42944 3956 42953
rect 3436 40340 3476 41140
rect 3436 39416 3476 40300
rect 3436 39367 3476 39376
rect 3532 42776 3572 42785
rect 3532 42104 3572 42736
rect 3916 42524 3956 42904
rect 3916 42475 3956 42484
rect 4492 42188 4532 43072
rect 4588 42692 4628 43180
rect 4588 42643 4628 42652
rect 4588 42524 4628 42533
rect 4588 42389 4628 42484
rect 4684 42272 4724 43576
rect 5356 43616 5396 43912
rect 5356 43567 5396 43576
rect 4780 43364 4820 43373
rect 4780 43280 4820 43324
rect 4780 43229 4820 43240
rect 4780 42944 4820 42953
rect 4780 42356 4820 42904
rect 5548 42944 5588 45172
rect 5644 44036 5684 45256
rect 5836 45212 5876 47280
rect 5836 45163 5876 45172
rect 6220 45212 6260 47280
rect 6220 45163 6260 45172
rect 6604 45212 6644 47280
rect 6604 45163 6644 45172
rect 6988 45212 7028 47280
rect 6988 45163 7028 45172
rect 7372 45212 7412 47280
rect 7372 45163 7412 45172
rect 7756 45212 7796 47280
rect 7756 45163 7796 45172
rect 8140 45212 8180 47280
rect 8140 45163 8180 45172
rect 8524 45212 8564 47280
rect 8524 45163 8564 45172
rect 8908 45212 8948 47280
rect 8908 45163 8948 45172
rect 9292 45212 9332 47280
rect 9292 45163 9332 45172
rect 9676 45212 9716 47280
rect 9676 45163 9716 45172
rect 10252 46304 10292 46313
rect 6124 45044 6164 45053
rect 5644 43987 5684 43996
rect 5740 44960 5780 44969
rect 5644 43868 5684 43877
rect 5644 43616 5684 43828
rect 5740 43784 5780 44920
rect 6124 44456 6164 45004
rect 6124 44407 6164 44416
rect 6508 44960 6548 44969
rect 6508 44456 6548 44920
rect 7276 44960 7316 44969
rect 6508 44407 6548 44416
rect 6796 44708 6836 44717
rect 6796 44456 6836 44668
rect 6796 44407 6836 44416
rect 7276 44456 7316 44920
rect 8044 44960 8084 44969
rect 7276 44407 7316 44416
rect 7756 44876 7796 44885
rect 7948 44876 7988 44885
rect 7756 44456 7796 44836
rect 7756 44407 7796 44416
rect 7852 44836 7948 44876
rect 6316 44288 6356 44297
rect 6316 44153 6356 44248
rect 6796 44288 6836 44297
rect 6412 44204 6452 44213
rect 5836 44120 5876 44131
rect 5836 44036 5876 44080
rect 5836 43987 5876 43996
rect 6220 44120 6260 44129
rect 5740 43735 5780 43744
rect 5644 43576 5780 43616
rect 5548 42895 5588 42904
rect 5644 43448 5684 43457
rect 5548 42692 5588 42701
rect 4780 42307 4820 42316
rect 4928 42356 5296 42365
rect 4968 42316 5010 42356
rect 5050 42316 5092 42356
rect 5132 42316 5174 42356
rect 5214 42316 5256 42356
rect 4928 42307 5296 42316
rect 4684 42223 4724 42232
rect 4492 42139 4532 42148
rect 3532 41096 3572 42064
rect 5548 42104 5588 42652
rect 5644 42188 5684 43408
rect 5644 42139 5684 42148
rect 4780 42020 4820 42029
rect 4588 41936 4628 41945
rect 3688 41600 4056 41609
rect 3728 41560 3770 41600
rect 3810 41560 3852 41600
rect 3892 41560 3934 41600
rect 3974 41560 4016 41600
rect 3688 41551 4056 41560
rect 3532 39248 3572 41056
rect 4108 40508 4148 40517
rect 3688 40088 4056 40097
rect 3728 40048 3770 40088
rect 3810 40048 3852 40088
rect 3892 40048 3934 40088
rect 3974 40048 4016 40088
rect 3688 40039 4056 40048
rect 4012 39920 4052 39929
rect 3436 39208 3572 39248
rect 3820 39332 3860 39341
rect 3436 36644 3476 39208
rect 3820 39080 3860 39292
rect 3820 39031 3860 39040
rect 3532 38996 3572 39005
rect 3532 36812 3572 38956
rect 4012 38996 4052 39880
rect 4012 38947 4052 38956
rect 4108 39752 4148 40468
rect 4396 40508 4436 40517
rect 3628 38912 3668 38921
rect 3628 38777 3668 38872
rect 3688 38576 4056 38585
rect 3728 38536 3770 38576
rect 3810 38536 3852 38576
rect 3892 38536 3934 38576
rect 3974 38536 4016 38576
rect 3688 38527 4056 38536
rect 3688 37064 4056 37073
rect 3728 37024 3770 37064
rect 3810 37024 3852 37064
rect 3892 37024 3934 37064
rect 3974 37024 4016 37064
rect 3688 37015 4056 37024
rect 3532 36763 3572 36772
rect 4012 36812 4052 36821
rect 4012 36644 4052 36772
rect 4108 36812 4148 39712
rect 4300 40424 4340 40433
rect 4300 40256 4340 40384
rect 4300 39668 4340 40216
rect 4300 39332 4340 39628
rect 4300 39283 4340 39292
rect 4396 39500 4436 40468
rect 4300 38996 4340 39005
rect 4204 38912 4244 38921
rect 4204 37316 4244 38872
rect 4300 38156 4340 38956
rect 4300 38107 4340 38116
rect 4204 37267 4244 37276
rect 4300 37400 4340 37409
rect 4108 36763 4148 36772
rect 4204 36644 4244 36653
rect 3436 36604 3668 36644
rect 4012 36604 4148 36644
rect 3532 36476 3572 36485
rect 3532 36341 3572 36436
rect 3532 35972 3572 35981
rect 3436 35888 3476 35897
rect 3436 34544 3476 35848
rect 3436 34495 3476 34504
rect 3532 34460 3572 35932
rect 3628 35972 3668 36604
rect 3628 35923 3668 35932
rect 3688 35552 4056 35561
rect 3728 35512 3770 35552
rect 3810 35512 3852 35552
rect 3892 35512 3934 35552
rect 3974 35512 4016 35552
rect 3688 35503 4056 35512
rect 3724 35384 3764 35393
rect 3436 34376 3476 34385
rect 3436 33788 3476 34336
rect 3436 33739 3476 33748
rect 3340 33655 3380 33664
rect 3436 33620 3476 33629
rect 3340 33452 3380 33461
rect 3340 32948 3380 33412
rect 3340 32899 3380 32908
rect 3244 32740 3380 32780
rect 3148 32311 3188 32320
rect 3244 32612 3284 32621
rect 2860 29716 2996 29756
rect 2860 29252 2900 29261
rect 2860 29000 2900 29212
rect 2860 28951 2900 28960
rect 2860 27572 2900 27667
rect 2860 27523 2900 27532
rect 2860 27320 2900 27329
rect 2860 27185 2900 27280
rect 2860 26984 2900 26993
rect 2860 26849 2900 26944
rect 2956 26900 2996 29716
rect 3052 29000 3092 29800
rect 3148 32192 3188 32201
rect 3148 31352 3188 32152
rect 3148 29252 3188 31312
rect 3244 30764 3284 32572
rect 3340 31352 3380 32740
rect 3436 31520 3476 33580
rect 3532 33536 3572 34420
rect 3628 35300 3668 35309
rect 3628 34376 3668 35260
rect 3724 35216 3764 35344
rect 3724 35167 3764 35176
rect 3916 34964 3956 34973
rect 3916 34829 3956 34924
rect 3628 34327 3668 34336
rect 3688 34040 4056 34049
rect 3728 34000 3770 34040
rect 3810 34000 3852 34040
rect 3892 34000 3934 34040
rect 3974 34000 4016 34040
rect 3688 33991 4056 34000
rect 3916 33872 3956 33881
rect 3532 33487 3572 33496
rect 3628 33704 3668 33713
rect 3628 33284 3668 33664
rect 3532 32864 3572 32873
rect 3532 32192 3572 32824
rect 3628 32696 3668 33244
rect 3916 33032 3956 33832
rect 3916 32983 3956 32992
rect 3628 32647 3668 32656
rect 3688 32528 4056 32537
rect 3728 32488 3770 32528
rect 3810 32488 3852 32528
rect 3892 32488 3934 32528
rect 3974 32488 4016 32528
rect 3688 32479 4056 32488
rect 3532 32143 3572 32152
rect 3628 32360 3668 32369
rect 3436 31471 3476 31480
rect 3532 31436 3572 31445
rect 3340 31312 3476 31352
rect 3244 30715 3284 30724
rect 3244 30428 3284 30437
rect 3244 30008 3284 30388
rect 3244 29959 3284 29968
rect 3340 30344 3380 30353
rect 3148 29203 3188 29212
rect 3244 29756 3284 29765
rect 3148 29084 3188 29093
rect 3148 29000 3188 29044
rect 3052 28960 3188 29000
rect 3244 29000 3284 29716
rect 3244 28832 3284 28960
rect 3148 28792 3284 28832
rect 2956 26851 2996 26860
rect 3052 28748 3092 28757
rect 2956 25388 2996 25397
rect 2956 24800 2996 25348
rect 2956 24751 2996 24760
rect 3052 24548 3092 28708
rect 3052 24499 3092 24508
rect 3148 25388 3188 28792
rect 3052 23960 3092 23969
rect 2956 23792 2996 23801
rect 2956 23540 2996 23752
rect 2668 22912 2804 22952
rect 2860 23500 2996 23540
rect 2668 22868 2708 22912
rect 2476 22828 2708 22868
rect 2476 16316 2516 22828
rect 2860 22700 2900 23500
rect 3052 23372 3092 23920
rect 2764 22660 2900 22700
rect 2956 23332 3092 23372
rect 2572 22364 2612 22373
rect 2572 19424 2612 22324
rect 2668 22280 2708 22291
rect 2668 22196 2708 22240
rect 2668 22147 2708 22156
rect 2764 21776 2804 22660
rect 2860 22532 2900 22541
rect 2860 22397 2900 22492
rect 2764 21727 2804 21736
rect 2860 22280 2900 22289
rect 2860 21608 2900 22240
rect 2956 22196 2996 23332
rect 3148 23204 3188 25348
rect 3244 28664 3284 28673
rect 3244 24716 3284 28624
rect 3340 28664 3380 30304
rect 3340 28615 3380 28624
rect 3436 28664 3476 31312
rect 3532 30260 3572 31396
rect 3628 31184 3668 32320
rect 4012 32360 4052 32369
rect 4012 32108 4052 32320
rect 4012 31520 4052 32068
rect 4012 31471 4052 31480
rect 3628 31135 3668 31144
rect 3688 31016 4056 31025
rect 3728 30976 3770 31016
rect 3810 30976 3852 31016
rect 3892 30976 3934 31016
rect 3974 30976 4016 31016
rect 3688 30967 4056 30976
rect 3916 30848 3956 30857
rect 3628 30680 3668 30775
rect 3628 30631 3668 30640
rect 3820 30596 3860 30605
rect 3628 30428 3668 30523
rect 3628 30379 3668 30388
rect 3532 30220 3668 30260
rect 3436 28615 3476 28624
rect 3532 30008 3572 30017
rect 3532 29000 3572 29968
rect 3628 29756 3668 30220
rect 3820 30008 3860 30556
rect 3820 29873 3860 29968
rect 3628 29707 3668 29716
rect 3724 29672 3764 29681
rect 3820 29672 3860 29681
rect 3764 29632 3820 29672
rect 3724 29623 3764 29632
rect 3820 29623 3860 29632
rect 3916 29672 3956 30808
rect 4012 30680 4052 30775
rect 4012 30631 4052 30640
rect 4012 30428 4052 30437
rect 4012 30176 4052 30388
rect 4108 30260 4148 36604
rect 4204 36140 4244 36604
rect 4300 36476 4340 37360
rect 4300 36427 4340 36436
rect 4204 36091 4244 36100
rect 4396 36392 4436 39460
rect 4204 35972 4244 35981
rect 4204 33872 4244 35932
rect 4204 33823 4244 33832
rect 4300 33956 4340 33965
rect 4300 33620 4340 33916
rect 4300 33368 4340 33580
rect 4300 33319 4340 33328
rect 4300 32948 4340 32957
rect 4204 32696 4244 32705
rect 4204 32192 4244 32656
rect 4204 32143 4244 32152
rect 4300 31940 4340 32908
rect 4300 31268 4340 31900
rect 4300 31219 4340 31228
rect 4204 30512 4244 30523
rect 4204 30428 4244 30472
rect 4204 30379 4244 30388
rect 4300 30428 4340 30437
rect 4108 30220 4244 30260
rect 4012 29924 4052 30136
rect 4052 29884 4148 29924
rect 4012 29875 4052 29884
rect 3916 29623 3956 29632
rect 3688 29504 4056 29513
rect 3728 29464 3770 29504
rect 3810 29464 3852 29504
rect 3892 29464 3934 29504
rect 3974 29464 4016 29504
rect 3688 29455 4056 29464
rect 4012 29252 4052 29261
rect 3436 28496 3476 28505
rect 3340 28412 3380 28421
rect 3340 26312 3380 28372
rect 3340 26060 3380 26272
rect 3340 26011 3380 26020
rect 3244 24667 3284 24676
rect 3244 24548 3284 24557
rect 3244 24044 3284 24508
rect 3244 23995 3284 24004
rect 3148 23120 3188 23164
rect 3052 23080 3188 23120
rect 3244 23288 3284 23297
rect 3052 22868 3092 23080
rect 3244 23036 3284 23248
rect 3052 22819 3092 22828
rect 3148 22996 3244 23036
rect 2956 22147 2996 22156
rect 3052 22700 3092 22709
rect 2764 21568 2900 21608
rect 2668 21440 2708 21449
rect 2668 19928 2708 21400
rect 2668 19879 2708 19888
rect 2612 19384 2708 19424
rect 2572 19375 2612 19384
rect 2572 19256 2612 19265
rect 2572 18416 2612 19216
rect 2572 18367 2612 18376
rect 2668 19088 2708 19384
rect 2764 19256 2804 21568
rect 3052 20936 3092 22660
rect 2956 20896 3092 20936
rect 2860 20264 2900 20273
rect 2860 20129 2900 20224
rect 2764 19207 2804 19216
rect 2476 16267 2516 16276
rect 2572 16652 2612 16661
rect 2572 16148 2612 16612
rect 2476 16108 2612 16148
rect 2476 11276 2516 16108
rect 2668 16064 2708 19048
rect 2956 18416 2996 20896
rect 3148 20852 3188 22996
rect 3244 22987 3284 22996
rect 2956 18367 2996 18376
rect 3052 20812 3148 20852
rect 3052 19676 3092 20812
rect 3148 20803 3188 20812
rect 3340 22952 3380 22961
rect 3340 20936 3380 22912
rect 3436 22700 3476 28456
rect 3532 27068 3572 28960
rect 3724 29000 3764 29009
rect 3724 28580 3764 28960
rect 3724 28531 3764 28540
rect 4012 28412 4052 29212
rect 4012 28160 4052 28372
rect 4108 29084 4148 29884
rect 4204 29252 4244 30220
rect 4204 29203 4244 29212
rect 4300 29168 4340 30388
rect 4396 29756 4436 36352
rect 4492 39584 4532 39593
rect 4492 34544 4532 39544
rect 4588 36812 4628 41896
rect 4684 41012 4724 41021
rect 4684 39668 4724 40972
rect 4684 39619 4724 39628
rect 4780 39500 4820 41980
rect 5452 41936 5492 41945
rect 4928 40844 5296 40853
rect 4968 40804 5010 40844
rect 5050 40804 5092 40844
rect 5132 40804 5174 40844
rect 5214 40804 5256 40844
rect 4928 40795 5296 40804
rect 4780 39451 4820 39460
rect 5356 40508 5396 40517
rect 4780 39332 4820 39341
rect 4780 37652 4820 39292
rect 4928 39332 5296 39341
rect 4968 39292 5010 39332
rect 5050 39292 5092 39332
rect 5132 39292 5174 39332
rect 5214 39292 5256 39332
rect 4928 39283 5296 39292
rect 5356 39332 5396 40468
rect 5356 39283 5396 39292
rect 5356 38576 5396 38585
rect 5356 38324 5396 38536
rect 5356 38275 5396 38284
rect 4928 37820 5296 37829
rect 4968 37780 5010 37820
rect 5050 37780 5092 37820
rect 5132 37780 5174 37820
rect 5214 37780 5256 37820
rect 4928 37771 5296 37780
rect 4780 37612 4916 37652
rect 4780 37400 4820 37409
rect 4588 36772 4724 36812
rect 4588 36644 4628 36653
rect 4588 35804 4628 36604
rect 4588 35755 4628 35764
rect 4532 34504 4628 34544
rect 4492 34495 4532 34504
rect 4396 29707 4436 29716
rect 4492 34208 4532 34217
rect 4300 29119 4340 29128
rect 4108 28328 4148 29044
rect 4492 29084 4532 34168
rect 4588 33620 4628 34504
rect 4588 33571 4628 33580
rect 4492 29035 4532 29044
rect 4588 33452 4628 33461
rect 4108 28279 4148 28288
rect 4204 29000 4244 29009
rect 4204 28580 4244 28960
rect 4012 28111 4052 28120
rect 3688 27992 4056 28001
rect 3728 27952 3770 27992
rect 3810 27952 3852 27992
rect 3892 27952 3934 27992
rect 3974 27952 4016 27992
rect 3688 27943 4056 27952
rect 3532 27019 3572 27028
rect 3688 26480 4056 26489
rect 3728 26440 3770 26480
rect 3810 26440 3852 26480
rect 3892 26440 3934 26480
rect 3974 26440 4016 26480
rect 3688 26431 4056 26440
rect 3916 26060 3956 26069
rect 3820 25892 3860 25901
rect 3820 25388 3860 25852
rect 3820 25136 3860 25348
rect 3916 25388 3956 26020
rect 4108 25892 4148 25901
rect 4108 25472 4148 25852
rect 4108 25423 4148 25432
rect 3916 25304 3956 25348
rect 3916 25253 3956 25264
rect 4108 25304 4148 25313
rect 4108 25136 4148 25264
rect 3820 25096 4148 25136
rect 3688 24968 4056 24977
rect 3728 24928 3770 24968
rect 3810 24928 3852 24968
rect 3892 24928 3934 24968
rect 3974 24928 4016 24968
rect 3688 24919 4056 24928
rect 3916 24380 3956 24389
rect 3916 24245 3956 24340
rect 4108 23792 4148 25096
rect 3688 23456 4056 23465
rect 3728 23416 3770 23456
rect 3810 23416 3852 23456
rect 3892 23416 3934 23456
rect 3974 23416 4016 23456
rect 3688 23407 4056 23416
rect 4012 23120 4052 23215
rect 4012 23071 4052 23080
rect 4012 22952 4052 22961
rect 3436 22651 3476 22660
rect 3724 22868 3764 22877
rect 3532 22364 3572 22373
rect 3436 22324 3532 22364
rect 3436 21692 3476 22324
rect 3532 22229 3572 22324
rect 3724 22112 3764 22828
rect 4012 22448 4052 22912
rect 4012 22399 4052 22408
rect 3724 22063 3764 22072
rect 3688 21944 4056 21953
rect 3728 21904 3770 21944
rect 3810 21904 3852 21944
rect 3892 21904 3934 21944
rect 3974 21904 4016 21944
rect 3688 21895 4056 21904
rect 3436 21643 3476 21652
rect 3148 20600 3188 20609
rect 3148 20180 3188 20560
rect 3340 20516 3380 20896
rect 3628 21608 3668 21617
rect 3628 21104 3668 21568
rect 4012 21608 4052 21617
rect 3628 20684 3668 21064
rect 3916 21272 3956 21281
rect 3916 20852 3956 21232
rect 3916 20717 3956 20812
rect 3628 20635 3668 20644
rect 4012 20684 4052 21568
rect 4108 21524 4148 23752
rect 4204 23288 4244 28540
rect 4396 29000 4436 29009
rect 4300 28244 4340 28253
rect 4300 27236 4340 28204
rect 4300 27187 4340 27196
rect 4396 27068 4436 28960
rect 4588 28748 4628 33412
rect 4684 33284 4724 36772
rect 4684 33235 4724 33244
rect 4780 35888 4820 37360
rect 4876 36896 4916 37612
rect 4876 36728 4916 36856
rect 5068 37484 5108 37493
rect 5068 36812 5108 37444
rect 5068 36763 5108 36772
rect 5356 37484 5396 37493
rect 4876 36679 4916 36688
rect 4928 36308 5296 36317
rect 4968 36268 5010 36308
rect 5050 36268 5092 36308
rect 5132 36268 5174 36308
rect 5214 36268 5256 36308
rect 4928 36259 5296 36268
rect 4780 31604 4820 35848
rect 5260 35888 5300 35897
rect 5164 35804 5204 35813
rect 5164 35384 5204 35764
rect 5260 35753 5300 35848
rect 5164 35335 5204 35344
rect 5356 35300 5396 37444
rect 5356 35251 5396 35260
rect 5356 35132 5396 35141
rect 4928 34796 5296 34805
rect 4968 34756 5010 34796
rect 5050 34756 5092 34796
rect 5132 34756 5174 34796
rect 5214 34756 5256 34796
rect 4928 34747 5296 34756
rect 4876 34544 4916 34553
rect 4876 33788 4916 34504
rect 5356 34460 5396 35092
rect 5356 34411 5396 34420
rect 4876 33739 4916 33748
rect 5356 34208 5396 34217
rect 4928 33284 5296 33293
rect 4968 33244 5010 33284
rect 5050 33244 5092 33284
rect 5132 33244 5174 33284
rect 5214 33244 5256 33284
rect 4928 33235 5296 33244
rect 5260 33032 5300 33041
rect 5260 32948 5300 32992
rect 5260 32897 5300 32908
rect 5356 32948 5396 34168
rect 5452 33452 5492 41896
rect 5548 39332 5588 42064
rect 5740 41180 5780 43576
rect 5836 43532 5876 43541
rect 5836 43364 5876 43492
rect 5836 43315 5876 43324
rect 5836 43196 5876 43205
rect 5836 42440 5876 43156
rect 5932 42944 5972 42953
rect 5932 42809 5972 42904
rect 5932 42692 5972 42701
rect 5932 42524 5972 42652
rect 6220 42608 6260 44080
rect 6220 42559 6260 42568
rect 6316 43952 6356 43961
rect 5932 42475 5972 42484
rect 5836 42391 5876 42400
rect 6220 42440 6260 42449
rect 5932 42188 5972 42197
rect 5548 37316 5588 39292
rect 5644 41140 5780 41180
rect 5836 41348 5876 41357
rect 5644 37484 5684 41140
rect 5740 41012 5780 41021
rect 5740 40877 5780 40972
rect 5836 40424 5876 41308
rect 5836 40375 5876 40384
rect 5932 39752 5972 42148
rect 6124 40928 6164 40937
rect 6124 40508 6164 40888
rect 6124 40340 6164 40468
rect 6124 40291 6164 40300
rect 5740 39712 5972 39752
rect 6028 39752 6068 39761
rect 5740 38324 5780 39712
rect 5836 38912 5876 38921
rect 5836 38777 5876 38872
rect 6028 38660 6068 39712
rect 6124 39668 6164 39677
rect 6124 39080 6164 39628
rect 6124 39031 6164 39040
rect 6028 38611 6068 38620
rect 5740 38275 5780 38284
rect 6124 38492 6164 38501
rect 5740 38156 5780 38165
rect 5740 37652 5780 38116
rect 6028 38156 6068 38165
rect 5740 37603 5780 37612
rect 5836 38072 5876 38081
rect 5644 37435 5684 37444
rect 5548 37267 5588 37276
rect 5644 37316 5684 37325
rect 5548 37148 5588 37157
rect 5548 36812 5588 37108
rect 5548 36763 5588 36772
rect 5644 36728 5684 37276
rect 5740 36812 5780 36907
rect 5740 36763 5780 36772
rect 5452 33403 5492 33412
rect 5548 36644 5588 36653
rect 5356 32899 5396 32908
rect 5452 33032 5492 33041
rect 4876 31940 4916 32035
rect 4876 31891 4916 31900
rect 4928 31772 5296 31781
rect 4968 31732 5010 31772
rect 5050 31732 5092 31772
rect 5132 31732 5174 31772
rect 5214 31732 5256 31772
rect 4928 31723 5296 31732
rect 4780 31555 4820 31564
rect 5356 31520 5396 31529
rect 4588 28699 4628 28708
rect 4684 31436 4724 31445
rect 4300 27028 4436 27068
rect 4588 27572 4628 27581
rect 4300 26312 4340 27028
rect 4300 26228 4340 26272
rect 4492 26984 4532 26993
rect 4300 26188 4436 26228
rect 4300 26060 4340 26069
rect 4300 25925 4340 26020
rect 4396 25556 4436 26188
rect 4300 25516 4396 25556
rect 4300 25472 4340 25516
rect 4396 25507 4436 25516
rect 4300 25423 4340 25432
rect 4396 25388 4436 25397
rect 4396 25253 4436 25348
rect 4396 24548 4436 24557
rect 4396 24044 4436 24508
rect 4396 23995 4436 24004
rect 4492 24464 4532 26944
rect 4588 26900 4628 27532
rect 4684 27068 4724 31396
rect 4780 31268 4820 31277
rect 4780 30092 4820 31228
rect 4928 30260 5296 30269
rect 4968 30220 5010 30260
rect 5050 30220 5092 30260
rect 5132 30220 5174 30260
rect 5214 30220 5256 30260
rect 4928 30211 5296 30220
rect 4876 30092 4916 30101
rect 4780 30052 4876 30092
rect 4876 30043 4916 30052
rect 4972 30008 5012 30017
rect 4780 29924 4820 29933
rect 4780 29789 4820 29884
rect 4972 29873 5012 29968
rect 5356 30008 5396 31480
rect 5452 31100 5492 32992
rect 5548 31520 5588 36604
rect 5644 36140 5684 36688
rect 5644 35804 5684 36100
rect 5740 36644 5780 36653
rect 5740 36056 5780 36604
rect 5740 36007 5780 36016
rect 5644 35764 5780 35804
rect 5644 35300 5684 35309
rect 5644 33704 5684 35260
rect 5644 33655 5684 33664
rect 5644 33368 5684 33377
rect 5644 33032 5684 33328
rect 5644 32983 5684 32992
rect 5548 31471 5588 31480
rect 5644 31940 5684 31949
rect 5548 31352 5588 31361
rect 5548 31217 5588 31312
rect 5452 31060 5588 31100
rect 5356 29959 5396 29968
rect 5452 30596 5492 30605
rect 4876 29840 4916 29849
rect 4684 27019 4724 27028
rect 4780 29168 4820 29177
rect 4780 28412 4820 29128
rect 4876 29000 4916 29800
rect 5164 29840 5204 29849
rect 5164 29252 5204 29800
rect 5452 29756 5492 30556
rect 5548 29924 5588 31060
rect 5548 29875 5588 29884
rect 5452 29707 5492 29716
rect 5548 29756 5588 29765
rect 5164 29203 5204 29212
rect 5452 29588 5492 29597
rect 4876 28951 4916 28960
rect 5356 29084 5396 29093
rect 4928 28748 5296 28757
rect 4968 28708 5010 28748
rect 5050 28708 5092 28748
rect 5132 28708 5174 28748
rect 5214 28708 5256 28748
rect 4928 28699 5296 28708
rect 4588 26732 4628 26860
rect 4588 26683 4628 26692
rect 4684 26648 4724 26657
rect 4204 23239 4244 23248
rect 4396 23204 4436 23213
rect 4108 21475 4148 21484
rect 4204 23120 4244 23129
rect 4012 20635 4052 20644
rect 4108 20600 4148 20609
rect 3340 20476 3438 20516
rect 3398 20348 3438 20476
rect 3688 20432 4056 20441
rect 3728 20392 3770 20432
rect 3810 20392 3852 20432
rect 3892 20392 3934 20432
rect 3974 20392 4016 20432
rect 3688 20383 4056 20392
rect 3398 20308 3476 20348
rect 3148 20131 3188 20140
rect 3340 20180 3380 20189
rect 3052 18500 3092 19636
rect 3148 20012 3188 20021
rect 3148 19172 3188 19972
rect 3148 19123 3188 19132
rect 2956 18248 2996 18257
rect 2956 17912 2996 18208
rect 2572 16024 2708 16064
rect 2764 17872 2996 17912
rect 2572 14804 2612 16024
rect 2764 14888 2804 17872
rect 3052 17828 3092 18460
rect 3052 17779 3092 17788
rect 3244 18500 3284 18509
rect 2956 17660 2996 17669
rect 2956 16988 2996 17620
rect 2956 16316 2996 16948
rect 2956 16267 2996 16276
rect 3052 17660 3092 17669
rect 2860 16232 2900 16241
rect 2860 14972 2900 16192
rect 2956 15812 2996 15821
rect 2956 15560 2996 15772
rect 3052 15644 3092 17620
rect 3052 15595 3092 15604
rect 2956 15511 2996 15520
rect 3148 15140 3188 15149
rect 2860 14923 2900 14932
rect 3052 15056 3092 15065
rect 2764 14839 2804 14848
rect 2956 14888 2996 14897
rect 2572 14720 2612 14764
rect 2860 14804 2900 14813
rect 2572 14671 2612 14680
rect 2668 14720 2708 14729
rect 2572 14132 2612 14141
rect 2572 12536 2612 14092
rect 2668 12620 2708 14680
rect 2764 14720 2804 14729
rect 2764 13964 2804 14680
rect 2860 14048 2900 14764
rect 2860 13999 2900 14008
rect 2764 12872 2804 13924
rect 2764 12823 2804 12832
rect 2860 13124 2900 13133
rect 2860 12704 2900 13084
rect 2860 12655 2900 12664
rect 2668 12571 2708 12580
rect 2572 12487 2612 12496
rect 2764 12452 2804 12461
rect 2476 11227 2516 11236
rect 2668 11780 2708 11789
rect 2476 11108 2516 11117
rect 2476 9176 2516 11068
rect 2476 9127 2516 9136
rect 2668 7916 2708 11740
rect 2764 10940 2804 12412
rect 2860 11948 2900 11957
rect 2860 11864 2900 11908
rect 2860 11813 2900 11824
rect 2860 11108 2900 11203
rect 2860 11059 2900 11068
rect 2956 11024 2996 14848
rect 3052 14720 3092 15016
rect 3052 13964 3092 14680
rect 3052 13915 3092 13924
rect 3052 13796 3092 13805
rect 3052 11948 3092 13756
rect 3052 11899 3092 11908
rect 2956 10975 2996 10984
rect 2860 10940 2900 10949
rect 2764 10900 2860 10940
rect 2860 10872 2900 10900
rect 2956 10016 2996 10025
rect 2956 9512 2996 9976
rect 2956 9463 2996 9472
rect 3052 9680 3092 9689
rect 2956 9344 2996 9353
rect 2860 8924 2900 8933
rect 2860 8789 2900 8884
rect 2764 8756 2804 8765
rect 2764 7916 2804 8716
rect 2860 8672 2900 8681
rect 2860 8537 2900 8632
rect 2860 7916 2900 7925
rect 2764 7876 2860 7916
rect 2668 7244 2708 7876
rect 2860 7848 2900 7876
rect 2668 7195 2708 7204
rect 2956 6992 2996 9304
rect 3052 7076 3092 9640
rect 3052 7027 3092 7036
rect 2956 6943 2996 6952
rect 2956 6404 2996 6413
rect 2476 6320 2516 6329
rect 2476 2120 2516 6280
rect 2956 6236 2996 6364
rect 2764 6196 2996 6236
rect 2764 5732 2804 6196
rect 2572 5648 2612 5657
rect 2572 4724 2612 5608
rect 2572 4675 2612 4684
rect 2668 4892 2708 4901
rect 2764 4892 2804 5692
rect 2860 4892 2900 4901
rect 2764 4852 2860 4892
rect 2668 4136 2708 4852
rect 2860 4824 2900 4852
rect 2668 4087 2708 4096
rect 2956 2792 2996 2801
rect 2572 2624 2612 2633
rect 2572 2489 2612 2584
rect 2476 2071 2516 2080
rect 2956 1952 2996 2752
rect 2956 1903 2996 1912
rect 2764 272 2804 281
rect 2764 80 2804 232
rect 3148 80 3188 15100
rect 3244 8168 3284 18460
rect 3340 17240 3380 20140
rect 3436 19844 3476 20308
rect 3916 20264 3956 20273
rect 3436 19795 3476 19804
rect 3532 20180 3572 20189
rect 3532 19676 3572 20140
rect 3436 19636 3572 19676
rect 3436 17996 3476 19636
rect 3532 19508 3572 19517
rect 3532 18752 3572 19468
rect 3628 19424 3668 19433
rect 3628 19289 3668 19384
rect 3724 19340 3764 19349
rect 3724 19205 3764 19300
rect 3916 19088 3956 20224
rect 4012 20096 4052 20105
rect 4012 19340 4052 20056
rect 4108 20012 4148 20560
rect 4108 19963 4148 19972
rect 4012 19291 4052 19300
rect 3916 19039 3956 19048
rect 3688 18920 4056 18929
rect 3728 18880 3770 18920
rect 3810 18880 3852 18920
rect 3892 18880 3934 18920
rect 3974 18880 4016 18920
rect 3688 18871 4056 18880
rect 3532 18703 3572 18712
rect 3436 17947 3476 17956
rect 3532 18332 3572 18341
rect 3532 17912 3572 18292
rect 3532 17863 3572 17872
rect 3340 17191 3380 17200
rect 3436 17828 3476 17837
rect 3340 16904 3380 16913
rect 3340 16316 3380 16864
rect 3340 16267 3380 16276
rect 3340 14636 3380 14645
rect 3340 13460 3380 14596
rect 3436 13796 3476 17788
rect 3532 17744 3572 17753
rect 3532 17156 3572 17704
rect 4108 17744 4148 17753
rect 3688 17408 4056 17417
rect 3728 17368 3770 17408
rect 3810 17368 3852 17408
rect 3892 17368 3934 17408
rect 3974 17368 4016 17408
rect 3688 17359 4056 17368
rect 3820 17240 3860 17249
rect 4108 17240 4148 17704
rect 3532 17107 3572 17116
rect 3628 17156 3668 17165
rect 3628 17072 3668 17116
rect 3628 17021 3668 17032
rect 3724 16988 3764 16997
rect 3628 16904 3668 16913
rect 3628 16484 3668 16864
rect 3724 16853 3764 16948
rect 3628 16435 3668 16444
rect 3436 13747 3476 13756
rect 3532 16232 3572 16241
rect 3340 13411 3380 13420
rect 3436 13628 3476 13637
rect 3340 13124 3380 13219
rect 3340 13075 3380 13084
rect 3340 12956 3380 12965
rect 3340 12452 3380 12916
rect 3436 12788 3476 13588
rect 3532 12956 3572 16192
rect 3820 16064 3860 17200
rect 3916 17200 4148 17240
rect 3916 17072 3956 17200
rect 3916 16820 3956 17032
rect 4108 16904 4148 16913
rect 3916 16316 3956 16780
rect 4012 16820 4052 16829
rect 4012 16400 4052 16780
rect 4012 16351 4052 16360
rect 3916 16267 3956 16276
rect 4108 16232 4148 16864
rect 4108 16183 4148 16192
rect 3820 16024 4148 16064
rect 3688 15896 4056 15905
rect 3728 15856 3770 15896
rect 3810 15856 3852 15896
rect 3892 15856 3934 15896
rect 3974 15856 4016 15896
rect 3688 15847 4056 15856
rect 4012 15728 4052 15737
rect 3628 15644 3668 15653
rect 3628 14888 3668 15604
rect 3820 15560 3860 15569
rect 3820 15425 3860 15520
rect 4012 15476 4052 15688
rect 4012 15427 4052 15436
rect 3628 14839 3668 14848
rect 3724 14804 3764 14813
rect 3724 14669 3764 14764
rect 3688 14384 4056 14393
rect 3728 14344 3770 14384
rect 3810 14344 3852 14384
rect 3892 14344 3934 14384
rect 3974 14344 4016 14384
rect 3688 14335 4056 14344
rect 4108 14216 4148 16024
rect 4012 14176 4148 14216
rect 3724 14132 3764 14141
rect 3628 13964 3668 13973
rect 3628 13829 3668 13924
rect 3724 13376 3764 14092
rect 3724 13040 3764 13336
rect 3724 12991 3764 13000
rect 3916 13040 3956 13135
rect 3916 12991 3956 13000
rect 4012 12980 4052 14176
rect 4204 14132 4244 23080
rect 4396 23036 4436 23164
rect 4396 22868 4436 22996
rect 4300 22828 4436 22868
rect 4300 22280 4340 22828
rect 4300 22231 4340 22240
rect 4396 22700 4436 22709
rect 4300 22112 4340 22121
rect 4300 21356 4340 22072
rect 4300 20768 4340 21316
rect 4396 20852 4436 22660
rect 4396 20803 4436 20812
rect 4300 20180 4340 20728
rect 4300 20140 4436 20180
rect 4396 17912 4436 20140
rect 4492 19424 4532 24424
rect 4492 19375 4532 19384
rect 4588 24632 4628 24641
rect 4492 19256 4532 19265
rect 4492 17996 4532 19216
rect 4492 17947 4532 17956
rect 4300 17576 4340 17585
rect 4300 16064 4340 17536
rect 4396 16988 4436 17872
rect 4396 16939 4436 16948
rect 4492 17744 4532 17753
rect 4396 16820 4436 16829
rect 4396 16568 4436 16780
rect 4396 16519 4436 16528
rect 4396 16400 4436 16409
rect 4396 16148 4436 16360
rect 4396 16099 4436 16108
rect 4300 16015 4340 16024
rect 4300 15644 4340 15655
rect 4300 15560 4340 15604
rect 4300 15511 4340 15520
rect 4300 15308 4340 15317
rect 4300 15173 4340 15268
rect 4492 14972 4532 17704
rect 4492 14923 4532 14932
rect 4108 14092 4244 14132
rect 4108 13124 4148 14092
rect 4204 13964 4244 13973
rect 4204 13208 4244 13924
rect 4492 13796 4532 13805
rect 4204 13168 4340 13208
rect 4108 13084 4244 13124
rect 4012 12940 4148 12980
rect 3532 12907 3572 12916
rect 3688 12872 4056 12881
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 3688 12823 4056 12832
rect 3436 12739 3476 12748
rect 3532 12788 3572 12797
rect 3340 12403 3380 12412
rect 3244 8119 3284 8128
rect 3340 12284 3380 12293
rect 3244 7832 3284 7841
rect 3244 3548 3284 7792
rect 3340 6488 3380 12244
rect 3532 11948 3572 12748
rect 3724 12704 3764 12713
rect 4108 12704 4148 12940
rect 4204 12872 4244 13084
rect 4204 12823 4244 12832
rect 4108 12664 4244 12704
rect 3532 11899 3572 11908
rect 3628 12452 3668 12461
rect 3628 11780 3668 12412
rect 3628 11731 3668 11740
rect 3532 11696 3572 11705
rect 3532 11612 3572 11656
rect 3724 11612 3764 12664
rect 3916 12620 3956 12629
rect 3532 11572 3764 11612
rect 3820 11696 3860 11705
rect 3820 11561 3860 11656
rect 3916 11528 3956 12580
rect 3916 11479 3956 11488
rect 4108 11780 4148 11789
rect 3532 11444 3572 11453
rect 3532 10268 3572 11404
rect 3688 11360 4056 11369
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 3688 11311 4056 11320
rect 4012 11192 4052 11201
rect 3820 11024 3860 11033
rect 3820 10772 3860 10984
rect 3820 10723 3860 10732
rect 3436 10228 3572 10268
rect 3436 7832 3476 10228
rect 3436 7783 3476 7792
rect 3532 10100 3572 10109
rect 4012 10100 4052 11152
rect 4108 10436 4148 11740
rect 4108 10387 4148 10396
rect 4012 10060 4148 10100
rect 3532 8756 3572 10060
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 3820 9428 3860 9437
rect 3820 9293 3860 9388
rect 3340 6439 3380 6448
rect 3436 7664 3476 7673
rect 3244 3499 3284 3508
rect 3340 4304 3380 4313
rect 3340 3464 3380 4264
rect 3436 3632 3476 7624
rect 3532 6572 3572 8716
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 3628 7412 3668 7421
rect 3628 7277 3668 7372
rect 3724 7160 3764 7169
rect 3724 7025 3764 7120
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 3532 6523 3572 6532
rect 3628 6656 3668 6665
rect 3628 6404 3668 6616
rect 4012 6656 4052 6665
rect 3436 3583 3476 3592
rect 3532 6364 3668 6404
rect 3820 6572 3860 6581
rect 3340 3415 3380 3424
rect 3436 3212 3476 3221
rect 3436 2876 3476 3172
rect 3436 1784 3476 2836
rect 3436 1735 3476 1744
rect 3532 80 3572 6364
rect 3820 5480 3860 6532
rect 4012 6152 4052 6616
rect 4012 5480 4052 6112
rect 4108 6320 4148 10060
rect 4108 5732 4148 6280
rect 4108 5683 4148 5692
rect 4012 5440 4148 5480
rect 3820 5431 3860 5440
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 3916 4892 3956 4901
rect 3916 4388 3956 4852
rect 3916 4339 3956 4348
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 4108 3464 4148 5440
rect 4108 3415 4148 3424
rect 4204 2900 4244 12664
rect 4300 11192 4340 13168
rect 4300 11143 4340 11152
rect 4396 12452 4436 12461
rect 4396 10940 4436 12412
rect 4492 11864 4532 13756
rect 4588 13208 4628 24592
rect 4684 24044 4724 26608
rect 4780 26312 4820 28372
rect 5356 28328 5396 29044
rect 5356 28279 5396 28288
rect 4928 27236 5296 27245
rect 4968 27196 5010 27236
rect 5050 27196 5092 27236
rect 5132 27196 5174 27236
rect 5214 27196 5256 27236
rect 4928 27187 5296 27196
rect 4780 26263 4820 26272
rect 4972 26900 5012 26909
rect 4972 26060 5012 26860
rect 5068 26564 5108 26573
rect 5068 26144 5108 26524
rect 5068 26095 5108 26104
rect 5260 26228 5300 26237
rect 4972 26011 5012 26020
rect 5260 25892 5300 26188
rect 5260 25843 5300 25852
rect 4928 25724 5296 25733
rect 4968 25684 5010 25724
rect 5050 25684 5092 25724
rect 5132 25684 5174 25724
rect 5214 25684 5256 25724
rect 4928 25675 5296 25684
rect 5356 25304 5396 25313
rect 4928 24212 5296 24221
rect 4968 24172 5010 24212
rect 5050 24172 5092 24212
rect 5132 24172 5174 24212
rect 5214 24172 5256 24212
rect 4928 24163 5296 24172
rect 4684 24004 4820 24044
rect 4684 23792 4724 23801
rect 4684 21356 4724 23752
rect 4780 23036 4820 24004
rect 4972 23960 5012 23969
rect 4780 22987 4820 22996
rect 4876 23120 4916 23129
rect 4876 22985 4916 23080
rect 4684 21307 4724 21316
rect 4780 22868 4820 22877
rect 4684 20684 4724 20693
rect 4684 19256 4724 20644
rect 4780 20012 4820 22828
rect 4972 22868 5012 23920
rect 5356 23876 5396 25264
rect 5356 23827 5396 23836
rect 5260 23792 5300 23801
rect 4972 22819 5012 22828
rect 5068 23708 5108 23717
rect 5068 22868 5108 23668
rect 5260 23120 5300 23752
rect 5452 23456 5492 29548
rect 5548 29168 5588 29716
rect 5548 29119 5588 29128
rect 5644 27320 5684 31900
rect 5740 27740 5780 35764
rect 5740 27691 5780 27700
rect 5644 27271 5684 27280
rect 5644 27152 5684 27161
rect 5644 24716 5684 27112
rect 5644 24667 5684 24676
rect 5740 25808 5780 25817
rect 5740 24044 5780 25768
rect 5740 23995 5780 24004
rect 5452 23407 5492 23416
rect 5260 22952 5300 23080
rect 5260 22903 5300 22912
rect 5356 23204 5396 23213
rect 5068 22819 5108 22828
rect 4928 22700 5296 22709
rect 4968 22660 5010 22700
rect 5050 22660 5092 22700
rect 5132 22660 5174 22700
rect 5214 22660 5256 22700
rect 4928 22651 5296 22660
rect 5260 22532 5300 22543
rect 5260 22448 5300 22492
rect 5260 22399 5300 22408
rect 5068 22364 5108 22373
rect 5108 22324 5204 22364
rect 5068 22229 5108 22324
rect 4972 22196 5012 22205
rect 4972 21608 5012 22156
rect 4972 21559 5012 21568
rect 5068 21692 5108 21701
rect 5068 21557 5108 21652
rect 5164 21608 5204 22324
rect 5164 21559 5204 21568
rect 4928 21188 5296 21197
rect 4968 21148 5010 21188
rect 5050 21148 5092 21188
rect 5132 21148 5174 21188
rect 5214 21148 5256 21188
rect 4928 21139 5296 21148
rect 4972 21020 5012 21029
rect 4780 19963 4820 19972
rect 4876 20852 4916 20861
rect 4876 19844 4916 20812
rect 4684 19207 4724 19216
rect 4780 19804 4916 19844
rect 4972 19844 5012 20980
rect 5260 20852 5300 20861
rect 5068 20096 5108 20105
rect 5260 20096 5300 20812
rect 5108 20056 5300 20096
rect 5068 20047 5108 20056
rect 5260 20012 5300 20056
rect 5356 20096 5396 23164
rect 5548 23036 5588 23045
rect 5452 22952 5492 22963
rect 5452 22868 5492 22912
rect 5452 22819 5492 22828
rect 5452 22700 5492 22709
rect 5452 22196 5492 22660
rect 5452 22147 5492 22156
rect 5452 21524 5492 21533
rect 5452 20852 5492 21484
rect 5452 20803 5492 20812
rect 5356 20047 5396 20056
rect 5452 20684 5492 20693
rect 5260 19963 5300 19972
rect 4684 18668 4724 18677
rect 4684 13292 4724 18628
rect 4780 17828 4820 19804
rect 4972 19795 5012 19804
rect 5452 19844 5492 20644
rect 5452 19795 5492 19804
rect 4928 19676 5296 19685
rect 4968 19636 5010 19676
rect 5050 19636 5092 19676
rect 5132 19636 5174 19676
rect 5214 19636 5256 19676
rect 4928 19627 5296 19636
rect 5548 19592 5588 22996
rect 5644 23036 5684 23047
rect 5644 22952 5684 22996
rect 5644 22903 5684 22912
rect 5740 22868 5780 22877
rect 5644 22700 5684 22709
rect 5644 21860 5684 22660
rect 5644 21440 5684 21820
rect 5740 21524 5780 22828
rect 5836 21608 5876 38032
rect 6028 38021 6068 38116
rect 6028 37652 6068 37661
rect 6028 36140 6068 37612
rect 6028 36091 6068 36100
rect 6124 37484 6164 38452
rect 6028 35972 6068 35981
rect 5932 35468 5972 35477
rect 5932 31436 5972 35428
rect 6028 35216 6068 35932
rect 6028 35167 6068 35176
rect 6124 33620 6164 37444
rect 6220 36224 6260 42400
rect 6316 42020 6356 43912
rect 6316 41348 6356 41980
rect 6316 41299 6356 41308
rect 6220 36175 6260 36184
rect 6316 37988 6356 37997
rect 6220 36056 6260 36065
rect 6220 34964 6260 36016
rect 6220 34915 6260 34924
rect 6220 34208 6260 34217
rect 6220 33704 6260 34168
rect 6220 33655 6260 33664
rect 6124 33571 6164 33580
rect 6220 33452 6260 33461
rect 6028 33116 6068 33125
rect 6028 32108 6068 33076
rect 6124 32864 6164 32873
rect 6124 32729 6164 32824
rect 6028 32059 6068 32068
rect 6124 32612 6164 32621
rect 6124 31940 6164 32572
rect 6124 31891 6164 31900
rect 6124 31436 6164 31445
rect 5932 31396 6124 31436
rect 6028 31268 6068 31277
rect 6028 30680 6068 31228
rect 6028 30631 6068 30640
rect 6028 30428 6068 30437
rect 6028 29924 6068 30388
rect 6028 29875 6068 29884
rect 5932 29840 5972 29849
rect 5932 29705 5972 29800
rect 5932 29168 5972 29177
rect 5932 28412 5972 29128
rect 6124 28916 6164 31396
rect 6220 29084 6260 33412
rect 6220 29035 6260 29044
rect 6124 28876 6260 28916
rect 5932 28363 5972 28372
rect 6028 28832 6068 28841
rect 6028 27572 6068 28792
rect 5932 27532 6068 27572
rect 5932 26144 5972 27532
rect 6124 27488 6164 27497
rect 5932 24716 5972 26104
rect 6028 27404 6068 27413
rect 6028 25388 6068 27364
rect 6028 25339 6068 25348
rect 5932 24676 6068 24716
rect 5932 24548 5972 24557
rect 5932 23960 5972 24508
rect 6028 24128 6068 24676
rect 6028 24079 6068 24088
rect 5932 22196 5972 23920
rect 6124 23876 6164 27448
rect 6124 23741 6164 23836
rect 5932 22147 5972 22156
rect 6028 23288 6068 23297
rect 5836 21568 5972 21608
rect 5740 21475 5780 21484
rect 5644 21391 5684 21400
rect 5836 21440 5876 21449
rect 5932 21440 5972 21568
rect 6028 21566 6068 23248
rect 6124 23120 6164 23129
rect 6124 22532 6164 23080
rect 6220 22868 6260 28876
rect 6220 22819 6260 22828
rect 6124 22483 6164 22492
rect 6220 22700 6260 22709
rect 6124 22196 6164 22205
rect 6124 22061 6164 22156
rect 6028 21517 6068 21526
rect 5932 21400 6068 21440
rect 5740 20936 5780 20945
rect 5644 20852 5684 20861
rect 5644 20180 5684 20812
rect 5644 20131 5684 20140
rect 5740 20096 5780 20896
rect 5836 20768 5876 21400
rect 5836 20719 5876 20728
rect 5932 21020 5972 21029
rect 5740 20047 5780 20056
rect 5836 20600 5876 20609
rect 5452 19552 5588 19592
rect 5164 19508 5204 19517
rect 5164 19340 5204 19468
rect 5164 18500 5204 19300
rect 5164 18451 5204 18460
rect 5260 18332 5300 18427
rect 5260 18283 5300 18292
rect 5356 18248 5396 18257
rect 4928 18164 5296 18173
rect 4968 18124 5010 18164
rect 5050 18124 5092 18164
rect 5132 18124 5174 18164
rect 5214 18124 5256 18164
rect 4928 18115 5296 18124
rect 4780 17693 4820 17788
rect 5068 17996 5108 18005
rect 5068 17744 5108 17956
rect 5356 17912 5396 18208
rect 5356 17863 5396 17872
rect 4972 17704 5068 17744
rect 4876 17408 4916 17417
rect 4780 17240 4820 17335
rect 4780 17191 4820 17200
rect 4876 17072 4916 17368
rect 4876 17023 4916 17032
rect 4780 16988 4820 16997
rect 4780 13460 4820 16948
rect 4972 16904 5012 17704
rect 5068 17695 5108 17704
rect 4972 16855 5012 16864
rect 5164 16988 5204 16997
rect 5164 16853 5204 16948
rect 5260 16820 5300 16915
rect 5260 16771 5300 16780
rect 5356 16736 5396 16745
rect 4928 16652 5296 16661
rect 4968 16612 5010 16652
rect 5050 16612 5092 16652
rect 5132 16612 5174 16652
rect 5214 16612 5256 16652
rect 4928 16603 5296 16612
rect 4972 16484 5012 16493
rect 4972 16349 5012 16444
rect 5356 16484 5396 16696
rect 5356 16435 5396 16444
rect 5356 16316 5396 16325
rect 4876 16232 4916 16241
rect 4876 16097 4916 16192
rect 5356 15728 5396 16276
rect 5260 15476 5300 15485
rect 5260 15341 5300 15436
rect 4928 15140 5296 15149
rect 4968 15100 5010 15140
rect 5050 15100 5092 15140
rect 5132 15100 5174 15140
rect 5214 15100 5256 15140
rect 4928 15091 5296 15100
rect 4876 14888 4916 14897
rect 4876 14132 4916 14848
rect 5356 14804 5396 15688
rect 5356 14755 5396 14764
rect 4876 14083 4916 14092
rect 5356 14636 5396 14645
rect 4928 13628 5296 13637
rect 4968 13588 5010 13628
rect 5050 13588 5092 13628
rect 5132 13588 5174 13628
rect 5214 13588 5256 13628
rect 4928 13579 5296 13588
rect 4780 13411 4820 13420
rect 4684 13252 4916 13292
rect 4588 13168 4820 13208
rect 4492 11815 4532 11824
rect 4684 13040 4724 13049
rect 4396 10891 4436 10900
rect 4492 11696 4532 11705
rect 4492 11108 4532 11656
rect 4396 10772 4436 10781
rect 4300 10184 4340 10193
rect 4300 8924 4340 10144
rect 4396 10016 4436 10732
rect 4492 10184 4532 11068
rect 4492 10135 4532 10144
rect 4588 10268 4628 10277
rect 4588 10133 4628 10228
rect 4396 9967 4436 9976
rect 4300 8875 4340 8884
rect 4396 9260 4436 9269
rect 4300 5732 4340 5741
rect 4300 5597 4340 5692
rect 4108 2860 4244 2900
rect 4300 4136 4340 4145
rect 3688 2288 4056 2297
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 3688 2239 4056 2248
rect 3724 1952 3764 1961
rect 3724 1817 3764 1912
rect 4108 188 4148 2860
rect 3916 148 4148 188
rect 3916 80 3956 148
rect 4300 80 4340 4096
rect 4396 3548 4436 9220
rect 4492 8588 4532 8597
rect 4492 7916 4532 8548
rect 4492 7867 4532 7876
rect 4396 3499 4436 3508
rect 4492 7748 4532 7757
rect 4492 3380 4532 7708
rect 4588 6488 4628 6497
rect 4588 5984 4628 6448
rect 4588 5900 4628 5944
rect 4588 5851 4628 5860
rect 4588 5732 4628 5741
rect 4588 5312 4628 5692
rect 4588 5263 4628 5272
rect 4588 4892 4628 4987
rect 4588 4843 4628 4852
rect 4588 4640 4628 4649
rect 4588 4472 4628 4600
rect 4588 3464 4628 4432
rect 4588 3415 4628 3424
rect 4396 3340 4532 3380
rect 4396 2900 4436 3340
rect 4588 3296 4628 3305
rect 4396 2860 4532 2900
rect 4492 2708 4532 2860
rect 4492 2659 4532 2668
rect 4396 2624 4436 2633
rect 4396 1952 4436 2584
rect 4588 2036 4628 3256
rect 4588 1987 4628 1996
rect 4396 1903 4436 1912
rect 4684 80 4724 13000
rect 4780 12536 4820 13168
rect 4780 12487 4820 12496
rect 4876 12284 4916 13252
rect 5068 12788 5108 12797
rect 5068 12536 5108 12748
rect 5068 12487 5108 12496
rect 4780 12244 4916 12284
rect 4780 9512 4820 12244
rect 4928 12116 5296 12125
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 4928 12067 5296 12076
rect 4876 11780 4916 11789
rect 4876 10772 4916 11740
rect 4972 11444 5012 11453
rect 4972 11024 5012 11404
rect 4972 10975 5012 10984
rect 4876 10723 4916 10732
rect 4928 10604 5296 10613
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 4928 10555 5296 10564
rect 5260 10436 5300 10445
rect 4876 10268 4916 10277
rect 4876 9848 4916 10228
rect 4876 9799 4916 9808
rect 5260 10100 5300 10396
rect 4780 9463 4820 9472
rect 5260 9428 5300 10060
rect 5260 9379 5300 9388
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 5260 7916 5300 7925
rect 5260 7781 5300 7876
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 4780 6404 4820 6413
rect 4780 5816 4820 6364
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 4780 5648 4820 5776
rect 4780 5608 4916 5648
rect 4780 5480 4820 5489
rect 4780 1868 4820 5440
rect 4876 4976 4916 5608
rect 4972 5480 5012 5489
rect 4972 5228 5012 5440
rect 4972 5179 5012 5188
rect 4876 4927 4916 4936
rect 4972 4892 5012 4901
rect 4972 4757 5012 4852
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 4780 1819 4820 1828
rect 4928 1532 5296 1541
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 4928 1483 5296 1492
rect 5356 1364 5396 14596
rect 5452 13124 5492 19552
rect 5548 19424 5588 19433
rect 5548 14720 5588 19384
rect 5644 18836 5684 18845
rect 5644 17996 5684 18796
rect 5644 17947 5684 17956
rect 5644 17828 5684 17837
rect 5644 16484 5684 17788
rect 5836 17324 5876 20560
rect 5932 19928 5972 20980
rect 6028 20096 6068 21400
rect 6124 20852 6164 20861
rect 6124 20264 6164 20812
rect 6124 20215 6164 20224
rect 6028 20056 6164 20096
rect 5932 19879 5972 19888
rect 5932 19760 5972 19769
rect 5932 19625 5972 19720
rect 6028 19676 6068 19685
rect 5932 18500 5972 18509
rect 5932 17660 5972 18460
rect 5932 17611 5972 17620
rect 5836 17275 5876 17284
rect 5740 17072 5780 17081
rect 5740 16937 5780 17032
rect 5932 16988 5972 16997
rect 5644 16435 5684 16444
rect 5836 16904 5876 16913
rect 5740 16316 5780 16325
rect 5740 16232 5780 16276
rect 5740 16181 5780 16192
rect 5548 14671 5588 14680
rect 5644 15896 5684 15905
rect 5452 13075 5492 13084
rect 5548 14552 5588 14561
rect 5068 1324 5396 1364
rect 5452 11948 5492 11957
rect 5068 80 5108 1324
rect 5452 80 5492 11908
rect 5548 10772 5588 14512
rect 5644 13208 5684 15856
rect 5740 15728 5780 15737
rect 5740 15560 5780 15688
rect 5740 15511 5780 15520
rect 5740 14804 5780 14813
rect 5740 14048 5780 14764
rect 5740 13999 5780 14008
rect 5644 13159 5684 13168
rect 5740 13880 5780 13889
rect 5644 12872 5684 12881
rect 5644 12116 5684 12832
rect 5644 12067 5684 12076
rect 5740 11948 5780 13840
rect 5836 12536 5876 16864
rect 5932 16568 5972 16948
rect 5932 16519 5972 16528
rect 6028 15896 6068 19636
rect 5932 15856 6068 15896
rect 5932 14636 5972 15856
rect 6028 15476 6068 15485
rect 6028 14804 6068 15436
rect 6028 14755 6068 14764
rect 5932 14587 5972 14596
rect 5836 12487 5876 12496
rect 6028 13544 6068 13553
rect 5740 11899 5780 11908
rect 5932 11864 5972 11873
rect 5548 10723 5588 10732
rect 5644 11780 5684 11789
rect 5548 10100 5588 10109
rect 5548 4136 5588 10060
rect 5644 7412 5684 11740
rect 5740 11780 5780 11789
rect 5740 11192 5780 11740
rect 5740 11143 5780 11152
rect 5740 10940 5780 10949
rect 5740 9764 5780 10900
rect 5932 10352 5972 11824
rect 5932 10303 5972 10312
rect 5740 9715 5780 9724
rect 5836 10268 5876 10277
rect 5836 9680 5876 10228
rect 6028 10268 6068 13504
rect 6124 12620 6164 20056
rect 6220 18164 6260 22660
rect 6220 18115 6260 18124
rect 6220 17996 6260 18005
rect 6220 17072 6260 17956
rect 6316 17828 6356 37948
rect 6412 32696 6452 44164
rect 6796 43784 6836 44248
rect 7276 44288 7316 44297
rect 6796 43735 6836 43744
rect 7180 44120 7220 44129
rect 7180 43280 7220 44080
rect 7276 43616 7316 44248
rect 7660 44288 7700 44297
rect 7660 43700 7700 44248
rect 7852 44036 7892 44836
rect 7948 44827 7988 44836
rect 7852 43987 7892 43996
rect 7948 44372 7988 44381
rect 7660 43651 7700 43660
rect 7276 43567 7316 43576
rect 7564 43616 7604 43625
rect 7180 43231 7220 43240
rect 7084 43196 7124 43205
rect 6988 42776 7028 42785
rect 6604 42692 6644 42701
rect 6508 42608 6548 42617
rect 6508 42524 6548 42568
rect 6508 42473 6548 42484
rect 6604 40340 6644 42652
rect 6700 42608 6740 42617
rect 6740 42568 6932 42608
rect 6700 42559 6740 42568
rect 6892 42524 6932 42568
rect 6892 42475 6932 42484
rect 6892 41012 6932 41021
rect 6604 40300 6740 40340
rect 6508 39500 6548 39509
rect 6508 35132 6548 39460
rect 6700 36056 6740 40300
rect 6892 39500 6932 40972
rect 6700 36007 6740 36016
rect 6796 39164 6836 39173
rect 6700 35888 6740 35897
rect 6700 35384 6740 35848
rect 6700 35335 6740 35344
rect 6796 35216 6836 39124
rect 6892 37652 6932 39460
rect 6892 37603 6932 37612
rect 6508 35083 6548 35092
rect 6700 35176 6836 35216
rect 6892 36224 6932 36233
rect 6412 32647 6452 32656
rect 6508 32864 6548 32873
rect 6412 32528 6452 32537
rect 6412 29840 6452 32488
rect 6412 29168 6452 29800
rect 6412 28244 6452 29128
rect 6412 28195 6452 28204
rect 6508 27068 6548 32824
rect 6604 31184 6644 31193
rect 6604 29924 6644 31144
rect 6604 29252 6644 29884
rect 6604 29203 6644 29212
rect 6604 28328 6644 28337
rect 6604 28193 6644 28288
rect 6700 28076 6740 35176
rect 6892 35132 6932 36184
rect 6796 35092 6932 35132
rect 6796 33620 6836 35092
rect 6796 33452 6836 33580
rect 6796 33403 6836 33412
rect 6892 34208 6932 34217
rect 6796 33284 6836 33293
rect 6796 33116 6836 33244
rect 6796 33067 6836 33076
rect 6796 32780 6836 32789
rect 6796 30596 6836 32740
rect 6892 32192 6932 34168
rect 6892 32143 6932 32152
rect 6796 30547 6836 30556
rect 6892 32024 6932 32033
rect 6796 28916 6836 28925
rect 6796 28781 6836 28876
rect 6892 28580 6932 31984
rect 6988 31772 7028 42736
rect 7084 40676 7124 43156
rect 7372 43028 7412 43037
rect 7276 42524 7316 42533
rect 7084 40627 7124 40636
rect 7180 42104 7220 42113
rect 7084 38156 7124 38165
rect 7084 37316 7124 38116
rect 7084 37267 7124 37276
rect 7180 36728 7220 42064
rect 7084 36688 7220 36728
rect 7276 39500 7316 42484
rect 7084 35636 7124 36688
rect 7180 36560 7220 36569
rect 7180 35804 7220 36520
rect 7180 35755 7220 35764
rect 7084 35596 7220 35636
rect 7084 35048 7124 35057
rect 7084 34460 7124 35008
rect 7084 34411 7124 34420
rect 7084 34292 7124 34301
rect 7084 32528 7124 34252
rect 7180 33704 7220 35596
rect 7180 33655 7220 33664
rect 7084 32479 7124 32488
rect 7180 33536 7220 33545
rect 6988 31723 7028 31732
rect 7084 32192 7124 32201
rect 7084 31604 7124 32152
rect 6412 27028 6508 27068
rect 6412 24548 6452 27028
rect 6508 27019 6548 27028
rect 6604 28036 6740 28076
rect 6796 28496 6836 28505
rect 6412 24499 6452 24508
rect 6508 25976 6548 25985
rect 6412 24296 6452 24305
rect 6412 23120 6452 24256
rect 6412 19676 6452 23080
rect 6508 22952 6548 25936
rect 6508 22903 6548 22912
rect 6412 19627 6452 19636
rect 6508 22784 6548 22793
rect 6508 20684 6548 22744
rect 6604 22364 6644 28036
rect 6700 27908 6740 27917
rect 6700 27320 6740 27868
rect 6700 26144 6740 27280
rect 6700 25556 6740 26104
rect 6700 25507 6740 25516
rect 6796 26228 6836 28456
rect 6796 24296 6836 26188
rect 6892 25808 6932 28540
rect 6988 31564 7124 31604
rect 6988 26228 7028 31564
rect 7084 31436 7124 31445
rect 7084 28580 7124 31396
rect 7180 30764 7220 33496
rect 7276 33284 7316 39460
rect 7372 36728 7412 42988
rect 7468 42860 7508 42869
rect 7468 39416 7508 42820
rect 7564 42608 7604 43576
rect 7564 39500 7604 42568
rect 7852 42692 7892 42701
rect 7852 42608 7892 42652
rect 7852 42557 7892 42568
rect 7948 42188 7988 44332
rect 8044 44120 8084 44920
rect 9580 44960 9620 44969
rect 9580 44456 9620 44920
rect 9580 44407 9620 44416
rect 9964 44960 10004 44969
rect 9964 44372 10004 44920
rect 10252 44456 10292 46264
rect 11020 45296 11060 45305
rect 10252 44407 10292 44416
rect 10348 44960 10388 44969
rect 9964 44323 10004 44332
rect 9004 44288 9044 44297
rect 8044 44071 8084 44080
rect 8236 44120 8276 44129
rect 8140 44036 8180 44045
rect 8140 43616 8180 43996
rect 8140 43567 8180 43576
rect 7948 42139 7988 42148
rect 8236 43448 8276 44080
rect 8236 42776 8276 43408
rect 9004 43700 9044 44248
rect 7756 41936 7796 41945
rect 7660 41896 7756 41936
rect 7660 41180 7700 41896
rect 7756 41887 7796 41896
rect 7660 40424 7700 41140
rect 7660 40375 7700 40384
rect 7852 41852 7892 41861
rect 7852 39668 7892 41812
rect 7852 39619 7892 39628
rect 7948 40508 7988 40517
rect 7948 40256 7988 40468
rect 7564 39460 7892 39500
rect 7468 39376 7796 39416
rect 7372 36679 7412 36688
rect 7468 39080 7508 39089
rect 7372 36560 7412 36569
rect 7372 34544 7412 36520
rect 7468 34628 7508 39040
rect 7660 38912 7700 38921
rect 7468 34579 7508 34588
rect 7564 38744 7604 38753
rect 7372 34495 7412 34504
rect 7564 34460 7604 38704
rect 7564 34411 7604 34420
rect 7660 37568 7700 38872
rect 7756 38240 7796 39376
rect 7756 38191 7796 38200
rect 7660 35132 7700 37528
rect 7756 37484 7796 37493
rect 7756 36476 7796 37444
rect 7756 36427 7796 36436
rect 7852 35804 7892 39460
rect 7948 39248 7988 40216
rect 7948 39199 7988 39208
rect 8044 39836 8084 39845
rect 7948 37484 7988 37493
rect 7948 37349 7988 37444
rect 8044 36476 8084 39796
rect 8140 39668 8180 39677
rect 8140 39533 8180 39628
rect 8140 38576 8180 38585
rect 8140 36644 8180 38536
rect 8140 36595 8180 36604
rect 8044 36436 8180 36476
rect 7852 35764 8084 35804
rect 7948 35636 7988 35645
rect 7756 35132 7796 35141
rect 7660 35092 7756 35132
rect 7660 34292 7700 35092
rect 7756 35083 7796 35092
rect 7852 34964 7892 34973
rect 7756 34880 7796 34889
rect 7756 34376 7796 34840
rect 7756 34327 7796 34336
rect 7276 33235 7316 33244
rect 7372 34252 7700 34292
rect 7180 30715 7220 30724
rect 7276 31688 7316 31697
rect 7276 31520 7316 31648
rect 7084 28531 7124 28540
rect 7180 30596 7220 30605
rect 7180 28496 7220 30556
rect 7276 28748 7316 31480
rect 7372 30512 7412 34252
rect 7756 33704 7796 33713
rect 7372 30463 7412 30472
rect 7468 33452 7508 33461
rect 7276 28699 7316 28708
rect 7372 29924 7412 29933
rect 7180 28447 7220 28456
rect 7276 28580 7316 28589
rect 7180 28328 7220 28337
rect 7180 27572 7220 28288
rect 6988 26179 7028 26188
rect 7084 27320 7124 27329
rect 7084 26900 7124 27280
rect 7180 27152 7220 27532
rect 7180 27103 7220 27112
rect 6892 25759 6932 25768
rect 6796 24247 6836 24256
rect 6892 25556 6932 25565
rect 6796 24128 6836 24137
rect 6700 24044 6740 24053
rect 6700 22868 6740 24004
rect 6700 22819 6740 22828
rect 6604 22315 6644 22324
rect 6508 19844 6548 20644
rect 6316 17779 6356 17788
rect 6412 18248 6452 18257
rect 6220 17023 6260 17032
rect 6316 17156 6356 17165
rect 6220 16820 6260 16829
rect 6220 14888 6260 16780
rect 6220 14839 6260 14848
rect 6124 11780 6164 12580
rect 6124 11731 6164 11740
rect 6220 14468 6260 14477
rect 6124 11192 6164 11201
rect 6124 10268 6164 11152
rect 6220 11024 6260 14428
rect 6316 14132 6356 17116
rect 6316 14083 6356 14092
rect 6412 12980 6452 18208
rect 6220 10975 6260 10984
rect 6316 12940 6452 12980
rect 6124 10228 6260 10268
rect 6028 10219 6068 10228
rect 5836 9631 5876 9640
rect 6124 10100 6164 10109
rect 5644 7363 5684 7372
rect 5740 9428 5780 9437
rect 5644 7244 5684 7253
rect 5644 6236 5684 7204
rect 5740 7244 5780 9388
rect 5740 7195 5780 7204
rect 5740 6992 5780 7001
rect 5740 6404 5780 6952
rect 5740 6355 5780 6364
rect 6028 6992 6068 7001
rect 5836 6236 5876 6245
rect 5644 6196 5780 6236
rect 5644 5648 5684 5657
rect 5644 5312 5684 5608
rect 5644 5263 5684 5272
rect 5548 4087 5588 4096
rect 5740 3548 5780 6196
rect 5836 5648 5876 6196
rect 5836 5599 5876 5608
rect 5932 4892 5972 4901
rect 5932 4304 5972 4852
rect 5932 4255 5972 4264
rect 5740 3499 5780 3508
rect 5548 3464 5588 3473
rect 5548 1868 5588 3424
rect 5548 1819 5588 1828
rect 5740 2876 5780 2885
rect 5740 1616 5780 2836
rect 6028 2120 6068 6952
rect 6124 2204 6164 10060
rect 6220 6656 6260 10228
rect 6220 6607 6260 6616
rect 6220 6404 6260 6413
rect 6220 4472 6260 6364
rect 6220 4220 6260 4432
rect 6220 4171 6260 4180
rect 6124 2155 6164 2164
rect 6028 2071 6068 2080
rect 5740 1567 5780 1576
rect 6316 188 6356 12940
rect 6412 12284 6452 12293
rect 6412 10856 6452 12244
rect 6508 11192 6548 19804
rect 6604 21524 6644 21533
rect 6604 20852 6644 21484
rect 6700 21020 6740 21029
rect 6700 20885 6740 20980
rect 6604 18500 6644 20812
rect 6700 20348 6740 20357
rect 6700 18668 6740 20308
rect 6700 18619 6740 18628
rect 6604 18451 6644 18460
rect 6604 18332 6644 18341
rect 6604 17912 6644 18292
rect 6796 18248 6836 24088
rect 6796 18199 6836 18208
rect 6796 18080 6836 18089
rect 6604 17863 6644 17872
rect 6700 17996 6740 18005
rect 6508 11143 6548 11152
rect 6604 17744 6644 17753
rect 6412 10807 6452 10816
rect 6508 10940 6548 10949
rect 6508 9428 6548 10900
rect 6508 8756 6548 9388
rect 6508 8707 6548 8716
rect 6412 8000 6452 8009
rect 6412 5564 6452 7960
rect 6412 5515 6452 5524
rect 5836 148 6356 188
rect 6412 5396 6452 5405
rect 5836 80 5876 148
rect 6412 104 6452 5356
rect 6508 2876 6548 2887
rect 6508 2792 6548 2836
rect 6508 2743 6548 2752
rect 6220 80 6452 104
rect 6604 80 6644 17704
rect 6700 11864 6740 17956
rect 6796 17408 6836 18040
rect 6796 17359 6836 17368
rect 6700 11815 6740 11824
rect 6796 17240 6836 17249
rect 6700 11360 6740 11369
rect 6700 10184 6740 11320
rect 6700 10135 6740 10144
rect 6700 5900 6740 5909
rect 6700 5765 6740 5860
rect 6700 5564 6740 5573
rect 6700 4388 6740 5524
rect 6700 4339 6740 4348
rect 6796 188 6836 17200
rect 6892 14468 6932 25516
rect 7084 24632 7124 26860
rect 7084 24583 7124 24592
rect 7180 26732 7220 26741
rect 7180 24884 7220 26692
rect 7276 25976 7316 28540
rect 7276 25927 7316 25936
rect 7372 26900 7412 29884
rect 7468 29168 7508 33412
rect 7756 31604 7796 33664
rect 7852 33620 7892 34924
rect 7852 33571 7892 33580
rect 7564 31268 7604 31277
rect 7564 31133 7604 31228
rect 7468 29119 7508 29128
rect 7564 30596 7604 30605
rect 6988 24464 7028 24473
rect 6988 17996 7028 24424
rect 7180 24464 7220 24844
rect 7180 24415 7220 24424
rect 7276 25724 7316 25733
rect 7276 24380 7316 25684
rect 7372 25220 7412 26860
rect 7468 29000 7508 29009
rect 7468 26144 7508 28960
rect 7468 26095 7508 26104
rect 7564 26144 7604 30556
rect 7660 30428 7700 30437
rect 7660 29924 7700 30388
rect 7660 29875 7700 29884
rect 7660 28580 7700 28589
rect 7660 26564 7700 28540
rect 7756 27656 7796 31564
rect 7852 33368 7892 33377
rect 7852 31604 7892 33328
rect 7852 28496 7892 31564
rect 7852 28447 7892 28456
rect 7756 27607 7796 27616
rect 7852 28328 7892 28337
rect 7660 26524 7796 26564
rect 7372 24548 7412 25180
rect 7372 24499 7412 24508
rect 7468 25976 7508 25985
rect 7276 24340 7412 24380
rect 7276 23036 7316 23045
rect 7180 22952 7220 22961
rect 6988 17947 7028 17956
rect 7084 22364 7124 22373
rect 7084 20012 7124 22324
rect 7084 18584 7124 19972
rect 6892 14419 6932 14428
rect 6988 17828 7028 17837
rect 6892 14300 6932 14309
rect 6892 5396 6932 14260
rect 6988 12980 7028 17788
rect 7084 17072 7124 18544
rect 7084 17023 7124 17032
rect 7180 16988 7220 22912
rect 7276 20348 7316 22996
rect 7276 20299 7316 20308
rect 7276 20180 7316 20189
rect 7276 19172 7316 20140
rect 7276 17912 7316 19132
rect 7276 17863 7316 17872
rect 7180 16853 7220 16948
rect 7276 17576 7316 17585
rect 7084 16316 7124 16325
rect 7084 14300 7124 16276
rect 7084 14251 7124 14260
rect 7180 15644 7220 15653
rect 7180 14216 7220 15604
rect 7180 14167 7220 14176
rect 7180 13964 7220 13973
rect 7180 13208 7220 13924
rect 7180 13159 7220 13168
rect 6988 12940 7220 12980
rect 7084 12788 7124 12797
rect 6988 10352 7028 10361
rect 6988 9428 7028 10312
rect 6988 9379 7028 9388
rect 6892 5347 6932 5356
rect 6988 8756 7028 8765
rect 6988 3464 7028 8716
rect 7084 5564 7124 12748
rect 7180 8756 7220 12940
rect 7180 8707 7220 8716
rect 7180 8588 7220 8597
rect 7180 7244 7220 8548
rect 7276 8000 7316 17536
rect 7276 7951 7316 7960
rect 7180 7195 7220 7204
rect 7276 6320 7316 6329
rect 7180 5984 7220 5993
rect 7180 5732 7220 5944
rect 7180 5683 7220 5692
rect 7276 5648 7316 6280
rect 7276 5599 7316 5608
rect 7084 5515 7124 5524
rect 6988 3415 7028 3424
rect 7372 2900 7412 24340
rect 7468 23960 7508 25936
rect 7468 23708 7508 23920
rect 7468 23659 7508 23668
rect 7564 25304 7604 26104
rect 7564 23540 7604 25264
rect 7468 23500 7604 23540
rect 7660 26396 7700 26405
rect 7468 23036 7508 23500
rect 7468 22987 7508 22996
rect 7564 23120 7604 23129
rect 7468 22784 7508 22793
rect 7468 22364 7508 22744
rect 7564 22532 7604 23080
rect 7564 22483 7604 22492
rect 7468 22324 7604 22364
rect 7564 22196 7604 22324
rect 7468 19256 7508 19265
rect 7468 19121 7508 19216
rect 7468 19004 7508 19013
rect 7468 18500 7508 18964
rect 7468 18451 7508 18460
rect 7468 18332 7508 18341
rect 7468 17744 7508 18292
rect 7468 17695 7508 17704
rect 7468 17408 7508 17417
rect 7468 16736 7508 17368
rect 7468 16687 7508 16696
rect 7564 16484 7604 22156
rect 7660 19340 7700 26356
rect 7756 25808 7796 26524
rect 7756 25759 7796 25768
rect 7852 24716 7892 28288
rect 7948 27740 7988 35596
rect 8044 30764 8084 35764
rect 8140 35216 8180 36436
rect 8140 35132 8180 35176
rect 8140 35052 8180 35092
rect 8044 30715 8084 30724
rect 8140 34544 8180 34553
rect 8140 33536 8180 34504
rect 8236 33704 8276 42736
rect 8716 43364 8756 43373
rect 8428 42608 8468 42617
rect 8428 42188 8468 42568
rect 8428 42139 8468 42148
rect 8716 42188 8756 43324
rect 9004 43220 9044 43660
rect 9388 44288 9428 44297
rect 9388 43700 9428 44248
rect 9196 43448 9236 43457
rect 9004 43180 9140 43220
rect 8716 42139 8756 42148
rect 8812 42524 8852 42533
rect 8620 40508 8660 40517
rect 8524 40424 8564 40433
rect 8236 33655 8276 33664
rect 8332 40340 8372 40349
rect 8332 33536 8372 40300
rect 8428 39752 8468 39761
rect 8428 39617 8468 39712
rect 8428 38912 8468 38921
rect 8428 38408 8468 38872
rect 8428 38359 8468 38368
rect 8524 38828 8564 40384
rect 8620 39668 8660 40468
rect 8620 38996 8660 39628
rect 8716 38996 8756 39005
rect 8620 38956 8716 38996
rect 8428 38240 8468 38249
rect 8428 35636 8468 38200
rect 8524 36980 8564 38788
rect 8620 38744 8660 38753
rect 8620 38156 8660 38704
rect 8716 38576 8756 38956
rect 8716 38527 8756 38536
rect 8620 38107 8660 38116
rect 8812 37988 8852 42484
rect 9100 42104 9140 43180
rect 9196 42608 9236 43408
rect 9388 42692 9428 43660
rect 10252 44288 10292 44297
rect 9388 42643 9428 42652
rect 9868 43112 9908 43121
rect 9196 42559 9236 42568
rect 9100 42055 9140 42064
rect 9388 42272 9428 42281
rect 9292 42020 9332 42029
rect 9100 41852 9140 41861
rect 8524 36931 8564 36940
rect 8620 37948 8852 37988
rect 8908 40508 8948 40517
rect 8908 40256 8948 40468
rect 8908 39668 8948 40216
rect 8908 38996 8948 39628
rect 8428 35587 8468 35596
rect 8524 35972 8564 35981
rect 8524 35048 8564 35932
rect 8524 34999 8564 35008
rect 7948 27691 7988 27700
rect 8044 30596 8084 30605
rect 7948 27572 7988 27581
rect 7948 25892 7988 27532
rect 7948 25757 7988 25852
rect 7756 24676 7892 24716
rect 7948 25304 7988 25313
rect 7756 23960 7796 24676
rect 7852 24548 7892 24557
rect 7852 24044 7892 24508
rect 7852 23995 7892 24004
rect 7756 23624 7796 23920
rect 7948 23876 7988 25264
rect 7756 23575 7796 23584
rect 7852 23836 7988 23876
rect 7660 18584 7700 19300
rect 7660 18535 7700 18544
rect 7756 23456 7796 23465
rect 7564 16435 7604 16444
rect 7660 17912 7700 17921
rect 7564 16316 7604 16325
rect 7468 16232 7508 16241
rect 7468 15476 7508 16192
rect 7564 15728 7604 16276
rect 7564 15679 7604 15688
rect 7468 14048 7508 15436
rect 7468 13999 7508 14008
rect 7564 14804 7604 14813
rect 7564 13124 7604 14764
rect 7660 13544 7700 17872
rect 7756 16400 7796 23416
rect 7852 23036 7892 23836
rect 8044 23792 8084 30556
rect 8140 28160 8180 33496
rect 8236 33496 8372 33536
rect 8428 34124 8468 34133
rect 8236 32864 8276 33496
rect 8332 33032 8372 33043
rect 8332 32948 8372 32992
rect 8332 32899 8372 32908
rect 8236 32192 8276 32824
rect 8236 32143 8276 32152
rect 8332 32108 8372 32117
rect 8236 31604 8276 31613
rect 8236 31469 8276 31564
rect 8332 31394 8372 32068
rect 8332 31268 8372 31354
rect 8332 31219 8372 31228
rect 8332 30764 8372 30773
rect 8236 29840 8276 29849
rect 8236 29705 8276 29800
rect 8332 29168 8372 30724
rect 8140 28111 8180 28120
rect 8236 29128 8372 29168
rect 8236 28328 8276 29128
rect 8236 27572 8276 28288
rect 8236 27523 8276 27532
rect 8332 29000 8372 29009
rect 8140 27488 8180 27497
rect 8140 26900 8180 27448
rect 8140 26851 8180 26860
rect 8236 27404 8276 27413
rect 7852 22987 7892 22996
rect 7948 23752 8084 23792
rect 8140 24884 8180 24893
rect 7852 22868 7892 22877
rect 7852 21020 7892 22828
rect 7948 22364 7988 23752
rect 8044 23624 8084 23633
rect 8044 22784 8084 23584
rect 8044 22735 8084 22744
rect 8044 22532 8084 22627
rect 8044 22483 8084 22492
rect 8044 22364 8084 22373
rect 7948 22324 8044 22364
rect 7852 18584 7892 20980
rect 8044 21524 8084 22324
rect 7852 18535 7892 18544
rect 7948 19928 7988 19937
rect 7756 16351 7796 16360
rect 7852 18416 7892 18425
rect 7756 16232 7796 16241
rect 7756 15056 7796 16192
rect 7756 15007 7796 15016
rect 7852 14804 7892 18376
rect 7948 17240 7988 19888
rect 7948 17191 7988 17200
rect 7948 16736 7988 16745
rect 7948 14972 7988 16696
rect 7948 14923 7988 14932
rect 7948 14804 7988 14813
rect 7852 14764 7948 14804
rect 7660 13495 7700 13504
rect 7564 12452 7604 13084
rect 7564 12403 7604 12412
rect 7756 13124 7796 13133
rect 7564 12284 7604 12293
rect 7564 11780 7604 12244
rect 7468 10940 7508 10949
rect 7468 9428 7508 10900
rect 7468 8924 7508 9388
rect 7564 9428 7604 11740
rect 7660 11528 7700 11537
rect 7660 10940 7700 11488
rect 7660 10891 7700 10900
rect 7564 9379 7604 9388
rect 7468 8875 7508 8884
rect 7756 8084 7796 13084
rect 7852 11948 7892 11957
rect 7852 11813 7892 11908
rect 7756 8044 7892 8084
rect 7660 8000 7700 8009
rect 7564 7076 7604 7085
rect 7564 6404 7604 7036
rect 7564 6355 7604 6364
rect 7660 5732 7700 7960
rect 7756 7916 7796 7925
rect 7756 7412 7796 7876
rect 7756 7363 7796 7372
rect 7756 5732 7796 5741
rect 7660 5692 7756 5732
rect 7756 4808 7796 5692
rect 7756 4759 7796 4768
rect 7852 2900 7892 8044
rect 7948 7916 7988 14764
rect 8044 13292 8084 21484
rect 8140 19256 8180 24844
rect 8140 18836 8180 19216
rect 8140 17744 8180 18796
rect 8236 24464 8276 27364
rect 8236 18752 8276 24424
rect 8332 25388 8372 28960
rect 8428 26732 8468 34084
rect 8524 33620 8564 33629
rect 8524 33116 8564 33580
rect 8524 33067 8564 33076
rect 8524 32780 8564 32789
rect 8524 32612 8564 32740
rect 8524 32563 8564 32572
rect 8620 32192 8660 37948
rect 8812 37400 8852 37409
rect 8716 37232 8756 37241
rect 8716 34544 8756 37192
rect 8812 37064 8852 37360
rect 8812 37015 8852 37024
rect 8716 34495 8756 34504
rect 8812 34880 8852 34889
rect 8716 34208 8756 34217
rect 8716 33788 8756 34168
rect 8716 33739 8756 33748
rect 8716 33620 8756 33629
rect 8716 32864 8756 33580
rect 8716 32815 8756 32824
rect 8620 32143 8660 32152
rect 8716 32612 8756 32621
rect 8524 32108 8564 32117
rect 8524 28832 8564 32068
rect 8524 28783 8564 28792
rect 8620 31520 8660 31529
rect 8428 26683 8468 26692
rect 8524 28160 8564 28169
rect 8332 23036 8372 25348
rect 8428 26144 8468 26153
rect 8428 23456 8468 26104
rect 8524 25304 8564 28120
rect 8620 26984 8660 31480
rect 8716 31436 8756 32572
rect 8716 30932 8756 31396
rect 8716 30883 8756 30892
rect 8812 30764 8852 34840
rect 8716 30724 8852 30764
rect 8716 30008 8756 30724
rect 8716 29959 8756 29968
rect 8812 30596 8852 30605
rect 8812 30344 8852 30556
rect 8716 29840 8756 29849
rect 8716 29705 8756 29800
rect 8716 29252 8756 29261
rect 8716 27068 8756 29212
rect 8812 29084 8852 30304
rect 8812 29035 8852 29044
rect 8716 27028 8852 27068
rect 8620 26944 8756 26984
rect 8620 26816 8660 26825
rect 8620 26732 8660 26776
rect 8620 26681 8660 26692
rect 8716 25388 8756 26944
rect 8812 26900 8852 27028
rect 8812 26851 8852 26860
rect 8524 25255 8564 25264
rect 8620 25348 8756 25388
rect 8620 23876 8660 25348
rect 8620 23827 8660 23836
rect 8716 25220 8756 25229
rect 8428 23120 8468 23416
rect 8428 23071 8468 23080
rect 8620 23708 8660 23717
rect 8620 23204 8660 23668
rect 8332 22952 8372 22996
rect 8332 22912 8468 22952
rect 8332 21608 8372 21617
rect 8332 21473 8372 21568
rect 8236 18712 8372 18752
rect 8332 18668 8372 18712
rect 8332 18619 8372 18628
rect 8236 18584 8276 18593
rect 8236 17828 8276 18544
rect 8236 17779 8276 17788
rect 8140 17695 8180 17704
rect 8044 13243 8084 13252
rect 8140 17492 8180 17501
rect 7948 7867 7988 7876
rect 8140 2900 8180 17452
rect 8332 16316 8372 16325
rect 8332 14804 8372 16276
rect 8428 16232 8468 22912
rect 8524 20096 8564 20105
rect 8524 18752 8564 20056
rect 8620 19928 8660 23164
rect 8620 19879 8660 19888
rect 8716 19424 8756 25180
rect 8908 25052 8948 38956
rect 9004 37904 9044 37913
rect 9004 37484 9044 37864
rect 9004 35972 9044 37444
rect 9004 35923 9044 35932
rect 9004 33704 9044 33713
rect 9004 32948 9044 33664
rect 9100 33032 9140 41812
rect 9196 41768 9236 41777
rect 9196 37568 9236 41728
rect 9292 41180 9332 41980
rect 9292 38744 9332 41140
rect 9292 38240 9332 38704
rect 9292 38191 9332 38200
rect 9196 37528 9332 37568
rect 9100 32983 9140 32992
rect 9196 35468 9236 35477
rect 9004 31436 9044 32908
rect 9100 32864 9140 32873
rect 9100 32108 9140 32824
rect 9100 32059 9140 32068
rect 9004 31387 9044 31396
rect 9100 31940 9140 31949
rect 9004 30008 9044 30017
rect 9004 29252 9044 29968
rect 9004 29203 9044 29212
rect 9100 28412 9140 31900
rect 9196 29168 9236 35428
rect 9292 32948 9332 37528
rect 9388 34880 9428 42232
rect 9484 41012 9524 41021
rect 9484 39668 9524 40972
rect 9484 39619 9524 39628
rect 9868 39752 9908 43072
rect 9964 42776 10004 42785
rect 9964 42641 10004 42736
rect 9964 42524 10004 42533
rect 9964 42020 10004 42484
rect 9964 41971 10004 41980
rect 10060 42104 10100 42113
rect 9964 41264 10004 41273
rect 9964 40424 10004 41224
rect 9964 40289 10004 40384
rect 10060 41012 10100 42064
rect 10060 40340 10100 40972
rect 10060 40291 10100 40300
rect 9772 38996 9812 39005
rect 9772 38408 9812 38956
rect 9772 38359 9812 38368
rect 9868 38156 9908 39712
rect 9868 37484 9908 38116
rect 9772 37444 9868 37484
rect 9580 37316 9620 37325
rect 9484 36476 9524 36485
rect 9484 36341 9524 36436
rect 9388 34831 9428 34840
rect 9484 36056 9524 36065
rect 9292 32899 9332 32908
rect 9388 34460 9428 34469
rect 9484 34460 9524 36016
rect 9428 34420 9524 34460
rect 9196 29119 9236 29128
rect 9292 32780 9332 32789
rect 9292 31352 9332 32740
rect 9292 29000 9332 31312
rect 8716 19375 8756 19384
rect 8812 25012 8948 25052
rect 9004 28372 9140 28412
rect 9196 28960 9332 29000
rect 8524 18703 8564 18712
rect 8716 19256 8756 19265
rect 8428 16183 8468 16192
rect 8524 18584 8564 18593
rect 8332 14755 8372 14764
rect 8428 14972 8468 14981
rect 8428 13964 8468 14932
rect 8428 13915 8468 13924
rect 8428 11948 8468 11957
rect 8332 9428 8372 9437
rect 8332 8756 8372 9388
rect 8236 8716 8332 8756
rect 8236 4892 8276 8716
rect 8332 8707 8372 8716
rect 8332 8084 8372 8093
rect 8332 7160 8372 8044
rect 8428 8000 8468 11908
rect 8428 7951 8468 7960
rect 8332 7111 8372 7120
rect 8332 5732 8372 5741
rect 8332 5144 8372 5692
rect 8332 5095 8372 5104
rect 8236 4220 8276 4852
rect 8236 4171 8276 4180
rect 7372 2860 7604 2900
rect 7564 2372 7604 2860
rect 7756 2860 7892 2900
rect 7948 2860 8180 2900
rect 7756 2540 7796 2860
rect 7756 2491 7796 2500
rect 7564 2332 7796 2372
rect 7372 1448 7412 1457
rect 6796 148 7124 188
rect 7084 104 7124 148
rect 6988 80 7124 104
rect 7372 80 7412 1408
rect 7756 80 7796 2332
rect 7948 1448 7988 2860
rect 7948 1399 7988 1408
rect 8140 1448 8180 1457
rect 8140 80 8180 1408
rect 8524 80 8564 18544
rect 8716 18500 8756 19216
rect 8716 18451 8756 18460
rect 8812 17828 8852 25012
rect 9004 24044 9044 28372
rect 9100 28244 9140 28253
rect 9100 28109 9140 28204
rect 9004 23995 9044 24004
rect 9100 26900 9140 26909
rect 9100 26144 9140 26860
rect 9004 23036 9044 23045
rect 8908 21440 8948 21449
rect 8908 20852 8948 21400
rect 8908 20803 8948 20812
rect 8908 20684 8948 20693
rect 8908 20549 8948 20644
rect 8812 17779 8852 17788
rect 8908 19424 8948 19433
rect 8812 17660 8852 17669
rect 8812 16988 8852 17620
rect 8812 16939 8852 16948
rect 8620 16400 8660 16409
rect 8620 15560 8660 16360
rect 8620 15511 8660 15520
rect 8812 16316 8852 16325
rect 8812 14720 8852 16276
rect 8812 14671 8852 14680
rect 8908 14804 8948 19384
rect 9004 16316 9044 22996
rect 9100 20936 9140 26104
rect 9196 23036 9236 28960
rect 9196 22987 9236 22996
rect 9292 28412 9332 28421
rect 9388 28412 9428 34420
rect 9332 28372 9428 28412
rect 9484 32948 9524 32957
rect 9484 30344 9524 32908
rect 9580 32192 9620 37276
rect 9580 32143 9620 32152
rect 9676 34292 9716 34301
rect 9484 29924 9524 30304
rect 9580 32024 9620 32033
rect 9580 31436 9620 31984
rect 9580 30176 9620 31396
rect 9580 30127 9620 30136
rect 9100 20012 9140 20896
rect 9100 19963 9140 19972
rect 9004 16267 9044 16276
rect 9100 19256 9140 19265
rect 8620 14552 8660 14561
rect 8620 13880 8660 14512
rect 8620 13831 8660 13840
rect 8812 13376 8852 13404
rect 8908 13376 8948 14764
rect 8852 13336 8948 13376
rect 8812 13327 8852 13336
rect 8908 12980 8948 13336
rect 8812 12940 8948 12980
rect 9004 15308 9044 15317
rect 8620 11780 8660 11789
rect 8620 10940 8660 11740
rect 8620 10891 8660 10900
rect 8812 11612 8852 12940
rect 8908 12620 8948 12629
rect 8908 11696 8948 12580
rect 8908 11647 8948 11656
rect 8716 10856 8756 10865
rect 8620 10184 8660 10193
rect 8620 9680 8660 10144
rect 8620 9631 8660 9640
rect 8716 9512 8756 10816
rect 8620 9472 8756 9512
rect 8620 7748 8660 9472
rect 8620 7699 8660 7708
rect 8716 8672 8756 8681
rect 8620 7244 8660 7253
rect 8620 5732 8660 7204
rect 8716 7076 8756 8632
rect 8716 7027 8756 7036
rect 8812 6908 8852 11572
rect 8908 10184 8948 10193
rect 8908 8168 8948 10144
rect 8908 8119 8948 8128
rect 8620 5060 8660 5692
rect 8620 5011 8660 5020
rect 8716 6868 8852 6908
rect 8716 2120 8756 6868
rect 8812 5732 8852 5741
rect 8812 5597 8852 5692
rect 9004 5312 9044 15268
rect 9100 13628 9140 19216
rect 9292 17996 9332 28372
rect 9484 26060 9524 29884
rect 9676 29084 9716 34252
rect 9580 29044 9716 29084
rect 9580 28244 9620 29044
rect 9676 28916 9716 28925
rect 9676 28781 9716 28876
rect 9580 28195 9620 28204
rect 9676 28496 9716 28505
rect 9388 26020 9524 26060
rect 9676 27488 9716 28456
rect 9388 24548 9428 26020
rect 9484 25892 9524 25901
rect 9484 25388 9524 25852
rect 9484 25339 9524 25348
rect 9580 25808 9620 25817
rect 9580 25220 9620 25768
rect 9388 24499 9428 24508
rect 9484 25180 9620 25220
rect 9388 24380 9428 24389
rect 9388 18164 9428 24340
rect 9484 19172 9524 25180
rect 9676 23960 9716 27448
rect 9676 23911 9716 23920
rect 9484 19123 9524 19132
rect 9580 23876 9620 23885
rect 9580 22364 9620 23836
rect 9580 20012 9620 22324
rect 9580 19340 9620 19972
rect 9388 18115 9428 18124
rect 9484 17996 9524 18005
rect 9292 17956 9428 17996
rect 9292 17828 9332 17837
rect 9100 13579 9140 13588
rect 9196 17744 9236 17753
rect 9100 13208 9140 13217
rect 9100 12704 9140 13168
rect 9100 12655 9140 12664
rect 9196 10856 9236 17704
rect 9292 17240 9332 17788
rect 9292 17191 9332 17200
rect 9292 16988 9332 16997
rect 9292 16736 9332 16948
rect 9388 16904 9428 17956
rect 9484 17072 9524 17956
rect 9484 17023 9524 17032
rect 9388 16864 9524 16904
rect 9292 16687 9332 16696
rect 9388 16316 9428 16325
rect 9388 15728 9428 16276
rect 9388 15679 9428 15688
rect 9388 14804 9428 14813
rect 9388 14216 9428 14764
rect 9388 14167 9428 14176
rect 9484 13796 9524 16864
rect 9580 16316 9620 19300
rect 9676 19844 9716 19853
rect 9676 18500 9716 19804
rect 9676 18451 9716 18460
rect 9676 16988 9716 16997
rect 9676 16568 9716 16948
rect 9676 16519 9716 16528
rect 9676 16316 9716 16325
rect 9580 16276 9676 16316
rect 9580 14048 9620 14057
rect 9580 13913 9620 14008
rect 9484 13756 9620 13796
rect 9484 13628 9524 13637
rect 9292 13292 9332 13301
rect 9292 12452 9332 13252
rect 9332 12412 9428 12452
rect 9292 12403 9332 12412
rect 9196 10807 9236 10816
rect 9292 11024 9332 11033
rect 9292 10100 9332 10984
rect 9292 10051 9332 10060
rect 9388 9512 9428 12412
rect 9388 7244 9428 9472
rect 9388 7195 9428 7204
rect 9004 5263 9044 5272
rect 9484 2900 9524 13588
rect 9580 11192 9620 13756
rect 9676 13712 9716 16276
rect 9676 13663 9716 13672
rect 9580 11143 9620 11152
rect 9676 13544 9716 13553
rect 8716 2071 8756 2080
rect 9292 2860 9524 2900
rect 8908 1448 8948 1457
rect 8908 80 8948 1408
rect 9292 80 9332 2860
rect 9676 80 9716 13504
rect 9772 9428 9812 37444
rect 9868 37435 9908 37444
rect 10156 39500 10196 39509
rect 10060 37064 10100 37073
rect 9964 36728 10004 36737
rect 9964 36593 10004 36688
rect 10060 36140 10100 37024
rect 10060 36091 10100 36100
rect 10060 35972 10100 35981
rect 9964 35132 10004 35141
rect 9868 34964 9908 34973
rect 9868 33620 9908 34924
rect 9868 33571 9908 33580
rect 9964 33368 10004 35092
rect 9868 33328 10004 33368
rect 9868 30596 9908 33328
rect 10060 33140 10100 35932
rect 9868 30547 9908 30556
rect 9964 33100 10100 33140
rect 9868 30428 9908 30437
rect 9868 30293 9908 30388
rect 9868 30176 9908 30185
rect 9868 28328 9908 30136
rect 9964 28412 10004 33100
rect 10060 32864 10100 32873
rect 10060 32729 10100 32824
rect 10156 32192 10196 39460
rect 10252 33200 10292 44248
rect 10348 43532 10388 44920
rect 11020 44456 11060 45256
rect 11020 44407 11060 44416
rect 11692 44792 11732 44801
rect 11692 44288 11732 44752
rect 11692 44239 11732 44248
rect 10348 43483 10388 43492
rect 10828 43784 10868 43793
rect 10540 43448 10580 43457
rect 10348 42776 10388 42785
rect 10348 42641 10388 42736
rect 10348 41936 10388 41945
rect 10348 41801 10388 41896
rect 10348 40424 10388 40433
rect 10348 36812 10388 40384
rect 10444 39500 10484 39509
rect 10444 39365 10484 39460
rect 10444 38912 10484 38921
rect 10444 38777 10484 38872
rect 10348 36772 10484 36812
rect 10252 33151 10292 33160
rect 10348 35216 10388 35225
rect 10156 32143 10196 32152
rect 10252 32108 10292 32117
rect 10156 31436 10196 31445
rect 9964 28363 10004 28372
rect 10060 30260 10100 30269
rect 10060 29924 10100 30220
rect 10156 30092 10196 31396
rect 10156 30043 10196 30052
rect 9868 28279 9908 28288
rect 9868 28076 9908 28085
rect 9868 20096 9908 28036
rect 9964 28076 10004 28085
rect 9964 24380 10004 28036
rect 10060 27572 10100 29884
rect 10252 29252 10292 32068
rect 10348 30848 10388 35176
rect 10348 30799 10388 30808
rect 10060 27523 10100 27532
rect 10156 29212 10292 29252
rect 9964 24331 10004 24340
rect 10060 24548 10100 24557
rect 9964 23960 10004 23969
rect 9964 20180 10004 23920
rect 10060 23876 10100 24508
rect 10060 21524 10100 23836
rect 10060 21475 10100 21484
rect 10060 20180 10100 20189
rect 9964 20140 10060 20180
rect 10060 20131 10100 20140
rect 9908 20056 10004 20096
rect 9868 20047 9908 20056
rect 9868 19508 9908 19517
rect 9868 18500 9908 19468
rect 9868 18451 9908 18460
rect 9964 18332 10004 20056
rect 10156 18752 10196 29212
rect 10348 29168 10388 29177
rect 10252 29084 10292 29093
rect 10252 28580 10292 29044
rect 10348 29033 10388 29128
rect 10252 28531 10292 28540
rect 10348 27404 10388 27413
rect 10348 26900 10388 27364
rect 10252 26860 10348 26900
rect 10252 24548 10292 26860
rect 10348 26851 10388 26860
rect 10252 24499 10292 24508
rect 10348 25388 10388 25397
rect 10252 22616 10292 22625
rect 10252 19508 10292 22576
rect 10348 21776 10388 25348
rect 10348 21727 10388 21736
rect 10348 21608 10388 21617
rect 10348 21440 10388 21568
rect 10348 21391 10388 21400
rect 10252 19468 10388 19508
rect 10156 18703 10196 18712
rect 10252 19340 10292 19349
rect 9868 18292 10004 18332
rect 10060 18584 10100 18593
rect 9868 16988 9908 18292
rect 9868 16939 9908 16948
rect 9964 18164 10004 18173
rect 9868 16820 9908 16829
rect 9868 15812 9908 16780
rect 9868 15763 9908 15772
rect 9964 13880 10004 18124
rect 10060 14048 10100 18544
rect 10156 16484 10196 16493
rect 10156 15560 10196 16444
rect 10156 15511 10196 15520
rect 10060 13999 10100 14008
rect 10252 13964 10292 19300
rect 9964 13840 10100 13880
rect 9964 13712 10004 13721
rect 9964 12620 10004 13672
rect 9964 12571 10004 12580
rect 10060 11948 10100 13840
rect 10252 12452 10292 13924
rect 10348 13796 10388 19468
rect 10348 13747 10388 13756
rect 10252 12403 10292 12412
rect 10348 13376 10388 13385
rect 10060 11899 10100 11908
rect 9772 8756 9812 9388
rect 9772 8707 9812 8716
rect 10156 11612 10196 11621
rect 10060 7748 10100 7757
rect 9964 6488 10004 6497
rect 9964 6353 10004 6448
rect 10060 4304 10100 7708
rect 10060 4255 10100 4264
rect 10156 2900 10196 11572
rect 10252 11024 10292 11033
rect 10252 10436 10292 10984
rect 10252 10387 10292 10396
rect 10348 10184 10388 13336
rect 10444 12980 10484 36772
rect 10540 28076 10580 43408
rect 10540 28027 10580 28036
rect 10636 41264 10676 41273
rect 10540 26648 10580 26657
rect 10540 18584 10580 26608
rect 10636 26312 10676 41224
rect 10732 40256 10772 40265
rect 10732 38240 10772 40216
rect 10732 38191 10772 38200
rect 10828 36140 10868 43744
rect 10924 43280 10964 43289
rect 10924 40256 10964 43240
rect 11692 42608 11732 42617
rect 11212 42524 11252 42533
rect 11116 41936 11156 41945
rect 10924 40207 10964 40216
rect 11020 41096 11060 41105
rect 11020 38240 11060 41056
rect 11020 38191 11060 38200
rect 10732 36100 10828 36140
rect 10732 32360 10772 36100
rect 10828 36091 10868 36100
rect 10924 38156 10964 38165
rect 10924 34628 10964 38116
rect 11116 37232 11156 41896
rect 11212 39248 11252 42484
rect 11692 42272 11732 42568
rect 11692 42223 11732 42232
rect 11212 39199 11252 39208
rect 11404 42020 11444 42029
rect 11116 37183 11156 37192
rect 11308 36728 11348 36737
rect 11020 36560 11060 36569
rect 11020 35216 11060 36520
rect 11020 35167 11060 35176
rect 11116 36476 11156 36485
rect 10828 34588 10924 34628
rect 10828 33116 10868 34588
rect 10924 34579 10964 34588
rect 10924 34376 10964 34385
rect 10924 33200 10964 34336
rect 11116 34208 11156 36436
rect 11116 34159 11156 34168
rect 11212 34964 11252 34973
rect 10924 33151 10964 33160
rect 11116 33452 11156 33461
rect 10828 33067 10868 33076
rect 10732 32311 10772 32320
rect 10828 32948 10868 32957
rect 10828 31688 10868 32908
rect 10828 31639 10868 31648
rect 10924 32864 10964 32873
rect 10828 29672 10868 29681
rect 10828 29168 10868 29632
rect 10828 29119 10868 29128
rect 10924 29000 10964 32824
rect 11020 32024 11060 32033
rect 11020 31184 11060 31984
rect 11020 31135 11060 31144
rect 10924 28951 10964 28960
rect 11020 29084 11060 29093
rect 10924 28664 10964 28673
rect 10924 28160 10964 28624
rect 10924 28111 10964 28120
rect 10636 26263 10676 26272
rect 10732 28076 10772 28085
rect 10636 23120 10676 23129
rect 10636 22532 10676 23080
rect 10636 22483 10676 22492
rect 10732 22448 10772 28036
rect 11020 27908 11060 29044
rect 10924 27868 11060 27908
rect 10732 22399 10772 22408
rect 10828 24548 10868 24557
rect 10732 21776 10772 21785
rect 10636 20852 10676 20861
rect 10636 19340 10676 20812
rect 10636 19291 10676 19300
rect 10540 18535 10580 18544
rect 10636 19088 10676 19097
rect 10540 18332 10580 18341
rect 10540 17324 10580 18292
rect 10636 17996 10676 19048
rect 10732 18248 10772 21736
rect 10732 18199 10772 18208
rect 10636 17947 10676 17956
rect 10732 18080 10772 18089
rect 10540 17275 10580 17284
rect 10636 17828 10676 17837
rect 10636 17156 10676 17788
rect 10732 17240 10772 18040
rect 10732 17191 10772 17200
rect 10540 17116 10676 17156
rect 10540 14300 10580 17116
rect 10732 16064 10772 16073
rect 10540 14251 10580 14260
rect 10636 15056 10676 15065
rect 10636 14216 10676 15016
rect 10732 14972 10772 16024
rect 10732 14923 10772 14932
rect 10636 14167 10676 14176
rect 10540 14132 10580 14143
rect 10540 14048 10580 14092
rect 10540 13999 10580 14008
rect 10444 12940 10772 12980
rect 10636 12032 10676 12041
rect 10636 10436 10676 11992
rect 10636 10387 10676 10396
rect 10348 10135 10388 10144
rect 10444 10100 10484 10109
rect 10348 9428 10388 9437
rect 10348 8756 10388 9388
rect 10252 8672 10292 8681
rect 10252 8000 10292 8632
rect 10252 7951 10292 7960
rect 10348 7832 10388 8716
rect 10444 8840 10484 10060
rect 10444 7916 10484 8800
rect 10636 9008 10676 9017
rect 10444 7867 10484 7876
rect 10540 8504 10580 8513
rect 10348 7783 10388 7792
rect 10540 7160 10580 8464
rect 10540 7111 10580 7120
rect 10636 7076 10676 8968
rect 10636 7027 10676 7036
rect 10732 6236 10772 12940
rect 10828 9428 10868 24508
rect 10924 17996 10964 27868
rect 10924 17947 10964 17956
rect 11020 27740 11060 27749
rect 10828 9379 10868 9388
rect 10924 17324 10964 17333
rect 10732 6187 10772 6196
rect 10924 3380 10964 17284
rect 11020 14720 11060 27700
rect 11020 14671 11060 14680
rect 11116 12788 11156 33412
rect 11212 33200 11252 34924
rect 11212 33151 11252 33160
rect 11212 31940 11252 31949
rect 11212 30176 11252 31900
rect 11212 30127 11252 30136
rect 11212 29000 11252 29009
rect 11212 17996 11252 28960
rect 11308 22616 11348 36688
rect 11404 33116 11444 41980
rect 11692 41852 11732 41861
rect 11692 41264 11732 41812
rect 11692 41215 11732 41224
rect 11500 41012 11540 41021
rect 11500 36224 11540 40972
rect 11500 36175 11540 36184
rect 11692 39920 11732 39929
rect 11404 28580 11444 33076
rect 11500 35972 11540 35981
rect 11500 29084 11540 35932
rect 11500 29035 11540 29044
rect 11596 35384 11636 35393
rect 11404 28531 11444 28540
rect 11500 28916 11540 28925
rect 11404 27740 11444 27749
rect 11404 26984 11444 27700
rect 11500 27152 11540 28876
rect 11500 27103 11540 27112
rect 11404 26944 11540 26984
rect 11404 25976 11444 25985
rect 11404 24128 11444 25936
rect 11404 24079 11444 24088
rect 11500 23060 11540 26944
rect 11596 25304 11636 35344
rect 11692 27740 11732 39880
rect 11692 27691 11732 27700
rect 11692 25976 11732 25985
rect 11732 25936 11828 25976
rect 11692 25927 11732 25936
rect 11596 25255 11636 25264
rect 11308 22567 11348 22576
rect 11404 23020 11540 23060
rect 11692 24716 11732 24725
rect 11404 22448 11444 23020
rect 11308 22408 11444 22448
rect 11596 22868 11636 22877
rect 11308 20852 11348 22408
rect 11308 20803 11348 20812
rect 11404 22280 11444 22289
rect 11212 17947 11252 17956
rect 11212 17072 11252 17081
rect 11212 15728 11252 17032
rect 11212 15679 11252 15688
rect 11116 12739 11156 12748
rect 11404 11444 11444 22240
rect 11404 11395 11444 11404
rect 11500 17996 11540 18005
rect 11500 11360 11540 17956
rect 11500 11311 11540 11320
rect 11596 3632 11636 22828
rect 11692 10268 11732 24676
rect 11788 12872 11828 25936
rect 11788 12823 11828 12832
rect 11692 10219 11732 10228
rect 11692 6320 11732 6329
rect 11692 5984 11732 6280
rect 11692 5935 11732 5944
rect 11692 5480 11732 5489
rect 11692 4976 11732 5440
rect 11692 4927 11732 4936
rect 11596 3583 11636 3592
rect 10924 3331 10964 3340
rect 11692 3212 11732 3221
rect 11692 2960 11732 3172
rect 11692 2911 11732 2920
rect 10156 2860 10292 2900
rect 10252 2624 10292 2860
rect 10252 2575 10292 2584
rect 11692 2456 11732 2465
rect 11692 1952 11732 2416
rect 11692 1903 11732 1912
rect 10444 1868 10484 1877
rect 10444 944 10484 1828
rect 10444 895 10484 904
rect 1976 0 2056 80
rect 2360 0 2440 80
rect 2744 0 2824 80
rect 3128 0 3208 80
rect 3512 0 3592 80
rect 3896 0 3976 80
rect 4280 0 4360 80
rect 4664 0 4744 80
rect 5048 0 5128 80
rect 5432 0 5512 80
rect 5816 0 5896 80
rect 6200 64 6452 80
rect 6200 0 6280 64
rect 6584 0 6664 80
rect 6968 64 7124 80
rect 6968 0 7048 64
rect 7352 0 7432 80
rect 7736 0 7816 80
rect 8120 0 8200 80
rect 8504 0 8584 80
rect 8888 0 8968 80
rect 9272 0 9352 80
rect 9656 0 9736 80
<< via3 >>
rect 1996 45172 2036 45212
rect 76 44248 116 44288
rect 364 38116 404 38156
rect 76 34168 116 34208
rect 460 24340 500 24380
rect 76 22408 116 22448
rect 172 22240 212 22280
rect 844 31984 884 32024
rect 844 24340 884 24380
rect 556 22240 596 22280
rect 1036 34504 1076 34544
rect 1612 40972 1652 41012
rect 1516 37192 1556 37232
rect 1132 33496 1172 33536
rect 1036 31480 1076 31520
rect 1132 31984 1172 32024
rect 1420 33496 1460 33536
rect 1516 33664 1556 33704
rect 1996 34588 2036 34628
rect 2764 44920 2804 44960
rect 2476 42652 2516 42692
rect 3148 43324 3188 43364
rect 3244 42988 3284 43028
rect 2956 42568 2996 42608
rect 3148 42148 3188 42188
rect 3052 41812 3092 41852
rect 2956 39712 2996 39752
rect 2860 39460 2900 39500
rect 2284 37444 2324 37484
rect 2284 35428 2324 35468
rect 2092 33916 2132 33956
rect 1708 33076 1748 33116
rect 1612 32824 1652 32864
rect 1900 32992 1940 33032
rect 1228 30976 1268 31016
rect 1420 31228 1460 31268
rect 1516 30892 1556 30932
rect 1420 29968 1460 30008
rect 1324 29800 1364 29840
rect 1420 27532 1460 27572
rect 940 19384 980 19424
rect 1132 20140 1172 20180
rect 1228 19300 1268 19340
rect 1516 20056 1556 20096
rect 1516 18628 1556 18668
rect 940 14512 980 14552
rect 1132 15016 1172 15056
rect 1228 14512 1268 14552
rect 1228 12412 1268 12452
rect 1420 11236 1460 11276
rect 1420 9472 1460 9512
rect 1324 7204 1364 7244
rect 1708 30220 1748 30260
rect 1804 32740 1844 32780
rect 1708 29884 1748 29924
rect 1708 27448 1748 27488
rect 1708 27280 1748 27320
rect 2188 35176 2228 35216
rect 2092 31564 2132 31604
rect 1996 30220 2036 30260
rect 1804 24676 1844 24716
rect 1708 22744 1748 22784
rect 1900 23080 1940 23120
rect 2668 36772 2708 36812
rect 2476 36604 2516 36644
rect 2476 34924 2516 34964
rect 2572 35428 2612 35468
rect 2284 31564 2324 31604
rect 2380 33160 2420 33200
rect 1612 16612 1652 16652
rect 1804 19804 1844 19844
rect 2092 21652 2132 21692
rect 1996 19468 2036 19508
rect 2092 18628 2132 18668
rect 1900 12664 1940 12704
rect 1900 12496 1940 12536
rect 1804 11488 1844 11528
rect 1804 9976 1844 10016
rect 1612 8548 1652 8588
rect 1612 6448 1652 6488
rect 1900 4768 1940 4808
rect 1900 4264 1940 4304
rect 2668 35092 2708 35132
rect 2572 33664 2612 33704
rect 2668 34924 2708 34964
rect 2572 33100 2612 33140
rect 2572 28792 2612 28832
rect 2668 28372 2708 28412
rect 2284 21652 2324 21692
rect 2284 14680 2324 14720
rect 2188 11908 2228 11948
rect 2284 12832 2324 12872
rect 2284 7204 2324 7244
rect 2092 4852 2132 4892
rect 2188 3424 2228 3464
rect 2188 2836 2228 2876
rect 2572 22996 2612 23036
rect 2860 37276 2900 37316
rect 3052 36016 3092 36056
rect 2860 35176 2900 35216
rect 2956 34588 2996 34628
rect 3244 37612 3284 37652
rect 2956 30556 2996 30596
rect 3148 33244 3188 33284
rect 3436 44248 3476 44288
rect 3436 43240 3476 43280
rect 4928 45340 4968 45380
rect 5010 45340 5050 45380
rect 5092 45340 5132 45380
rect 5174 45340 5214 45380
rect 5256 45340 5296 45380
rect 5164 45172 5204 45212
rect 4588 44920 4628 44960
rect 3688 44584 3728 44624
rect 3770 44584 3810 44624
rect 3852 44584 3892 44624
rect 3934 44584 3974 44624
rect 4016 44584 4056 44624
rect 4492 44080 4532 44120
rect 4204 43408 4244 43448
rect 4928 43828 4968 43868
rect 5010 43828 5050 43868
rect 5092 43828 5132 43868
rect 5174 43828 5214 43868
rect 5256 43828 5296 43868
rect 4396 43324 4436 43364
rect 3688 43072 3728 43112
rect 3770 43072 3810 43112
rect 3852 43072 3892 43112
rect 3934 43072 3974 43112
rect 4016 43072 4056 43112
rect 3916 42904 3956 42944
rect 4588 42484 4628 42524
rect 4780 43240 4820 43280
rect 5644 43996 5684 44036
rect 6316 44248 6356 44288
rect 5836 44080 5876 44120
rect 5644 43408 5684 43448
rect 4928 42316 4968 42356
rect 5010 42316 5050 42356
rect 5092 42316 5132 42356
rect 5174 42316 5214 42356
rect 5256 42316 5296 42356
rect 3688 41560 3728 41600
rect 3770 41560 3810 41600
rect 3852 41560 3892 41600
rect 3934 41560 3974 41600
rect 4016 41560 4056 41600
rect 3688 40048 3728 40088
rect 3770 40048 3810 40088
rect 3852 40048 3892 40088
rect 3934 40048 3974 40088
rect 4016 40048 4056 40088
rect 3628 38872 3668 38912
rect 3688 38536 3728 38576
rect 3770 38536 3810 38576
rect 3852 38536 3892 38576
rect 3934 38536 3974 38576
rect 4016 38536 4056 38576
rect 3688 37024 3728 37064
rect 3770 37024 3810 37064
rect 3852 37024 3892 37064
rect 3934 37024 3974 37064
rect 4016 37024 4056 37064
rect 4012 36772 4052 36812
rect 3532 36436 3572 36476
rect 3628 35932 3668 35972
rect 3688 35512 3728 35552
rect 3770 35512 3810 35552
rect 3852 35512 3892 35552
rect 3934 35512 3974 35552
rect 4016 35512 4056 35552
rect 3436 33748 3476 33788
rect 3148 32320 3188 32360
rect 2860 29212 2900 29252
rect 2860 27532 2900 27572
rect 2860 27280 2900 27320
rect 2860 26944 2900 26984
rect 3628 35260 3668 35300
rect 3916 34924 3956 34964
rect 3688 34000 3728 34040
rect 3770 34000 3810 34040
rect 3852 34000 3892 34040
rect 3934 34000 3974 34040
rect 4016 34000 4056 34040
rect 3916 33832 3956 33872
rect 3688 32488 3728 32528
rect 3770 32488 3810 32528
rect 3852 32488 3892 32528
rect 3934 32488 3974 32528
rect 4016 32488 4056 32528
rect 3628 32320 3668 32360
rect 3148 29212 3188 29252
rect 3244 29716 3284 29756
rect 3052 28708 3092 28748
rect 2956 25348 2996 25388
rect 2668 22156 2708 22196
rect 2860 22492 2900 22532
rect 3244 28624 3284 28664
rect 3688 30976 3728 31016
rect 3770 30976 3810 31016
rect 3852 30976 3892 31016
rect 3934 30976 3974 31016
rect 4016 30976 4056 31016
rect 3916 30808 3956 30848
rect 3628 30640 3668 30680
rect 3628 30388 3668 30428
rect 3436 28624 3476 28664
rect 3532 29968 3572 30008
rect 3820 29968 3860 30008
rect 3628 29716 3668 29756
rect 3724 29632 3764 29672
rect 4012 30640 4052 30680
rect 4012 30388 4052 30428
rect 4204 35932 4244 35972
rect 4204 33832 4244 33872
rect 4300 33916 4340 33956
rect 4300 33328 4340 33368
rect 4204 30388 4244 30428
rect 3916 29632 3956 29672
rect 3688 29464 3728 29504
rect 3770 29464 3810 29504
rect 3852 29464 3892 29504
rect 3934 29464 3974 29504
rect 4016 29464 4056 29504
rect 4012 29212 4052 29252
rect 3244 24676 3284 24716
rect 3148 23164 3188 23204
rect 3244 23248 3284 23288
rect 3052 22660 3092 22700
rect 2860 20224 2900 20264
rect 2476 16276 2516 16316
rect 2572 16612 2612 16652
rect 4204 29212 4244 29252
rect 4928 40804 4968 40844
rect 5010 40804 5050 40844
rect 5092 40804 5132 40844
rect 5174 40804 5214 40844
rect 5256 40804 5296 40844
rect 4928 39292 4968 39332
rect 5010 39292 5050 39332
rect 5092 39292 5132 39332
rect 5174 39292 5214 39332
rect 5256 39292 5296 39332
rect 4928 37780 4968 37820
rect 5010 37780 5050 37820
rect 5092 37780 5132 37820
rect 5174 37780 5214 37820
rect 5256 37780 5296 37820
rect 4588 33412 4628 33452
rect 4012 28120 4052 28160
rect 3688 27952 3728 27992
rect 3770 27952 3810 27992
rect 3852 27952 3892 27992
rect 3934 27952 3974 27992
rect 4016 27952 4056 27992
rect 3688 26440 3728 26480
rect 3770 26440 3810 26480
rect 3852 26440 3892 26480
rect 3934 26440 3974 26480
rect 4016 26440 4056 26480
rect 3916 25348 3956 25388
rect 3688 24928 3728 24968
rect 3770 24928 3810 24968
rect 3852 24928 3892 24968
rect 3934 24928 3974 24968
rect 4016 24928 4056 24968
rect 3916 24340 3956 24380
rect 3688 23416 3728 23456
rect 3770 23416 3810 23456
rect 3852 23416 3892 23456
rect 3934 23416 3974 23456
rect 4016 23416 4056 23456
rect 4012 23080 4052 23120
rect 3436 22660 3476 22700
rect 3532 22324 3572 22364
rect 4012 22408 4052 22448
rect 3688 21904 3728 21944
rect 3770 21904 3810 21944
rect 3852 21904 3892 21944
rect 3934 21904 3974 21944
rect 4016 21904 4056 21944
rect 3916 20812 3956 20852
rect 4684 33244 4724 33284
rect 5068 36772 5108 36812
rect 5356 37444 5396 37484
rect 4928 36268 4968 36308
rect 5010 36268 5050 36308
rect 5092 36268 5132 36308
rect 5174 36268 5214 36308
rect 5256 36268 5296 36308
rect 5260 35848 5300 35888
rect 5356 35260 5396 35300
rect 4928 34756 4968 34796
rect 5010 34756 5050 34796
rect 5092 34756 5132 34796
rect 5174 34756 5214 34796
rect 5256 34756 5296 34796
rect 4876 34504 4916 34544
rect 4928 33244 4968 33284
rect 5010 33244 5050 33284
rect 5092 33244 5132 33284
rect 5174 33244 5214 33284
rect 5256 33244 5296 33284
rect 5260 32908 5300 32948
rect 5836 43324 5876 43364
rect 5932 42904 5972 42944
rect 5932 42652 5972 42692
rect 5932 42148 5972 42188
rect 5740 40972 5780 41012
rect 5836 38872 5876 38912
rect 6028 38116 6068 38156
rect 5644 37444 5684 37484
rect 5548 37276 5588 37316
rect 5740 36772 5780 36812
rect 5452 33412 5492 33452
rect 5452 32992 5492 33032
rect 4876 31900 4916 31940
rect 4928 31732 4968 31772
rect 5010 31732 5050 31772
rect 5092 31732 5132 31772
rect 5174 31732 5214 31772
rect 5256 31732 5296 31772
rect 5356 31480 5396 31520
rect 4588 28708 4628 28748
rect 4300 26020 4340 26060
rect 4396 25516 4436 25556
rect 4396 25348 4436 25388
rect 4928 30220 4968 30260
rect 5010 30220 5050 30260
rect 5092 30220 5132 30260
rect 5174 30220 5214 30260
rect 5256 30220 5296 30260
rect 4972 29968 5012 30008
rect 4780 29884 4820 29924
rect 5644 35260 5684 35300
rect 5644 33328 5684 33368
rect 5548 31480 5588 31520
rect 5644 31900 5684 31940
rect 5548 31312 5588 31352
rect 5356 29968 5396 30008
rect 5452 30556 5492 30596
rect 5548 29884 5588 29924
rect 5452 29716 5492 29756
rect 5452 29548 5492 29588
rect 4876 28960 4916 29000
rect 4928 28708 4968 28748
rect 5010 28708 5050 28748
rect 5092 28708 5132 28748
rect 5174 28708 5214 28748
rect 5256 28708 5296 28748
rect 4396 23164 4436 23204
rect 4204 23080 4244 23120
rect 3688 20392 3728 20432
rect 3770 20392 3810 20432
rect 3852 20392 3892 20432
rect 3934 20392 3974 20432
rect 4016 20392 4056 20432
rect 3340 20140 3380 20180
rect 2956 17620 2996 17660
rect 2956 15772 2996 15812
rect 3148 15100 3188 15140
rect 2860 14932 2900 14972
rect 3052 15016 3092 15056
rect 2764 14848 2804 14888
rect 2956 14848 2996 14888
rect 2572 14680 2612 14720
rect 2764 14680 2804 14720
rect 2764 12832 2804 12872
rect 2572 12496 2612 12536
rect 2476 11068 2516 11108
rect 2860 11908 2900 11948
rect 2860 11068 2900 11108
rect 3052 13756 3092 13796
rect 2860 8884 2900 8924
rect 2860 8632 2900 8672
rect 2956 2752 2996 2792
rect 2572 2584 2612 2624
rect 2764 232 2804 272
rect 3436 19804 3476 19844
rect 3532 20140 3572 20180
rect 3628 19384 3668 19424
rect 3724 19300 3764 19340
rect 4012 20056 4052 20096
rect 3916 19048 3956 19088
rect 3688 18880 3728 18920
rect 3770 18880 3810 18920
rect 3852 18880 3892 18920
rect 3934 18880 3974 18920
rect 4016 18880 4056 18920
rect 3436 17956 3476 17996
rect 3340 17200 3380 17240
rect 3688 17368 3728 17408
rect 3770 17368 3810 17408
rect 3852 17368 3892 17408
rect 3934 17368 3974 17408
rect 4016 17368 4056 17408
rect 3820 17200 3860 17240
rect 3628 17116 3668 17156
rect 3724 16948 3764 16988
rect 3628 16444 3668 16484
rect 3436 13756 3476 13796
rect 3436 13588 3476 13628
rect 3340 13084 3380 13124
rect 4108 16864 4148 16904
rect 3916 16780 3956 16820
rect 3688 15856 3728 15896
rect 3770 15856 3810 15896
rect 3852 15856 3892 15896
rect 3934 15856 3974 15896
rect 4016 15856 4056 15896
rect 3820 15520 3860 15560
rect 3724 14764 3764 14804
rect 3688 14344 3728 14384
rect 3770 14344 3810 14384
rect 3852 14344 3892 14384
rect 3934 14344 3974 14384
rect 4016 14344 4056 14384
rect 3628 13924 3668 13964
rect 3916 13000 3956 13040
rect 3532 12916 3572 12956
rect 4396 20812 4436 20852
rect 4492 19384 4532 19424
rect 4492 19216 4532 19256
rect 4396 16948 4436 16988
rect 4396 16360 4436 16400
rect 4300 15604 4340 15644
rect 4300 15268 4340 15308
rect 3688 12832 3728 12872
rect 3770 12832 3810 12872
rect 3852 12832 3892 12872
rect 3934 12832 3974 12872
rect 4016 12832 4056 12872
rect 3436 12748 3476 12788
rect 3340 12244 3380 12284
rect 3244 7792 3284 7832
rect 4204 12832 4244 12872
rect 3820 11656 3860 11696
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 4012 11152 4052 11192
rect 3820 10984 3860 11024
rect 3436 7792 3476 7832
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 3820 9388 3860 9428
rect 3340 4264 3380 4304
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 3628 7372 3668 7412
rect 3724 7120 3764 7160
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 3628 6616 3668 6656
rect 3820 6532 3860 6572
rect 3820 5440 3860 5480
rect 4108 5692 4148 5732
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 4928 27196 4968 27236
rect 5010 27196 5050 27236
rect 5092 27196 5132 27236
rect 5174 27196 5214 27236
rect 5256 27196 5296 27236
rect 4928 25684 4968 25724
rect 5010 25684 5050 25724
rect 5092 25684 5132 25724
rect 5174 25684 5214 25724
rect 5256 25684 5296 25724
rect 4928 24172 4968 24212
rect 5010 24172 5050 24212
rect 5092 24172 5132 24212
rect 5174 24172 5214 24212
rect 5256 24172 5296 24212
rect 4780 22996 4820 23036
rect 4876 23080 4916 23120
rect 4684 20644 4724 20684
rect 5644 27112 5684 27152
rect 5644 24676 5684 24716
rect 5452 23416 5492 23456
rect 5260 23080 5300 23120
rect 5260 22912 5300 22952
rect 5068 22828 5108 22868
rect 4928 22660 4968 22700
rect 5010 22660 5050 22700
rect 5092 22660 5132 22700
rect 5174 22660 5214 22700
rect 5256 22660 5296 22700
rect 5260 22492 5300 22532
rect 5068 22324 5108 22364
rect 5068 21652 5108 21692
rect 4928 21148 4968 21188
rect 5010 21148 5050 21188
rect 5092 21148 5132 21188
rect 5174 21148 5214 21188
rect 5256 21148 5296 21188
rect 4972 20980 5012 21020
rect 4876 20812 4916 20852
rect 4684 19216 4724 19256
rect 5548 22996 5588 23036
rect 5452 22828 5492 22868
rect 4972 19804 5012 19844
rect 4928 19636 4968 19676
rect 5010 19636 5050 19676
rect 5092 19636 5132 19676
rect 5174 19636 5214 19676
rect 5256 19636 5296 19676
rect 5644 22912 5684 22952
rect 5644 22660 5684 22700
rect 6028 36100 6068 36140
rect 5932 35428 5972 35468
rect 6220 36016 6260 36056
rect 6220 34924 6260 34964
rect 6220 34168 6260 34208
rect 6124 32824 6164 32864
rect 6124 32572 6164 32612
rect 5932 29800 5972 29840
rect 6124 27448 6164 27488
rect 6124 23836 6164 23876
rect 5932 22156 5972 22196
rect 5740 21484 5780 21524
rect 6220 22660 6260 22700
rect 6124 22156 6164 22196
rect 5164 19468 5204 19508
rect 5260 18292 5300 18332
rect 4928 18124 4968 18164
rect 5010 18124 5050 18164
rect 5092 18124 5132 18164
rect 5174 18124 5214 18164
rect 5256 18124 5296 18164
rect 4780 17788 4820 17828
rect 5068 17956 5108 17996
rect 4780 17200 4820 17240
rect 4780 16948 4820 16988
rect 4972 16864 5012 16904
rect 5164 16948 5204 16988
rect 5260 16780 5300 16820
rect 4928 16612 4968 16652
rect 5010 16612 5050 16652
rect 5092 16612 5132 16652
rect 5174 16612 5214 16652
rect 5256 16612 5296 16652
rect 4972 16444 5012 16484
rect 5356 16444 5396 16484
rect 4876 16192 4916 16232
rect 5260 15436 5300 15476
rect 4928 15100 4968 15140
rect 5010 15100 5050 15140
rect 5092 15100 5132 15140
rect 5174 15100 5214 15140
rect 5256 15100 5296 15140
rect 4876 14848 4916 14888
rect 5356 14596 5396 14636
rect 4928 13588 4968 13628
rect 5010 13588 5050 13628
rect 5092 13588 5132 13628
rect 5174 13588 5214 13628
rect 5256 13588 5296 13628
rect 4492 11824 4532 11864
rect 4396 10732 4436 10772
rect 4588 10228 4628 10268
rect 4300 5692 4340 5732
rect 4300 4096 4340 4136
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 3724 1912 3764 1952
rect 4396 3508 4436 3548
rect 4588 5944 4628 5984
rect 4588 4852 4628 4892
rect 4588 3256 4628 3296
rect 4928 12076 4968 12116
rect 5010 12076 5050 12116
rect 5092 12076 5132 12116
rect 5174 12076 5214 12116
rect 5256 12076 5296 12116
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 5260 7876 5300 7916
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 4972 5440 5012 5480
rect 4972 4852 5012 4892
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 5548 19384 5588 19424
rect 5932 19720 5972 19760
rect 6028 19636 6068 19676
rect 5932 17620 5972 17660
rect 5740 17032 5780 17072
rect 5740 16276 5780 16316
rect 5548 14680 5588 14720
rect 5452 13084 5492 13124
rect 5452 11908 5492 11948
rect 5740 15688 5780 15728
rect 5644 13168 5684 13208
rect 5740 13840 5780 13880
rect 5644 12832 5684 12872
rect 6028 15436 6068 15476
rect 5932 14596 5972 14636
rect 5740 11908 5780 11948
rect 5644 11740 5684 11780
rect 5548 10060 5588 10100
rect 6220 18124 6260 18164
rect 6604 42652 6644 42692
rect 6508 42568 6548 42608
rect 6700 36016 6740 36056
rect 6700 35344 6740 35384
rect 6412 32656 6452 32696
rect 6412 32488 6452 32528
rect 6604 28288 6644 28328
rect 6796 33412 6836 33452
rect 6796 33244 6836 33284
rect 6892 32152 6932 32192
rect 6796 28876 6836 28916
rect 7084 32488 7124 32528
rect 7180 33496 7220 33536
rect 6988 31732 7028 31772
rect 7084 32152 7124 32192
rect 6796 28456 6836 28496
rect 6412 24256 6452 24296
rect 6508 22912 6548 22952
rect 6412 19636 6452 19676
rect 6700 27868 6740 27908
rect 6700 27280 6740 27320
rect 7852 42652 7892 42692
rect 7372 36688 7412 36728
rect 7756 38200 7796 38240
rect 7948 37444 7988 37484
rect 8140 39628 8180 39668
rect 7948 35596 7988 35636
rect 7276 33244 7316 33284
rect 7180 28456 7220 28496
rect 6796 24256 6836 24296
rect 6316 17788 6356 17828
rect 6412 18208 6452 18248
rect 6220 16780 6260 16820
rect 6220 14848 6260 14888
rect 5644 7204 5684 7244
rect 5548 4096 5588 4136
rect 6220 6616 6260 6656
rect 6220 6364 6260 6404
rect 6700 20980 6740 21020
rect 6700 20308 6740 20348
rect 6796 18208 6836 18248
rect 6796 18040 6836 18080
rect 6700 17956 6740 17996
rect 6412 5356 6452 5396
rect 6508 2836 6548 2876
rect 6796 17368 6836 17408
rect 6700 5860 6740 5900
rect 7564 31228 7604 31268
rect 7468 26104 7508 26144
rect 7852 31564 7892 31604
rect 7276 22996 7316 23036
rect 6988 17956 7028 17996
rect 6892 14428 6932 14468
rect 6988 17788 7028 17828
rect 6892 14260 6932 14300
rect 7276 20308 7316 20348
rect 7276 20140 7316 20180
rect 7180 16948 7220 16988
rect 7084 14260 7124 14300
rect 7084 12748 7124 12788
rect 6892 5356 6932 5396
rect 6988 8716 7028 8756
rect 7180 8716 7220 8756
rect 7180 5944 7220 5984
rect 7564 23080 7604 23120
rect 7468 22744 7508 22784
rect 7468 19216 7508 19256
rect 7468 17368 7508 17408
rect 8140 35092 8180 35132
rect 8044 30724 8084 30764
rect 8428 42568 8468 42608
rect 8428 39712 8468 39752
rect 8428 38200 8468 38240
rect 8428 35596 8468 35636
rect 7948 27532 7988 27572
rect 7948 25852 7988 25892
rect 8332 32908 8372 32948
rect 8236 31564 8276 31604
rect 8332 31228 8372 31268
rect 8332 30724 8372 30764
rect 8236 29800 8276 29840
rect 8236 27532 8276 27572
rect 8332 28960 8372 29000
rect 7852 22996 7892 23036
rect 8044 22744 8084 22784
rect 8044 22492 8084 22532
rect 7852 18544 7892 18584
rect 7756 15016 7796 15056
rect 7564 9388 7604 9428
rect 7852 11908 7892 11948
rect 8812 34840 8852 34880
rect 8428 26104 8468 26144
rect 8716 30892 8756 30932
rect 8812 30304 8852 30344
rect 8716 29800 8756 29840
rect 8620 26692 8660 26732
rect 8332 21568 8372 21608
rect 8140 17452 8180 17492
rect 9100 32992 9140 33032
rect 9100 32068 9140 32108
rect 9964 42736 10004 42776
rect 9964 40384 10004 40424
rect 10060 40300 10100 40340
rect 9484 36436 9524 36476
rect 9388 34840 9428 34880
rect 9292 32908 9332 32948
rect 8716 19384 8756 19424
rect 8716 19216 8756 19256
rect 8524 18544 8564 18584
rect 8332 9388 8372 9428
rect 7372 1408 7412 1448
rect 8140 1408 8180 1448
rect 9100 28204 9140 28244
rect 8908 20644 8948 20684
rect 8908 19384 8948 19424
rect 8812 17620 8852 17660
rect 9484 32908 9524 32948
rect 9580 31984 9620 32024
rect 9580 30136 9620 30176
rect 8812 5692 8852 5732
rect 9676 28876 9716 28916
rect 9580 28204 9620 28244
rect 9388 24340 9428 24380
rect 9388 18124 9428 18164
rect 9100 13588 9140 13628
rect 9580 14008 9620 14048
rect 9484 13588 9524 13628
rect 9676 13672 9716 13712
rect 9676 13504 9716 13544
rect 9964 36688 10004 36728
rect 9868 30388 9908 30428
rect 9868 30136 9908 30176
rect 10060 32824 10100 32864
rect 10348 42736 10388 42776
rect 10348 41896 10388 41936
rect 10444 39460 10484 39500
rect 10444 38872 10484 38912
rect 9964 28372 10004 28412
rect 10060 30220 10100 30260
rect 9868 28036 9908 28076
rect 9964 24340 10004 24380
rect 10060 20140 10100 20180
rect 10348 29128 10388 29168
rect 10252 22576 10292 22616
rect 10348 21736 10388 21776
rect 10348 21400 10388 21440
rect 10156 18712 10196 18752
rect 10060 18544 10100 18584
rect 9964 18124 10004 18164
rect 9964 13672 10004 13712
rect 10156 11572 10196 11612
rect 9964 6448 10004 6488
rect 10540 28036 10580 28076
rect 10732 40216 10772 40256
rect 10924 33160 10964 33200
rect 10828 33076 10868 33116
rect 10828 32908 10868 32948
rect 10924 32824 10964 32864
rect 10924 28960 10964 29000
rect 11020 29044 11060 29084
rect 10732 28036 10772 28076
rect 10732 21736 10772 21776
rect 10540 18544 10580 18584
rect 10732 18208 10772 18248
rect 10636 17788 10676 17828
rect 10540 14092 10580 14132
rect 10444 10060 10484 10100
rect 10924 17956 10964 17996
rect 11020 27700 11060 27740
rect 11212 28960 11252 29000
rect 11500 29044 11540 29084
rect 11692 27700 11732 27740
rect 11308 22576 11348 22616
rect 11212 17956 11252 17996
rect 11500 17956 11540 17996
<< metal4 >>
rect 4919 45340 4928 45380
rect 4968 45340 5010 45380
rect 5050 45340 5092 45380
rect 5132 45340 5174 45380
rect 5214 45340 5256 45380
rect 5296 45340 5305 45380
rect 1987 45172 1996 45212
rect 2036 45172 5164 45212
rect 5204 45172 5213 45212
rect 2755 44920 2764 44960
rect 2804 44920 4588 44960
rect 4628 44920 4637 44960
rect 3679 44584 3688 44624
rect 3728 44584 3770 44624
rect 3810 44584 3852 44624
rect 3892 44584 3934 44624
rect 3974 44584 4016 44624
rect 4056 44584 4065 44624
rect 67 44248 76 44288
rect 116 44248 3436 44288
rect 3476 44248 3485 44288
rect 6307 44248 6316 44288
rect 6356 44248 6412 44288
rect 6452 44248 6461 44288
rect 4483 44080 4492 44120
rect 4532 44080 5836 44120
rect 5876 44080 5885 44120
rect 5635 43996 5644 44036
rect 5684 43996 5693 44036
rect 4919 43828 4928 43868
rect 4968 43828 5010 43868
rect 5050 43828 5092 43868
rect 5132 43828 5174 43868
rect 5214 43828 5256 43868
rect 5296 43828 5305 43868
rect 5644 43448 5684 43996
rect 4195 43408 4204 43448
rect 4244 43408 4532 43448
rect 5635 43408 5644 43448
rect 5684 43408 5693 43448
rect 4492 43364 4532 43408
rect 3139 43324 3148 43364
rect 3188 43324 4396 43364
rect 4436 43324 4445 43364
rect 4492 43324 5836 43364
rect 5876 43324 5885 43364
rect 3427 43240 3436 43280
rect 3476 43240 4780 43280
rect 4820 43240 4829 43280
rect 3679 43072 3688 43112
rect 3728 43072 3770 43112
rect 3810 43072 3852 43112
rect 3892 43072 3934 43112
rect 3974 43072 4016 43112
rect 4056 43072 4065 43112
rect 3235 42988 3244 43028
rect 3284 42988 6508 43028
rect 6548 42988 6557 43028
rect 3907 42904 3916 42944
rect 3956 42904 5932 42944
rect 5972 42904 5981 42944
rect 9763 42736 9772 42776
rect 9812 42736 9964 42776
rect 10004 42736 10013 42776
rect 10147 42736 10156 42776
rect 10196 42736 10348 42776
rect 10388 42736 10397 42776
rect 2467 42652 2476 42692
rect 2516 42652 5932 42692
rect 5972 42652 6604 42692
rect 6644 42652 7852 42692
rect 7892 42652 7901 42692
rect 2947 42568 2956 42608
rect 2996 42568 6508 42608
rect 6548 42568 8428 42608
rect 8468 42568 8477 42608
rect 4493 42484 4588 42524
rect 4628 42484 4637 42524
rect 4919 42316 4928 42356
rect 4968 42316 5010 42356
rect 5050 42316 5092 42356
rect 5132 42316 5174 42356
rect 5214 42316 5256 42356
rect 5296 42316 5305 42356
rect 3139 42148 3148 42188
rect 3188 42148 5932 42188
rect 5972 42148 5981 42188
rect 10253 41896 10348 41936
rect 10388 41896 10397 41936
rect 2957 41812 3052 41852
rect 3092 41812 3101 41852
rect 3679 41560 3688 41600
rect 3728 41560 3770 41600
rect 3810 41560 3852 41600
rect 3892 41560 3934 41600
rect 3974 41560 4016 41600
rect 4056 41560 4065 41600
rect 1517 40972 1612 41012
rect 1652 40972 1661 41012
rect 5645 40972 5740 41012
rect 5780 40972 5789 41012
rect 4919 40804 4928 40844
rect 4968 40804 5010 40844
rect 5050 40804 5092 40844
rect 5132 40804 5174 40844
rect 5214 40804 5256 40844
rect 5296 40804 5305 40844
rect 9869 40384 9964 40424
rect 10004 40384 10013 40424
rect 10051 40300 10060 40340
rect 10100 40300 10109 40340
rect 10060 40256 10100 40300
rect 10060 40216 10732 40256
rect 10772 40216 10781 40256
rect 3679 40048 3688 40088
rect 3728 40048 3770 40088
rect 3810 40048 3852 40088
rect 3892 40048 3934 40088
rect 3974 40048 4016 40088
rect 4056 40048 4065 40088
rect 2947 39712 2956 39752
rect 2996 39712 3091 39752
rect 7075 39712 7084 39752
rect 7124 39712 8428 39752
rect 8468 39712 8477 39752
rect 8131 39628 8140 39668
rect 8180 39628 8524 39668
rect 8564 39628 8573 39668
rect 2851 39460 2860 39500
rect 2900 39460 2995 39500
rect 10349 39460 10444 39500
rect 10484 39460 10493 39500
rect 4919 39292 4928 39332
rect 4968 39292 5010 39332
rect 5050 39292 5092 39332
rect 5132 39292 5174 39332
rect 5214 39292 5256 39332
rect 5296 39292 5305 39332
rect 3427 38872 3436 38912
rect 3476 38872 3628 38912
rect 3668 38872 3677 38912
rect 5741 38872 5836 38912
rect 5876 38872 5885 38912
rect 10243 38872 10252 38912
rect 10292 38872 10444 38912
rect 10484 38872 10493 38912
rect 3679 38536 3688 38576
rect 3728 38536 3770 38576
rect 3810 38536 3852 38576
rect 3892 38536 3934 38576
rect 3974 38536 4016 38576
rect 4056 38536 4065 38576
rect 7747 38200 7756 38240
rect 7796 38200 8428 38240
rect 8468 38200 8477 38240
rect 355 38116 364 38156
rect 404 38116 6028 38156
rect 6068 38116 6077 38156
rect 4919 37780 4928 37820
rect 4968 37780 5010 37820
rect 5050 37780 5092 37820
rect 5132 37780 5174 37820
rect 5214 37780 5256 37820
rect 5296 37780 5305 37820
rect 3149 37612 3244 37652
rect 3284 37612 3293 37652
rect 2860 37528 5452 37568
rect 5492 37528 5501 37568
rect 2860 37484 2900 37528
rect 2275 37444 2284 37484
rect 2324 37444 2900 37484
rect 5347 37444 5356 37484
rect 5396 37444 5644 37484
rect 5684 37444 5693 37484
rect 7853 37444 7948 37484
rect 7988 37444 7997 37484
rect 2851 37276 2860 37316
rect 2900 37276 5548 37316
rect 5588 37276 5597 37316
rect 1421 37192 1516 37232
rect 1556 37192 1565 37232
rect 3679 37024 3688 37064
rect 3728 37024 3770 37064
rect 3810 37024 3852 37064
rect 3892 37024 3934 37064
rect 3974 37024 4016 37064
rect 4056 37024 4065 37064
rect 2659 36772 2668 36812
rect 2708 36772 4012 36812
rect 4052 36772 4061 36812
rect 5059 36772 5068 36812
rect 5108 36772 5548 36812
rect 5588 36772 5740 36812
rect 5780 36772 5789 36812
rect 7171 36688 7180 36728
rect 7220 36688 7372 36728
rect 7412 36688 7421 36728
rect 9571 36688 9580 36728
rect 9620 36688 9964 36728
rect 10004 36688 10013 36728
rect 2371 36604 2380 36644
rect 2420 36604 2476 36644
rect 2516 36604 2525 36644
rect 3437 36436 3532 36476
rect 3572 36436 3581 36476
rect 9389 36436 9484 36476
rect 9524 36436 9533 36476
rect 4919 36268 4928 36308
rect 4968 36268 5010 36308
rect 5050 36268 5092 36308
rect 5132 36268 5174 36308
rect 5214 36268 5256 36308
rect 5296 36268 5305 36308
rect 5932 36100 6028 36140
rect 6068 36100 6077 36140
rect 3043 36016 3052 36056
rect 3092 36016 3244 36056
rect 3284 36016 3293 36056
rect 3619 35932 3628 35972
rect 3668 35932 4204 35972
rect 4244 35932 4253 35972
rect 5251 35848 5260 35888
rect 5300 35848 5548 35888
rect 5588 35848 5597 35888
rect 3679 35512 3688 35552
rect 3728 35512 3770 35552
rect 3810 35512 3852 35552
rect 3892 35512 3934 35552
rect 3974 35512 4016 35552
rect 4056 35512 4065 35552
rect 5932 35468 5972 36100
rect 6211 36016 6220 36056
rect 6260 36016 6700 36056
rect 6740 36016 6749 36056
rect 7939 35596 7948 35636
rect 7988 35596 8428 35636
rect 8468 35596 8477 35636
rect 2275 35428 2284 35468
rect 2324 35428 2572 35468
rect 2612 35428 2621 35468
rect 5923 35428 5932 35468
rect 5972 35428 5981 35468
rect 2275 35344 2284 35384
rect 2324 35344 6700 35384
rect 6740 35344 6749 35384
rect 2947 35260 2956 35300
rect 2996 35260 3628 35300
rect 3668 35260 3677 35300
rect 5347 35260 5356 35300
rect 5396 35260 5644 35300
rect 5684 35260 5693 35300
rect 2179 35176 2188 35216
rect 2228 35176 2860 35216
rect 2900 35176 2909 35216
rect 2659 35092 2668 35132
rect 2708 35092 8140 35132
rect 8180 35092 8189 35132
rect 2467 34924 2476 34964
rect 2516 34924 2668 34964
rect 2708 34924 2717 34964
rect 3907 34924 3916 34964
rect 3956 34924 5644 34964
rect 5684 34924 6220 34964
rect 6260 34924 6269 34964
rect 8803 34840 8812 34880
rect 8852 34840 9388 34880
rect 9428 34840 9437 34880
rect 4919 34756 4928 34796
rect 4968 34756 5010 34796
rect 5050 34756 5092 34796
rect 5132 34756 5174 34796
rect 5214 34756 5256 34796
rect 5296 34756 5305 34796
rect 1987 34588 1996 34628
rect 2036 34588 2956 34628
rect 2996 34588 3005 34628
rect 1027 34504 1036 34544
rect 1076 34504 4876 34544
rect 4916 34504 4925 34544
rect 67 34168 76 34208
rect 116 34168 6220 34208
rect 6260 34168 6269 34208
rect 3679 34000 3688 34040
rect 3728 34000 3770 34040
rect 3810 34000 3852 34040
rect 3892 34000 3934 34040
rect 3974 34000 4016 34040
rect 4056 34000 4065 34040
rect 2083 33916 2092 33956
rect 2132 33916 4300 33956
rect 4340 33916 4349 33956
rect 3907 33832 3916 33872
rect 3956 33832 4204 33872
rect 4244 33832 4253 33872
rect 3148 33748 3436 33788
rect 3476 33748 3485 33788
rect 1507 33664 1516 33704
rect 1556 33664 2572 33704
rect 2612 33664 2621 33704
rect 1123 33496 1132 33536
rect 1172 33496 1420 33536
rect 1460 33496 1469 33536
rect 3148 33284 3188 33748
rect 7085 33496 7180 33536
rect 7220 33496 7229 33536
rect 4579 33412 4588 33452
rect 4628 33412 5452 33452
rect 5492 33412 5501 33452
rect 6691 33412 6700 33452
rect 6740 33412 6796 33452
rect 6836 33412 6845 33452
rect 4291 33328 4300 33368
rect 4340 33328 5644 33368
rect 5684 33328 5693 33368
rect 3139 33244 3148 33284
rect 3188 33244 3197 33284
rect 4675 33244 4684 33284
rect 4724 33244 4733 33284
rect 4919 33244 4928 33284
rect 4968 33244 5010 33284
rect 5050 33244 5092 33284
rect 5132 33244 5174 33284
rect 5214 33244 5256 33284
rect 5296 33244 5305 33284
rect 6787 33244 6796 33284
rect 6836 33244 7276 33284
rect 7316 33244 7325 33284
rect 2285 33160 2380 33200
rect 2420 33160 2429 33200
rect 1613 33076 1708 33116
rect 1748 33076 1757 33116
rect 2563 33100 2572 33140
rect 2612 33100 2621 33140
rect 4684 33116 4724 33244
rect 10915 33160 10924 33200
rect 10964 33160 10973 33200
rect 2572 33032 2612 33100
rect 4684 33076 5492 33116
rect 10819 33076 10828 33116
rect 10868 33076 10877 33116
rect 5452 33032 5492 33076
rect 1891 32992 1900 33032
rect 1940 32992 2612 33032
rect 5443 32992 5452 33032
rect 5492 32992 5501 33032
rect 9005 32992 9100 33032
rect 9140 32992 9149 33032
rect 10828 32948 10868 33076
rect 5251 32908 5260 32948
rect 5300 32908 8332 32948
rect 8372 32908 8381 32948
rect 9283 32908 9292 32948
rect 9332 32908 9484 32948
rect 9524 32908 9533 32948
rect 10819 32908 10828 32948
rect 10868 32908 10877 32948
rect 10924 32864 10964 33160
rect 1603 32824 1612 32864
rect 1652 32824 1661 32864
rect 6115 32824 6124 32864
rect 6164 32824 6220 32864
rect 6260 32824 6269 32864
rect 9965 32824 10060 32864
rect 10100 32824 10109 32864
rect 10915 32824 10924 32864
rect 10964 32824 10973 32864
rect 1612 32780 1652 32824
rect 1612 32740 1804 32780
rect 1844 32740 1853 32780
rect 6403 32656 6412 32696
rect 6452 32656 7852 32696
rect 7892 32656 7901 32696
rect 5635 32572 5644 32612
rect 5684 32572 6124 32612
rect 6164 32572 6173 32612
rect 3679 32488 3688 32528
rect 3728 32488 3770 32528
rect 3810 32488 3852 32528
rect 3892 32488 3934 32528
rect 3974 32488 4016 32528
rect 4056 32488 4065 32528
rect 6403 32488 6412 32528
rect 6452 32488 7084 32528
rect 7124 32488 7133 32528
rect 3139 32320 3148 32360
rect 3188 32320 3628 32360
rect 3668 32320 3677 32360
rect 6883 32152 6892 32192
rect 6932 32152 7084 32192
rect 7124 32152 7133 32192
rect 9091 32068 9100 32108
rect 9140 32068 9149 32108
rect 9100 32024 9140 32068
rect 835 31984 844 32024
rect 884 31984 1132 32024
rect 1172 31984 1181 32024
rect 9100 31984 9580 32024
rect 9620 31984 9629 32024
rect 4675 31900 4684 31940
rect 4724 31900 4876 31940
rect 4916 31900 4925 31940
rect 5539 31900 5548 31940
rect 5588 31900 5644 31940
rect 5684 31900 5693 31940
rect 4919 31732 4928 31772
rect 4968 31732 5010 31772
rect 5050 31732 5092 31772
rect 5132 31732 5174 31772
rect 5214 31732 5256 31772
rect 5296 31732 5305 31772
rect 6979 31732 6988 31772
rect 7028 31732 7372 31772
rect 7412 31732 7421 31772
rect 2083 31564 2092 31604
rect 2132 31564 2284 31604
rect 2324 31564 2333 31604
rect 7843 31564 7852 31604
rect 7892 31564 8236 31604
rect 8276 31564 8285 31604
rect 1027 31480 1036 31520
rect 1076 31480 1085 31520
rect 5347 31480 5356 31520
rect 5396 31480 5548 31520
rect 5588 31480 5597 31520
rect 1036 31016 1076 31480
rect 5453 31312 5548 31352
rect 5588 31312 5597 31352
rect 1325 31228 1420 31268
rect 1460 31228 1469 31268
rect 7469 31228 7564 31268
rect 7604 31228 8332 31268
rect 8372 31228 8381 31268
rect 1036 30976 1228 31016
rect 1268 30976 1277 31016
rect 3679 30976 3688 31016
rect 3728 30976 3770 31016
rect 3810 30976 3852 31016
rect 3892 30976 3934 31016
rect 3974 30976 4016 31016
rect 4056 30976 4065 31016
rect 1507 30892 1516 30932
rect 1556 30892 8716 30932
rect 8756 30892 8765 30932
rect 3916 30848 3956 30892
rect 3907 30808 3916 30848
rect 3956 30808 3965 30848
rect 8035 30724 8044 30764
rect 8084 30724 8332 30764
rect 8372 30724 8381 30764
rect 3523 30640 3532 30680
rect 3572 30640 3628 30680
rect 3668 30640 3677 30680
rect 4003 30640 4012 30680
rect 4052 30640 7084 30680
rect 7124 30640 7133 30680
rect 3628 30596 3668 30640
rect 2947 30556 2956 30596
rect 2996 30556 3091 30596
rect 3628 30556 5452 30596
rect 5492 30556 5501 30596
rect 3619 30388 3628 30428
rect 3668 30388 4012 30428
rect 4052 30388 4204 30428
rect 4244 30388 4253 30428
rect 9773 30388 9868 30428
rect 9908 30388 9917 30428
rect 8803 30304 8812 30344
rect 8852 30304 10100 30344
rect 10060 30260 10100 30304
rect 1699 30220 1708 30260
rect 1748 30220 1996 30260
rect 2036 30220 2045 30260
rect 4919 30220 4928 30260
rect 4968 30220 5010 30260
rect 5050 30220 5092 30260
rect 5132 30220 5174 30260
rect 5214 30220 5256 30260
rect 5296 30220 5305 30260
rect 10051 30220 10060 30260
rect 10100 30220 10109 30260
rect 9571 30136 9580 30176
rect 9620 30136 9868 30176
rect 9908 30136 9917 30176
rect 1325 29968 1420 30008
rect 1460 29968 1469 30008
rect 3523 29968 3532 30008
rect 3572 29968 3820 30008
rect 3860 29968 3869 30008
rect 4771 29968 4780 30008
rect 4820 29968 4972 30008
rect 5012 29968 5356 30008
rect 5396 29968 5405 30008
rect 1699 29884 1708 29924
rect 1748 29884 4780 29924
rect 4820 29884 4829 29924
rect 5539 29884 5548 29924
rect 5588 29884 5644 29924
rect 5684 29884 5693 29924
rect 1315 29800 1324 29840
rect 1364 29800 5932 29840
rect 5972 29800 5981 29840
rect 8141 29800 8236 29840
rect 8276 29800 8285 29840
rect 8621 29800 8716 29840
rect 8756 29800 8765 29840
rect 3235 29716 3244 29756
rect 3284 29716 3628 29756
rect 3668 29716 3677 29756
rect 4387 29716 4396 29756
rect 4436 29716 5452 29756
rect 5492 29716 5501 29756
rect 3715 29632 3724 29672
rect 3764 29632 3773 29672
rect 3907 29632 3916 29672
rect 3956 29632 4204 29672
rect 4244 29632 4253 29672
rect 3724 29588 3764 29632
rect 3724 29548 5452 29588
rect 5492 29548 5501 29588
rect 3679 29464 3688 29504
rect 3728 29464 3770 29504
rect 3810 29464 3852 29504
rect 3892 29464 3934 29504
rect 3974 29464 4016 29504
rect 4056 29464 4065 29504
rect 2851 29212 2860 29252
rect 2900 29212 3148 29252
rect 3188 29212 3197 29252
rect 4003 29212 4012 29252
rect 4052 29212 4204 29252
rect 4244 29212 4253 29252
rect 1603 29128 1612 29168
rect 1652 29128 10348 29168
rect 10388 29128 10397 29168
rect 11011 29044 11020 29084
rect 11060 29044 11500 29084
rect 11540 29044 11549 29084
rect 4867 28960 4876 29000
rect 4916 28960 8332 29000
rect 8372 28960 8381 29000
rect 10915 28960 10924 29000
rect 10964 28960 11212 29000
rect 11252 28960 11261 29000
rect 6701 28876 6796 28916
rect 6836 28876 6845 28916
rect 9581 28876 9676 28916
rect 9716 28876 9725 28916
rect 1699 28792 1708 28832
rect 1748 28792 2572 28832
rect 2612 28792 2621 28832
rect 2755 28708 2764 28748
rect 2804 28708 3052 28748
rect 3092 28708 3101 28748
rect 3148 28708 4588 28748
rect 4628 28708 4637 28748
rect 4919 28708 4928 28748
rect 4968 28708 5010 28748
rect 5050 28708 5092 28748
rect 5132 28708 5174 28748
rect 5214 28708 5256 28748
rect 5296 28708 5305 28748
rect 3148 28664 3188 28708
rect 2563 28624 2572 28664
rect 2612 28624 3188 28664
rect 3235 28624 3244 28664
rect 3284 28624 3436 28664
rect 3476 28624 3485 28664
rect 6787 28456 6796 28496
rect 6836 28456 7180 28496
rect 7220 28456 7229 28496
rect 2659 28372 2668 28412
rect 2708 28372 9100 28412
rect 9140 28372 9149 28412
rect 9955 28372 9964 28412
rect 10004 28372 10013 28412
rect 6509 28288 6604 28328
rect 6644 28288 6653 28328
rect 9005 28204 9100 28244
rect 9140 28204 9580 28244
rect 9620 28204 9629 28244
rect 3235 28120 3244 28160
rect 3284 28120 4012 28160
rect 4052 28120 4061 28160
rect 9964 28076 10004 28372
rect 9859 28036 9868 28076
rect 9908 28036 10004 28076
rect 10531 28036 10540 28076
rect 10580 28036 10732 28076
rect 10772 28036 10781 28076
rect 3679 27952 3688 27992
rect 3728 27952 3770 27992
rect 3810 27952 3852 27992
rect 3892 27952 3934 27992
rect 3974 27952 4016 27992
rect 4056 27952 4065 27992
rect 6605 27868 6700 27908
rect 6740 27868 6749 27908
rect 11011 27700 11020 27740
rect 11060 27700 11692 27740
rect 11732 27700 11741 27740
rect 1411 27532 1420 27572
rect 1460 27532 1469 27572
rect 2851 27532 2860 27572
rect 2900 27532 2956 27572
rect 2996 27532 3005 27572
rect 7939 27532 7948 27572
rect 7988 27532 8236 27572
rect 8276 27532 8285 27572
rect 1420 27320 1460 27532
rect 1699 27448 1708 27488
rect 1748 27448 6124 27488
rect 6164 27448 6173 27488
rect 1420 27280 1708 27320
rect 1748 27280 1757 27320
rect 2851 27280 2860 27320
rect 2900 27280 6700 27320
rect 6740 27280 6749 27320
rect 4919 27196 4928 27236
rect 4968 27196 5010 27236
rect 5050 27196 5092 27236
rect 5132 27196 5174 27236
rect 5214 27196 5256 27236
rect 5296 27196 5305 27236
rect 5549 27112 5644 27152
rect 5684 27112 5693 27152
rect 2851 26944 2860 26984
rect 2900 26944 9772 26984
rect 9812 26944 9821 26984
rect 1603 26692 1612 26732
rect 1652 26692 8620 26732
rect 8660 26692 8669 26732
rect 3679 26440 3688 26480
rect 3728 26440 3770 26480
rect 3810 26440 3852 26480
rect 3892 26440 3934 26480
rect 3974 26440 4016 26480
rect 4056 26440 4065 26480
rect 7459 26104 7468 26144
rect 7508 26104 8428 26144
rect 8468 26104 8477 26144
rect 4291 26020 4300 26060
rect 4340 26020 4780 26060
rect 4820 26020 4829 26060
rect 7651 25852 7660 25892
rect 7700 25852 7948 25892
rect 7988 25852 7997 25892
rect 4919 25684 4928 25724
rect 4968 25684 5010 25724
rect 5050 25684 5092 25724
rect 5132 25684 5174 25724
rect 5214 25684 5256 25724
rect 5296 25684 5305 25724
rect 4387 25516 4396 25556
rect 4436 25516 5644 25556
rect 5684 25516 5693 25556
rect 2947 25348 2956 25388
rect 2996 25348 3916 25388
rect 3956 25348 3965 25388
rect 4301 25348 4396 25388
rect 4436 25348 4445 25388
rect 3679 24928 3688 24968
rect 3728 24928 3770 24968
rect 3810 24928 3852 24968
rect 3892 24928 3934 24968
rect 3974 24928 4016 24968
rect 4056 24928 4065 24968
rect 1795 24676 1804 24716
rect 1844 24676 3244 24716
rect 3284 24676 3293 24716
rect 5635 24676 5644 24716
rect 5684 24676 5693 24716
rect 5644 24464 5684 24676
rect 5644 24424 8140 24464
rect 8180 24424 8189 24464
rect 451 24340 460 24380
rect 500 24340 844 24380
rect 884 24340 893 24380
rect 3523 24340 3532 24380
rect 3572 24340 3916 24380
rect 3956 24340 3965 24380
rect 9379 24340 9388 24380
rect 9428 24340 9964 24380
rect 10004 24340 10013 24380
rect 6403 24256 6412 24296
rect 6452 24256 6796 24296
rect 6836 24256 6845 24296
rect 4919 24172 4928 24212
rect 4968 24172 5010 24212
rect 5050 24172 5092 24212
rect 5132 24172 5174 24212
rect 5214 24172 5256 24212
rect 5296 24172 5305 24212
rect 6115 23836 6124 23876
rect 6164 23836 6316 23876
rect 6356 23836 6365 23876
rect 3679 23416 3688 23456
rect 3728 23416 3770 23456
rect 3810 23416 3852 23456
rect 3892 23416 3934 23456
rect 3974 23416 4016 23456
rect 4056 23416 4065 23456
rect 5443 23416 5452 23456
rect 5492 23416 9772 23456
rect 9812 23416 9821 23456
rect 3149 23248 3244 23288
rect 3284 23248 3293 23288
rect 3139 23164 3148 23204
rect 3188 23164 4396 23204
rect 4436 23164 4445 23204
rect 1891 23080 1900 23120
rect 1940 23080 4012 23120
rect 4052 23080 4061 23120
rect 4109 23080 4204 23120
rect 4244 23080 4253 23120
rect 4771 23080 4780 23120
rect 4820 23080 4876 23120
rect 4916 23080 4925 23120
rect 5251 23080 5260 23120
rect 5300 23080 7564 23120
rect 7604 23080 7660 23120
rect 7700 23080 7728 23120
rect 2563 22996 2572 23036
rect 2612 22996 3340 23036
rect 3380 22996 3389 23036
rect 4771 22996 4780 23036
rect 4820 22996 5548 23036
rect 5588 22996 5597 23036
rect 7267 22996 7276 23036
rect 7316 22996 7852 23036
rect 7892 22996 7901 23036
rect 3235 22912 3244 22952
rect 3284 22912 5260 22952
rect 5300 22912 5309 22952
rect 5635 22912 5644 22952
rect 5684 22912 5932 22952
rect 5972 22912 5981 22952
rect 6499 22912 6508 22952
rect 6548 22912 6557 22952
rect 3139 22828 3148 22868
rect 3188 22828 5068 22868
rect 5108 22828 5117 22868
rect 5443 22828 5452 22868
rect 5492 22828 5684 22868
rect 1699 22744 1708 22784
rect 1748 22744 4396 22784
rect 4436 22744 4445 22784
rect 5644 22700 5684 22828
rect 6508 22700 6548 22912
rect 7459 22744 7468 22784
rect 7508 22744 8044 22784
rect 8084 22744 8093 22784
rect 3043 22660 3052 22700
rect 3092 22660 3436 22700
rect 3476 22660 3485 22700
rect 4919 22660 4928 22700
rect 4968 22660 5010 22700
rect 5050 22660 5092 22700
rect 5132 22660 5174 22700
rect 5214 22660 5256 22700
rect 5296 22660 5305 22700
rect 5635 22660 5644 22700
rect 5684 22660 5693 22700
rect 6211 22660 6220 22700
rect 6260 22660 6548 22700
rect 10243 22576 10252 22616
rect 10292 22576 11308 22616
rect 11348 22576 11357 22616
rect 2851 22492 2860 22532
rect 2900 22492 5260 22532
rect 5300 22492 5309 22532
rect 6499 22492 6508 22532
rect 6548 22492 8044 22532
rect 8084 22492 8093 22532
rect 67 22408 76 22448
rect 116 22408 4012 22448
rect 4052 22408 4061 22448
rect 3331 22324 3340 22364
rect 3380 22324 3532 22364
rect 3572 22324 3581 22364
rect 5059 22324 5068 22364
rect 5108 22324 5644 22364
rect 5684 22324 5693 22364
rect 163 22240 172 22280
rect 212 22240 556 22280
rect 596 22240 605 22280
rect 2659 22156 2668 22196
rect 2708 22156 5644 22196
rect 5684 22156 5932 22196
rect 5972 22156 6124 22196
rect 6164 22156 6173 22196
rect 3679 21904 3688 21944
rect 3728 21904 3770 21944
rect 3810 21904 3852 21944
rect 3892 21904 3934 21944
rect 3974 21904 4016 21944
rect 4056 21904 4065 21944
rect 10339 21736 10348 21776
rect 10388 21736 10732 21776
rect 10772 21736 10781 21776
rect 2083 21652 2092 21692
rect 2132 21652 2284 21692
rect 2324 21652 2333 21692
rect 4387 21652 4396 21692
rect 4436 21652 5068 21692
rect 5108 21652 5117 21692
rect 8237 21568 8332 21608
rect 8372 21568 8381 21608
rect 2179 21484 2188 21524
rect 2228 21484 5740 21524
rect 5780 21484 5789 21524
rect 1891 21400 1900 21440
rect 1940 21400 10348 21440
rect 10388 21400 10397 21440
rect 4919 21148 4928 21188
rect 4968 21148 5010 21188
rect 5050 21148 5092 21188
rect 5132 21148 5174 21188
rect 5214 21148 5256 21188
rect 5296 21148 5305 21188
rect 4771 20980 4780 21020
rect 4820 20980 4972 21020
rect 5012 20980 5021 21020
rect 6691 20980 6700 21020
rect 6740 20980 9292 21020
rect 9332 20980 9341 21020
rect 3907 20812 3916 20852
rect 3956 20812 4396 20852
rect 4436 20812 4876 20852
rect 4916 20812 4925 20852
rect 4387 20644 4396 20684
rect 4436 20644 4684 20684
rect 4724 20644 4733 20684
rect 5923 20644 5932 20684
rect 5972 20644 8908 20684
rect 8948 20644 8957 20684
rect 3679 20392 3688 20432
rect 3728 20392 3770 20432
rect 3810 20392 3852 20432
rect 3892 20392 3934 20432
rect 3974 20392 4016 20432
rect 4056 20392 4065 20432
rect 6691 20308 6700 20348
rect 6740 20308 7276 20348
rect 7316 20308 7325 20348
rect 2851 20224 2860 20264
rect 2900 20224 3148 20264
rect 3188 20224 3197 20264
rect 3244 20224 7564 20264
rect 7604 20224 7613 20264
rect 3244 20180 3284 20224
rect 1037 20140 1132 20180
rect 1172 20140 1181 20180
rect 2947 20140 2956 20180
rect 2996 20140 3284 20180
rect 3331 20140 3340 20180
rect 3380 20140 3475 20180
rect 3523 20140 3532 20180
rect 3572 20140 3667 20180
rect 7267 20140 7276 20180
rect 7316 20140 8524 20180
rect 8564 20140 8573 20180
rect 10051 20140 10060 20180
rect 10100 20140 10109 20180
rect 10060 20096 10100 20140
rect 1507 20056 1516 20096
rect 1556 20056 4012 20096
rect 4052 20056 4061 20096
rect 9379 20056 9388 20096
rect 9428 20056 10100 20096
rect 1795 19804 1804 19844
rect 1844 19804 3436 19844
rect 3476 19804 4204 19844
rect 4244 19804 4253 19844
rect 4771 19804 4780 19844
rect 4820 19804 4972 19844
rect 5012 19804 5021 19844
rect 5837 19720 5932 19760
rect 5972 19720 5981 19760
rect 4919 19636 4928 19676
rect 4968 19636 5010 19676
rect 5050 19636 5092 19676
rect 5132 19636 5174 19676
rect 5214 19636 5256 19676
rect 5296 19636 5305 19676
rect 6019 19636 6028 19676
rect 6068 19636 6412 19676
rect 6452 19636 6461 19676
rect 1987 19468 1996 19508
rect 2036 19468 5164 19508
rect 5204 19468 5213 19508
rect 931 19384 940 19424
rect 980 19384 3628 19424
rect 3668 19384 3677 19424
rect 4483 19384 4492 19424
rect 4532 19384 5548 19424
rect 5588 19384 5597 19424
rect 8707 19384 8716 19424
rect 8756 19384 8908 19424
rect 8948 19384 8957 19424
rect 1219 19300 1228 19340
rect 1268 19300 3724 19340
rect 3764 19300 3773 19340
rect 4483 19216 4492 19256
rect 4532 19216 4684 19256
rect 4724 19216 4733 19256
rect 7075 19216 7084 19256
rect 7124 19216 7468 19256
rect 7508 19216 8716 19256
rect 8756 19216 8765 19256
rect 3907 19048 3916 19088
rect 3956 19048 4492 19088
rect 4532 19048 4541 19088
rect 3679 18880 3688 18920
rect 3728 18880 3770 18920
rect 3810 18880 3852 18920
rect 3892 18880 3934 18920
rect 3974 18880 4016 18920
rect 4056 18880 4065 18920
rect 4291 18880 4300 18920
rect 4340 18880 8716 18920
rect 8756 18880 8765 18920
rect 6499 18796 6508 18836
rect 6548 18796 9964 18836
rect 10004 18796 10013 18836
rect 8803 18712 8812 18752
rect 8852 18712 10156 18752
rect 10196 18712 10205 18752
rect 1507 18628 1516 18668
rect 1556 18628 2092 18668
rect 2132 18628 2141 18668
rect 7843 18544 7852 18584
rect 7892 18544 8524 18584
rect 8564 18544 8573 18584
rect 10051 18544 10060 18584
rect 10100 18544 10540 18584
rect 10580 18544 10589 18584
rect 4579 18460 4588 18500
rect 4628 18460 7468 18500
rect 7508 18460 7517 18500
rect 5251 18292 5260 18332
rect 5300 18292 9388 18332
rect 9428 18292 9437 18332
rect 6403 18208 6412 18248
rect 6452 18208 6796 18248
rect 6836 18208 6845 18248
rect 10636 18208 10732 18248
rect 10772 18208 10781 18248
rect 4919 18124 4928 18164
rect 4968 18124 5010 18164
rect 5050 18124 5092 18164
rect 5132 18124 5174 18164
rect 5214 18124 5256 18164
rect 5296 18124 5305 18164
rect 6211 18124 6220 18164
rect 6260 18124 6269 18164
rect 9379 18124 9388 18164
rect 9428 18124 9964 18164
rect 10004 18124 10013 18164
rect 6220 18080 6260 18124
rect 6220 18040 6796 18080
rect 6836 18040 6845 18080
rect 3427 17956 3436 17996
rect 3476 17956 3532 17996
rect 3572 17956 3581 17996
rect 4771 17956 4780 17996
rect 4820 17956 5068 17996
rect 5108 17956 5117 17996
rect 6691 17956 6700 17996
rect 6740 17956 6988 17996
rect 7028 17956 7037 17996
rect 10636 17828 10676 18208
rect 10829 17956 10924 17996
rect 10964 17956 10973 17996
rect 11203 17956 11212 17996
rect 11252 17956 11500 17996
rect 11540 17956 11549 17996
rect 4685 17788 4780 17828
rect 4820 17788 4829 17828
rect 6307 17788 6316 17828
rect 6356 17788 6988 17828
rect 7028 17788 7037 17828
rect 10627 17788 10636 17828
rect 10676 17788 10685 17828
rect 2947 17620 2956 17660
rect 2996 17620 5932 17660
rect 5972 17620 8812 17660
rect 8852 17620 8861 17660
rect 8035 17452 8044 17492
rect 8084 17452 8140 17492
rect 8180 17452 8189 17492
rect 3679 17368 3688 17408
rect 3728 17368 3770 17408
rect 3810 17368 3852 17408
rect 3892 17368 3934 17408
rect 3974 17368 4016 17408
rect 4056 17368 4065 17408
rect 6787 17368 6796 17408
rect 6836 17368 7468 17408
rect 7508 17368 7517 17408
rect 3331 17200 3340 17240
rect 3380 17200 3820 17240
rect 3860 17200 3869 17240
rect 4771 17200 4780 17240
rect 4820 17200 4829 17240
rect 4780 17156 4820 17200
rect 3619 17116 3628 17156
rect 3668 17116 4820 17156
rect 4483 17032 4492 17072
rect 4532 17032 5740 17072
rect 5780 17032 5789 17072
rect 3715 16948 3724 16988
rect 3764 16948 4396 16988
rect 4436 16948 4445 16988
rect 4771 16948 4780 16988
rect 4820 16948 5164 16988
rect 5204 16948 5213 16988
rect 6019 16948 6028 16988
rect 6068 16948 7180 16988
rect 7220 16948 7229 16988
rect 4099 16864 4108 16904
rect 4148 16864 4972 16904
rect 5012 16864 5021 16904
rect 3907 16780 3916 16820
rect 3956 16780 5260 16820
rect 5300 16780 5309 16820
rect 5635 16780 5644 16820
rect 5684 16780 6220 16820
rect 6260 16780 6269 16820
rect 1603 16612 1612 16652
rect 1652 16612 2572 16652
rect 2612 16612 2621 16652
rect 4919 16612 4928 16652
rect 4968 16612 5010 16652
rect 5050 16612 5092 16652
rect 5132 16612 5174 16652
rect 5214 16612 5256 16652
rect 5296 16612 5305 16652
rect 3619 16444 3628 16484
rect 3668 16444 4972 16484
rect 5012 16444 5021 16484
rect 5347 16444 5356 16484
rect 5396 16444 5405 16484
rect 5356 16400 5396 16444
rect 4387 16360 4396 16400
rect 4436 16360 5396 16400
rect 2467 16276 2476 16316
rect 2516 16276 5740 16316
rect 5780 16276 5789 16316
rect 4195 16192 4204 16232
rect 4244 16192 4876 16232
rect 4916 16192 4925 16232
rect 3679 15856 3688 15896
rect 3728 15856 3770 15896
rect 3810 15856 3852 15896
rect 3892 15856 3934 15896
rect 3974 15856 4016 15896
rect 4056 15856 4065 15896
rect 2947 15772 2956 15812
rect 2996 15772 6220 15812
rect 6260 15772 6269 15812
rect 5731 15688 5740 15728
rect 5780 15688 10444 15728
rect 10484 15688 10493 15728
rect 4291 15604 4300 15644
rect 4340 15604 8236 15644
rect 8276 15604 8285 15644
rect 3811 15520 3820 15560
rect 3860 15520 5740 15560
rect 5780 15520 5789 15560
rect 4771 15436 4780 15476
rect 4820 15436 5260 15476
rect 5300 15436 5309 15476
rect 5443 15436 5452 15476
rect 5492 15436 6028 15476
rect 6068 15436 6077 15476
rect 2851 15268 2860 15308
rect 2900 15268 4300 15308
rect 4340 15268 4349 15308
rect 2947 15100 2956 15140
rect 2996 15100 3148 15140
rect 3188 15100 3197 15140
rect 4919 15100 4928 15140
rect 4968 15100 5010 15140
rect 5050 15100 5092 15140
rect 5132 15100 5174 15140
rect 5214 15100 5256 15140
rect 5296 15100 5305 15140
rect 1123 15016 1132 15056
rect 1172 15016 3052 15056
rect 3092 15016 7756 15056
rect 7796 15016 7805 15056
rect 2851 14932 2860 14972
rect 2900 14932 4588 14972
rect 4628 14932 4637 14972
rect 2755 14848 2764 14888
rect 2804 14848 2956 14888
rect 2996 14848 3005 14888
rect 4867 14848 4876 14888
rect 4916 14848 6220 14888
rect 6260 14848 6269 14888
rect 3715 14764 3724 14804
rect 3764 14764 4204 14804
rect 4244 14764 4253 14804
rect 2189 14680 2284 14720
rect 2324 14680 2333 14720
rect 2563 14680 2572 14720
rect 2612 14680 2764 14720
rect 2804 14680 2813 14720
rect 5539 14680 5548 14720
rect 5588 14680 5644 14720
rect 5684 14680 5693 14720
rect 5347 14596 5356 14636
rect 5396 14596 5932 14636
rect 5972 14596 5981 14636
rect 931 14512 940 14552
rect 980 14512 1228 14552
rect 1268 14512 1277 14552
rect 5740 14428 6892 14468
rect 6932 14428 6941 14468
rect 3679 14344 3688 14384
rect 3728 14344 3770 14384
rect 3810 14344 3852 14384
rect 3892 14344 3934 14384
rect 3974 14344 4016 14384
rect 4056 14344 4065 14384
rect 3619 13924 3628 13964
rect 3668 13924 4204 13964
rect 4244 13924 4253 13964
rect 5740 13880 5780 14428
rect 6883 14260 6892 14300
rect 6932 14260 7084 14300
rect 7124 14260 7133 14300
rect 7459 14092 7468 14132
rect 7508 14092 10540 14132
rect 10580 14092 10589 14132
rect 9485 14008 9580 14048
rect 9620 14008 9629 14048
rect 5731 13840 5740 13880
rect 5780 13840 5789 13880
rect 3043 13756 3052 13796
rect 3092 13756 3436 13796
rect 3476 13756 3485 13796
rect 9667 13672 9676 13712
rect 9716 13672 9964 13712
rect 10004 13672 10013 13712
rect 3427 13588 3436 13628
rect 3476 13588 3532 13628
rect 3572 13588 3581 13628
rect 4919 13588 4928 13628
rect 4968 13588 5010 13628
rect 5050 13588 5092 13628
rect 5132 13588 5174 13628
rect 5214 13588 5256 13628
rect 5296 13588 5305 13628
rect 9091 13588 9100 13628
rect 9140 13588 9484 13628
rect 9524 13588 9533 13628
rect 9379 13504 9388 13544
rect 9428 13504 9676 13544
rect 9716 13504 9725 13544
rect 5635 13168 5644 13208
rect 5684 13168 5740 13208
rect 5780 13168 5789 13208
rect 3043 13084 3052 13124
rect 3092 13084 3340 13124
rect 3380 13084 3389 13124
rect 5443 13084 5452 13124
rect 5492 13084 5836 13124
rect 5876 13084 5885 13124
rect 3139 13000 3148 13040
rect 3188 13000 3916 13040
rect 3956 13000 3965 13040
rect 3523 12916 3532 12956
rect 3572 12916 5108 12956
rect 2275 12832 2284 12872
rect 2324 12832 2764 12872
rect 2804 12832 2813 12872
rect 3679 12832 3688 12872
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 4056 12832 4065 12872
rect 4195 12832 4204 12872
rect 4244 12832 4339 12872
rect 5068 12788 5108 12916
rect 5635 12832 5644 12872
rect 5684 12832 5836 12872
rect 5876 12832 5885 12872
rect 3427 12748 3436 12788
rect 3476 12748 3532 12788
rect 3572 12748 3581 12788
rect 5068 12748 7084 12788
rect 7124 12748 7133 12788
rect 1795 12664 1804 12704
rect 1844 12664 1900 12704
rect 1940 12664 1949 12704
rect 1891 12496 1900 12536
rect 1940 12496 2572 12536
rect 2612 12496 2621 12536
rect 1123 12412 1132 12452
rect 1172 12412 1228 12452
rect 1268 12412 1277 12452
rect 3331 12244 3340 12284
rect 3380 12244 4492 12284
rect 4532 12244 4541 12284
rect 4919 12076 4928 12116
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 5296 12076 5305 12116
rect 2179 11908 2188 11948
rect 2228 11908 2860 11948
rect 2900 11908 2909 11948
rect 5443 11908 5452 11948
rect 5492 11908 5740 11948
rect 5780 11908 5789 11948
rect 7757 11908 7852 11948
rect 7892 11908 7901 11948
rect 4397 11824 4492 11864
rect 4532 11824 4541 11864
rect 5549 11740 5644 11780
rect 5684 11740 5693 11780
rect 3811 11656 3820 11696
rect 3860 11656 10252 11696
rect 10292 11656 10301 11696
rect 9283 11572 9292 11612
rect 9332 11572 10156 11612
rect 10196 11572 10205 11612
rect 1795 11488 1804 11528
rect 1844 11488 9868 11528
rect 9908 11488 9917 11528
rect 3679 11320 3688 11360
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 4056 11320 4065 11360
rect 1411 11236 1420 11276
rect 1460 11236 9676 11276
rect 9716 11236 9725 11276
rect 4003 11152 4012 11192
rect 4052 11152 4204 11192
rect 4244 11152 4253 11192
rect 1123 11068 1132 11108
rect 1172 11068 2476 11108
rect 2516 11068 2525 11108
rect 2765 11068 2860 11108
rect 2900 11068 2909 11108
rect 3811 10984 3820 11024
rect 3860 10984 6124 11024
rect 6164 10984 6173 11024
rect 4387 10732 4396 10772
rect 4436 10732 4492 10772
rect 4532 10732 4541 10772
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 4579 10228 4588 10268
rect 4628 10228 4780 10268
rect 4820 10228 4829 10268
rect 5539 10060 5548 10100
rect 5588 10060 6412 10100
rect 6452 10060 6461 10100
rect 10435 10060 10444 10100
rect 10484 10060 10924 10100
rect 10964 10060 10973 10100
rect 1709 9976 1804 10016
rect 1844 9976 1853 10016
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 1411 9472 1420 9512
rect 1460 9472 9484 9512
rect 9524 9472 9533 9512
rect 3811 9388 3820 9428
rect 3860 9388 7564 9428
rect 7604 9388 8332 9428
rect 8372 9388 8381 9428
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 2851 8884 2860 8924
rect 2900 8884 6508 8924
rect 6548 8884 6557 8924
rect 6979 8716 6988 8756
rect 7028 8716 7180 8756
rect 7220 8716 7229 8756
rect 2851 8632 2860 8672
rect 2900 8632 10156 8672
rect 10196 8632 10205 8672
rect 1603 8548 1612 8588
rect 1652 8548 3436 8588
rect 3476 8548 3485 8588
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 4579 7876 4588 7916
rect 4628 7876 5260 7916
rect 5300 7876 5309 7916
rect 3235 7792 3244 7832
rect 3284 7792 3436 7832
rect 3476 7792 3485 7832
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 3619 7372 3628 7412
rect 3668 7372 10348 7412
rect 10388 7372 10397 7412
rect 1315 7204 1324 7244
rect 1364 7204 1516 7244
rect 1556 7204 2284 7244
rect 2324 7204 2333 7244
rect 5635 7204 5644 7244
rect 5684 7204 5740 7244
rect 5780 7204 5789 7244
rect 3715 7120 3724 7160
rect 3764 7120 10060 7160
rect 10100 7120 10109 7160
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 3619 6616 3628 6656
rect 3668 6616 6220 6656
rect 6260 6616 6269 6656
rect 3523 6532 3532 6572
rect 3572 6532 3820 6572
rect 3860 6532 3869 6572
rect 1517 6448 1612 6488
rect 1652 6448 1661 6488
rect 9763 6448 9772 6488
rect 9812 6448 9964 6488
rect 10004 6448 10013 6488
rect 6211 6364 6220 6404
rect 6260 6364 6316 6404
rect 6356 6364 6365 6404
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 4579 5944 4588 5984
rect 4628 5944 7180 5984
rect 7220 5944 7229 5984
rect 4579 5860 4588 5900
rect 4628 5860 6700 5900
rect 6740 5860 6749 5900
rect 4099 5692 4108 5732
rect 4148 5692 4300 5732
rect 4340 5692 4349 5732
rect 8717 5692 8812 5732
rect 8852 5692 8861 5732
rect 3811 5440 3820 5480
rect 3860 5440 4972 5480
rect 5012 5440 5021 5480
rect 6403 5356 6412 5396
rect 6452 5356 6892 5396
rect 6932 5356 6941 5396
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 2083 4852 2092 4892
rect 2132 4852 4300 4892
rect 4340 4852 4349 4892
rect 4493 4852 4588 4892
rect 4628 4852 4637 4892
rect 4963 4852 4972 4892
rect 5012 4852 9100 4892
rect 9140 4852 9149 4892
rect 1891 4768 1900 4808
rect 1940 4768 8332 4808
rect 8372 4768 8381 4808
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 1805 4264 1900 4304
rect 1940 4264 1949 4304
rect 3331 4264 3340 4304
rect 3380 4264 6604 4304
rect 6644 4264 6653 4304
rect 4291 4096 4300 4136
rect 4340 4096 5548 4136
rect 5588 4096 5597 4136
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 4387 3508 4396 3548
rect 4436 3508 4445 3548
rect 2093 3424 2188 3464
rect 2228 3424 2237 3464
rect 4396 3296 4436 3508
rect 4396 3256 4588 3296
rect 4628 3256 4637 3296
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 2179 2836 2188 2876
rect 2228 2836 5548 2876
rect 5588 2836 5597 2876
rect 6499 2836 6508 2876
rect 6548 2836 7948 2876
rect 7988 2836 7997 2876
rect 2947 2752 2956 2792
rect 2996 2752 6796 2792
rect 6836 2752 6845 2792
rect 2477 2584 2572 2624
rect 2612 2584 2621 2624
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 3715 1912 3724 1952
rect 3764 1912 4684 1952
rect 4724 1912 4733 1952
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 7277 1408 7372 1448
rect 7412 1408 7421 1448
rect 8045 1408 8140 1448
rect 8180 1408 8189 1448
rect 2755 232 2764 272
rect 2804 232 6028 272
rect 6068 232 6077 272
<< via4 >>
rect 4928 45340 4968 45380
rect 5010 45340 5050 45380
rect 5092 45340 5132 45380
rect 5174 45340 5214 45380
rect 5256 45340 5296 45380
rect 3688 44584 3728 44624
rect 3770 44584 3810 44624
rect 3852 44584 3892 44624
rect 3934 44584 3974 44624
rect 4016 44584 4056 44624
rect 6412 44248 6452 44288
rect 4928 43828 4968 43868
rect 5010 43828 5050 43868
rect 5092 43828 5132 43868
rect 5174 43828 5214 43868
rect 5256 43828 5296 43868
rect 3688 43072 3728 43112
rect 3770 43072 3810 43112
rect 3852 43072 3892 43112
rect 3934 43072 3974 43112
rect 4016 43072 4056 43112
rect 6508 42988 6548 43028
rect 9772 42736 9812 42776
rect 10156 42736 10196 42776
rect 4588 42484 4628 42524
rect 4928 42316 4968 42356
rect 5010 42316 5050 42356
rect 5092 42316 5132 42356
rect 5174 42316 5214 42356
rect 5256 42316 5296 42356
rect 10348 41896 10388 41936
rect 3052 41812 3092 41852
rect 3688 41560 3728 41600
rect 3770 41560 3810 41600
rect 3852 41560 3892 41600
rect 3934 41560 3974 41600
rect 4016 41560 4056 41600
rect 1612 40972 1652 41012
rect 5740 40972 5780 41012
rect 4928 40804 4968 40844
rect 5010 40804 5050 40844
rect 5092 40804 5132 40844
rect 5174 40804 5214 40844
rect 5256 40804 5296 40844
rect 9964 40384 10004 40424
rect 3688 40048 3728 40088
rect 3770 40048 3810 40088
rect 3852 40048 3892 40088
rect 3934 40048 3974 40088
rect 4016 40048 4056 40088
rect 2956 39712 2996 39752
rect 7084 39712 7124 39752
rect 8524 39628 8564 39668
rect 2860 39460 2900 39500
rect 10444 39460 10484 39500
rect 4928 39292 4968 39332
rect 5010 39292 5050 39332
rect 5092 39292 5132 39332
rect 5174 39292 5214 39332
rect 5256 39292 5296 39332
rect 3436 38872 3476 38912
rect 5836 38872 5876 38912
rect 10252 38872 10292 38912
rect 3688 38536 3728 38576
rect 3770 38536 3810 38576
rect 3852 38536 3892 38576
rect 3934 38536 3974 38576
rect 4016 38536 4056 38576
rect 4928 37780 4968 37820
rect 5010 37780 5050 37820
rect 5092 37780 5132 37820
rect 5174 37780 5214 37820
rect 5256 37780 5296 37820
rect 3244 37612 3284 37652
rect 5452 37528 5492 37568
rect 7948 37444 7988 37484
rect 1516 37192 1556 37232
rect 3688 37024 3728 37064
rect 3770 37024 3810 37064
rect 3852 37024 3892 37064
rect 3934 37024 3974 37064
rect 4016 37024 4056 37064
rect 5548 36772 5588 36812
rect 7180 36688 7220 36728
rect 9580 36688 9620 36728
rect 2380 36604 2420 36644
rect 3532 36436 3572 36476
rect 9484 36436 9524 36476
rect 4928 36268 4968 36308
rect 5010 36268 5050 36308
rect 5092 36268 5132 36308
rect 5174 36268 5214 36308
rect 5256 36268 5296 36308
rect 3244 36016 3284 36056
rect 5548 35848 5588 35888
rect 3688 35512 3728 35552
rect 3770 35512 3810 35552
rect 3852 35512 3892 35552
rect 3934 35512 3974 35552
rect 4016 35512 4056 35552
rect 2284 35344 2324 35384
rect 2956 35260 2996 35300
rect 5644 34924 5684 34964
rect 4928 34756 4968 34796
rect 5010 34756 5050 34796
rect 5092 34756 5132 34796
rect 5174 34756 5214 34796
rect 5256 34756 5296 34796
rect 3688 34000 3728 34040
rect 3770 34000 3810 34040
rect 3852 34000 3892 34040
rect 3934 34000 3974 34040
rect 4016 34000 4056 34040
rect 7180 33496 7220 33536
rect 6700 33412 6740 33452
rect 4928 33244 4968 33284
rect 5010 33244 5050 33284
rect 5092 33244 5132 33284
rect 5174 33244 5214 33284
rect 5256 33244 5296 33284
rect 2380 33160 2420 33200
rect 1708 33076 1748 33116
rect 9100 32992 9140 33032
rect 6220 32824 6260 32864
rect 10060 32824 10100 32864
rect 7852 32656 7892 32696
rect 5644 32572 5684 32612
rect 3688 32488 3728 32528
rect 3770 32488 3810 32528
rect 3852 32488 3892 32528
rect 3934 32488 3974 32528
rect 4016 32488 4056 32528
rect 4684 31900 4724 31940
rect 5548 31900 5588 31940
rect 4928 31732 4968 31772
rect 5010 31732 5050 31772
rect 5092 31732 5132 31772
rect 5174 31732 5214 31772
rect 5256 31732 5296 31772
rect 7372 31732 7412 31772
rect 5548 31312 5588 31352
rect 1420 31228 1460 31268
rect 7564 31228 7604 31268
rect 3688 30976 3728 31016
rect 3770 30976 3810 31016
rect 3852 30976 3892 31016
rect 3934 30976 3974 31016
rect 4016 30976 4056 31016
rect 3532 30640 3572 30680
rect 7084 30640 7124 30680
rect 2956 30556 2996 30596
rect 9868 30388 9908 30428
rect 4928 30220 4968 30260
rect 5010 30220 5050 30260
rect 5092 30220 5132 30260
rect 5174 30220 5214 30260
rect 5256 30220 5296 30260
rect 1420 29968 1460 30008
rect 4780 29968 4820 30008
rect 5644 29884 5684 29924
rect 8236 29800 8276 29840
rect 8716 29800 8756 29840
rect 4396 29716 4436 29756
rect 4204 29632 4244 29672
rect 3688 29464 3728 29504
rect 3770 29464 3810 29504
rect 3852 29464 3892 29504
rect 3934 29464 3974 29504
rect 4016 29464 4056 29504
rect 1612 29128 1652 29168
rect 6796 28876 6836 28916
rect 9676 28876 9716 28916
rect 1708 28792 1748 28832
rect 2764 28708 2804 28748
rect 4928 28708 4968 28748
rect 5010 28708 5050 28748
rect 5092 28708 5132 28748
rect 5174 28708 5214 28748
rect 5256 28708 5296 28748
rect 2572 28624 2612 28664
rect 9100 28372 9140 28412
rect 6604 28288 6644 28328
rect 9100 28204 9140 28244
rect 3244 28120 3284 28160
rect 3688 27952 3728 27992
rect 3770 27952 3810 27992
rect 3852 27952 3892 27992
rect 3934 27952 3974 27992
rect 4016 27952 4056 27992
rect 6700 27868 6740 27908
rect 2956 27532 2996 27572
rect 4928 27196 4968 27236
rect 5010 27196 5050 27236
rect 5092 27196 5132 27236
rect 5174 27196 5214 27236
rect 5256 27196 5296 27236
rect 5644 27112 5684 27152
rect 9772 26944 9812 26984
rect 1612 26692 1652 26732
rect 3688 26440 3728 26480
rect 3770 26440 3810 26480
rect 3852 26440 3892 26480
rect 3934 26440 3974 26480
rect 4016 26440 4056 26480
rect 4780 26020 4820 26060
rect 7660 25852 7700 25892
rect 4928 25684 4968 25724
rect 5010 25684 5050 25724
rect 5092 25684 5132 25724
rect 5174 25684 5214 25724
rect 5256 25684 5296 25724
rect 5644 25516 5684 25556
rect 4396 25348 4436 25388
rect 3688 24928 3728 24968
rect 3770 24928 3810 24968
rect 3852 24928 3892 24968
rect 3934 24928 3974 24968
rect 4016 24928 4056 24968
rect 8140 24424 8180 24464
rect 3532 24340 3572 24380
rect 4928 24172 4968 24212
rect 5010 24172 5050 24212
rect 5092 24172 5132 24212
rect 5174 24172 5214 24212
rect 5256 24172 5296 24212
rect 6316 23836 6356 23876
rect 3688 23416 3728 23456
rect 3770 23416 3810 23456
rect 3852 23416 3892 23456
rect 3934 23416 3974 23456
rect 4016 23416 4056 23456
rect 9772 23416 9812 23456
rect 3244 23248 3284 23288
rect 4204 23080 4244 23120
rect 4780 23080 4820 23120
rect 7660 23080 7700 23120
rect 3340 22996 3380 23036
rect 3244 22912 3284 22952
rect 5932 22912 5972 22952
rect 3148 22828 3188 22868
rect 4396 22744 4436 22784
rect 4928 22660 4968 22700
rect 5010 22660 5050 22700
rect 5092 22660 5132 22700
rect 5174 22660 5214 22700
rect 5256 22660 5296 22700
rect 6508 22492 6548 22532
rect 8044 22492 8084 22532
rect 3340 22324 3380 22364
rect 5644 22324 5684 22364
rect 5644 22156 5684 22196
rect 3688 21904 3728 21944
rect 3770 21904 3810 21944
rect 3852 21904 3892 21944
rect 3934 21904 3974 21944
rect 4016 21904 4056 21944
rect 4396 21652 4436 21692
rect 8332 21568 8372 21608
rect 2188 21484 2228 21524
rect 1900 21400 1940 21440
rect 4928 21148 4968 21188
rect 5010 21148 5050 21188
rect 5092 21148 5132 21188
rect 5174 21148 5214 21188
rect 5256 21148 5296 21188
rect 4780 20980 4820 21020
rect 9292 20980 9332 21020
rect 4396 20644 4436 20684
rect 5932 20644 5972 20684
rect 3688 20392 3728 20432
rect 3770 20392 3810 20432
rect 3852 20392 3892 20432
rect 3934 20392 3974 20432
rect 4016 20392 4056 20432
rect 3148 20224 3188 20264
rect 7564 20224 7604 20264
rect 1132 20140 1172 20180
rect 2956 20140 2996 20180
rect 3340 20140 3380 20180
rect 3532 20140 3572 20180
rect 8524 20140 8564 20180
rect 9388 20056 9428 20096
rect 4204 19804 4244 19844
rect 4780 19804 4820 19844
rect 5932 19720 5972 19760
rect 4928 19636 4968 19676
rect 5010 19636 5050 19676
rect 5092 19636 5132 19676
rect 5174 19636 5214 19676
rect 5256 19636 5296 19676
rect 7084 19216 7124 19256
rect 4492 19048 4532 19088
rect 3688 18880 3728 18920
rect 3770 18880 3810 18920
rect 3852 18880 3892 18920
rect 3934 18880 3974 18920
rect 4016 18880 4056 18920
rect 4300 18880 4340 18920
rect 8716 18880 8756 18920
rect 6508 18796 6548 18836
rect 9964 18796 10004 18836
rect 8812 18712 8852 18752
rect 4588 18460 4628 18500
rect 7468 18460 7508 18500
rect 9388 18292 9428 18332
rect 4928 18124 4968 18164
rect 5010 18124 5050 18164
rect 5092 18124 5132 18164
rect 5174 18124 5214 18164
rect 5256 18124 5296 18164
rect 3532 17956 3572 17996
rect 4780 17956 4820 17996
rect 10924 17956 10964 17996
rect 4780 17788 4820 17828
rect 8044 17452 8084 17492
rect 3688 17368 3728 17408
rect 3770 17368 3810 17408
rect 3852 17368 3892 17408
rect 3934 17368 3974 17408
rect 4016 17368 4056 17408
rect 4492 17032 4532 17072
rect 6028 16948 6068 16988
rect 5644 16780 5684 16820
rect 4928 16612 4968 16652
rect 5010 16612 5050 16652
rect 5092 16612 5132 16652
rect 5174 16612 5214 16652
rect 5256 16612 5296 16652
rect 4204 16192 4244 16232
rect 3688 15856 3728 15896
rect 3770 15856 3810 15896
rect 3852 15856 3892 15896
rect 3934 15856 3974 15896
rect 4016 15856 4056 15896
rect 6220 15772 6260 15812
rect 10444 15688 10484 15728
rect 8236 15604 8276 15644
rect 5740 15520 5780 15560
rect 4780 15436 4820 15476
rect 5452 15436 5492 15476
rect 2860 15268 2900 15308
rect 2956 15100 2996 15140
rect 4928 15100 4968 15140
rect 5010 15100 5050 15140
rect 5092 15100 5132 15140
rect 5174 15100 5214 15140
rect 5256 15100 5296 15140
rect 4588 14932 4628 14972
rect 4204 14764 4244 14804
rect 2284 14680 2324 14720
rect 5644 14680 5684 14720
rect 3688 14344 3728 14384
rect 3770 14344 3810 14384
rect 3852 14344 3892 14384
rect 3934 14344 3974 14384
rect 4016 14344 4056 14384
rect 4204 13924 4244 13964
rect 7468 14092 7508 14132
rect 9580 14008 9620 14048
rect 3532 13588 3572 13628
rect 4928 13588 4968 13628
rect 5010 13588 5050 13628
rect 5092 13588 5132 13628
rect 5174 13588 5214 13628
rect 5256 13588 5296 13628
rect 9388 13504 9428 13544
rect 5740 13168 5780 13208
rect 3052 13084 3092 13124
rect 5836 13084 5876 13124
rect 3148 13000 3188 13040
rect 3688 12832 3728 12872
rect 3770 12832 3810 12872
rect 3852 12832 3892 12872
rect 3934 12832 3974 12872
rect 4016 12832 4056 12872
rect 4204 12832 4244 12872
rect 5836 12832 5876 12872
rect 3532 12748 3572 12788
rect 1804 12664 1844 12704
rect 1132 12412 1172 12452
rect 4492 12244 4532 12284
rect 4928 12076 4968 12116
rect 5010 12076 5050 12116
rect 5092 12076 5132 12116
rect 5174 12076 5214 12116
rect 5256 12076 5296 12116
rect 7852 11908 7892 11948
rect 4492 11824 4532 11864
rect 5644 11740 5684 11780
rect 10252 11656 10292 11696
rect 9292 11572 9332 11612
rect 9868 11488 9908 11528
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 9676 11236 9716 11276
rect 4204 11152 4244 11192
rect 1132 11068 1172 11108
rect 2860 11068 2900 11108
rect 6124 10984 6164 11024
rect 4492 10732 4532 10772
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 4780 10228 4820 10268
rect 6412 10060 6452 10100
rect 10924 10060 10964 10100
rect 1804 9976 1844 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 9484 9472 9524 9512
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 6508 8884 6548 8924
rect 10156 8632 10196 8672
rect 3436 8548 3476 8588
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 4588 7876 4628 7916
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 10348 7372 10388 7412
rect 1516 7204 1556 7244
rect 5740 7204 5780 7244
rect 10060 7120 10100 7160
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 3532 6532 3572 6572
rect 1612 6448 1652 6488
rect 9772 6448 9812 6488
rect 6316 6364 6356 6404
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 4588 5860 4628 5900
rect 8812 5692 8852 5732
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 4300 4852 4340 4892
rect 4588 4852 4628 4892
rect 9100 4852 9140 4892
rect 8332 4768 8372 4808
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 1900 4264 1940 4304
rect 6604 4264 6644 4304
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 2188 3424 2228 3464
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 5548 2836 5588 2876
rect 7948 2836 7988 2876
rect 6796 2752 6836 2792
rect 2572 2584 2612 2624
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 4684 1912 4724 1952
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 7372 1408 7412 1448
rect 8140 1408 8180 1448
rect 6028 232 6068 272
<< metal5 >>
rect 3652 44624 4092 47360
rect 3652 44584 3688 44624
rect 3728 44584 3770 44624
rect 3810 44584 3852 44624
rect 3892 44584 3934 44624
rect 3974 44584 4016 44624
rect 4056 44584 4092 44624
rect 3652 43112 4092 44584
rect 3652 43072 3688 43112
rect 3728 43072 3770 43112
rect 3810 43072 3852 43112
rect 3892 43072 3934 43112
rect 3974 43072 4016 43112
rect 4056 43072 4092 43112
rect 3052 41852 3092 41861
rect 1612 41012 1652 41021
rect 1516 37232 1556 37241
rect 1420 31268 1460 31277
rect 1420 30008 1460 31228
rect 1420 29959 1460 29968
rect 1132 20180 1172 20189
rect 1132 12452 1172 20140
rect 1132 11108 1172 12412
rect 1132 11059 1172 11068
rect 1516 7244 1556 37192
rect 1612 29168 1652 40972
rect 2956 39752 2996 39761
rect 2764 39500 2900 39528
rect 2764 39488 2860 39500
rect 2380 36644 2420 36653
rect 2284 35384 2324 35393
rect 1612 29119 1652 29128
rect 1708 33116 1748 33125
rect 1708 28832 1748 33076
rect 1708 28783 1748 28792
rect 1516 7195 1556 7204
rect 1612 26732 1652 26741
rect 1612 6488 1652 26692
rect 2188 21524 2228 21533
rect 1900 21440 1940 21449
rect 1804 12704 1844 12713
rect 1804 10016 1844 12664
rect 1804 9967 1844 9976
rect 1612 6439 1652 6448
rect 1900 4304 1940 21400
rect 1900 4255 1940 4264
rect 2188 3464 2228 21484
rect 2284 14720 2324 35344
rect 2380 33200 2420 36604
rect 2380 33151 2420 33160
rect 2764 28748 2804 39488
rect 2860 39451 2900 39460
rect 2956 35300 2996 39712
rect 2956 35251 2996 35260
rect 2764 28699 2804 28708
rect 2956 30596 2996 30605
rect 2284 14671 2324 14680
rect 2572 28664 2612 28673
rect 2188 3415 2228 3424
rect 2572 2624 2612 28624
rect 2956 27572 2996 30556
rect 2956 27523 2996 27532
rect 2956 20180 2996 20189
rect 2860 15308 2900 15317
rect 2860 11108 2900 15268
rect 2956 15140 2996 20140
rect 2956 15091 2996 15100
rect 3052 13124 3092 41812
rect 3652 41600 4092 43072
rect 4892 45380 5332 47360
rect 4892 45340 4928 45380
rect 4968 45340 5010 45380
rect 5050 45340 5092 45380
rect 5132 45340 5174 45380
rect 5214 45340 5256 45380
rect 5296 45340 5332 45380
rect 4892 43868 5332 45340
rect 4892 43828 4928 43868
rect 4968 43828 5010 43868
rect 5050 43828 5092 43868
rect 5132 43828 5174 43868
rect 5214 43828 5256 43868
rect 5296 43828 5332 43868
rect 3652 41560 3688 41600
rect 3728 41560 3770 41600
rect 3810 41560 3852 41600
rect 3892 41560 3934 41600
rect 3974 41560 4016 41600
rect 4056 41560 4092 41600
rect 3652 40088 4092 41560
rect 3652 40048 3688 40088
rect 3728 40048 3770 40088
rect 3810 40048 3852 40088
rect 3892 40048 3934 40088
rect 3974 40048 4016 40088
rect 4056 40048 4092 40088
rect 3436 38912 3476 38921
rect 3244 37652 3284 37661
rect 3244 36056 3284 37612
rect 3244 36007 3284 36016
rect 3244 28160 3284 28169
rect 3244 23288 3284 28120
rect 3244 23239 3284 23248
rect 3340 23036 3380 23045
rect 3244 22952 3284 22961
rect 3052 13075 3092 13084
rect 3148 22868 3188 22877
rect 3148 20264 3188 22828
rect 3148 13040 3188 20224
rect 3244 20180 3284 22912
rect 3340 22364 3380 22996
rect 3340 22315 3380 22324
rect 3340 20180 3380 20189
rect 3244 20140 3340 20180
rect 3340 20131 3380 20140
rect 3148 12991 3188 13000
rect 2860 11059 2900 11068
rect 3436 8588 3476 38872
rect 3652 38576 4092 40048
rect 3652 38536 3688 38576
rect 3728 38536 3770 38576
rect 3810 38536 3852 38576
rect 3892 38536 3934 38576
rect 3974 38536 4016 38576
rect 4056 38536 4092 38576
rect 3652 37064 4092 38536
rect 3652 37024 3688 37064
rect 3728 37024 3770 37064
rect 3810 37024 3852 37064
rect 3892 37024 3934 37064
rect 3974 37024 4016 37064
rect 4056 37024 4092 37064
rect 3532 36476 3572 36485
rect 3532 30680 3572 36436
rect 3532 30631 3572 30640
rect 3652 35552 4092 37024
rect 3652 35512 3688 35552
rect 3728 35512 3770 35552
rect 3810 35512 3852 35552
rect 3892 35512 3934 35552
rect 3974 35512 4016 35552
rect 4056 35512 4092 35552
rect 3652 34040 4092 35512
rect 3652 34000 3688 34040
rect 3728 34000 3770 34040
rect 3810 34000 3852 34040
rect 3892 34000 3934 34040
rect 3974 34000 4016 34040
rect 4056 34000 4092 34040
rect 3652 32528 4092 34000
rect 3652 32488 3688 32528
rect 3728 32488 3770 32528
rect 3810 32488 3852 32528
rect 3892 32488 3934 32528
rect 3974 32488 4016 32528
rect 4056 32488 4092 32528
rect 3652 31016 4092 32488
rect 3652 30976 3688 31016
rect 3728 30976 3770 31016
rect 3810 30976 3852 31016
rect 3892 30976 3934 31016
rect 3974 30976 4016 31016
rect 4056 30976 4092 31016
rect 3652 29504 4092 30976
rect 4588 42524 4628 42533
rect 4396 29756 4436 29765
rect 3652 29464 3688 29504
rect 3728 29464 3770 29504
rect 3810 29464 3852 29504
rect 3892 29464 3934 29504
rect 3974 29464 4016 29504
rect 4056 29464 4092 29504
rect 3652 27992 4092 29464
rect 3652 27952 3688 27992
rect 3728 27952 3770 27992
rect 3810 27952 3852 27992
rect 3892 27952 3934 27992
rect 3974 27952 4016 27992
rect 4056 27952 4092 27992
rect 3652 26480 4092 27952
rect 3652 26440 3688 26480
rect 3728 26440 3770 26480
rect 3810 26440 3852 26480
rect 3892 26440 3934 26480
rect 3974 26440 4016 26480
rect 4056 26440 4092 26480
rect 3652 24968 4092 26440
rect 3652 24928 3688 24968
rect 3728 24928 3770 24968
rect 3810 24928 3852 24968
rect 3892 24928 3934 24968
rect 3974 24928 4016 24968
rect 4056 24928 4092 24968
rect 3532 24380 3572 24389
rect 3532 20180 3572 24340
rect 3532 20131 3572 20140
rect 3652 23456 4092 24928
rect 3652 23416 3688 23456
rect 3728 23416 3770 23456
rect 3810 23416 3852 23456
rect 3892 23416 3934 23456
rect 3974 23416 4016 23456
rect 4056 23416 4092 23456
rect 3652 21944 4092 23416
rect 4204 29672 4244 29681
rect 4204 23120 4244 29632
rect 4204 23071 4244 23080
rect 4396 25388 4436 29716
rect 3652 21904 3688 21944
rect 3728 21904 3770 21944
rect 3810 21904 3852 21944
rect 3892 21904 3934 21944
rect 3974 21904 4016 21944
rect 4056 21904 4092 21944
rect 3652 20432 4092 21904
rect 4396 22784 4436 25348
rect 4396 21692 4436 22744
rect 4396 20684 4436 21652
rect 4396 20635 4436 20644
rect 3652 20392 3688 20432
rect 3728 20392 3770 20432
rect 3810 20392 3852 20432
rect 3892 20392 3934 20432
rect 3974 20392 4016 20432
rect 4056 20392 4092 20432
rect 3652 18920 4092 20392
rect 3652 18880 3688 18920
rect 3728 18880 3770 18920
rect 3810 18880 3852 18920
rect 3892 18880 3934 18920
rect 3974 18880 4016 18920
rect 4056 18880 4092 18920
rect 3532 17996 3572 18005
rect 3532 13628 3572 17956
rect 3532 13579 3572 13588
rect 3652 17408 4092 18880
rect 3652 17368 3688 17408
rect 3728 17368 3770 17408
rect 3810 17368 3852 17408
rect 3892 17368 3934 17408
rect 3974 17368 4016 17408
rect 4056 17368 4092 17408
rect 3652 15896 4092 17368
rect 3652 15856 3688 15896
rect 3728 15856 3770 15896
rect 3810 15856 3852 15896
rect 3892 15856 3934 15896
rect 3974 15856 4016 15896
rect 4056 15856 4092 15896
rect 3652 14384 4092 15856
rect 3652 14344 3688 14384
rect 3728 14344 3770 14384
rect 3810 14344 3852 14384
rect 3892 14344 3934 14384
rect 3974 14344 4016 14384
rect 4056 14344 4092 14384
rect 3652 12872 4092 14344
rect 4204 19844 4244 19853
rect 4204 16232 4244 19804
rect 4492 19088 4532 19097
rect 4300 18920 4340 18929
rect 4300 18096 4340 18880
rect 4300 18056 4436 18096
rect 4204 14804 4244 16192
rect 4396 15816 4436 18056
rect 4204 13964 4244 14764
rect 4204 13915 4244 13924
rect 4300 15776 4436 15816
rect 4492 17072 4532 19048
rect 4588 18500 4628 42484
rect 4892 42356 5332 43828
rect 4892 42316 4928 42356
rect 4968 42316 5010 42356
rect 5050 42316 5092 42356
rect 5132 42316 5174 42356
rect 5214 42316 5256 42356
rect 5296 42316 5332 42356
rect 4892 40844 5332 42316
rect 6412 44288 6452 44297
rect 4892 40804 4928 40844
rect 4968 40804 5010 40844
rect 5050 40804 5092 40844
rect 5132 40804 5174 40844
rect 5214 40804 5256 40844
rect 5296 40804 5332 40844
rect 4892 39332 5332 40804
rect 4892 39292 4928 39332
rect 4968 39292 5010 39332
rect 5050 39292 5092 39332
rect 5132 39292 5174 39332
rect 5214 39292 5256 39332
rect 5296 39292 5332 39332
rect 4892 37820 5332 39292
rect 4892 37780 4928 37820
rect 4968 37780 5010 37820
rect 5050 37780 5092 37820
rect 5132 37780 5174 37820
rect 5214 37780 5256 37820
rect 5296 37780 5332 37820
rect 4892 36308 5332 37780
rect 5740 41012 5780 41021
rect 4892 36268 4928 36308
rect 4968 36268 5010 36308
rect 5050 36268 5092 36308
rect 5132 36268 5174 36308
rect 5214 36268 5256 36308
rect 5296 36268 5332 36308
rect 4892 34796 5332 36268
rect 4892 34756 4928 34796
rect 4968 34756 5010 34796
rect 5050 34756 5092 34796
rect 5132 34756 5174 34796
rect 5214 34756 5256 34796
rect 5296 34756 5332 34796
rect 4892 33284 5332 34756
rect 4892 33244 4928 33284
rect 4968 33244 5010 33284
rect 5050 33244 5092 33284
rect 5132 33244 5174 33284
rect 5214 33244 5256 33284
rect 5296 33244 5332 33284
rect 4588 18451 4628 18460
rect 4684 31940 4724 31949
rect 3652 12832 3688 12872
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 4056 12832 4092 12872
rect 3436 8539 3476 8548
rect 3532 12788 3572 12797
rect 3532 6572 3572 12748
rect 3532 6523 3572 6532
rect 3652 11360 4092 12832
rect 3652 11320 3688 11360
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 4056 11320 4092 11360
rect 3652 9848 4092 11320
rect 4204 12872 4244 12881
rect 4204 11192 4244 12832
rect 4204 11143 4244 11152
rect 3652 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4092 9848
rect 3652 8336 4092 9808
rect 3652 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4092 8336
rect 3652 6824 4092 8296
rect 3652 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4092 6824
rect 2572 2575 2612 2584
rect 3652 5312 4092 6784
rect 3652 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4092 5312
rect 3652 3800 4092 5272
rect 4300 4892 4340 15776
rect 4492 12284 4532 17032
rect 4492 12235 4532 12244
rect 4588 14972 4628 14981
rect 4492 11864 4532 11873
rect 4492 10772 4532 11824
rect 4492 10723 4532 10732
rect 4300 4843 4340 4852
rect 4588 7916 4628 14932
rect 4588 5900 4628 7876
rect 4588 4892 4628 5860
rect 4588 4843 4628 4852
rect 3652 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4092 3800
rect 3652 2288 4092 3760
rect 3652 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4092 2288
rect 3652 0 4092 2248
rect 4684 1952 4724 31900
rect 4892 31772 5332 33244
rect 4892 31732 4928 31772
rect 4968 31732 5010 31772
rect 5050 31732 5092 31772
rect 5132 31732 5174 31772
rect 5214 31732 5256 31772
rect 5296 31732 5332 31772
rect 4892 30260 5332 31732
rect 4892 30220 4928 30260
rect 4968 30220 5010 30260
rect 5050 30220 5092 30260
rect 5132 30220 5174 30260
rect 5214 30220 5256 30260
rect 5296 30220 5332 30260
rect 4780 30008 4820 30017
rect 4780 26060 4820 29968
rect 4780 23120 4820 26020
rect 4780 21020 4820 23080
rect 4780 20971 4820 20980
rect 4892 28748 5332 30220
rect 4892 28708 4928 28748
rect 4968 28708 5010 28748
rect 5050 28708 5092 28748
rect 5132 28708 5174 28748
rect 5214 28708 5256 28748
rect 5296 28708 5332 28748
rect 4892 27236 5332 28708
rect 4892 27196 4928 27236
rect 4968 27196 5010 27236
rect 5050 27196 5092 27236
rect 5132 27196 5174 27236
rect 5214 27196 5256 27236
rect 5296 27196 5332 27236
rect 4892 25724 5332 27196
rect 4892 25684 4928 25724
rect 4968 25684 5010 25724
rect 5050 25684 5092 25724
rect 5132 25684 5174 25724
rect 5214 25684 5256 25724
rect 5296 25684 5332 25724
rect 4892 24212 5332 25684
rect 4892 24172 4928 24212
rect 4968 24172 5010 24212
rect 5050 24172 5092 24212
rect 5132 24172 5174 24212
rect 5214 24172 5256 24212
rect 5296 24172 5332 24212
rect 4892 22700 5332 24172
rect 4892 22660 4928 22700
rect 4968 22660 5010 22700
rect 5050 22660 5092 22700
rect 5132 22660 5174 22700
rect 5214 22660 5256 22700
rect 5296 22660 5332 22700
rect 4892 21188 5332 22660
rect 4892 21148 4928 21188
rect 4968 21148 5010 21188
rect 5050 21148 5092 21188
rect 5132 21148 5174 21188
rect 5214 21148 5256 21188
rect 5296 21148 5332 21188
rect 4780 19844 4820 19853
rect 4780 17996 4820 19804
rect 4780 17947 4820 17956
rect 4892 19676 5332 21148
rect 4892 19636 4928 19676
rect 4968 19636 5010 19676
rect 5050 19636 5092 19676
rect 5132 19636 5174 19676
rect 5214 19636 5256 19676
rect 5296 19636 5332 19676
rect 4892 18164 5332 19636
rect 4892 18124 4928 18164
rect 4968 18124 5010 18164
rect 5050 18124 5092 18164
rect 5132 18124 5174 18164
rect 5214 18124 5256 18164
rect 5296 18124 5332 18164
rect 4780 17828 4820 17837
rect 4780 15476 4820 17788
rect 4780 10268 4820 15436
rect 4780 10219 4820 10228
rect 4892 16652 5332 18124
rect 4892 16612 4928 16652
rect 4968 16612 5010 16652
rect 5050 16612 5092 16652
rect 5132 16612 5174 16652
rect 5214 16612 5256 16652
rect 5296 16612 5332 16652
rect 4892 15140 5332 16612
rect 5452 37568 5492 37577
rect 5452 15476 5492 37528
rect 5548 36812 5588 36821
rect 5548 35888 5588 36772
rect 5548 31940 5588 35848
rect 5644 34964 5684 34973
rect 5644 32612 5684 34924
rect 5644 32563 5684 32572
rect 5548 31891 5588 31900
rect 5452 15427 5492 15436
rect 5548 31352 5588 31361
rect 4892 15100 4928 15140
rect 4968 15100 5010 15140
rect 5050 15100 5092 15140
rect 5132 15100 5174 15140
rect 5214 15100 5256 15140
rect 5296 15100 5332 15140
rect 4892 13628 5332 15100
rect 4892 13588 4928 13628
rect 4968 13588 5010 13628
rect 5050 13588 5092 13628
rect 5132 13588 5174 13628
rect 5214 13588 5256 13628
rect 5296 13588 5332 13628
rect 4892 12116 5332 13588
rect 4892 12076 4928 12116
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 5296 12076 5332 12116
rect 4892 10604 5332 12076
rect 4892 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5332 10604
rect 4684 1903 4724 1912
rect 4892 9092 5332 10564
rect 4892 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5332 9092
rect 4892 7580 5332 9052
rect 4892 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5332 7580
rect 4892 6068 5332 7540
rect 4892 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5332 6068
rect 4892 4556 5332 6028
rect 4892 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5332 4556
rect 4892 3044 5332 4516
rect 4892 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5332 3044
rect 4892 1532 5332 3004
rect 5548 2876 5588 31312
rect 5644 29924 5684 29933
rect 5644 27152 5684 29884
rect 5644 27103 5684 27112
rect 5644 25556 5684 25565
rect 5644 22364 5684 25516
rect 5644 22315 5684 22324
rect 5644 22196 5684 22205
rect 5644 16820 5684 22156
rect 5644 16771 5684 16780
rect 5740 15560 5780 40972
rect 5836 38912 5876 38921
rect 5836 18096 5876 38872
rect 6220 32864 6260 32873
rect 5932 22952 5972 22961
rect 5932 20684 5972 22912
rect 5932 19760 5972 20644
rect 5932 19711 5972 19720
rect 5836 18056 6164 18096
rect 5740 15511 5780 15520
rect 6028 16988 6068 16997
rect 5644 14720 5684 14729
rect 5644 11780 5684 14680
rect 5644 11731 5684 11740
rect 5740 13208 5780 13217
rect 5740 7244 5780 13168
rect 5836 13124 5876 13133
rect 5836 12872 5876 13084
rect 5836 12823 5876 12832
rect 5740 7195 5780 7204
rect 5548 2827 5588 2836
rect 4892 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5332 1532
rect 4892 0 5332 1492
rect 6028 272 6068 16948
rect 6124 11024 6164 18056
rect 6220 15812 6260 32824
rect 6220 15763 6260 15772
rect 6316 23876 6356 23885
rect 6124 10975 6164 10984
rect 6316 6404 6356 23836
rect 6412 10100 6452 44248
rect 6508 43028 6548 43037
rect 6508 22532 6548 42988
rect 9772 42776 9812 42785
rect 7084 39752 7124 39761
rect 6700 33452 6740 33461
rect 6508 22483 6548 22492
rect 6604 28328 6644 28337
rect 6412 10051 6452 10060
rect 6508 18836 6548 18845
rect 6508 8924 6548 18796
rect 6508 8875 6548 8884
rect 6316 6355 6356 6364
rect 6604 4304 6644 28288
rect 6700 27908 6740 33412
rect 7084 30680 7124 39712
rect 8524 39668 8564 39677
rect 7948 37484 7988 37493
rect 7180 36728 7220 36737
rect 7180 33536 7220 36688
rect 7180 33487 7220 33496
rect 7852 32696 7892 32705
rect 6700 27859 6740 27868
rect 6796 28916 6836 28925
rect 6604 4255 6644 4264
rect 6796 2792 6836 28876
rect 7084 19256 7124 30640
rect 7084 19207 7124 19216
rect 7372 31772 7412 31781
rect 6796 2743 6836 2752
rect 7372 1448 7412 31732
rect 7564 31268 7604 31277
rect 7564 20264 7604 31228
rect 7660 25892 7700 25901
rect 7660 23120 7700 25852
rect 7660 23071 7700 23080
rect 7564 20215 7604 20224
rect 7468 18500 7508 18509
rect 7468 14132 7508 18460
rect 7468 14083 7508 14092
rect 7852 11948 7892 32656
rect 7852 11899 7892 11908
rect 7948 2876 7988 37444
rect 8236 29840 8276 29849
rect 8140 24464 8180 24473
rect 8044 22532 8084 22541
rect 8044 17492 8084 22492
rect 8044 17443 8084 17452
rect 7948 2827 7988 2836
rect 7372 1399 7412 1408
rect 8140 1448 8180 24424
rect 8236 15644 8276 29800
rect 8236 15595 8276 15604
rect 8332 21608 8372 21617
rect 8332 4808 8372 21568
rect 8524 20180 8564 39628
rect 9580 36728 9620 36737
rect 9484 36476 9524 36485
rect 9100 33032 9140 33041
rect 8524 20131 8564 20140
rect 8716 29840 8756 29849
rect 8716 18920 8756 29800
rect 9100 28412 9140 32992
rect 9100 28363 9140 28372
rect 8716 18871 8756 18880
rect 9100 28244 9140 28253
rect 8812 18752 8852 18761
rect 8812 5732 8852 18712
rect 8812 5683 8852 5692
rect 9100 4892 9140 28204
rect 9292 21020 9332 21029
rect 9292 11612 9332 20980
rect 9388 20096 9428 20105
rect 9388 18332 9428 20056
rect 9388 13544 9428 18292
rect 9388 13495 9428 13504
rect 9292 11563 9332 11572
rect 9484 9512 9524 36436
rect 9580 14048 9620 36688
rect 9580 13999 9620 14008
rect 9676 28916 9716 28925
rect 9676 11276 9716 28876
rect 9772 26984 9812 42736
rect 10156 42776 10196 42785
rect 9964 40424 10004 40433
rect 9772 26935 9812 26944
rect 9868 30428 9908 30437
rect 9676 11227 9716 11236
rect 9772 23456 9812 23465
rect 9484 9463 9524 9472
rect 9772 6488 9812 23416
rect 9868 11528 9908 30388
rect 9964 18836 10004 40384
rect 9964 18787 10004 18796
rect 10060 32864 10100 32873
rect 9868 11479 9908 11488
rect 10060 7160 10100 32824
rect 10156 8672 10196 42736
rect 10348 41936 10388 41945
rect 10252 38912 10292 38921
rect 10252 11696 10292 38872
rect 10252 11647 10292 11656
rect 10156 8623 10196 8632
rect 10348 7412 10388 41896
rect 10444 39500 10484 39509
rect 10444 15728 10484 39460
rect 10444 15679 10484 15688
rect 10924 17996 10964 18005
rect 10924 10100 10964 17956
rect 10924 10051 10964 10060
rect 10348 7363 10388 7372
rect 10060 7111 10100 7120
rect 9772 6439 9812 6448
rect 9100 4843 9140 4852
rect 8332 4759 8372 4768
rect 8140 1399 8180 1408
rect 6028 223 6068 232
use sg13g2_inv_1  _053_
timestamp 1676382929
transform -1 0 5760 0 -1 25704
box -48 -56 336 834
use sg13g2_inv_1  _054_
timestamp 1676382929
transform -1 0 5376 0 1 15120
box -48 -56 336 834
use sg13g2_inv_1  _055_
timestamp 1676382929
transform 1 0 5568 0 1 22680
box -48 -56 336 834
use sg13g2_inv_1  _056_
timestamp 1676382929
transform 1 0 2880 0 -1 27216
box -48 -56 336 834
use sg13g2_mux4_1  _057_
timestamp 1677257233
transform 1 0 2784 0 1 21168
box -48 -56 2064 834
use sg13g2_nor2_1  _058_
timestamp 1676627187
transform -1 0 4992 0 -1 24192
box -48 -56 432 834
use sg13g2_nor2_1  _059_
timestamp 1676627187
transform 1 0 3936 0 1 25704
box -48 -56 432 834
use sg13g2_nor2b_1  _060_
timestamp 1685181386
transform 1 0 2880 0 -1 25704
box -54 -56 528 834
use sg13g2_nor3_1  _061_
timestamp 1676639442
transform -1 0 3840 0 -1 25704
box -48 -56 528 834
use sg13g2_mux2_1  _062_
timestamp 1677247768
transform 1 0 3840 0 -1 25704
box -48 -56 1008 834
use sg13g2_a21o_1  _063_
timestamp 1677175127
transform -1 0 5472 0 -1 25704
box -48 -56 720 834
use sg13g2_o21ai_1  _064_
timestamp 1685175443
transform 1 0 3456 0 1 24192
box -48 -56 538 834
use sg13g2_mux2_1  _065_
timestamp 1677247768
transform 1 0 1824 0 1 21168
box -48 -56 1008 834
use sg13g2_mux2_1  _066_
timestamp 1677247768
transform -1 0 3744 0 -1 22680
box -48 -56 1008 834
use sg13g2_mux2_1  _067_
timestamp 1677247768
transform 1 0 2592 0 1 22680
box -48 -56 1008 834
use sg13g2_mux2_1  _068_
timestamp 1677247768
transform 1 0 1152 0 -1 24192
box -48 -56 1008 834
use sg13g2_mux4_1  _069_
timestamp 1677257233
transform 1 0 2112 0 -1 24192
box -48 -56 2064 834
use sg13g2_nand2b_1  _070_
timestamp 1676567195
transform 1 0 2976 0 1 24192
box -48 -56 528 834
use sg13g2_o21ai_1  _071_
timestamp 1685175443
transform -1 0 4512 0 1 24192
box -48 -56 538 834
use sg13g2_mux4_1  _072_
timestamp 1677257233
transform 1 0 3648 0 -1 21168
box -48 -56 2064 834
use sg13g2_nor2_1  _073_
timestamp 1676627187
transform -1 0 6240 0 1 19656
box -48 -56 432 834
use sg13g2_nor2_1  _074_
timestamp 1676627187
transform -1 0 5376 0 1 22680
box -48 -56 432 834
use sg13g2_nor2b_1  _075_
timestamp 1685181386
transform -1 0 4992 0 1 22680
box -54 -56 528 834
use sg13g2_nor3_1  _076_
timestamp 1676639442
transform -1 0 5376 0 1 19656
box -48 -56 528 834
use sg13g2_mux2_1  _077_
timestamp 1677247768
transform 1 0 4800 0 1 21168
box -48 -56 1008 834
use sg13g2_a21o_1  _078_
timestamp 1677175127
transform -1 0 6432 0 1 21168
box -48 -56 720 834
use sg13g2_o21ai_1  _079_
timestamp 1685175443
transform 1 0 5664 0 -1 21168
box -48 -56 538 834
use sg13g2_mux2_1  _080_
timestamp 1677247768
transform 1 0 1920 0 1 19656
box -48 -56 1008 834
use sg13g2_mux2_1  _081_
timestamp 1677247768
transform 1 0 2016 0 -1 19656
box -48 -56 1008 834
use sg13g2_mux2_1  _082_
timestamp 1677247768
transform 1 0 2688 0 -1 21168
box -48 -56 1008 834
use sg13g2_mux2_1  _083_
timestamp 1677247768
transform 1 0 1728 0 -1 21168
box -48 -56 1008 834
use sg13g2_mux4_1  _084_
timestamp 1677257233
transform 1 0 2880 0 1 19656
box -48 -56 2064 834
use sg13g2_nand2b_1  _085_
timestamp 1676567195
transform -1 0 5856 0 1 19656
box -48 -56 528 834
use sg13g2_o21ai_1  _086_
timestamp 1685175443
transform 1 0 6144 0 -1 21168
box -48 -56 538 834
use sg13g2_mux4_1  _087_
timestamp 1677257233
transform 1 0 6240 0 1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _088_
timestamp 1677257233
transform 1 0 6528 0 -1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _089_
timestamp 1677257233
transform 1 0 4512 0 -1 36288
box -48 -56 2064 834
use sg13g2_mux4_1  _090_
timestamp 1677257233
transform 1 0 3552 0 -1 33264
box -48 -56 2064 834
use sg13g2_mux4_1  _091_
timestamp 1677257233
transform 1 0 6048 0 1 10584
box -48 -56 2064 834
use sg13g2_mux4_1  _092_
timestamp 1677257233
transform 1 0 4224 0 1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _093_
timestamp 1677257233
transform 1 0 7584 0 -1 18144
box -48 -56 2064 834
use sg13g2_mux4_1  _094_
timestamp 1677257233
transform 1 0 7680 0 -1 15120
box -48 -56 2064 834
use sg13g2_mux4_1  _095_
timestamp 1677257233
transform 1 0 3648 0 -1 40824
box -48 -56 2064 834
use sg13g2_mux4_1  _096_
timestamp 1677257233
transform 1 0 5952 0 -1 30240
box -48 -56 2064 834
use sg13g2_mux4_1  _097_
timestamp 1677257233
transform 1 0 7776 0 1 39312
box -48 -56 2064 834
use sg13g2_mux4_1  _098_
timestamp 1677257233
transform 1 0 7776 0 -1 25704
box -48 -56 2064 834
use sg13g2_mux4_1  _099_
timestamp 1677257233
transform 1 0 2304 0 -1 15120
box -48 -56 2064 834
use sg13g2_mux4_1  _100_
timestamp 1677257233
transform 1 0 1728 0 -1 18144
box -48 -56 2064 834
use sg13g2_mux4_1  _101_
timestamp 1677257233
transform 1 0 8352 0 -1 28728
box -48 -56 2064 834
use sg13g2_mux4_1  _102_
timestamp 1677257233
transform 1 0 8448 0 -1 31752
box -48 -56 2064 834
use sg13g2_mux4_1  _103_
timestamp 1677257233
transform 1 0 8064 0 -1 39312
box -48 -56 2064 834
use sg13g2_mux4_1  _104_
timestamp 1677257233
transform 1 0 6144 0 1 24192
box -48 -56 2064 834
use sg13g2_mux4_1  _105_
timestamp 1677257233
transform 1 0 8064 0 1 33264
box -48 -56 2064 834
use sg13g2_mux4_1  _106_
timestamp 1677257233
transform 1 0 7104 0 1 36288
box -48 -56 2064 834
use sg13g2_mux4_1  _107_
timestamp 1677257233
transform 1 0 2400 0 1 13608
box -48 -56 2064 834
use sg13g2_mux4_1  _108_
timestamp 1677257233
transform 1 0 1824 0 1 18144
box -48 -56 2064 834
use sg13g2_mux4_1  _109_
timestamp 1677257233
transform 1 0 3840 0 -1 22680
box -48 -56 2064 834
use sg13g2_mux4_1  _110_
timestamp 1677257233
transform 1 0 4320 0 -1 18144
box -48 -56 2064 834
use sg13g2_mux4_1  _111_
timestamp 1677257233
transform 1 0 7872 0 -1 34776
box -48 -56 2064 834
use sg13g2_mux4_1  _112_
timestamp 1677257233
transform 1 0 7872 0 -1 33264
box -48 -56 2064 834
use sg13g2_mux4_1  _113_
timestamp 1677257233
transform 1 0 7680 0 -1 40824
box -48 -56 2064 834
use sg13g2_mux4_1  _114_
timestamp 1677257233
transform 1 0 6432 0 -1 27216
box -48 -56 2064 834
use sg13g2_mux4_1  _115_
timestamp 1677257233
transform 1 0 4128 0 -1 10584
box -48 -56 2064 834
use sg13g2_mux4_1  _116_
timestamp 1677257233
transform 1 0 3936 0 1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _117_
timestamp 1677257233
transform 1 0 7872 0 1 18144
box -48 -56 2064 834
use sg13g2_mux4_1  _118_
timestamp 1677257233
transform 1 0 7872 0 1 22680
box -48 -56 2064 834
use sg13g2_mux4_1  _119_
timestamp 1677257233
transform 1 0 4992 0 1 36288
box -48 -56 2064 834
use sg13g2_mux4_1  _120_
timestamp 1677257233
transform 1 0 3264 0 -1 31752
box -48 -56 2064 834
use sg13g2_mux4_1  _121_
timestamp 1677257233
transform 1 0 2880 0 1 36288
box -48 -56 2064 834
use sg13g2_mux4_1  _122_
timestamp 1677257233
transform 1 0 4512 0 1 28728
box -48 -56 2064 834
use sg13g2_mux4_1  _123_
timestamp 1677257233
transform 1 0 4032 0 -1 12096
box -48 -56 2064 834
use sg13g2_mux4_1  _124_
timestamp 1677257233
transform 1 0 2976 0 -1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _125_
timestamp 1677257233
transform 1 0 6720 0 -1 19656
box -48 -56 2064 834
use sg13g2_mux4_1  _126_
timestamp 1677257233
transform 1 0 7680 0 -1 16632
box -48 -56 2064 834
use sg13g2_mux4_1  _127_
timestamp 1677257233
transform 1 0 3840 0 -1 37800
box -48 -56 2064 834
use sg13g2_mux4_1  _128_
timestamp 1677257233
transform 1 0 2784 0 1 31752
box -48 -56 2064 834
use sg13g2_mux4_1  _129_
timestamp 1677257233
transform 1 0 3072 0 1 39312
box -48 -56 2064 834
use sg13g2_mux4_1  _130_
timestamp 1677257233
transform 1 0 4320 0 -1 28728
box -48 -56 2064 834
use sg13g2_mux2_1  _131_
timestamp 1677247768
transform 1 0 5760 0 -1 9072
box -48 -56 1008 834
use sg13g2_mux2_1  _132_
timestamp 1677247768
transform 1 0 4800 0 1 7560
box -48 -56 1008 834
use sg13g2_mux2_1  _133_
timestamp 1677247768
transform 1 0 7584 0 1 7560
box -48 -56 1008 834
use sg13g2_mux2_1  _134_
timestamp 1677247768
transform 1 0 6816 0 -1 13608
box -48 -56 1008 834
use sg13g2_nand2b_1  _135_
timestamp 1676567195
transform 1 0 5664 0 1 16632
box -48 -56 528 834
use sg13g2_o21ai_1  _136_
timestamp 1685175443
transform 1 0 4704 0 -1 16632
box -48 -56 538 834
use sg13g2_nor2b_1  _137_
timestamp 1685181386
transform 1 0 4224 0 1 16632
box -54 -56 528 834
use sg13g2_a21oi_1  _138_
timestamp 1683973020
transform 1 0 5184 0 1 16632
box -48 -56 528 834
use sg13g2_o21ai_1  _139_
timestamp 1685175443
transform 1 0 3264 0 1 16632
box -48 -56 538 834
use sg13g2_nor3_1  _140_
timestamp 1676639442
transform 1 0 3840 0 -1 18144
box -48 -56 528 834
use sg13g2_o21ai_1  _141_
timestamp 1685175443
transform 1 0 3744 0 1 16632
box -48 -56 538 834
use sg13g2_nand2_1  _142_
timestamp 1676557249
transform 1 0 3840 0 -1 16632
box -48 -56 432 834
use sg13g2_nand3_1  _143_
timestamp 1683988354
transform 1 0 4704 0 1 16632
box -48 -56 528 834
use sg13g2_o21ai_1  _144_
timestamp 1685175443
transform 1 0 4224 0 -1 16632
box -48 -56 538 834
use sg13g2_nor2_1  _145_
timestamp 1676627187
transform 1 0 3936 0 -1 28728
box -48 -56 432 834
use sg13g2_a21oi_1  _146_
timestamp 1683973020
transform -1 0 3936 0 -1 28728
box -48 -56 528 834
use sg13g2_nor2_1  _147_
timestamp 1676627187
transform -1 0 4512 0 1 30240
box -48 -56 432 834
use sg13g2_a221oi_1  _148_
timestamp 1685197497
transform 1 0 3072 0 1 28728
box -48 -56 816 834
use sg13g2_nor2b_1  _149_
timestamp 1685181386
transform 1 0 3840 0 1 28728
box -54 -56 528 834
use sg13g2_a22oi_1  _150_
timestamp 1685173987
transform -1 0 4704 0 -1 30240
box -48 -56 624 834
use sg13g2_o21ai_1  _151_
timestamp 1685175443
transform -1 0 3648 0 1 30240
box -48 -56 538 834
use sg13g2_nand3_1  _152_
timestamp 1683988354
transform -1 0 3360 0 -1 30240
box -48 -56 528 834
use sg13g2_nand2b_2  _153_
timestamp 1685211885
transform 1 0 3360 0 -1 30240
box -48 -56 816 834
use sg13g2_dlhq_1  _154_
timestamp 1678805552
transform 1 0 6240 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _155_
timestamp 1678805552
transform 1 0 8448 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _156_
timestamp 1678805552
transform 1 0 9024 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _157_
timestamp 1678805552
transform -1 0 10560 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _158_
timestamp 1678805552
transform 1 0 9024 0 1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _159_
timestamp 1678805552
transform 1 0 8736 0 -1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _160_
timestamp 1678805552
transform -1 0 10656 0 1 12096
box -50 -56 1692 834
use sg13g2_dlhq_1  _161_
timestamp 1678805552
transform 1 0 9024 0 -1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _162_
timestamp 1678805552
transform 1 0 4608 0 -1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _163_
timestamp 1678805552
transform 1 0 6048 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _164_
timestamp 1678805552
transform 1 0 3072 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _165_
timestamp 1678805552
transform 1 0 3936 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _166_
timestamp 1678805552
transform 1 0 2400 0 1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _167_
timestamp 1678805552
transform 1 0 4416 0 1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _168_
timestamp 1678805552
transform 1 0 1536 0 1 40824
box -50 -56 1692 834
use sg13g2_dlhq_1  _169_
timestamp 1678805552
transform 1 0 3744 0 1 40824
box -50 -56 1692 834
use sg13g2_dlhq_1  _170_
timestamp 1678805552
transform 1 0 1152 0 1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _171_
timestamp 1678805552
transform 1 0 1920 0 -1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _172_
timestamp 1678805552
transform 1 0 2304 0 1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _173_
timestamp 1678805552
transform 1 0 4128 0 1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _174_
timestamp 1678805552
transform 1 0 6048 0 1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _175_
timestamp 1678805552
transform 1 0 8256 0 1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _176_
timestamp 1678805552
transform 1 0 5088 0 -1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _177_
timestamp 1678805552
transform 1 0 6528 0 1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _178_
timestamp 1678805552
transform 1 0 1344 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _179_
timestamp 1678805552
transform 1 0 2496 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _180_
timestamp 1678805552
transform 1 0 2208 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _181_
timestamp 1678805552
transform 1 0 4320 0 1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _182_
timestamp 1678805552
transform 1 0 1920 0 -1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _183_
timestamp 1678805552
transform 1 0 4704 0 1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _184_
timestamp 1678805552
transform 1 0 1248 0 1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _185_
timestamp 1678805552
transform 1 0 2592 0 -1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _186_
timestamp 1678805552
transform 1 0 1344 0 -1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _187_
timestamp 1678805552
transform 1 0 3168 0 -1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _188_
timestamp 1678805552
transform -1 0 10464 0 -1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _189_
timestamp 1678805552
transform -1 0 10368 0 -1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _190_
timestamp 1678805552
transform -1 0 10464 0 -1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _191_
timestamp 1678805552
transform 1 0 8352 0 -1 22680
box -50 -56 1692 834
use sg13g2_dlhq_1  _192_
timestamp 1678805552
transform -1 0 10656 0 -1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _193_
timestamp 1678805552
transform 1 0 8832 0 1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _194_
timestamp 1678805552
transform 1 0 1728 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _195_
timestamp 1678805552
transform 1 0 4224 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _196_
timestamp 1678805552
transform 1 0 2208 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _197_
timestamp 1678805552
transform 1 0 3936 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _198_
timestamp 1678805552
transform 1 0 6144 0 1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _199_
timestamp 1678805552
transform 1 0 4800 0 -1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _200_
timestamp 1678805552
transform 1 0 6336 0 1 40824
box -50 -56 1692 834
use sg13g2_dlhq_1  _201_
timestamp 1678805552
transform 1 0 6048 0 -1 40824
box -50 -56 1692 834
use sg13g2_dlhq_1  _202_
timestamp 1678805552
transform 1 0 6336 0 1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _203_
timestamp 1678805552
transform 1 0 6240 0 -1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _204_
timestamp 1678805552
transform 1 0 6048 0 -1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _205_
timestamp 1678805552
transform 1 0 6048 0 -1 39312
box -50 -56 1692 834
use sg13g2_dlhq_1  _206_
timestamp 1678805552
transform -1 0 6048 0 -1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _207_
timestamp 1678805552
transform -1 0 7008 0 -1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _208_
timestamp 1678805552
transform 1 0 1152 0 -1 22680
box -50 -56 1692 834
use sg13g2_dlhq_1  _209_
timestamp 1678805552
transform -1 0 7680 0 -1 22680
box -50 -56 1692 834
use sg13g2_dlhq_1  _210_
timestamp 1678805552
transform 1 0 1440 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _211_
timestamp 1678805552
transform 1 0 1152 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _212_
timestamp 1678805552
transform 1 0 2112 0 1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _213_
timestamp 1678805552
transform -1 0 4416 0 1 12096
box -50 -56 1692 834
use sg13g2_dlhq_1  _214_
timestamp 1678805552
transform 1 0 7104 0 -1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _215_
timestamp 1678805552
transform 1 0 5856 0 -1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _216_
timestamp 1678805552
transform 1 0 8640 0 1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _217_
timestamp 1678805552
transform 1 0 6336 0 1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _218_
timestamp 1678805552
transform 1 0 5856 0 -1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _219_
timestamp 1678805552
transform 1 0 4512 0 1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _220_
timestamp 1678805552
transform 1 0 8736 0 1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _221_
timestamp 1678805552
transform 1 0 6912 0 1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _222_
timestamp 1678805552
transform 1 0 9024 0 -1 30240
box -50 -56 1692 834
use sg13g2_dlhq_1  _223_
timestamp 1678805552
transform 1 0 7776 0 1 30240
box -50 -56 1692 834
use sg13g2_dlhq_1  _224_
timestamp 1678805552
transform 1 0 8832 0 1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _225_
timestamp 1678805552
transform 1 0 7488 0 1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _226_
timestamp 1678805552
transform 1 0 1440 0 -1 12096
box -50 -56 1692 834
use sg13g2_dlhq_1  _227_
timestamp 1678805552
transform 1 0 1152 0 1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _228_
timestamp 1678805552
transform 1 0 1344 0 -1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _229_
timestamp 1678805552
transform 1 0 1152 0 1 12096
box -50 -56 1692 834
use sg13g2_dlhq_1  _230_
timestamp 1678805552
transform 1 0 5952 0 -1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _231_
timestamp 1678805552
transform 1 0 7680 0 1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _232_
timestamp 1678805552
transform 1 0 6336 0 -1 42336
box -50 -56 1692 834
use sg13g2_dlhq_1  _233_
timestamp 1678805552
transform 1 0 7968 0 1 40824
box -50 -56 1692 834
use sg13g2_dlhq_1  _234_
timestamp 1678805552
transform 1 0 4512 0 1 30240
box -50 -56 1692 834
use sg13g2_dlhq_1  _235_
timestamp 1678805552
transform 1 0 6144 0 1 30240
box -50 -56 1692 834
use sg13g2_dlhq_1  _236_
timestamp 1678805552
transform 1 0 2016 0 -1 40824
box -50 -56 1692 834
use sg13g2_dlhq_1  _237_
timestamp 1678805552
transform 1 0 3936 0 -1 39312
box -50 -56 1692 834
use sg13g2_dlhq_1  _238_
timestamp 1678805552
transform 1 0 6048 0 -1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _239_
timestamp 1678805552
transform 1 0 7680 0 1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _240_
timestamp 1678805552
transform 1 0 5376 0 1 18144
box -50 -56 1692 834
use sg13g2_dlhq_1  _241_
timestamp 1678805552
transform 1 0 7776 0 1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _242_
timestamp 1678805552
transform 1 0 2112 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _243_
timestamp 1678805552
transform 1 0 3936 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _244_
timestamp 1678805552
transform 1 0 1920 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _245_
timestamp 1678805552
transform 1 0 6144 0 -1 12096
box -50 -56 1692 834
use sg13g2_dlhq_1  _246_
timestamp 1678805552
transform 1 0 1632 0 1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _247_
timestamp 1678805552
transform 1 0 3840 0 -1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _248_
timestamp 1678805552
transform 1 0 1536 0 1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _249_
timestamp 1678805552
transform 1 0 3936 0 1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _250_
timestamp 1678805552
transform 1 0 5664 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _251_
timestamp 1678805552
transform 1 0 6912 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _252_
timestamp 1678805552
transform -1 0 9888 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _253_
timestamp 1678805552
transform 1 0 6912 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _254_
timestamp 1678805552
transform -1 0 10272 0 1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _255_
timestamp 1678805552
transform -1 0 8256 0 1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _256_
timestamp 1678805552
transform -1 0 10464 0 -1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _257_
timestamp 1678805552
transform -1 0 8832 0 -1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _258_
timestamp 1678805552
transform 1 0 2976 0 -1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _259_
timestamp 1678805552
transform 1 0 1632 0 1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _260_
timestamp 1678805552
transform 1 0 1728 0 -1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _261_
timestamp 1678805552
transform 1 0 1152 0 1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _262_
timestamp 1678805552
transform 1 0 1728 0 1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _263_
timestamp 1678805552
transform 1 0 1152 0 -1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _264_
timestamp 1678805552
transform 1 0 1344 0 1 39312
box -50 -56 1692 834
use sg13g2_dlhq_1  _265_
timestamp 1678805552
transform 1 0 1344 0 -1 39312
box -50 -56 1692 834
use sg13g2_dlhq_1  _266_
timestamp 1678805552
transform 1 0 1152 0 -1 30240
box -50 -56 1692 834
use sg13g2_dlhq_1  _267_
timestamp 1678805552
transform 1 0 1344 0 1 30240
box -50 -56 1692 834
use sg13g2_tiehi  _268__196
timestamp 1680000651
transform 1 0 8640 0 1 12096
box -48 -56 432 834
use sg13g2_dfrbp_1  _268_
timestamp 1678705109
transform 1 0 8160 0 -1 12096
box -60 -56 2556 834
use sg13g2_dfrbp_1  _269_
timestamp 1678705109
transform 1 0 8160 0 1 10584
box -60 -56 2556 834
use sg13g2_tiehi  _269__197
timestamp 1680000651
transform -1 0 9600 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  _272_
timestamp 1676381911
transform 1 0 5472 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  _273_
timestamp 1676381911
transform 1 0 5952 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  _274_
timestamp 1676381911
transform 1 0 1632 0 -1 19656
box -48 -56 432 834
use sg13g2_buf_1  _275_
timestamp 1676381911
transform 1 0 7008 0 1 18144
box -48 -56 432 834
use sg13g2_buf_2  _276_
timestamp 1676381867
transform 1 0 1344 0 1 4536
box -48 -56 528 834
use sg13g2_buf_2  _277_
timestamp 1676381867
transform -1 0 2112 0 -1 4536
box -48 -56 528 834
use sg13g2_buf_1  _278_
timestamp 1676381911
transform 1 0 3744 0 1 10584
box -48 -56 432 834
use sg13g2_buf_2  _279_
timestamp 1676381867
transform 1 0 3072 0 -1 12096
box -48 -56 528 834
use sg13g2_buf_1  _280_
timestamp 1676381911
transform 1 0 5952 0 1 34776
box -48 -56 432 834
use sg13g2_buf_1  _281_
timestamp 1676381911
transform 1 0 5472 0 -1 34776
box -48 -56 432 834
use sg13g2_buf_1  _282_
timestamp 1676381911
transform 1 0 1152 0 1 40824
box -48 -56 432 834
use sg13g2_buf_1  _283_
timestamp 1676381911
transform 1 0 5568 0 1 34776
box -48 -56 432 834
use sg13g2_buf_2  _284_
timestamp 1676381867
transform -1 0 2304 0 1 4536
box -48 -56 528 834
use sg13g2_buf_2  _285_
timestamp 1676381867
transform -1 0 9024 0 -1 6048
box -48 -56 528 834
use sg13g2_buf_1  _286_
timestamp 1676381911
transform 1 0 9792 0 1 39312
box -48 -56 432 834
use sg13g2_buf_1  _287_
timestamp 1676381911
transform 1 0 8448 0 -1 37800
box -48 -56 432 834
use sg13g2_buf_1  _288_
timestamp 1676381911
transform 1 0 10080 0 1 30240
box -48 -56 432 834
use sg13g2_buf_2  _289_
timestamp 1676381867
transform -1 0 7680 0 1 13608
box -48 -56 528 834
use sg13g2_buf_2  _290_
timestamp 1676381867
transform -1 0 9792 0 1 13608
box -48 -56 528 834
use sg13g2_buf_1  _291_
timestamp 1676381911
transform 1 0 9312 0 1 25704
box -48 -56 432 834
use sg13g2_buf_2  _292_
timestamp 1676381867
transform -1 0 3264 0 -1 7560
box -48 -56 528 834
use sg13g2_buf_2  _293_
timestamp 1676381867
transform -1 0 1728 0 -1 9072
box -48 -56 528 834
use sg13g2_buf_2  _294_
timestamp 1676381867
transform -1 0 2208 0 -1 9072
box -48 -56 528 834
use sg13g2_buf_2  _295_
timestamp 1676381867
transform -1 0 2592 0 1 22680
box -48 -56 528 834
use sg13g2_buf_2  _296_
timestamp 1676381867
transform -1 0 2400 0 -1 27216
box -48 -56 528 834
use sg13g2_buf_2  _297_
timestamp 1676381867
transform -1 0 2880 0 -1 27216
box -48 -56 528 834
use sg13g2_buf_1  _298_
timestamp 1676381911
transform 1 0 5664 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  _299_
timestamp 1676381911
transform 1 0 3552 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_2  _300_
timestamp 1676381867
transform -1 0 3744 0 1 33264
box -48 -56 528 834
use sg13g2_buf_2  _301_
timestamp 1676381867
transform -1 0 4704 0 1 33264
box -48 -56 528 834
use sg13g2_buf_1  _302_
timestamp 1676381911
transform 1 0 1152 0 1 34776
box -48 -56 432 834
use sg13g2_buf_1  _303_
timestamp 1676381911
transform -1 0 9984 0 -1 42336
box -48 -56 432 834
use sg13g2_buf_1  _304_
timestamp 1676381911
transform -1 0 8352 0 -1 42336
box -48 -56 432 834
use sg13g2_buf_1  _305_
timestamp 1676381911
transform -1 0 5184 0 1 42336
box -48 -56 432 834
use sg13g2_buf_1  _306_
timestamp 1676381911
transform -1 0 7392 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  _307_
timestamp 1676381911
transform -1 0 6528 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  _308_
timestamp 1676381911
transform 1 0 2400 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  _309_
timestamp 1676381911
transform 1 0 3552 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  _310_
timestamp 1676381911
transform 1 0 2784 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  _311_
timestamp 1676381911
transform 1 0 4800 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  _312_
timestamp 1676381911
transform -1 0 6912 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  _313_
timestamp 1676381911
transform -1 0 8160 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  _314_
timestamp 1676381911
transform -1 0 7776 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  _315_
timestamp 1676381911
transform 1 0 5184 0 1 42336
box -48 -56 432 834
use sg13g2_buf_1  _316_
timestamp 1676381911
transform 1 0 3168 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  _317_
timestamp 1676381911
transform 1 0 4416 0 -1 42336
box -48 -56 432 834
use sg13g2_buf_1  _318_
timestamp 1676381911
transform 1 0 3936 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  _319_
timestamp 1676381911
transform 1 0 3072 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  _320_
timestamp 1676381911
transform 1 0 8928 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  _321_
timestamp 1676381911
transform 1 0 9312 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  _322_
timestamp 1676381911
transform -1 0 8160 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  _323_
timestamp 1676381911
transform -1 0 8160 0 -1 13608
box -48 -56 432 834
use sg13g2_buf_1  _324_
timestamp 1676381911
transform -1 0 8448 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _325_
timestamp 1676381911
transform -1 0 6144 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _326_
timestamp 1676381911
transform -1 0 6240 0 1 9072
box -48 -56 432 834
use sg13g2_buf_2  _327_
timestamp 1676381867
transform -1 0 6816 0 -1 28728
box -48 -56 528 834
use sg13g2_buf_2  _328_
timestamp 1676381867
transform -1 0 5568 0 -1 42336
box -48 -56 528 834
use sg13g2_buf_2  _329_
timestamp 1676381867
transform -1 0 5280 0 1 31752
box -48 -56 528 834
use sg13g2_buf_2  _330_
timestamp 1676381867
transform -1 0 6336 0 1 37800
box -48 -56 528 834
use sg13g2_buf_1  _331_
timestamp 1676381911
transform -1 0 10272 0 1 15120
box -48 -56 432 834
use sg13g2_buf_2  _332_
timestamp 1676381867
transform -1 0 10368 0 1 18144
box -48 -56 528 834
use sg13g2_buf_1  _333_
timestamp 1676381911
transform -1 0 5376 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _334_
timestamp 1676381911
transform -1 0 6432 0 1 12096
box -48 -56 432 834
use sg13g2_buf_2  _335_
timestamp 1676381867
transform -1 0 7008 0 1 28728
box -48 -56 528 834
use sg13g2_buf_2  _336_
timestamp 1676381867
transform 1 0 3360 0 -1 37800
box -48 -56 528 834
use sg13g2_buf_2  _337_
timestamp 1676381867
transform -1 0 5760 0 -1 31752
box -48 -56 528 834
use sg13g2_buf_2  _338_
timestamp 1676381867
transform -1 0 8160 0 -1 37800
box -48 -56 528 834
use sg13g2_buf_2  _339_
timestamp 1676381867
transform -1 0 10368 0 1 22680
box -48 -56 528 834
use sg13g2_buf_1  _340_
timestamp 1676381911
transform -1 0 9984 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  _341_
timestamp 1676381911
transform 1 0 5760 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _342_
timestamp 1676381911
transform -1 0 6528 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_2  _343_
timestamp 1676381867
transform -1 0 10272 0 -1 25704
box -48 -56 528 834
use sg13g2_buf_2  _344_
timestamp 1676381867
transform -1 0 10656 0 1 39312
box -48 -56 528 834
use sg13g2_buf_2  _345_
timestamp 1676381867
transform -1 0 8448 0 -1 30240
box -48 -56 528 834
use sg13g2_buf_2  _346_
timestamp 1676381867
transform -1 0 6048 0 1 40824
box -48 -56 528 834
use sg13g2_buf_1  _347_
timestamp 1676381911
transform -1 0 10080 0 -1 15120
box -48 -56 432 834
use sg13g2_buf_1  _348_
timestamp 1676381911
transform -1 0 10272 0 1 16632
box -48 -56 432 834
use sg13g2_buf_1  _349_
timestamp 1676381911
transform -1 0 6624 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _350_
timestamp 1676381911
transform -1 0 8352 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_2  _351_
timestamp 1676381867
transform -1 0 6048 0 -1 33264
box -48 -56 528 834
use sg13g2_buf_2  _352_
timestamp 1676381867
transform -1 0 7008 0 -1 36288
box -48 -56 528 834
use sg13g2_buf_1  _353_
timestamp 1676381911
transform -1 0 9408 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _354_
timestamp 1676381911
transform -1 0 8736 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_2  _355_
timestamp 1676381867
transform -1 0 8928 0 -1 27216
box -48 -56 528 834
use sg13g2_buf_2  _356_
timestamp 1676381867
transform -1 0 10656 0 -1 40824
box -48 -56 528 834
use sg13g2_buf_2  _357_
timestamp 1676381867
transform -1 0 10368 0 -1 33264
box -48 -56 528 834
use sg13g2_buf_2  _358_
timestamp 1676381867
transform -1 0 10368 0 -1 34776
box -48 -56 528 834
use sg13g2_buf_1  _359_
timestamp 1676381911
transform -1 0 6624 0 1 16632
box -48 -56 432 834
use sg13g2_buf_1  _360_
timestamp 1676381911
transform -1 0 6240 0 1 22680
box -48 -56 432 834
use sg13g2_buf_1  _361_
timestamp 1676381911
transform -1 0 4704 0 1 18144
box -48 -56 432 834
use sg13g2_buf_1  _362_
timestamp 1676381911
transform -1 0 4800 0 1 13608
box -48 -56 432 834
use sg13g2_buf_2  _363_
timestamp 1676381867
transform -1 0 9696 0 1 36288
box -48 -56 528 834
use sg13g2_buf_2  _364_
timestamp 1676381867
transform -1 0 10560 0 1 33264
box -48 -56 528 834
use sg13g2_buf_2  _365_
timestamp 1676381867
transform -1 0 8640 0 1 24192
box -48 -56 528 834
use sg13g2_buf_2  _366_
timestamp 1676381867
transform -1 0 10560 0 -1 39312
box -48 -56 528 834
use sg13g2_buf_2  _367_
timestamp 1676381867
transform 1 0 9600 0 1 30240
box -48 -56 528 834
use sg13g2_buf_2  _368_
timestamp 1676381867
transform 1 0 9600 0 1 28728
box -48 -56 528 834
use sg13g2_buf_1  _369_
timestamp 1676381911
transform -1 0 5088 0 1 18144
box -48 -56 432 834
use sg13g2_buf_1  _370_
timestamp 1676381911
transform -1 0 4704 0 1 15120
box -48 -56 432 834
use sg13g2_buf_2  _371_
timestamp 1676381867
transform -1 0 4800 0 1 42336
box -48 -56 528 834
use sg13g2_buf_2  _372_
timestamp 1676381867
transform -1 0 5952 0 1 39312
box -48 -56 528 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform 1 0 9888 0 -1 40824
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_2
timestamp 1679999689
transform 1 0 9216 0 1 31752
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_3
timestamp 1679999689
transform 1 0 8352 0 1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_4
timestamp 1679999689
transform 1 0 8928 0 1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_5
timestamp 1679999689
transform 1 0 4800 0 -1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_6
timestamp 1679999689
transform 1 0 6432 0 1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_7
timestamp 1679999689
transform 1 0 10368 0 1 37800
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_8
timestamp 1679999689
transform 1 0 8640 0 1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_9
timestamp 1679999689
transform 1 0 6048 0 1 40824
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_10
timestamp 1679999689
transform 1 0 7008 0 1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_11
timestamp 1679999689
transform 1 0 5856 0 1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_12
timestamp 1679999689
transform 1 0 6144 0 1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_13
timestamp 1679999689
transform 1 0 5568 0 1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_14
timestamp 1679999689
transform 1 0 5568 0 -1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_15
timestamp 1679999689
transform 1 0 4128 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_16
timestamp 1679999689
transform -1 0 5280 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_17
timestamp 1679999689
transform -1 0 4704 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_18
timestamp 1679999689
transform 1 0 5952 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_19
timestamp 1679999689
transform 1 0 10368 0 -1 36288
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_20
timestamp 1679999689
transform 1 0 7776 0 1 33264
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_21
timestamp 1679999689
transform 1 0 8928 0 1 31752
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_22
timestamp 1679999689
transform 1 0 6720 0 1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_23
timestamp 1679999689
transform 1 0 7296 0 1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_24
timestamp 1679999689
transform 1 0 9600 0 1 40824
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_25
timestamp 1679999689
transform 1 0 9312 0 1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_26
timestamp 1679999689
transform 1 0 6720 0 1 39312
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_27
timestamp 1679999689
transform 1 0 8064 0 -1 28728
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_28
timestamp 1679999689
transform 1 0 7872 0 1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_29
timestamp 1679999689
transform 1 0 8352 0 -1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_30
timestamp 1679999689
transform 1 0 7584 0 1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_31
timestamp 1679999689
transform 1 0 5856 0 -1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_32
timestamp 1679999689
transform -1 0 4992 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_33
timestamp 1679999689
transform 1 0 4416 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_34
timestamp 1679999689
transform 1 0 4608 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_35
timestamp 1679999689
transform 1 0 6144 0 -1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_36
timestamp 1679999689
transform 1 0 8448 0 1 31752
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_37
timestamp 1679999689
transform 1 0 6912 0 -1 31752
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_38
timestamp 1679999689
transform 1 0 9600 0 1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_39
timestamp 1679999689
transform 1 0 7008 0 1 39312
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_40
timestamp 1679999689
transform 1 0 7296 0 1 39312
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_41
timestamp 1679999689
transform 1 0 8928 0 -1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_42
timestamp 1679999689
transform 1 0 9984 0 -1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_43
timestamp 1679999689
transform 1 0 8160 0 -1 37800
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_44
timestamp 1679999689
transform 1 0 7392 0 1 25704
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_45
timestamp 1679999689
transform 1 0 3648 0 1 34776
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_46
timestamp 1679999689
transform 1 0 3552 0 -1 34776
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_47
timestamp 1679999689
transform 1 0 4224 0 -1 36288
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_48
timestamp 1679999689
transform 1 0 8640 0 -1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_49
timestamp 1679999689
transform 1 0 4992 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_50
timestamp 1679999689
transform 1 0 4704 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_51
timestamp 1679999689
transform 1 0 4320 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_52
timestamp 1679999689
transform -1 0 5856 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_53
timestamp 1679999689
transform 1 0 7776 0 -1 28728
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_54
timestamp 1679999689
transform 1 0 8064 0 1 27216
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_55
timestamp 1679999689
transform 1 0 10368 0 1 22680
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_56
timestamp 1679999689
transform -1 0 1920 0 -1 34776
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_57
timestamp 1679999689
transform 1 0 5760 0 1 31752
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_58
timestamp 1679999689
transform 1 0 10368 0 -1 34776
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_59
timestamp 1679999689
transform 1 0 10368 0 -1 33264
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_60
timestamp 1679999689
transform 1 0 6432 0 -1 31752
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_61
timestamp 1679999689
transform 1 0 5280 0 -1 24192
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_62
timestamp 1679999689
transform 1 0 6048 0 1 31752
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_63
timestamp 1679999689
transform 1 0 6144 0 -1 31752
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_64
timestamp 1679999689
transform 1 0 7392 0 1 33264
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_65
timestamp 1679999689
transform 1 0 7104 0 1 33264
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_66
timestamp 1679999689
transform 1 0 5280 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_67
timestamp 1679999689
transform 1 0 1152 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_68
timestamp 1679999689
transform -1 0 4416 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_69
timestamp 1679999689
transform -1 0 6144 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_70
timestamp 1679999689
transform 1 0 9984 0 -1 22680
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_71
timestamp 1679999689
transform 1 0 8640 0 1 24192
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_72
timestamp 1679999689
transform 1 0 8256 0 -1 24192
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_73
timestamp 1679999689
transform -1 0 1920 0 1 27216
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_74
timestamp 1679999689
transform 1 0 6816 0 -1 28728
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_75
timestamp 1679999689
transform 1 0 7200 0 -1 31752
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_76
timestamp 1679999689
transform 1 0 10368 0 -1 28728
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_77
timestamp 1679999689
transform 1 0 6240 0 1 22680
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_78
timestamp 1679999689
transform 1 0 7680 0 -1 22680
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_79
timestamp 1679999689
transform 1 0 7104 0 -1 28728
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_80
timestamp 1679999689
transform 1 0 5088 0 1 25704
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_81
timestamp 1679999689
transform -1 0 1920 0 -1 27216
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_82
timestamp 1679999689
transform 1 0 7008 0 1 28728
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_83
timestamp 1679999689
transform 1 0 4896 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_84
timestamp 1679999689
transform 1 0 5568 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_85
timestamp 1679999689
transform 1 0 5184 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_86
timestamp 1679999689
transform -1 0 4128 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_87
timestamp 1679999689
transform 1 0 7776 0 -1 24192
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_88
timestamp 1679999689
transform 1 0 7392 0 1 18144
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_89
timestamp 1679999689
transform 1 0 8160 0 1 19656
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_90
timestamp 1679999689
transform 1 0 5664 0 1 25704
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_91
timestamp 1679999689
transform 1 0 5952 0 1 25704
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_92
timestamp 1679999689
transform 1 0 7488 0 -1 28728
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_93
timestamp 1679999689
transform 1 0 7776 0 1 27216
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_94
timestamp 1679999689
transform 1 0 6624 0 -1 21168
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_95
timestamp 1679999689
transform 1 0 8160 0 1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_96
timestamp 1679999689
transform 1 0 6528 0 1 25704
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_97
timestamp 1679999689
transform 1 0 6816 0 1 25704
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_98
timestamp 1679999689
transform 1 0 6240 0 1 25704
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_99
timestamp 1679999689
transform 1 0 5376 0 1 25704
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_100
timestamp 1679999689
transform 1 0 6144 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_101
timestamp 1679999689
transform 1 0 5856 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_102
timestamp 1679999689
transform 1 0 5472 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_103
timestamp 1679999689
transform 1 0 3552 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_104
timestamp 1679999689
transform -1 0 4320 0 -1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_105
timestamp 1679999689
transform 1 0 8448 0 1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_106
timestamp 1679999689
transform 1 0 8448 0 -1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_107
timestamp 1679999689
transform 1 0 5568 0 -1 24192
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_108
timestamp 1679999689
transform -1 0 7392 0 1 25704
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_109
timestamp 1679999689
transform 1 0 8544 0 -1 24192
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_110
timestamp 1679999689
transform 1 0 6240 0 1 19656
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_111
timestamp 1679999689
transform 1 0 5664 0 -1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_112
timestamp 1679999689
transform 1 0 7488 0 -1 24192
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_113
timestamp 1679999689
transform 1 0 6528 0 1 22680
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_114
timestamp 1679999689
transform 1 0 4992 0 -1 24192
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_115
timestamp 1679999689
transform 1 0 5760 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_116
timestamp 1679999689
transform 1 0 6432 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_117
timestamp 1679999689
transform -1 0 5568 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_118
timestamp 1679999689
transform 1 0 3840 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_119
timestamp 1679999689
transform 1 0 5952 0 -1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_120
timestamp 1679999689
transform 1 0 8160 0 -1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_121
timestamp 1679999689
transform 1 0 7872 0 -1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_122
timestamp 1679999689
transform 1 0 7392 0 1 22680
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_123
timestamp 1679999689
transform 1 0 7968 0 -1 22680
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_124
timestamp 1679999689
transform 1 0 8736 0 -1 19656
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_125
timestamp 1679999689
transform 1 0 5088 0 1 18144
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_126
timestamp 1679999689
transform -1 0 3456 0 1 40824
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_127
timestamp 1679999689
transform 1 0 7584 0 -1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_128
timestamp 1679999689
transform -1 0 1920 0 1 19656
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_129
timestamp 1679999689
transform 1 0 6720 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_130
timestamp 1679999689
transform 1 0 7296 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_131
timestamp 1679999689
transform 1 0 6048 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_132
timestamp 1679999689
transform 1 0 3840 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_133
timestamp 1679999689
transform 1 0 6240 0 -1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_134
timestamp 1679999689
transform 1 0 6912 0 -1 21168
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_135
timestamp 1679999689
transform 1 0 6336 0 -1 18144
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_136
timestamp 1679999689
transform 1 0 9600 0 -1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_137
timestamp 1679999689
transform -1 0 3456 0 1 42336
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_138
timestamp 1679999689
transform 1 0 3456 0 1 40824
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_139
timestamp 1679999689
transform 1 0 7296 0 -1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_140
timestamp 1679999689
transform -1 0 3072 0 1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_141
timestamp 1679999689
transform 1 0 7008 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_142
timestamp 1679999689
transform 1 0 6624 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_143
timestamp 1679999689
transform 1 0 6336 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_144
timestamp 1679999689
transform -1 0 3648 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_145
timestamp 1679999689
transform 1 0 6528 0 -1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_146
timestamp 1679999689
transform 1 0 3072 0 1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_147
timestamp 1679999689
transform 1 0 8928 0 -1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_148
timestamp 1679999689
transform 1 0 9312 0 -1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_149
timestamp 1679999689
transform 1 0 7008 0 -1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_150
timestamp 1679999689
transform 1 0 2400 0 -1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_151
timestamp 1679999689
transform 1 0 4800 0 -1 43848
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_152
timestamp 1679999689
transform 1 0 1152 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_153
timestamp 1679999689
transform 1 0 1152 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_154
timestamp 1679999689
transform 1 0 1536 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_155
timestamp 1679999689
transform 1 0 3648 0 1 6048
box -48 -56 336 834
use sg13g2_buf_2  fanout59
timestamp 1676381867
transform 1 0 9888 0 1 9072
box -48 -56 528 834
use sg13g2_buf_2  fanout60
timestamp 1676381867
transform -1 0 8832 0 1 27216
box -48 -56 528 834
use sg13g2_buf_2  fanout61
timestamp 1676381867
transform -1 0 3936 0 -1 42336
box -48 -56 528 834
use sg13g2_buf_2  fanout62
timestamp 1676381867
transform 1 0 6816 0 1 12096
box -48 -56 528 834
use sg13g2_buf_4  fanout63
timestamp 1676384057
transform 1 0 9696 0 -1 16632
box -48 -56 816 834
use sg13g2_buf_2  fanout64
timestamp 1676381867
transform -1 0 7968 0 -1 31752
box -48 -56 528 834
use sg13g2_buf_2  fanout65
timestamp 1676381867
transform 1 0 7968 0 -1 31752
box -48 -56 528 834
use sg13g2_buf_2  fanout66
timestamp 1676381867
transform 1 0 7968 0 1 31752
box -48 -56 528 834
use sg13g2_buf_2  fanout67
timestamp 1676381867
transform 1 0 6816 0 1 16632
box -48 -56 528 834
use sg13g2_buf_2  fanout68
timestamp 1676381867
transform -1 0 7776 0 1 16632
box -48 -56 528 834
use sg13g2_buf_2  fanout69
timestamp 1676381867
transform 1 0 8160 0 1 34776
box -48 -56 528 834
use sg13g2_buf_1  fanout70
timestamp 1676381911
transform 1 0 7680 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_2  fanout71
timestamp 1676381867
transform -1 0 7392 0 1 22680
box -48 -56 528 834
use sg13g2_buf_2  fanout72
timestamp 1676381867
transform -1 0 8544 0 1 12096
box -48 -56 528 834
use sg13g2_buf_2  fanout73
timestamp 1676381867
transform -1 0 9888 0 1 16632
box -48 -56 528 834
use sg13g2_buf_2  fanout74
timestamp 1676381867
transform -1 0 3936 0 1 25704
box -48 -56 528 834
use sg13g2_buf_2  fanout75
timestamp 1676381867
transform 1 0 1920 0 1 27216
box -48 -56 528 834
use sg13g2_buf_2  fanout76
timestamp 1676381867
transform 1 0 2208 0 1 28728
box -48 -56 528 834
use sg13g2_buf_2  fanout77
timestamp 1676381867
transform 1 0 2976 0 -1 28728
box -48 -56 528 834
use sg13g2_decap_8  FILLER_0_52
timestamp 1679581782
transform 1 0 6144 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_59
timestamp 1679581782
transform 1 0 6816 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_66
timestamp 1679581782
transform 1 0 7488 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_73
timestamp 1679581782
transform 1 0 8160 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_80
timestamp 1679581782
transform 1 0 8832 0 1 1512
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_87
timestamp 1679577901
transform 1 0 9504 0 1 1512
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_7
timestamp 1677579658
transform 1 0 1824 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_24
timestamp 1677579658
transform 1 0 3456 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_31
timestamp 1677580104
transform 1 0 4128 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_57
timestamp 1679581782
transform 1 0 6624 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_64
timestamp 1679581782
transform 1 0 7296 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_71
timestamp 1679581782
transform 1 0 7968 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_78
timestamp 1679581782
transform 1 0 8640 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_85
timestamp 1679581782
transform 1 0 9312 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_92
timestamp 1677580104
transform 1 0 9984 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_94
timestamp 1677579658
transform 1 0 10176 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_3
timestamp 1677579658
transform 1 0 1440 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_64
timestamp 1679581782
transform 1 0 7296 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_71
timestamp 1679581782
transform 1 0 7968 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_78
timestamp 1679581782
transform 1 0 8640 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_85
timestamp 1679581782
transform 1 0 9312 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_92
timestamp 1677580104
transform 1 0 9984 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_94
timestamp 1677579658
transform 1 0 10176 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_3
timestamp 1677580104
transform 1 0 1440 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_27
timestamp 1677580104
transform 1 0 3744 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_46
timestamp 1677579658
transform 1 0 5568 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_67
timestamp 1679581782
transform 1 0 7584 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_74
timestamp 1679581782
transform 1 0 8256 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_81
timestamp 1679581782
transform 1 0 8928 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_88
timestamp 1677580104
transform 1 0 9600 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_90
timestamp 1677579658
transform 1 0 9792 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_0
timestamp 1677580104
transform 1 0 1152 0 1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_12
timestamp 1677580104
transform 1 0 2304 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_31
timestamp 1677579658
transform 1 0 4128 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_77
timestamp 1679581782
transform 1 0 8544 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_84
timestamp 1679581782
transform 1 0 9216 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_91
timestamp 1679581782
transform 1 0 9888 0 1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_98
timestamp 1677579658
transform 1 0 10560 0 1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_0
timestamp 1677580104
transform 1 0 1152 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_55
timestamp 1677579658
transform 1 0 6432 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_86
timestamp 1679581782
transform 1 0 9408 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_93
timestamp 1677580104
transform 1 0 10080 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_0
timestamp 1677580104
transform 1 0 1152 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_70
timestamp 1679581782
transform 1 0 7872 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_77
timestamp 1679581782
transform 1 0 8544 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_84
timestamp 1679581782
transform 1 0 9216 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_30
timestamp 1677580104
transform 1 0 4032 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_49
timestamp 1677580104
transform 1 0 5856 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_68
timestamp 1679577901
transform 1 0 7680 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_93
timestamp 1677580104
transform 1 0 10080 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_37
timestamp 1677579658
transform 1 0 4704 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_60
timestamp 1679581782
transform 1 0 6912 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_77
timestamp 1679577901
transform 1 0 8544 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_98
timestamp 1677579658
transform 1 0 10560 0 1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_0
timestamp 1677579658
transform 1 0 1152 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_28
timestamp 1677579658
transform 1 0 3840 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_46
timestamp 1677580104
transform 1 0 5568 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_58
timestamp 1677580104
transform 1 0 6720 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_77
timestamp 1677579658
transform 1 0 8544 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_46
timestamp 1677580104
transform 1 0 5568 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_48
timestamp 1677579658
transform 1 0 5760 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_96
timestamp 1677580104
transform 1 0 10368 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_98
timestamp 1677579658
transform 1 0 10560 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_8
timestamp 1677580104
transform 1 0 1920 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_10
timestamp 1677579658
transform 1 0 2112 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_28
timestamp 1677580104
transform 1 0 3840 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_30
timestamp 1677579658
transform 1 0 4032 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_60
timestamp 1679581782
transform 1 0 6912 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_67
timestamp 1679577901
transform 1 0 7584 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_79
timestamp 1677579658
transform 1 0 8736 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_88
timestamp 1677580104
transform 1 0 9600 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_90
timestamp 1677579658
transform 1 0 9792 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_8
timestamp 1677580104
transform 1 0 1920 0 1 10584
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_31
timestamp 1677580104
transform 1 0 4128 0 1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_50
timestamp 1677579658
transform 1 0 5952 0 1 10584
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_72
timestamp 1677579658
transform 1 0 8064 0 1 10584
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_0
timestamp 1677580104
transform 1 0 1152 0 -1 12096
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_2
timestamp 1677579658
transform 1 0 1344 0 -1 12096
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_29
timestamp 1677579658
transform 1 0 3936 0 -1 12096
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_51
timestamp 1677579658
transform 1 0 6048 0 -1 12096
box -48 -56 144 834
use sg13g2_decap_4  FILLER_14_46
timestamp 1679577901
transform 1 0 5568 0 1 12096
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_50
timestamp 1677579658
transform 1 0 5952 0 1 12096
box -48 -56 144 834
use sg13g2_decap_4  FILLER_14_55
timestamp 1679577901
transform 1 0 6432 0 1 12096
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_64
timestamp 1679581782
transform 1 0 7296 0 1 12096
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_71
timestamp 1677579658
transform 1 0 7968 0 1 12096
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_77
timestamp 1677579658
transform 1 0 8544 0 1 12096
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_0
timestamp 1677580104
transform 1 0 1152 0 -1 13608
box -48 -56 240 834
use sg13g2_decap_4  FILLER_15_53
timestamp 1679577901
transform 1 0 6240 0 -1 13608
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_57
timestamp 1677580104
transform 1 0 6624 0 -1 13608
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_73
timestamp 1677580104
transform 1 0 8160 0 -1 13608
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_96
timestamp 1677580104
transform 1 0 10368 0 -1 13608
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_98
timestamp 1677579658
transform 1 0 10560 0 -1 13608
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_12
timestamp 1677579658
transform 1 0 2304 0 1 13608
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_42
timestamp 1677580104
transform 1 0 5184 0 1 13608
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_44
timestamp 1677579658
transform 1 0 5376 0 1 13608
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_49
timestamp 1677579658
transform 1 0 5856 0 1 13608
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_54
timestamp 1679581782
transform 1 0 6336 0 1 13608
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_61
timestamp 1677580104
transform 1 0 7008 0 1 13608
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_90
timestamp 1677579658
transform 1 0 9792 0 1 13608
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_33
timestamp 1677579658
transform 1 0 4320 0 -1 15120
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_93
timestamp 1677580104
transform 1 0 10080 0 -1 15120
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_44
timestamp 1679581782
transform 1 0 5376 0 1 15120
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_68
timestamp 1679577901
transform 1 0 7680 0 1 15120
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_72
timestamp 1677580104
transform 1 0 8064 0 1 15120
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_5
timestamp 1677579658
transform 1 0 1632 0 -1 16632
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_27
timestamp 1677579658
transform 1 0 3744 0 -1 16632
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_42
timestamp 1677580104
transform 1 0 5184 0 -1 16632
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_61
timestamp 1679581782
transform 1 0 7008 0 -1 16632
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_97
timestamp 1677580104
transform 1 0 10464 0 -1 16632
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_52
timestamp 1677579658
transform 1 0 6144 0 1 16632
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_57
timestamp 1677580104
transform 1 0 6624 0 1 16632
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_5
timestamp 1677579658
transform 1 0 1632 0 -1 18144
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_27
timestamp 1677579658
transform 1 0 3744 0 -1 18144
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_57
timestamp 1679581782
transform 1 0 6624 0 -1 18144
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_64
timestamp 1677580104
transform 1 0 7296 0 -1 18144
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_66
timestamp 1677579658
transform 1 0 7488 0 -1 18144
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_92
timestamp 1677580104
transform 1 0 9984 0 -1 18144
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_94
timestamp 1677579658
transform 1 0 10176 0 -1 18144
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_5
timestamp 1677580104
transform 1 0 1632 0 1 18144
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_68
timestamp 1677580104
transform 1 0 7680 0 1 18144
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_96
timestamp 1677580104
transform 1 0 10368 0 1 18144
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_98
timestamp 1677579658
transform 1 0 10560 0 1 18144
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_39
timestamp 1677580104
transform 1 0 4896 0 -1 19656
box -48 -56 240 834
use sg13g2_fill_2  FILLER_24_97
timestamp 1677580104
transform 1 0 10464 0 1 19656
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_5
timestamp 1677579658
transform 1 0 1632 0 -1 21168
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_97
timestamp 1677580104
transform 1 0 10464 0 -1 21168
box -48 -56 240 834
use sg13g2_fill_2  FILLER_26_5
timestamp 1677580104
transform 1 0 1632 0 1 21168
box -48 -56 240 834
use sg13g2_fill_2  FILLER_26_55
timestamp 1677580104
transform 1 0 6432 0 1 21168
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_27
timestamp 1677579658
transform 1 0 3744 0 -1 22680
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_49
timestamp 1677580104
transform 1 0 5856 0 -1 22680
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_74
timestamp 1677579658
transform 1 0 8256 0 -1 22680
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_44
timestamp 1677580104
transform 1 0 5376 0 1 22680
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_59
timestamp 1677579658
transform 1 0 6816 0 1 22680
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_68
timestamp 1677580104
transform 1 0 7680 0 1 22680
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_72
timestamp 1677580104
transform 1 0 8064 0 -1 24192
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_97
timestamp 1677580104
transform 1 0 10464 0 -1 24192
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_17
timestamp 1677580104
transform 1 0 2784 0 1 24192
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_29
timestamp 1677579658
transform 1 0 3936 0 1 24192
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_81
timestamp 1677579658
transform 1 0 8928 0 1 24192
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_17
timestamp 1677579658
transform 1 0 2784 0 -1 25704
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_48
timestamp 1677580104
transform 1 0 5760 0 -1 25704
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_67
timestamp 1677580104
transform 1 0 7584 0 -1 25704
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_5
timestamp 1677579658
transform 1 0 1632 0 1 25704
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_23
timestamp 1677579658
transform 1 0 3360 0 1 25704
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_89
timestamp 1677580104
transform 1 0 9696 0 1 25704
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_81
timestamp 1677579658
transform 1 0 8928 0 -1 27216
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_51
timestamp 1677579658
transform 1 0 6048 0 1 27216
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_97
timestamp 1677580104
transform 1 0 10464 0 1 27216
box -48 -56 240 834
use sg13g2_fill_2  FILLER_35_0
timestamp 1677580104
transform 1 0 1152 0 -1 28728
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_65
timestamp 1677579658
transform 1 0 7392 0 -1 28728
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_10
timestamp 1677579658
transform 1 0 2112 0 1 28728
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_33
timestamp 1677580104
transform 1 0 4320 0 1 28728
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_64
timestamp 1677580104
transform 1 0 7296 0 1 28728
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_83
timestamp 1677579658
transform 1 0 9120 0 1 28728
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_93
timestamp 1677580104
transform 1 0 10080 0 1 28728
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_17
timestamp 1677579658
transform 1 0 2784 0 -1 30240
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_76
timestamp 1677580104
transform 1 0 8448 0 -1 30240
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_0
timestamp 1677580104
transform 1 0 1152 0 1 30240
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_19
timestamp 1677580104
transform 1 0 2976 0 1 30240
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_86
timestamp 1677580104
transform 1 0 9408 0 1 30240
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_97
timestamp 1677580104
transform 1 0 10464 0 1 30240
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_58
timestamp 1677580104
transform 1 0 6720 0 -1 31752
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_97
timestamp 1677580104
transform 1 0 10464 0 -1 31752
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_79
timestamp 1677580104
transform 1 0 8736 0 1 31752
box -48 -56 240 834
use sg13g2_fill_2  FILLER_41_51
timestamp 1677580104
transform 1 0 6048 0 -1 33264
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_68
timestamp 1677579658
transform 1 0 7680 0 1 33264
box -48 -56 144 834
use sg13g2_fill_1  FILLER_42_98
timestamp 1677579658
transform 1 0 10560 0 1 33264
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_71
timestamp 1677580104
transform 1 0 7968 0 1 34776
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_61
timestamp 1677579658
transform 1 0 7008 0 -1 36288
box -48 -56 144 834
use sg13g2_fill_1  FILLER_46_0
timestamp 1677579658
transform 1 0 1152 0 1 36288
box -48 -56 144 834
use sg13g2_fill_1  FILLER_46_39
timestamp 1677579658
transform 1 0 4896 0 1 36288
box -48 -56 144 834
use sg13g2_fill_1  FILLER_46_61
timestamp 1677579658
transform 1 0 7008 0 1 36288
box -48 -56 144 834
use sg13g2_fill_1  FILLER_46_83
timestamp 1677579658
transform 1 0 9120 0 1 36288
box -48 -56 144 834
use sg13g2_fill_2  FILLER_46_89
timestamp 1677580104
transform 1 0 9696 0 1 36288
box -48 -56 240 834
use sg13g2_fill_2  FILLER_47_49
timestamp 1677580104
transform 1 0 5856 0 -1 37800
box -48 -56 240 834
use sg13g2_fill_2  FILLER_47_97
timestamp 1677580104
transform 1 0 10464 0 -1 37800
box -48 -56 240 834
use sg13g2_fill_2  FILLER_48_29
timestamp 1677580104
transform 1 0 3936 0 1 37800
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_48
timestamp 1677579658
transform 1 0 5760 0 1 37800
box -48 -56 144 834
use sg13g2_fill_1  FILLER_48_59
timestamp 1677579658
transform 1 0 6816 0 1 37800
box -48 -56 144 834
use sg13g2_fill_2  FILLER_48_77
timestamp 1677580104
transform 1 0 8544 0 1 37800
box -48 -56 240 834
use sg13g2_fill_2  FILLER_49_0
timestamp 1677580104
transform 1 0 1152 0 -1 39312
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_98
timestamp 1677579658
transform 1 0 10560 0 -1 39312
box -48 -56 144 834
use sg13g2_fill_2  FILLER_50_0
timestamp 1677580104
transform 1 0 1152 0 1 39312
box -48 -56 240 834
use sg13g2_fill_1  FILLER_50_19
timestamp 1677579658
transform 1 0 2976 0 1 39312
box -48 -56 144 834
use sg13g2_fill_2  FILLER_50_67
timestamp 1677580104
transform 1 0 7584 0 1 39312
box -48 -56 240 834
use sg13g2_fill_1  FILLER_51_8
timestamp 1677579658
transform 1 0 1920 0 -1 40824
box -48 -56 144 834
use sg13g2_fill_2  FILLER_51_89
timestamp 1677580104
transform 1 0 9696 0 -1 40824
box -48 -56 240 834
use sg13g2_fill_2  FILLER_52_44
timestamp 1677580104
transform 1 0 5376 0 1 40824
box -48 -56 240 834
use sg13g2_fill_2  FILLER_53_52
timestamp 1677580104
transform 1 0 6144 0 -1 42336
box -48 -56 240 834
use sg13g2_fill_1  FILLER_54_20
timestamp 1677579658
transform 1 0 3072 0 1 42336
box -48 -56 144 834
use sg13g2_fill_2  FILLER_54_73
timestamp 1677580104
transform 1 0 8160 0 1 42336
box -48 -56 240 834
use sg13g2_fill_1  FILLER_54_84
timestamp 1677579658
transform 1 0 9216 0 1 42336
box -48 -56 144 834
use sg13g2_fill_1  FILLER_55_16
timestamp 1677579658
transform 1 0 2688 0 -1 43848
box -48 -56 144 834
use sg13g2_fill_1  FILLER_55_29
timestamp 1677579658
transform 1 0 3936 0 -1 43848
box -48 -56 144 834
use sg13g2_fill_1  FILLER_55_37
timestamp 1677579658
transform 1 0 4704 0 -1 43848
box -48 -56 144 834
use sg13g2_fill_2  FILLER_55_45
timestamp 1677580104
transform 1 0 5472 0 -1 43848
box -48 -56 240 834
use sg13g2_fill_2  FILLER_55_59
timestamp 1677580104
transform 1 0 6816 0 -1 43848
box -48 -56 240 834
use sg13g2_fill_2  FILLER_55_79
timestamp 1677580104
transform 1 0 8736 0 -1 43848
box -48 -56 240 834
use sg13g2_fill_1  FILLER_55_84
timestamp 1677579658
transform 1 0 9216 0 -1 43848
box -48 -56 144 834
use sg13g2_fill_2  FILLER_56_23
timestamp 1677580104
transform 1 0 3360 0 1 43848
box -48 -56 240 834
use sg13g2_fill_1  FILLER_56_37
timestamp 1677579658
transform 1 0 4704 0 1 43848
box -48 -56 144 834
use sg13g2_fill_2  FILLER_56_50
timestamp 1677580104
transform 1 0 5952 0 1 43848
box -48 -56 240 834
use sg13g2_fill_1  FILLER_56_60
timestamp 1677579658
transform 1 0 6912 0 1 43848
box -48 -56 144 834
use sg13g2_fill_2  FILLER_56_79
timestamp 1677580104
transform 1 0 8736 0 1 43848
box -48 -56 240 834
use sg13g2_fill_2  FILLER_56_89
timestamp 1677580104
transform 1 0 9696 0 1 43848
box -48 -56 240 834
use sg13g2_fill_2  FILLER_57_8
timestamp 1677580104
transform 1 0 1920 0 -1 45360
box -48 -56 240 834
use sg13g2_fill_1  FILLER_57_28
timestamp 1677579658
transform 1 0 3840 0 -1 45360
box -48 -56 144 834
use sg13g2_fill_2  FILLER_57_93
timestamp 1677580104
transform 1 0 10080 0 -1 45360
box -48 -56 240 834
use sg13g2_buf_4  input1
timestamp 1676384057
transform 1 0 9888 0 1 1512
box -48 -56 816 834
use sg13g2_buf_4  input2
timestamp 1676384057
transform 1 0 9888 0 -1 4536
box -48 -56 816 834
use sg13g2_buf_1  input3
timestamp 1676381911
transform 1 0 1152 0 -1 15120
box -48 -56 432 834
use sg13g2_buf_2  input4
timestamp 1676381867
transform -1 0 1632 0 -1 16632
box -48 -56 528 834
use sg13g2_buf_2  input5
timestamp 1676381867
transform -1 0 4320 0 1 18144
box -48 -56 528 834
use sg13g2_buf_2  input6
timestamp 1676381867
transform -1 0 4896 0 -1 19656
box -48 -56 528 834
use sg13g2_buf_2  input7
timestamp 1676381867
transform -1 0 4512 0 1 22680
box -48 -56 528 834
use sg13g2_buf_2  input8
timestamp 1676381867
transform -1 0 1632 0 -1 21168
box -48 -56 528 834
use sg13g2_buf_2  input9
timestamp 1676381867
transform -1 0 4032 0 1 22680
box -48 -56 528 834
use sg13g2_buf_2  input10
timestamp 1676381867
transform -1 0 4608 0 -1 24192
box -48 -56 528 834
use sg13g2_buf_2  input11
timestamp 1676381867
transform -1 0 1632 0 1 21168
box -48 -56 528 834
use sg13g2_buf_2  input12
timestamp 1676381867
transform -1 0 2112 0 1 22680
box -48 -56 528 834
use sg13g2_buf_2  input13
timestamp 1676381867
transform -1 0 1632 0 1 22680
box -48 -56 528 834
use sg13g2_buf_2  input14
timestamp 1676381867
transform -1 0 1632 0 1 25704
box -48 -56 528 834
use sg13g2_buf_2  input15
timestamp 1676381867
transform -1 0 1632 0 1 16632
box -48 -56 528 834
use sg13g2_buf_2  input16
timestamp 1676381867
transform -1 0 4416 0 -1 19656
box -48 -56 528 834
use sg13g2_buf_2  input17
timestamp 1676381867
transform -1 0 3936 0 -1 19656
box -48 -56 528 834
use sg13g2_buf_2  input18
timestamp 1676381867
transform -1 0 1632 0 -1 18144
box -48 -56 528 834
use sg13g2_buf_2  input19
timestamp 1676381867
transform -1 0 3456 0 -1 19656
box -48 -56 528 834
use sg13g2_buf_2  input20
timestamp 1676381867
transform -1 0 1632 0 1 18144
box -48 -56 528 834
use sg13g2_buf_2  input21
timestamp 1676381867
transform -1 0 1632 0 -1 19656
box -48 -56 528 834
use sg13g2_buf_2  input22
timestamp 1676381867
transform -1 0 1632 0 1 19656
box -48 -56 528 834
use sg13g2_buf_2  input23
timestamp 1676381867
transform -1 0 1632 0 1 33264
box -48 -56 528 834
use sg13g2_buf_1  input24
timestamp 1676381911
transform 1 0 1920 0 1 37800
box -48 -56 432 834
use sg13g2_buf_1  input25
timestamp 1676381911
transform 1 0 6336 0 1 33264
box -48 -56 432 834
use sg13g2_buf_4  input26
timestamp 1676384057
transform -1 0 1920 0 -1 31752
box -48 -56 816 834
use sg13g2_buf_2  input27
timestamp 1676381867
transform -1 0 1632 0 -1 34776
box -48 -56 528 834
use sg13g2_buf_2  input28
timestamp 1676381867
transform -1 0 4224 0 1 33264
box -48 -56 528 834
use sg13g2_buf_2  input29
timestamp 1676381867
transform -1 0 5760 0 1 31752
box -48 -56 528 834
use sg13g2_buf_2  input30
timestamp 1676381867
transform -1 0 1632 0 -1 36288
box -48 -56 528 834
use sg13g2_buf_2  input31
timestamp 1676381867
transform -1 0 2112 0 -1 36288
box -48 -56 528 834
use sg13g2_buf_2  input32
timestamp 1676381867
transform -1 0 2592 0 -1 36288
box -48 -56 528 834
use sg13g2_buf_4  input33
timestamp 1676384057
transform -1 0 1920 0 -1 33264
box -48 -56 816 834
use sg13g2_buf_2  input34
timestamp 1676381867
transform -1 0 3648 0 1 34776
box -48 -56 528 834
use sg13g2_buf_2  input35
timestamp 1676381867
transform -1 0 1632 0 -1 27216
box -48 -56 528 834
use sg13g2_buf_2  input36
timestamp 1676381867
transform -1 0 4128 0 1 30240
box -48 -56 528 834
use sg13g2_buf_2  input37
timestamp 1676381867
transform -1 0 5184 0 -1 30240
box -48 -56 528 834
use sg13g2_buf_1  input38
timestamp 1676381911
transform 1 0 2880 0 -1 31752
box -48 -56 432 834
use sg13g2_buf_1  input39
timestamp 1676381911
transform -1 0 5568 0 -1 30240
box -48 -56 432 834
use sg13g2_buf_1  input40
timestamp 1676381911
transform -1 0 5952 0 -1 30240
box -48 -56 432 834
use sg13g2_buf_1  input41
timestamp 1676381911
transform 1 0 5760 0 -1 31752
box -48 -56 432 834
use sg13g2_buf_2  input42
timestamp 1676381867
transform -1 0 1632 0 1 27216
box -48 -56 528 834
use sg13g2_buf_1  input43
timestamp 1676381911
transform 1 0 4320 0 1 25704
box -48 -56 432 834
use sg13g2_buf_2  input44
timestamp 1676381867
transform -1 0 1632 0 1 28728
box -48 -56 528 834
use sg13g2_buf_1  input45
timestamp 1676381911
transform 1 0 4032 0 1 27216
box -48 -56 432 834
use sg13g2_buf_1  input46
timestamp 1676381911
transform 1 0 2688 0 1 28728
box -48 -56 432 834
use sg13g2_buf_2  input47
timestamp 1676381867
transform -1 0 2112 0 1 28728
box -48 -56 528 834
use sg13g2_buf_1  input48
timestamp 1676381911
transform 1 0 4704 0 1 25704
box -48 -56 432 834
use sg13g2_buf_2  input49
timestamp 1676381867
transform -1 0 2400 0 -1 31752
box -48 -56 528 834
use sg13g2_buf_2  input50
timestamp 1676381867
transform -1 0 2880 0 -1 31752
box -48 -56 528 834
use sg13g2_buf_1  input51
timestamp 1676381911
transform -1 0 7104 0 1 33264
box -48 -56 432 834
use sg13g2_buf_1  input52
timestamp 1676381911
transform 1 0 2688 0 1 42336
box -48 -56 432 834
use sg13g2_buf_1  input53
timestamp 1676381911
transform 1 0 5088 0 1 39312
box -48 -56 432 834
use sg13g2_buf_1  input54
timestamp 1676381911
transform 1 0 5952 0 1 39312
box -48 -56 432 834
use sg13g2_buf_1  input55
timestamp 1676381911
transform -1 0 6720 0 1 39312
box -48 -56 432 834
use sg13g2_buf_4  input56
timestamp 1676384057
transform -1 0 1920 0 -1 40824
box -48 -56 816 834
use sg13g2_buf_4  input57
timestamp 1676384057
transform -1 0 1920 0 1 37800
box -48 -56 816 834
use sg13g2_buf_4  input58
timestamp 1676384057
transform -1 0 1920 0 -1 42336
box -48 -56 816 834
use sg13g2_buf_4  input59
timestamp 1676384057
transform -1 0 2688 0 -1 42336
box -48 -56 816 834
use sg13g2_buf_2  input60
timestamp 1676381867
transform -1 0 4416 0 -1 42336
box -48 -56 528 834
use sg13g2_buf_4  input61
timestamp 1676384057
transform -1 0 1920 0 1 42336
box -48 -56 816 834
use sg13g2_buf_1  input62
timestamp 1676381911
transform -1 0 7872 0 -1 34776
box -48 -56 432 834
use sg13g2_buf_4  input63
timestamp 1676384057
transform -1 0 2688 0 1 42336
box -48 -56 816 834
use sg13g2_buf_2  input64
timestamp 1676381867
transform -1 0 4320 0 1 42336
box -48 -56 528 834
use sg13g2_buf_4  input65
timestamp 1676384057
transform -1 0 3456 0 -1 42336
box -48 -56 816 834
use sg13g2_buf_4  input66
timestamp 1676384057
transform -1 0 1920 0 1 43848
box -48 -56 816 834
use sg13g2_buf_4  input67
timestamp 1676384057
transform -1 0 2400 0 -1 43848
box -48 -56 816 834
use sg13g2_buf_4  input68
timestamp 1676384057
transform -1 0 1920 0 -1 45360
box -48 -56 816 834
use sg13g2_buf_2  input69
timestamp 1676381867
transform -1 0 2400 0 1 43848
box -48 -56 528 834
use sg13g2_buf_2  input70
timestamp 1676381867
transform -1 0 1632 0 -1 43848
box -48 -56 528 834
use sg13g2_buf_1  input71
timestamp 1676381911
transform 1 0 4320 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  input72
timestamp 1676381911
transform 1 0 4320 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_2  input73
timestamp 1676381867
transform -1 0 2400 0 -1 37800
box -48 -56 528 834
use sg13g2_buf_2  input74
timestamp 1676381867
transform -1 0 3072 0 -1 45360
box -48 -56 528 834
use sg13g2_buf_2  input75
timestamp 1676381867
transform -1 0 2592 0 -1 45360
box -48 -56 528 834
use sg13g2_buf_2  input76
timestamp 1676381867
transform -1 0 2880 0 -1 37800
box -48 -56 528 834
use sg13g2_buf_2  input77
timestamp 1676381867
transform -1 0 3360 0 -1 37800
box -48 -56 528 834
use sg13g2_buf_2  input78
timestamp 1676381867
transform -1 0 3456 0 -1 39312
box -48 -56 528 834
use sg13g2_buf_2  input79
timestamp 1676381867
transform -1 0 3936 0 -1 39312
box -48 -56 528 834
use sg13g2_buf_4  input80
timestamp 1676384057
transform -1 0 1920 0 -1 37800
box -48 -56 816 834
use sg13g2_buf_2  input81
timestamp 1676381867
transform -1 0 6048 0 -1 39312
box -48 -56 528 834
use sg13g2_buf_2  input82
timestamp 1676381867
transform -1 0 6816 0 1 37800
box -48 -56 528 834
use sg13g2_buf_1  output83
timestamp 1676381911
transform 1 0 10272 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output84
timestamp 1676381911
transform 1 0 10272 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output85
timestamp 1676381911
transform 1 0 10272 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output86
timestamp 1676381911
transform 1 0 8640 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output87
timestamp 1676381911
transform 1 0 10272 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output88
timestamp 1676381911
transform 1 0 8832 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output89
timestamp 1676381911
transform 1 0 10272 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output90
timestamp 1676381911
transform 1 0 9888 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output91
timestamp 1676381911
transform 1 0 9888 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output92
timestamp 1676381911
transform 1 0 10272 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output93
timestamp 1676381911
transform 1 0 8352 0 -1 13608
box -48 -56 432 834
use sg13g2_buf_1  output94
timestamp 1676381911
transform 1 0 9888 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  output95
timestamp 1676381911
transform 1 0 10272 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  output96
timestamp 1676381911
transform 1 0 10272 0 -1 25704
box -48 -56 432 834
use sg13g2_buf_1  output97
timestamp 1676381911
transform 1 0 9888 0 1 25704
box -48 -56 432 834
use sg13g2_buf_1  output98
timestamp 1676381911
transform 1 0 10272 0 1 28728
box -48 -56 432 834
use sg13g2_buf_1  output99
timestamp 1676381911
transform 1 0 9216 0 1 28728
box -48 -56 432 834
use sg13g2_buf_1  output100
timestamp 1676381911
transform 1 0 8640 0 -1 30240
box -48 -56 432 834
use sg13g2_buf_1  output101
timestamp 1676381911
transform 1 0 10272 0 1 31752
box -48 -56 432 834
use sg13g2_buf_1  output102
timestamp 1676381911
transform 1 0 9888 0 1 31752
box -48 -56 432 834
use sg13g2_buf_1  output103
timestamp 1676381911
transform 1 0 9504 0 1 31752
box -48 -56 432 834
use sg13g2_buf_1  output104
timestamp 1676381911
transform 1 0 10272 0 1 34776
box -48 -56 432 834
use sg13g2_buf_1  output105
timestamp 1676381911
transform 1 0 10272 0 1 36288
box -48 -56 432 834
use sg13g2_buf_1  output106
timestamp 1676381911
transform 1 0 10272 0 -1 15120
box -48 -56 432 834
use sg13g2_buf_1  output107
timestamp 1676381911
transform 1 0 9888 0 1 36288
box -48 -56 432 834
use sg13g2_buf_1  output108
timestamp 1676381911
transform 1 0 10272 0 1 40824
box -48 -56 432 834
use sg13g2_buf_1  output109
timestamp 1676381911
transform 1 0 10272 0 -1 42336
box -48 -56 432 834
use sg13g2_buf_1  output110
timestamp 1676381911
transform 1 0 9888 0 1 40824
box -48 -56 432 834
use sg13g2_buf_1  output111
timestamp 1676381911
transform 1 0 10272 0 1 42336
box -48 -56 432 834
use sg13g2_buf_1  output112
timestamp 1676381911
transform 1 0 10272 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  output113
timestamp 1676381911
transform 1 0 9216 0 -1 42336
box -48 -56 432 834
use sg13g2_buf_1  output114
timestamp 1676381911
transform 1 0 9888 0 1 42336
box -48 -56 432 834
use sg13g2_buf_1  output115
timestamp 1676381911
transform 1 0 9888 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  output116
timestamp 1676381911
transform 1 0 10272 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output117
timestamp 1676381911
transform 1 0 10272 0 1 15120
box -48 -56 432 834
use sg13g2_buf_1  output118
timestamp 1676381911
transform 1 0 10272 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  output119
timestamp 1676381911
transform 1 0 9888 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  output120
timestamp 1676381911
transform 1 0 10272 0 1 16632
box -48 -56 432 834
use sg13g2_buf_1  output121
timestamp 1676381911
transform 1 0 10272 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  output122
timestamp 1676381911
transform 1 0 8448 0 1 19656
box -48 -56 432 834
use sg13g2_buf_1  output123
timestamp 1676381911
transform 1 0 8256 0 1 21168
box -48 -56 432 834
use sg13g2_buf_1  output124
timestamp 1676381911
transform 1 0 10272 0 1 21168
box -48 -56 432 834
use sg13g2_buf_1  output125
timestamp 1676381911
transform 1 0 10272 0 -1 22680
box -48 -56 432 834
use sg13g2_buf_1  output126
timestamp 1676381911
transform 1 0 10272 0 1 25704
box -48 -56 432 834
use sg13g2_buf_1  output127
timestamp 1676381911
transform -1 0 3840 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output128
timestamp 1676381911
transform -1 0 6624 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output129
timestamp 1676381911
transform -1 0 7008 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output130
timestamp 1676381911
transform -1 0 7392 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output131
timestamp 1676381911
transform -1 0 7776 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output132
timestamp 1676381911
transform -1 0 8160 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output133
timestamp 1676381911
transform -1 0 8544 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output134
timestamp 1676381911
transform -1 0 8928 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output135
timestamp 1676381911
transform -1 0 9312 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output136
timestamp 1676381911
transform -1 0 9696 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output137
timestamp 1676381911
transform -1 0 10080 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output138
timestamp 1676381911
transform -1 0 5472 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  output139
timestamp 1676381911
transform -1 0 5952 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  output140
timestamp 1676381911
transform -1 0 3840 0 1 42336
box -48 -56 432 834
use sg13g2_buf_1  output141
timestamp 1676381911
transform -1 0 4320 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output142
timestamp 1676381911
transform -1 0 4704 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output143
timestamp 1676381911
transform -1 0 5088 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output144
timestamp 1676381911
transform -1 0 5472 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output145
timestamp 1676381911
transform -1 0 5856 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output146
timestamp 1676381911
transform -1 0 6240 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output147
timestamp 1676381911
transform -1 0 5568 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  output148
timestamp 1676381911
transform -1 0 3456 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output149
timestamp 1676381911
transform -1 0 2688 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output150
timestamp 1676381911
transform -1 0 3072 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output151
timestamp 1676381911
transform -1 0 3456 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output152
timestamp 1676381911
transform -1 0 3456 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output153
timestamp 1676381911
transform -1 0 2688 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output154
timestamp 1676381911
transform -1 0 3840 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output155
timestamp 1676381911
transform -1 0 1536 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output156
timestamp 1676381911
transform -1 0 5760 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output157
timestamp 1676381911
transform -1 0 3072 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output158
timestamp 1676381911
transform -1 0 2304 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output159
timestamp 1676381911
transform -1 0 2688 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output160
timestamp 1676381911
transform -1 0 3072 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output161
timestamp 1676381911
transform -1 0 1536 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output162
timestamp 1676381911
transform -1 0 2304 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output163
timestamp 1676381911
transform -1 0 1920 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output164
timestamp 1676381911
transform -1 0 3840 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output165
timestamp 1676381911
transform -1 0 6912 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output166
timestamp 1676381911
transform -1 0 6528 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output167
timestamp 1676381911
transform -1 0 1920 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output168
timestamp 1676381911
transform -1 0 5184 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  output169
timestamp 1676381911
transform -1 0 3744 0 -1 16632
box -48 -56 432 834
use sg13g2_buf_1  output170
timestamp 1676381911
transform -1 0 1920 0 -1 15120
box -48 -56 432 834
use sg13g2_buf_1  output171
timestamp 1676381911
transform -1 0 5088 0 1 15120
box -48 -56 432 834
use sg13g2_buf_1  output172
timestamp 1676381911
transform -1 0 4320 0 1 15120
box -48 -56 432 834
use sg13g2_buf_1  output173
timestamp 1676381911
transform -1 0 3936 0 1 15120
box -48 -56 432 834
use sg13g2_buf_1  output174
timestamp 1676381911
transform -1 0 2304 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  output175
timestamp 1676381911
transform -1 0 3552 0 1 15120
box -48 -56 432 834
use sg13g2_buf_1  output176
timestamp 1676381911
transform -1 0 1920 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  output177
timestamp 1676381911
transform -1 0 1536 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  output178
timestamp 1676381911
transform -1 0 3168 0 1 15120
box -48 -56 432 834
use sg13g2_buf_1  output179
timestamp 1676381911
transform -1 0 2304 0 -1 15120
box -48 -56 432 834
use sg13g2_buf_1  output180
timestamp 1676381911
transform -1 0 1728 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output181
timestamp 1676381911
transform -1 0 4800 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  output182
timestamp 1676381911
transform -1 0 3936 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  output183
timestamp 1676381911
transform -1 0 1920 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output184
timestamp 1676381911
transform -1 0 1536 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output185
timestamp 1676381911
transform -1 0 1920 0 1 10584
box -48 -56 432 834
use sg13g2_buf_1  output186
timestamp 1676381911
transform -1 0 1536 0 1 10584
box -48 -56 432 834
use sg13g2_buf_1  output187
timestamp 1676381911
transform -1 0 4032 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output188
timestamp 1676381911
transform -1 0 3648 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output189
timestamp 1676381911
transform -1 0 6912 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output190
timestamp 1676381911
transform -1 0 5568 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  output191
timestamp 1676381911
transform -1 0 2304 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output192
timestamp 1676381911
transform -1 0 3936 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output193
timestamp 1676381911
transform -1 0 1920 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output194
timestamp 1676381911
transform -1 0 1536 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output195
timestamp 1676381911
transform -1 0 5184 0 1 12096
box -48 -56 432 834
<< labels >>
flabel metal2 s 11750 1892 11840 1972 0 FreeSans 320 0 0 0 A_I_top
port 0 nsew signal output
flabel metal2 s 11750 884 11840 964 0 FreeSans 320 0 0 0 A_O_top
port 1 nsew signal input
flabel metal2 s 11750 2900 11840 2980 0 FreeSans 320 0 0 0 A_T_top
port 2 nsew signal output
flabel metal2 s 11750 6932 11840 7012 0 FreeSans 320 0 0 0 A_config_C_bit0
port 3 nsew signal output
flabel metal2 s 11750 7940 11840 8020 0 FreeSans 320 0 0 0 A_config_C_bit1
port 4 nsew signal output
flabel metal2 s 11750 8948 11840 9028 0 FreeSans 320 0 0 0 A_config_C_bit2
port 5 nsew signal output
flabel metal2 s 11750 9956 11840 10036 0 FreeSans 320 0 0 0 A_config_C_bit3
port 6 nsew signal output
flabel metal2 s 11750 4916 11840 4996 0 FreeSans 320 0 0 0 B_I_top
port 7 nsew signal output
flabel metal2 s 11750 3908 11840 3988 0 FreeSans 320 0 0 0 B_O_top
port 8 nsew signal input
flabel metal2 s 11750 5924 11840 6004 0 FreeSans 320 0 0 0 B_T_top
port 9 nsew signal output
flabel metal2 s 11750 10964 11840 11044 0 FreeSans 320 0 0 0 B_config_C_bit0
port 10 nsew signal output
flabel metal2 s 11750 11972 11840 12052 0 FreeSans 320 0 0 0 B_config_C_bit1
port 11 nsew signal output
flabel metal2 s 11750 12980 11840 13060 0 FreeSans 320 0 0 0 B_config_C_bit2
port 12 nsew signal output
flabel metal2 s 11750 13988 11840 14068 0 FreeSans 320 0 0 0 B_config_C_bit3
port 13 nsew signal output
flabel metal2 s 0 18356 90 18436 0 FreeSans 320 0 0 0 E1END[0]
port 14 nsew signal input
flabel metal2 s 0 18692 90 18772 0 FreeSans 320 0 0 0 E1END[1]
port 15 nsew signal input
flabel metal2 s 0 19028 90 19108 0 FreeSans 320 0 0 0 E1END[2]
port 16 nsew signal input
flabel metal2 s 0 19364 90 19444 0 FreeSans 320 0 0 0 E1END[3]
port 17 nsew signal input
flabel metal2 s 0 22388 90 22468 0 FreeSans 320 0 0 0 E2END[0]
port 18 nsew signal input
flabel metal2 s 0 22724 90 22804 0 FreeSans 320 0 0 0 E2END[1]
port 19 nsew signal input
flabel metal2 s 0 23060 90 23140 0 FreeSans 320 0 0 0 E2END[2]
port 20 nsew signal input
flabel metal2 s 0 23396 90 23476 0 FreeSans 320 0 0 0 E2END[3]
port 21 nsew signal input
flabel metal2 s 0 23732 90 23812 0 FreeSans 320 0 0 0 E2END[4]
port 22 nsew signal input
flabel metal2 s 0 24068 90 24148 0 FreeSans 320 0 0 0 E2END[5]
port 23 nsew signal input
flabel metal2 s 0 24404 90 24484 0 FreeSans 320 0 0 0 E2END[6]
port 24 nsew signal input
flabel metal2 s 0 24740 90 24820 0 FreeSans 320 0 0 0 E2END[7]
port 25 nsew signal input
flabel metal2 s 0 19700 90 19780 0 FreeSans 320 0 0 0 E2MID[0]
port 26 nsew signal input
flabel metal2 s 0 20036 90 20116 0 FreeSans 320 0 0 0 E2MID[1]
port 27 nsew signal input
flabel metal2 s 0 20372 90 20452 0 FreeSans 320 0 0 0 E2MID[2]
port 28 nsew signal input
flabel metal2 s 0 20708 90 20788 0 FreeSans 320 0 0 0 E2MID[3]
port 29 nsew signal input
flabel metal2 s 0 21044 90 21124 0 FreeSans 320 0 0 0 E2MID[4]
port 30 nsew signal input
flabel metal2 s 0 21380 90 21460 0 FreeSans 320 0 0 0 E2MID[5]
port 31 nsew signal input
flabel metal2 s 0 21716 90 21796 0 FreeSans 320 0 0 0 E2MID[6]
port 32 nsew signal input
flabel metal2 s 0 22052 90 22132 0 FreeSans 320 0 0 0 E2MID[7]
port 33 nsew signal input
flabel metal2 s 0 30452 90 30532 0 FreeSans 320 0 0 0 E6END[0]
port 34 nsew signal input
flabel metal2 s 0 33812 90 33892 0 FreeSans 320 0 0 0 E6END[10]
port 35 nsew signal input
flabel metal2 s 0 34148 90 34228 0 FreeSans 320 0 0 0 E6END[11]
port 36 nsew signal input
flabel metal2 s 0 30788 90 30868 0 FreeSans 320 0 0 0 E6END[1]
port 37 nsew signal input
flabel metal2 s 0 31124 90 31204 0 FreeSans 320 0 0 0 E6END[2]
port 38 nsew signal input
flabel metal2 s 0 31460 90 31540 0 FreeSans 320 0 0 0 E6END[3]
port 39 nsew signal input
flabel metal2 s 0 31796 90 31876 0 FreeSans 320 0 0 0 E6END[4]
port 40 nsew signal input
flabel metal2 s 0 32132 90 32212 0 FreeSans 320 0 0 0 E6END[5]
port 41 nsew signal input
flabel metal2 s 0 32468 90 32548 0 FreeSans 320 0 0 0 E6END[6]
port 42 nsew signal input
flabel metal2 s 0 32804 90 32884 0 FreeSans 320 0 0 0 E6END[7]
port 43 nsew signal input
flabel metal2 s 0 33140 90 33220 0 FreeSans 320 0 0 0 E6END[8]
port 44 nsew signal input
flabel metal2 s 0 33476 90 33556 0 FreeSans 320 0 0 0 E6END[9]
port 45 nsew signal input
flabel metal2 s 0 25076 90 25156 0 FreeSans 320 0 0 0 EE4END[0]
port 46 nsew signal input
flabel metal2 s 0 28436 90 28516 0 FreeSans 320 0 0 0 EE4END[10]
port 47 nsew signal input
flabel metal2 s 0 28772 90 28852 0 FreeSans 320 0 0 0 EE4END[11]
port 48 nsew signal input
flabel metal2 s 0 29108 90 29188 0 FreeSans 320 0 0 0 EE4END[12]
port 49 nsew signal input
flabel metal2 s 0 29444 90 29524 0 FreeSans 320 0 0 0 EE4END[13]
port 50 nsew signal input
flabel metal2 s 0 29780 90 29860 0 FreeSans 320 0 0 0 EE4END[14]
port 51 nsew signal input
flabel metal2 s 0 30116 90 30196 0 FreeSans 320 0 0 0 EE4END[15]
port 52 nsew signal input
flabel metal2 s 0 25412 90 25492 0 FreeSans 320 0 0 0 EE4END[1]
port 53 nsew signal input
flabel metal2 s 0 25748 90 25828 0 FreeSans 320 0 0 0 EE4END[2]
port 54 nsew signal input
flabel metal2 s 0 26084 90 26164 0 FreeSans 320 0 0 0 EE4END[3]
port 55 nsew signal input
flabel metal2 s 0 26420 90 26500 0 FreeSans 320 0 0 0 EE4END[4]
port 56 nsew signal input
flabel metal2 s 0 26756 90 26836 0 FreeSans 320 0 0 0 EE4END[5]
port 57 nsew signal input
flabel metal2 s 0 27092 90 27172 0 FreeSans 320 0 0 0 EE4END[6]
port 58 nsew signal input
flabel metal2 s 0 27428 90 27508 0 FreeSans 320 0 0 0 EE4END[7]
port 59 nsew signal input
flabel metal2 s 0 27764 90 27844 0 FreeSans 320 0 0 0 EE4END[8]
port 60 nsew signal input
flabel metal2 s 0 28100 90 28180 0 FreeSans 320 0 0 0 EE4END[9]
port 61 nsew signal input
flabel metal2 s 0 34484 90 34564 0 FreeSans 320 0 0 0 FrameData[0]
port 62 nsew signal input
flabel metal2 s 0 37844 90 37924 0 FreeSans 320 0 0 0 FrameData[10]
port 63 nsew signal input
flabel metal2 s 0 38180 90 38260 0 FreeSans 320 0 0 0 FrameData[11]
port 64 nsew signal input
flabel metal2 s 0 38516 90 38596 0 FreeSans 320 0 0 0 FrameData[12]
port 65 nsew signal input
flabel metal2 s 0 38852 90 38932 0 FreeSans 320 0 0 0 FrameData[13]
port 66 nsew signal input
flabel metal2 s 0 39188 90 39268 0 FreeSans 320 0 0 0 FrameData[14]
port 67 nsew signal input
flabel metal2 s 0 39524 90 39604 0 FreeSans 320 0 0 0 FrameData[15]
port 68 nsew signal input
flabel metal2 s 0 39860 90 39940 0 FreeSans 320 0 0 0 FrameData[16]
port 69 nsew signal input
flabel metal2 s 0 40196 90 40276 0 FreeSans 320 0 0 0 FrameData[17]
port 70 nsew signal input
flabel metal2 s 0 40532 90 40612 0 FreeSans 320 0 0 0 FrameData[18]
port 71 nsew signal input
flabel metal2 s 0 40868 90 40948 0 FreeSans 320 0 0 0 FrameData[19]
port 72 nsew signal input
flabel metal2 s 0 34820 90 34900 0 FreeSans 320 0 0 0 FrameData[1]
port 73 nsew signal input
flabel metal2 s 0 41204 90 41284 0 FreeSans 320 0 0 0 FrameData[20]
port 74 nsew signal input
flabel metal2 s 0 41540 90 41620 0 FreeSans 320 0 0 0 FrameData[21]
port 75 nsew signal input
flabel metal2 s 0 41876 90 41956 0 FreeSans 320 0 0 0 FrameData[22]
port 76 nsew signal input
flabel metal2 s 0 42212 90 42292 0 FreeSans 320 0 0 0 FrameData[23]
port 77 nsew signal input
flabel metal2 s 0 42548 90 42628 0 FreeSans 320 0 0 0 FrameData[24]
port 78 nsew signal input
flabel metal2 s 0 42884 90 42964 0 FreeSans 320 0 0 0 FrameData[25]
port 79 nsew signal input
flabel metal2 s 0 43220 90 43300 0 FreeSans 320 0 0 0 FrameData[26]
port 80 nsew signal input
flabel metal2 s 0 43556 90 43636 0 FreeSans 320 0 0 0 FrameData[27]
port 81 nsew signal input
flabel metal2 s 0 43892 90 43972 0 FreeSans 320 0 0 0 FrameData[28]
port 82 nsew signal input
flabel metal2 s 0 44228 90 44308 0 FreeSans 320 0 0 0 FrameData[29]
port 83 nsew signal input
flabel metal2 s 0 35156 90 35236 0 FreeSans 320 0 0 0 FrameData[2]
port 84 nsew signal input
flabel metal2 s 0 44564 90 44644 0 FreeSans 320 0 0 0 FrameData[30]
port 85 nsew signal input
flabel metal2 s 0 44900 90 44980 0 FreeSans 320 0 0 0 FrameData[31]
port 86 nsew signal input
flabel metal2 s 0 35492 90 35572 0 FreeSans 320 0 0 0 FrameData[3]
port 87 nsew signal input
flabel metal2 s 0 35828 90 35908 0 FreeSans 320 0 0 0 FrameData[4]
port 88 nsew signal input
flabel metal2 s 0 36164 90 36244 0 FreeSans 320 0 0 0 FrameData[5]
port 89 nsew signal input
flabel metal2 s 0 36500 90 36580 0 FreeSans 320 0 0 0 FrameData[6]
port 90 nsew signal input
flabel metal2 s 0 36836 90 36916 0 FreeSans 320 0 0 0 FrameData[7]
port 91 nsew signal input
flabel metal2 s 0 37172 90 37252 0 FreeSans 320 0 0 0 FrameData[8]
port 92 nsew signal input
flabel metal2 s 0 37508 90 37588 0 FreeSans 320 0 0 0 FrameData[9]
port 93 nsew signal input
flabel metal2 s 11750 14996 11840 15076 0 FreeSans 320 0 0 0 FrameData_O[0]
port 94 nsew signal output
flabel metal2 s 11750 25076 11840 25156 0 FreeSans 320 0 0 0 FrameData_O[10]
port 95 nsew signal output
flabel metal2 s 11750 26084 11840 26164 0 FreeSans 320 0 0 0 FrameData_O[11]
port 96 nsew signal output
flabel metal2 s 11750 27092 11840 27172 0 FreeSans 320 0 0 0 FrameData_O[12]
port 97 nsew signal output
flabel metal2 s 11750 28100 11840 28180 0 FreeSans 320 0 0 0 FrameData_O[13]
port 98 nsew signal output
flabel metal2 s 11750 29108 11840 29188 0 FreeSans 320 0 0 0 FrameData_O[14]
port 99 nsew signal output
flabel metal2 s 11750 30116 11840 30196 0 FreeSans 320 0 0 0 FrameData_O[15]
port 100 nsew signal output
flabel metal2 s 11750 31124 11840 31204 0 FreeSans 320 0 0 0 FrameData_O[16]
port 101 nsew signal output
flabel metal2 s 11750 32132 11840 32212 0 FreeSans 320 0 0 0 FrameData_O[17]
port 102 nsew signal output
flabel metal2 s 11750 33140 11840 33220 0 FreeSans 320 0 0 0 FrameData_O[18]
port 103 nsew signal output
flabel metal2 s 11750 34148 11840 34228 0 FreeSans 320 0 0 0 FrameData_O[19]
port 104 nsew signal output
flabel metal2 s 11750 16004 11840 16084 0 FreeSans 320 0 0 0 FrameData_O[1]
port 105 nsew signal output
flabel metal2 s 11750 35156 11840 35236 0 FreeSans 320 0 0 0 FrameData_O[20]
port 106 nsew signal output
flabel metal2 s 11750 36164 11840 36244 0 FreeSans 320 0 0 0 FrameData_O[21]
port 107 nsew signal output
flabel metal2 s 11750 37172 11840 37252 0 FreeSans 320 0 0 0 FrameData_O[22]
port 108 nsew signal output
flabel metal2 s 11750 38180 11840 38260 0 FreeSans 320 0 0 0 FrameData_O[23]
port 109 nsew signal output
flabel metal2 s 11750 39188 11840 39268 0 FreeSans 320 0 0 0 FrameData_O[24]
port 110 nsew signal output
flabel metal2 s 11750 40196 11840 40276 0 FreeSans 320 0 0 0 FrameData_O[25]
port 111 nsew signal output
flabel metal2 s 11750 41204 11840 41284 0 FreeSans 320 0 0 0 FrameData_O[26]
port 112 nsew signal output
flabel metal2 s 11750 42212 11840 42292 0 FreeSans 320 0 0 0 FrameData_O[27]
port 113 nsew signal output
flabel metal2 s 11750 43220 11840 43300 0 FreeSans 320 0 0 0 FrameData_O[28]
port 114 nsew signal output
flabel metal2 s 11750 44228 11840 44308 0 FreeSans 320 0 0 0 FrameData_O[29]
port 115 nsew signal output
flabel metal2 s 11750 17012 11840 17092 0 FreeSans 320 0 0 0 FrameData_O[2]
port 116 nsew signal output
flabel metal2 s 11750 45236 11840 45316 0 FreeSans 320 0 0 0 FrameData_O[30]
port 117 nsew signal output
flabel metal2 s 11750 46244 11840 46324 0 FreeSans 320 0 0 0 FrameData_O[31]
port 118 nsew signal output
flabel metal2 s 11750 18020 11840 18100 0 FreeSans 320 0 0 0 FrameData_O[3]
port 119 nsew signal output
flabel metal2 s 11750 19028 11840 19108 0 FreeSans 320 0 0 0 FrameData_O[4]
port 120 nsew signal output
flabel metal2 s 11750 20036 11840 20116 0 FreeSans 320 0 0 0 FrameData_O[5]
port 121 nsew signal output
flabel metal2 s 11750 21044 11840 21124 0 FreeSans 320 0 0 0 FrameData_O[6]
port 122 nsew signal output
flabel metal2 s 11750 22052 11840 22132 0 FreeSans 320 0 0 0 FrameData_O[7]
port 123 nsew signal output
flabel metal2 s 11750 23060 11840 23140 0 FreeSans 320 0 0 0 FrameData_O[8]
port 124 nsew signal output
flabel metal2 s 11750 24068 11840 24148 0 FreeSans 320 0 0 0 FrameData_O[9]
port 125 nsew signal output
flabel metal3 s 2360 0 2440 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 126 nsew signal input
flabel metal3 s 6200 0 6280 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 127 nsew signal input
flabel metal3 s 6584 0 6664 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 128 nsew signal input
flabel metal3 s 6968 0 7048 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 129 nsew signal input
flabel metal3 s 7352 0 7432 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 130 nsew signal input
flabel metal3 s 7736 0 7816 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 131 nsew signal input
flabel metal3 s 8120 0 8200 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 132 nsew signal input
flabel metal3 s 8504 0 8584 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 133 nsew signal input
flabel metal3 s 8888 0 8968 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 134 nsew signal input
flabel metal3 s 9272 0 9352 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 135 nsew signal input
flabel metal3 s 9656 0 9736 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 136 nsew signal input
flabel metal3 s 2744 0 2824 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 137 nsew signal input
flabel metal3 s 3128 0 3208 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 138 nsew signal input
flabel metal3 s 3512 0 3592 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 139 nsew signal input
flabel metal3 s 3896 0 3976 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 140 nsew signal input
flabel metal3 s 4280 0 4360 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 141 nsew signal input
flabel metal3 s 4664 0 4744 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 142 nsew signal input
flabel metal3 s 5048 0 5128 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 143 nsew signal input
flabel metal3 s 5432 0 5512 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 144 nsew signal input
flabel metal3 s 5816 0 5896 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 145 nsew signal input
flabel metal3 s 2360 47280 2440 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 146 nsew signal output
flabel metal3 s 6200 47280 6280 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 147 nsew signal output
flabel metal3 s 6584 47280 6664 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 148 nsew signal output
flabel metal3 s 6968 47280 7048 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 149 nsew signal output
flabel metal3 s 7352 47280 7432 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 150 nsew signal output
flabel metal3 s 7736 47280 7816 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 151 nsew signal output
flabel metal3 s 8120 47280 8200 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 152 nsew signal output
flabel metal3 s 8504 47280 8584 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 153 nsew signal output
flabel metal3 s 8888 47280 8968 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 154 nsew signal output
flabel metal3 s 9272 47280 9352 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 155 nsew signal output
flabel metal3 s 9656 47280 9736 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 156 nsew signal output
flabel metal3 s 2744 47280 2824 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 157 nsew signal output
flabel metal3 s 3128 47280 3208 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 158 nsew signal output
flabel metal3 s 3512 47280 3592 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 159 nsew signal output
flabel metal3 s 3896 47280 3976 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 160 nsew signal output
flabel metal3 s 4280 47280 4360 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 161 nsew signal output
flabel metal3 s 4664 47280 4744 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 162 nsew signal output
flabel metal3 s 5048 47280 5128 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 163 nsew signal output
flabel metal3 s 5432 47280 5512 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 164 nsew signal output
flabel metal3 s 5816 47280 5896 47360 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 165 nsew signal output
flabel metal3 s 1976 0 2056 80 0 FreeSans 320 0 0 0 UserCLK
port 166 nsew signal input
flabel metal3 s 1976 47280 2056 47360 0 FreeSans 320 0 0 0 UserCLKo
port 167 nsew signal output
flabel metal5 s 4892 0 5332 47360 0 FreeSans 2560 90 0 0 VGND
port 168 nsew ground bidirectional
flabel metal5 s 4892 0 5332 40 0 FreeSans 320 0 0 0 VGND
port 168 nsew ground bidirectional
flabel metal5 s 4892 47320 5332 47360 0 FreeSans 320 0 0 0 VGND
port 168 nsew ground bidirectional
flabel metal5 s 3652 0 4092 47360 0 FreeSans 2560 90 0 0 VPWR
port 169 nsew power bidirectional
flabel metal5 s 3652 0 4092 40 0 FreeSans 320 0 0 0 VPWR
port 169 nsew power bidirectional
flabel metal5 s 3652 47320 4092 47360 0 FreeSans 320 0 0 0 VPWR
port 169 nsew power bidirectional
flabel metal2 s 0 2228 90 2308 0 FreeSans 320 0 0 0 W1BEG[0]
port 170 nsew signal output
flabel metal2 s 0 2564 90 2644 0 FreeSans 320 0 0 0 W1BEG[1]
port 171 nsew signal output
flabel metal2 s 0 2900 90 2980 0 FreeSans 320 0 0 0 W1BEG[2]
port 172 nsew signal output
flabel metal2 s 0 3236 90 3316 0 FreeSans 320 0 0 0 W1BEG[3]
port 173 nsew signal output
flabel metal2 s 0 3572 90 3652 0 FreeSans 320 0 0 0 W2BEG[0]
port 174 nsew signal output
flabel metal2 s 0 3908 90 3988 0 FreeSans 320 0 0 0 W2BEG[1]
port 175 nsew signal output
flabel metal2 s 0 4244 90 4324 0 FreeSans 320 0 0 0 W2BEG[2]
port 176 nsew signal output
flabel metal2 s 0 4580 90 4660 0 FreeSans 320 0 0 0 W2BEG[3]
port 177 nsew signal output
flabel metal2 s 0 4916 90 4996 0 FreeSans 320 0 0 0 W2BEG[4]
port 178 nsew signal output
flabel metal2 s 0 5252 90 5332 0 FreeSans 320 0 0 0 W2BEG[5]
port 179 nsew signal output
flabel metal2 s 0 5588 90 5668 0 FreeSans 320 0 0 0 W2BEG[6]
port 180 nsew signal output
flabel metal2 s 0 5924 90 6004 0 FreeSans 320 0 0 0 W2BEG[7]
port 181 nsew signal output
flabel metal2 s 0 6260 90 6340 0 FreeSans 320 0 0 0 W2BEGb[0]
port 182 nsew signal output
flabel metal2 s 0 6596 90 6676 0 FreeSans 320 0 0 0 W2BEGb[1]
port 183 nsew signal output
flabel metal2 s 0 6932 90 7012 0 FreeSans 320 0 0 0 W2BEGb[2]
port 184 nsew signal output
flabel metal2 s 0 7268 90 7348 0 FreeSans 320 0 0 0 W2BEGb[3]
port 185 nsew signal output
flabel metal2 s 0 7604 90 7684 0 FreeSans 320 0 0 0 W2BEGb[4]
port 186 nsew signal output
flabel metal2 s 0 7940 90 8020 0 FreeSans 320 0 0 0 W2BEGb[5]
port 187 nsew signal output
flabel metal2 s 0 8276 90 8356 0 FreeSans 320 0 0 0 W2BEGb[6]
port 188 nsew signal output
flabel metal2 s 0 8612 90 8692 0 FreeSans 320 0 0 0 W2BEGb[7]
port 189 nsew signal output
flabel metal2 s 0 14324 90 14404 0 FreeSans 320 0 0 0 W6BEG[0]
port 190 nsew signal output
flabel metal2 s 0 17684 90 17764 0 FreeSans 320 0 0 0 W6BEG[10]
port 191 nsew signal output
flabel metal2 s 0 18020 90 18100 0 FreeSans 320 0 0 0 W6BEG[11]
port 192 nsew signal output
flabel metal2 s 0 14660 90 14740 0 FreeSans 320 0 0 0 W6BEG[1]
port 193 nsew signal output
flabel metal2 s 0 14996 90 15076 0 FreeSans 320 0 0 0 W6BEG[2]
port 194 nsew signal output
flabel metal2 s 0 15332 90 15412 0 FreeSans 320 0 0 0 W6BEG[3]
port 195 nsew signal output
flabel metal2 s 0 15668 90 15748 0 FreeSans 320 0 0 0 W6BEG[4]
port 196 nsew signal output
flabel metal2 s 0 16004 90 16084 0 FreeSans 320 0 0 0 W6BEG[5]
port 197 nsew signal output
flabel metal2 s 0 16340 90 16420 0 FreeSans 320 0 0 0 W6BEG[6]
port 198 nsew signal output
flabel metal2 s 0 16676 90 16756 0 FreeSans 320 0 0 0 W6BEG[7]
port 199 nsew signal output
flabel metal2 s 0 17012 90 17092 0 FreeSans 320 0 0 0 W6BEG[8]
port 200 nsew signal output
flabel metal2 s 0 17348 90 17428 0 FreeSans 320 0 0 0 W6BEG[9]
port 201 nsew signal output
flabel metal2 s 0 8948 90 9028 0 FreeSans 320 0 0 0 WW4BEG[0]
port 202 nsew signal output
flabel metal2 s 0 12308 90 12388 0 FreeSans 320 0 0 0 WW4BEG[10]
port 203 nsew signal output
flabel metal2 s 0 12644 90 12724 0 FreeSans 320 0 0 0 WW4BEG[11]
port 204 nsew signal output
flabel metal2 s 0 12980 90 13060 0 FreeSans 320 0 0 0 WW4BEG[12]
port 205 nsew signal output
flabel metal2 s 0 13316 90 13396 0 FreeSans 320 0 0 0 WW4BEG[13]
port 206 nsew signal output
flabel metal2 s 0 13652 90 13732 0 FreeSans 320 0 0 0 WW4BEG[14]
port 207 nsew signal output
flabel metal2 s 0 13988 90 14068 0 FreeSans 320 0 0 0 WW4BEG[15]
port 208 nsew signal output
flabel metal2 s 0 9284 90 9364 0 FreeSans 320 0 0 0 WW4BEG[1]
port 209 nsew signal output
flabel metal2 s 0 9620 90 9700 0 FreeSans 320 0 0 0 WW4BEG[2]
port 210 nsew signal output
flabel metal2 s 0 9956 90 10036 0 FreeSans 320 0 0 0 WW4BEG[3]
port 211 nsew signal output
flabel metal2 s 0 10292 90 10372 0 FreeSans 320 0 0 0 WW4BEG[4]
port 212 nsew signal output
flabel metal2 s 0 10628 90 10708 0 FreeSans 320 0 0 0 WW4BEG[5]
port 213 nsew signal output
flabel metal2 s 0 10964 90 11044 0 FreeSans 320 0 0 0 WW4BEG[6]
port 214 nsew signal output
flabel metal2 s 0 11300 90 11380 0 FreeSans 320 0 0 0 WW4BEG[7]
port 215 nsew signal output
flabel metal2 s 0 11636 90 11716 0 FreeSans 320 0 0 0 WW4BEG[8]
port 216 nsew signal output
flabel metal2 s 0 11972 90 12052 0 FreeSans 320 0 0 0 WW4BEG[9]
port 217 nsew signal output
rlabel metal1 5904 45360 5904 45360 0 VGND
rlabel metal1 5904 44604 5904 44604 0 VPWR
rlabel metal2 11750 1932 11750 1932 0 A_I_top
rlabel metal2 11126 924 11126 924 0 A_O_top
rlabel metal2 11750 2940 11750 2940 0 A_T_top
rlabel metal2 10608 6804 10608 6804 0 A_config_C_bit0
rlabel metal2 11030 7980 11030 7980 0 A_config_C_bit1
rlabel metal2 10632 7056 10632 7056 0 A_config_C_bit2
rlabel metal2 11270 9996 11270 9996 0 A_config_C_bit3
rlabel metal2 11750 4956 11750 4956 0 B_I_top
rlabel metal2 10848 4200 10848 4200 0 B_O_top
rlabel metal2 11750 5964 11750 5964 0 B_T_top
rlabel metal2 10248 10416 10248 10416 0 B_config_C_bit0
rlabel metal2 10632 10416 10632 10416 0 B_config_C_bit1
rlabel metal2 11078 13020 11078 13020 0 B_config_C_bit2
rlabel metal2 11414 14028 11414 14028 0 B_config_C_bit3
rlabel metal2 512 18396 512 18396 0 E1END[0]
rlabel metal2 416 18732 416 18732 0 E1END[1]
rlabel metal2 752 19068 752 19068 0 E1END[2]
rlabel metal2 512 19404 512 19404 0 E1END[3]
rlabel via2 80 22428 80 22428 0 E2END[0]
rlabel metal2 656 22764 656 22764 0 E2END[1]
rlabel metal2 368 23100 368 23100 0 E2END[2]
rlabel metal2 1472 23436 1472 23436 0 E2END[3]
rlabel metal2 840 21504 840 21504 0 E2END[4]
rlabel metal2 416 24108 416 24108 0 E2END[5]
rlabel metal2 936 23016 936 23016 0 E2END[6]
rlabel metal2 368 24780 368 24780 0 E2END[7]
rlabel metal2 320 19740 320 19740 0 E2MID[0]
rlabel metal2 800 20076 800 20076 0 E2MID[1]
rlabel metal2 656 20412 656 20412 0 E2MID[2]
rlabel metal2 272 20748 272 20748 0 E2MID[3]
rlabel metal2 176 21084 176 21084 0 E2MID[4]
rlabel metal2 368 21420 368 21420 0 E2MID[5]
rlabel metal2 224 21756 224 21756 0 E2MID[6]
rlabel metal2 320 22092 320 22092 0 E2MID[7]
rlabel metal2 984 33600 984 33600 0 E6END[0]
rlabel metal2 800 33852 800 33852 0 E6END[10]
rlabel via2 80 34188 80 34188 0 E6END[11]
rlabel metal2 704 30828 704 30828 0 E6END[1]
rlabel metal2 656 31164 656 31164 0 E6END[2]
rlabel metal2 992 31500 992 31500 0 E6END[3]
rlabel metal2 2624 31836 2624 31836 0 E6END[4]
rlabel metal2 864 35952 864 35952 0 E6END[5]
rlabel metal2 1536 35952 1536 35952 0 E6END[6]
rlabel metal2 2016 35952 2016 35952 0 E6END[7]
rlabel metal2 80 33180 80 33180 0 E6END[8]
rlabel metal2 944 33516 944 33516 0 E6END[9]
rlabel metal2 656 25116 656 25116 0 EE4END[0]
rlabel metal2 80 28476 80 28476 0 EE4END[10]
rlabel metal2 896 28812 896 28812 0 EE4END[11]
rlabel metal2 800 29148 800 29148 0 EE4END[12]
rlabel metal2 1472 29484 1472 29484 0 EE4END[13]
rlabel metal2 704 29820 704 29820 0 EE4END[14]
rlabel metal2 752 30156 752 30156 0 EE4END[15]
rlabel metal2 224 25452 224 25452 0 EE4END[1]
rlabel metal2 800 25788 800 25788 0 EE4END[2]
rlabel metal2 416 26124 416 26124 0 EE4END[3]
rlabel metal2 800 26460 800 26460 0 EE4END[4]
rlabel metal2 176 26796 176 26796 0 EE4END[5]
rlabel metal2 704 27132 704 27132 0 EE4END[6]
rlabel metal2 560 27468 560 27468 0 EE4END[7]
rlabel metal2 560 27804 560 27804 0 EE4END[8]
rlabel metal2 272 28140 272 28140 0 EE4END[9]
rlabel metal2 560 34524 560 34524 0 FrameData[0]
rlabel metal2 1040 37884 1040 37884 0 FrameData[10]
rlabel metal2 800 38220 800 38220 0 FrameData[11]
rlabel metal2 1472 38556 1472 38556 0 FrameData[12]
rlabel metal2 800 38892 800 38892 0 FrameData[13]
rlabel metal2 704 39228 704 39228 0 FrameData[14]
rlabel metal2 464 39564 464 39564 0 FrameData[15]
rlabel metal2 176 39900 176 39900 0 FrameData[16]
rlabel metal2 560 40236 560 40236 0 FrameData[17]
rlabel metal2 944 40572 944 40572 0 FrameData[18]
rlabel metal2 704 40908 704 40908 0 FrameData[19]
rlabel metal2 3264 34944 3264 34944 0 FrameData[1]
rlabel metal2 560 41244 560 41244 0 FrameData[20]
rlabel metal2 1136 41580 1136 41580 0 FrameData[21]
rlabel metal2 1472 41916 1472 41916 0 FrameData[22]
rlabel metal2 368 42252 368 42252 0 FrameData[23]
rlabel metal2 944 42588 944 42588 0 FrameData[24]
rlabel metal2 704 42924 704 42924 0 FrameData[25]
rlabel metal2 464 43260 464 43260 0 FrameData[26]
rlabel metal2 656 43596 656 43596 0 FrameData[27]
rlabel via2 80 43932 80 43932 0 FrameData[28]
rlabel via2 80 44268 80 44268 0 FrameData[29]
rlabel metal2 560 35196 560 35196 0 FrameData[2]
rlabel metal2 1376 44604 1376 44604 0 FrameData[30]
rlabel metal2 752 44940 752 44940 0 FrameData[31]
rlabel metal2 656 35532 656 35532 0 FrameData[3]
rlabel metal2 128 35868 128 35868 0 FrameData[4]
rlabel metal3 3072 37590 3072 37590 0 FrameData[5]
rlabel metal2 800 36540 800 36540 0 FrameData[6]
rlabel metal2 704 36876 704 36876 0 FrameData[7]
rlabel metal2 128 37212 128 37212 0 FrameData[8]
rlabel metal2 224 37548 224 37548 0 FrameData[9]
rlabel metal2 10632 14196 10632 14196 0 FrameData_O[0]
rlabel metal2 11198 25116 11198 25116 0 FrameData_O[10]
rlabel metal2 11414 26124 11414 26124 0 FrameData_O[11]
rlabel metal2 11654 27132 11654 27132 0 FrameData_O[12]
rlabel metal2 9600 28770 9600 28770 0 FrameData_O[13]
rlabel metal2 11318 29148 11318 29148 0 FrameData_O[14]
rlabel metal2 11510 30156 11510 30156 0 FrameData_O[15]
rlabel metal2 11414 31164 11414 31164 0 FrameData_O[16]
rlabel metal2 11318 32172 11318 32172 0 FrameData_O[17]
rlabel metal2 11510 33180 11510 33180 0 FrameData_O[18]
rlabel metal2 11462 34188 11462 34188 0 FrameData_O[19]
rlabel metal2 10680 14952 10680 14952 0 FrameData_O[1]
rlabel metal2 11414 35196 11414 35196 0 FrameData_O[20]
rlabel metal2 11654 36204 11654 36204 0 FrameData_O[21]
rlabel metal2 11462 37212 11462 37212 0 FrameData_O[22]
rlabel metal2 11414 38220 11414 38220 0 FrameData_O[23]
rlabel metal2 11510 39228 11510 39228 0 FrameData_O[24]
rlabel metal2 11366 40236 11366 40236 0 FrameData_O[25]
rlabel metal2 11750 41244 11750 41244 0 FrameData_O[26]
rlabel metal2 11750 42252 11750 42252 0 FrameData_O[27]
rlabel metal2 11414 43260 11414 43260 0 FrameData_O[28]
rlabel metal2 11750 44268 11750 44268 0 FrameData_O[29]
rlabel metal2 10920 15708 10920 15708 0 FrameData_O[2]
rlabel metal2 10824 44436 10824 44436 0 FrameData_O[30]
rlabel metal2 10248 44436 10248 44436 0 FrameData_O[31]
rlabel metal2 10680 17220 10680 17220 0 FrameData_O[3]
rlabel metal2 10632 17976 10632 17976 0 FrameData_O[4]
rlabel metal2 11030 20076 11030 20076 0 FrameData_O[5]
rlabel metal2 10214 21084 10214 21084 0 FrameData_O[6]
rlabel metal2 10608 21924 10608 21924 0 FrameData_O[7]
rlabel metal2 10632 22512 10632 22512 0 FrameData_O[8]
rlabel metal2 11606 24108 11606 24108 0 FrameData_O[9]
rlabel metal3 2400 11550 2400 11550 0 FrameStrobe[0]
rlabel metal3 6240 72 6240 72 0 FrameStrobe[10]
rlabel metal3 7488 18018 7488 18018 0 FrameStrobe[11]
rlabel metal3 7008 72 7008 72 0 FrameStrobe[12]
rlabel metal3 7392 744 7392 744 0 FrameStrobe[13]
rlabel metal3 7776 1206 7776 1206 0 FrameStrobe[14]
rlabel metal3 8160 744 8160 744 0 FrameStrobe[15]
rlabel metal2 7488 21000 7488 21000 0 FrameStrobe[16]
rlabel metal3 8928 744 8928 744 0 FrameStrobe[17]
rlabel metal2 8976 19236 8976 19236 0 FrameStrobe[18]
rlabel metal2 10752 42000 10752 42000 0 FrameStrobe[19]
rlabel metal3 2784 156 2784 156 0 FrameStrobe[1]
rlabel metal4 5424 20244 5424 20244 0 FrameStrobe[2]
rlabel metal2 6480 19824 6480 19824 0 FrameStrobe[3]
rlabel metal3 3936 114 3936 114 0 FrameStrobe[4]
rlabel metal4 4944 4116 4944 4116 0 FrameStrobe[5]
rlabel metal3 1824 20076 1824 20076 0 FrameStrobe[6]
rlabel metal3 5088 702 5088 702 0 FrameStrobe[7]
rlabel metal2 1728 27174 1728 27174 0 FrameStrobe[8]
rlabel metal3 5856 114 5856 114 0 FrameStrobe[9]
rlabel metal3 2400 46246 2400 46246 0 FrameStrobe_O[0]
rlabel metal2 6264 45192 6264 45192 0 FrameStrobe_O[10]
rlabel metal2 6648 45192 6648 45192 0 FrameStrobe_O[11]
rlabel metal2 7032 45192 7032 45192 0 FrameStrobe_O[12]
rlabel metal2 7416 45192 7416 45192 0 FrameStrobe_O[13]
rlabel metal2 7800 45192 7800 45192 0 FrameStrobe_O[14]
rlabel metal2 8184 45192 8184 45192 0 FrameStrobe_O[15]
rlabel metal2 8568 45192 8568 45192 0 FrameStrobe_O[16]
rlabel metal2 8952 45192 8952 45192 0 FrameStrobe_O[17]
rlabel metal2 9336 45192 9336 45192 0 FrameStrobe_O[18]
rlabel metal2 9720 45192 9720 45192 0 FrameStrobe_O[19]
rlabel metal3 2784 46120 2784 46120 0 FrameStrobe_O[1]
rlabel metal2 5544 44436 5544 44436 0 FrameStrobe_O[2]
rlabel metal2 3528 42924 3528 42924 0 FrameStrobe_O[3]
rlabel metal2 3960 45192 3960 45192 0 FrameStrobe_O[4]
rlabel metal2 4344 45192 4344 45192 0 FrameStrobe_O[5]
rlabel metal2 4728 45192 4728 45192 0 FrameStrobe_O[6]
rlabel metal2 5256 45192 5256 45192 0 FrameStrobe_O[7]
rlabel metal2 5496 45108 5496 45108 0 FrameStrobe_O[8]
rlabel metal2 5880 45192 5880 45192 0 FrameStrobe_O[9]
rlabel metal4 9696 18144 9696 18144 0 Inst_A_IO_1_bidirectional_frame_config_pass.Q
rlabel metal3 9360 17976 9360 17976 0 Inst_B_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 3840 40530 3840 40530 0 Inst_E_IO_ConfigMem.Inst_frame0_bit0.Q
rlabel metal3 5376 39900 5376 39900 0 Inst_E_IO_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 3264 33432 3264 33432 0 Inst_E_IO_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 5328 32928 5328 32928 0 Inst_E_IO_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 3024 35364 3024 35364 0 Inst_E_IO_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 5328 35364 5328 35364 0 Inst_E_IO_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 6960 4368 6960 4368 0 Inst_E_IO_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 8304 5712 8304 5712 0 Inst_E_IO_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 6432 9366 6432 9366 0 Inst_E_IO_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 8352 8904 8352 8904 0 Inst_E_IO_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 4992 21462 4992 21462 0 Inst_E_IO_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 5952 21588 5952 21588 0 Inst_E_IO_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 7872 14826 7872 14826 0 Inst_E_IO_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 6144 19908 6144 19908 0 Inst_E_IO_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 5952 20874 5952 20874 0 Inst_E_IO_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 5225 16968 5225 16968 0 Inst_E_IO_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 4032 17052 4032 17052 0 Inst_E_IO_ConfigMem.Inst_frame0_bit23.Q
rlabel metal3 3936 16926 3936 16926 0 Inst_E_IO_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 4032 25326 4032 25326 0 Inst_E_IO_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 3840 23814 3840 23814 0 Inst_E_IO_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 5136 23856 5136 23856 0 Inst_E_IO_ConfigMem.Inst_frame0_bit27.Q
rlabel metal5 2784 34118 2784 34118 0 Inst_E_IO_ConfigMem.Inst_frame0_bit28.Q
rlabel metal3 3120 33432 3120 33432 0 Inst_E_IO_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 9312 14196 9312 14196 0 Inst_E_IO_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 3360 30156 3360 30156 0 Inst_E_IO_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 2928 30408 2928 30408 0 Inst_E_IO_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 7200 17808 7200 17808 0 Inst_E_IO_ConfigMem.Inst_frame0_bit4.Q
rlabel metal3 9312 17514 9312 17514 0 Inst_E_IO_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 3792 4368 3792 4368 0 Inst_E_IO_ConfigMem.Inst_frame0_bit6.Q
rlabel via2 5960 4872 5960 4872 0 Inst_E_IO_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 3456 9702 3456 9702 0 Inst_E_IO_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 7736 10920 7736 10920 0 Inst_E_IO_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 9600 34482 9600 34482 0 Inst_E_IO_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 7824 34440 7824 34440 0 Inst_E_IO_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 8744 36624 8744 36624 0 Inst_E_IO_ConfigMem.Inst_frame1_bit10.Q
rlabel metal3 7392 35532 7392 35532 0 Inst_E_IO_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 9864 33600 9864 33600 0 Inst_E_IO_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 8064 33600 8064 33600 0 Inst_E_IO_ConfigMem.Inst_frame1_bit13.Q
rlabel via2 7880 24528 7880 24528 0 Inst_E_IO_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 6192 24528 6192 24528 0 Inst_E_IO_ConfigMem.Inst_frame1_bit15.Q
rlabel metal3 9792 38682 9792 38682 0 Inst_E_IO_ConfigMem.Inst_frame1_bit16.Q
rlabel metal3 8448 38640 8448 38640 0 Inst_E_IO_ConfigMem.Inst_frame1_bit17.Q
rlabel metal3 10176 30744 10176 30744 0 Inst_E_IO_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 8976 30828 8976 30828 0 Inst_E_IO_ConfigMem.Inst_frame1_bit19.Q
rlabel metal3 4512 16338 4512 16338 0 Inst_E_IO_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 10080 28350 10080 28350 0 Inst_E_IO_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 8544 28434 8544 28434 0 Inst_E_IO_ConfigMem.Inst_frame1_bit21.Q
rlabel metal4 3264 13776 3264 13776 0 Inst_E_IO_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 2304 15708 2304 15708 0 Inst_E_IO_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 3120 13440 3120 13440 0 Inst_E_IO_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 2592 14700 2592 14700 0 Inst_E_IO_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 7728 25368 7728 25368 0 Inst_E_IO_ConfigMem.Inst_frame1_bit26.Q
rlabel metal3 9504 25620 9504 25620 0 Inst_E_IO_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 7905 39648 7905 39648 0 Inst_E_IO_ConfigMem.Inst_frame1_bit28.Q
rlabel via2 9512 39648 9512 39648 0 Inst_E_IO_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 5568 16464 5568 16464 0 Inst_E_IO_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 6096 29904 6096 29904 0 Inst_E_IO_ConfigMem.Inst_frame1_bit30.Q
rlabel metal3 7680 30156 7680 30156 0 Inst_E_IO_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 4032 22386 4032 22386 0 Inst_E_IO_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 5856 22344 5856 22344 0 Inst_E_IO_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 3416 18480 3416 18480 0 Inst_E_IO_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 1776 18480 1776 18480 0 Inst_E_IO_ConfigMem.Inst_frame1_bit7.Q
rlabel metal3 4272 13188 4272 13188 0 Inst_E_IO_ConfigMem.Inst_frame1_bit8.Q
rlabel metal3 2304 13482 2304 13482 0 Inst_E_IO_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 4032 37506 4032 37506 0 Inst_E_IO_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 5616 37464 5616 37464 0 Inst_E_IO_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 3984 34188 3984 34188 0 Inst_E_IO_ConfigMem.Inst_frame2_bit10.Q
rlabel via2 6248 29064 6248 29064 0 Inst_E_IO_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 3072 36582 3072 36582 0 Inst_E_IO_ConfigMem.Inst_frame2_bit12.Q
rlabel via2 4616 36624 4616 36624 0 Inst_E_IO_ConfigMem.Inst_frame2_bit13.Q
rlabel metal3 2688 29988 2688 29988 0 Inst_E_IO_ConfigMem.Inst_frame2_bit14.Q
rlabel metal3 4704 29232 4704 29232 0 Inst_E_IO_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 5184 36666 5184 36666 0 Inst_E_IO_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 8016 35784 8016 35784 0 Inst_E_IO_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 8064 23058 8064 23058 0 Inst_E_IO_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 9792 22512 9792 22512 0 Inst_E_IO_ConfigMem.Inst_frame2_bit19.Q
rlabel metal3 7584 16002 7584 16002 0 Inst_E_IO_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 7776 18480 7776 18480 0 Inst_E_IO_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 9672 18480 9672 18480 0 Inst_E_IO_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 3696 6384 3696 6384 0 Inst_E_IO_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 5736 6384 5736 6384 0 Inst_E_IO_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 4032 8904 4032 8904 0 Inst_E_IO_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 5664 9660 5664 9660 0 Inst_E_IO_ConfigMem.Inst_frame2_bit25.Q
rlabel metal3 8160 27174 8160 27174 0 Inst_E_IO_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 6624 26922 6624 26922 0 Inst_E_IO_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 9216 40488 9216 40488 0 Inst_E_IO_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 7872 40530 7872 40530 0 Inst_E_IO_ConfigMem.Inst_frame2_bit29.Q
rlabel metal3 9408 16002 9408 16002 0 Inst_E_IO_ConfigMem.Inst_frame2_bit3.Q
rlabel metal2 8736 32340 8736 32340 0 Inst_E_IO_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 8064 32970 8064 32970 0 Inst_E_IO_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 6768 19320 6768 19320 0 Inst_E_IO_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 8256 19320 8256 19320 0 Inst_E_IO_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 3168 5754 3168 5754 0 Inst_E_IO_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 4032 5166 4032 5166 0 Inst_E_IO_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 3936 10416 3936 10416 0 Inst_E_IO_ConfigMem.Inst_frame2_bit8.Q
rlabel metal3 5760 11466 5760 11466 0 Inst_E_IO_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 7008 13314 7008 13314 0 Inst_E_IO_ConfigMem.Inst_frame3_bit22.Q
rlabel metal3 7776 7644 7776 7644 0 Inst_E_IO_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 4992 7854 4992 7854 0 Inst_E_IO_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 5952 8778 5952 8778 0 Inst_E_IO_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 4224 27804 4224 27804 0 Inst_E_IO_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 6000 27804 6000 27804 0 Inst_E_IO_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 3168 39648 3168 39648 0 Inst_E_IO_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 4760 39648 4760 39648 0 Inst_E_IO_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 2784 32004 2784 32004 0 Inst_E_IO_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 4328 32088 4328 32088 0 Inst_E_IO_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 8064 13104 8064 13104 0 Inst_E_IO_switch_matrix.W1BEG0
rlabel metal3 8352 7602 8352 7602 0 Inst_E_IO_switch_matrix.W1BEG1
rlabel metal2 6048 8022 6048 8022 0 Inst_E_IO_switch_matrix.W1BEG2
rlabel metal2 6408 8904 6408 8904 0 Inst_E_IO_switch_matrix.W1BEG3
rlabel metal2 6336 28392 6336 28392 0 Inst_E_IO_switch_matrix.W2BEG0
rlabel metal2 4896 39480 4896 39480 0 Inst_E_IO_switch_matrix.W2BEG1
rlabel metal2 4776 32088 4776 32088 0 Inst_E_IO_switch_matrix.W2BEG2
rlabel metal2 5832 38136 5832 38136 0 Inst_E_IO_switch_matrix.W2BEG3
rlabel metal2 9888 16464 9888 16464 0 Inst_E_IO_switch_matrix.W2BEG4
rlabel metal2 9264 19488 9264 19488 0 Inst_E_IO_switch_matrix.W2BEG5
rlabel metal2 5112 5628 5112 5628 0 Inst_E_IO_switch_matrix.W2BEG6
rlabel metal2 6144 12516 6144 12516 0 Inst_E_IO_switch_matrix.W2BEG7
rlabel metal2 6528 29064 6528 29064 0 Inst_E_IO_switch_matrix.W2BEGb0
rlabel metal2 3817 37464 3817 37464 0 Inst_E_IO_switch_matrix.W2BEGb1
rlabel metal2 5376 31500 5376 31500 0 Inst_E_IO_switch_matrix.W2BEGb2
rlabel metal2 7344 36456 7344 36456 0 Inst_E_IO_switch_matrix.W2BEGb3
rlabel metal2 9840 22848 9840 22848 0 Inst_E_IO_switch_matrix.W2BEGb4
rlabel metal2 9840 17724 9840 17724 0 Inst_E_IO_switch_matrix.W2BEGb5
rlabel metal3 5856 5922 5856 5922 0 Inst_E_IO_switch_matrix.W2BEGb6
rlabel metal2 6264 10164 6264 10164 0 Inst_E_IO_switch_matrix.W2BEGb7
rlabel metal2 9888 25452 9888 25452 0 Inst_E_IO_switch_matrix.W6BEG0
rlabel metal2 10224 39606 10224 39606 0 Inst_E_IO_switch_matrix.W6BEG1
rlabel metal2 9168 5628 9168 5628 0 Inst_E_IO_switch_matrix.W6BEG10
rlabel metal2 8424 9660 8424 9660 0 Inst_E_IO_switch_matrix.W6BEG11
rlabel metal2 7968 29904 7968 29904 0 Inst_E_IO_switch_matrix.W6BEG2
rlabel metal2 5599 41160 5599 41160 0 Inst_E_IO_switch_matrix.W6BEG3
rlabel metal2 9816 14700 9816 14700 0 Inst_E_IO_switch_matrix.W6BEG4
rlabel metal3 9504 17514 9504 17514 0 Inst_E_IO_switch_matrix.W6BEG5
rlabel metal2 6360 4956 6360 4956 0 Inst_E_IO_switch_matrix.W6BEG6
rlabel metal2 8112 10164 8112 10164 0 Inst_E_IO_switch_matrix.W6BEG7
rlabel metal2 5568 32928 5568 32928 0 Inst_E_IO_switch_matrix.W6BEG8
rlabel metal2 6552 35952 6552 35952 0 Inst_E_IO_switch_matrix.W6BEG9
rlabel metal2 8448 26880 8448 26880 0 Inst_E_IO_switch_matrix.WW4BEG0
rlabel metal2 9936 40488 9936 40488 0 Inst_E_IO_switch_matrix.WW4BEG1
rlabel metal2 8160 24528 8160 24528 0 Inst_E_IO_switch_matrix.WW4BEG10
rlabel metal2 10176 39060 10176 39060 0 Inst_E_IO_switch_matrix.WW4BEG11
rlabel metal2 10056 30618 10056 30618 0 Inst_E_IO_switch_matrix.WW4BEG12
rlabel metal2 10153 29064 10153 29064 0 Inst_E_IO_switch_matrix.WW4BEG13
rlabel metal2 4992 18396 4992 18396 0 Inst_E_IO_switch_matrix.WW4BEG14
rlabel metal2 4560 15540 4560 15540 0 Inst_E_IO_switch_matrix.WW4BEG15
rlabel metal2 9888 32928 9888 32928 0 Inst_E_IO_switch_matrix.WW4BEG2
rlabel metal2 9912 34440 9912 34440 0 Inst_E_IO_switch_matrix.WW4BEG3
rlabel metal3 6240 17514 6240 17514 0 Inst_E_IO_switch_matrix.WW4BEG4
rlabel metal2 5952 22512 5952 22512 0 Inst_E_IO_switch_matrix.WW4BEG5
rlabel metal2 4608 18480 4608 18480 0 Inst_E_IO_switch_matrix.WW4BEG6
rlabel metal2 4536 14028 4536 14028 0 Inst_E_IO_switch_matrix.WW4BEG7
rlabel metal2 9144 36624 9144 36624 0 Inst_E_IO_switch_matrix.WW4BEG8
rlabel metal2 10056 33600 10056 33600 0 Inst_E_IO_switch_matrix.WW4BEG9
rlabel metal3 2016 5826 2016 5826 0 UserCLK
rlabel metal3 2016 46246 2016 46246 0 UserCLKo
rlabel metal2 800 2268 800 2268 0 W1BEG[0]
rlabel metal2 608 2604 608 2604 0 W1BEG[1]
rlabel metal2 2040 2856 2040 2856 0 W1BEG[2]
rlabel metal2 1584 1848 1584 1848 0 W1BEG[3]
rlabel metal2 128 3612 128 3612 0 W2BEG[0]
rlabel metal2 1752 2772 1752 2772 0 W2BEG[1]
rlabel metal2 1872 1596 1872 1596 0 W2BEG[2]
rlabel metal2 840 2100 840 2100 0 W2BEG[3]
rlabel metal2 1472 4956 1472 4956 0 W2BEG[4]
rlabel metal2 704 5292 704 5292 0 W2BEG[5]
rlabel metal2 1464 1764 1464 1764 0 W2BEG[6]
rlabel metal2 656 5964 656 5964 0 W2BEG[7]
rlabel metal2 2616 2100 2616 2100 0 W2BEGb[0]
rlabel metal2 696 2856 696 2856 0 W2BEGb[1]
rlabel metal2 1896 2604 1896 2604 0 W2BEGb[2]
rlabel metal2 752 7308 752 7308 0 W2BEGb[3]
rlabel metal2 3480 3612 3480 3612 0 W2BEGb[4]
rlabel metal2 128 7980 128 7980 0 W2BEGb[5]
rlabel metal2 1472 8316 1472 8316 0 W2BEGb[6]
rlabel metal2 1080 2016 1080 2016 0 W2BEGb[7]
rlabel metal2 128 14364 128 14364 0 W6BEG[0]
rlabel via2 80 17724 80 17724 0 W6BEG[10]
rlabel metal2 224 18060 224 18060 0 W6BEG[11]
rlabel metal2 128 14700 128 14700 0 W6BEG[1]
rlabel via2 80 15036 80 15036 0 W6BEG[2]
rlabel metal2 416 15372 416 15372 0 W6BEG[3]
rlabel metal2 704 15708 704 15708 0 W6BEG[4]
rlabel metal2 128 16044 128 16044 0 W6BEG[5]
rlabel metal2 560 16380 560 16380 0 W6BEG[6]
rlabel metal2 368 16716 368 16716 0 W6BEG[7]
rlabel metal2 752 17052 752 17052 0 W6BEG[8]
rlabel metal2 272 17388 272 17388 0 W6BEG[9]
rlabel metal2 416 8988 416 8988 0 WW4BEG[0]
rlabel metal2 128 12348 128 12348 0 WW4BEG[10]
rlabel metal2 752 12684 752 12684 0 WW4BEG[11]
rlabel metal2 416 13020 416 13020 0 WW4BEG[12]
rlabel metal2 368 13356 368 13356 0 WW4BEG[13]
rlabel metal2 704 13692 704 13692 0 WW4BEG[14]
rlabel metal2 320 14028 320 14028 0 WW4BEG[15]
rlabel metal2 3336 6972 3336 6972 0 WW4BEG[1]
rlabel metal2 3192 7056 3192 7056 0 WW4BEG[2]
rlabel metal2 560 9996 560 9996 0 WW4BEG[3]
rlabel metal2 272 10332 272 10332 0 WW4BEG[4]
rlabel metal2 560 10668 560 10668 0 WW4BEG[5]
rlabel metal2 608 11004 608 11004 0 WW4BEG[6]
rlabel metal2 656 11340 656 11340 0 WW4BEG[7]
rlabel metal2 128 11676 128 11676 0 WW4BEG[8]
rlabel metal2 464 12012 464 12012 0 WW4BEG[9]
rlabel metal2 5304 25368 5304 25368 0 _000_
rlabel metal2 3744 17808 3744 17808 0 _001_
rlabel metal2 5928 23268 5928 23268 0 _002_
rlabel metal2 4032 30576 4032 30576 0 _003_
rlabel metal2 4704 23814 4704 23814 0 _004_
rlabel metal2 4608 24024 4608 24024 0 _005_
rlabel metal2 3619 25368 3619 25368 0 _006_
rlabel metal2 3456 25410 3456 25410 0 _007_
rlabel metal2 3486 24528 3486 24528 0 _008_
rlabel metal2 4809 25536 4809 25536 0 _009_
rlabel metal2 3648 24654 3648 24654 0 _010_
rlabel metal2 4091 24612 4091 24612 0 _011_
rlabel metal3 2784 22218 2784 22218 0 _012_
rlabel metal2 2400 23898 2400 23898 0 _013_
rlabel metal2 3407 23856 3407 23856 0 _014_
rlabel metal2 2640 23856 2640 23856 0 _015_
rlabel metal2 3243 24528 3243 24528 0 _016_
rlabel metal2 3600 24360 3600 24360 0 _017_
rlabel metal2 5760 21000 5760 21000 0 _018_
rlabel metal2 6048 20244 6048 20244 0 _019_
rlabel metal2 5155 19992 5155 19992 0 _020_
rlabel metal2 4896 19992 4896 19992 0 _021_
rlabel metal2 5685 20832 5685 20832 0 _022_
rlabel metal2 5784 21336 5784 21336 0 _023_
rlabel metal3 5856 21084 5856 21084 0 _024_
rlabel metal2 6192 20748 6192 20748 0 _025_
rlabel metal2 3514 19992 3514 19992 0 _026_
rlabel metal2 3024 19152 3024 19152 0 _027_
rlabel metal3 4128 20286 4128 20286 0 _028_
rlabel metal2 3552 20118 3552 20118 0 _029_
rlabel metal2 5592 19992 5592 19992 0 _030_
rlabel metal2 6432 20748 6432 20748 0 _031_
rlabel metal2 4992 16338 4992 16338 0 _032_
rlabel metal2 5040 16464 5040 16464 0 _033_
rlabel metal2 5472 16968 5472 16968 0 _034_
rlabel metal2 3552 17010 3552 17010 0 _035_
rlabel metal2 4512 16338 4512 16338 0 _036_
rlabel via1 4296 16285 4296 16285 0 _037_
rlabel via1 4913 16968 4913 16968 0 _038_
rlabel metal2 4224 16464 4224 16464 0 _039_
rlabel metal2 4440 16212 4440 16212 0 _040_
rlabel metal2 3991 28476 3991 28476 0 _041_
rlabel metal3 3744 28770 3744 28770 0 _042_
rlabel metal2 3869 29148 3869 29148 0 _043_
rlabel metal2 3456 29820 3456 29820 0 _044_
rlabel metal2 4272 29316 4272 29316 0 _045_
rlabel via1 3126 29904 3126 29904 0 _046_
rlabel metal2 3243 29988 3243 29988 0 _047_
rlabel metal2 3696 29904 3696 29904 0 _048_
rlabel metal2 9408 2100 9408 2100 0 net1
rlabel metal2 4752 22344 4752 22344 0 net10
rlabel metal3 2304 9828 2304 9828 0 net100
rlabel metal3 5904 21588 5904 21588 0 net101
rlabel metal2 10320 2604 10320 2604 0 net102
rlabel metal4 5712 7224 5712 7224 0 net103
rlabel metal2 10368 6510 10368 6510 0 net104
rlabel metal2 9360 7056 9360 7056 0 net105
rlabel metal2 10464 7140 10464 7140 0 net106
rlabel metal2 8976 8148 8976 8148 0 net107
rlabel metal4 3504 13608 3504 13608 0 net108
rlabel metal4 9888 6468 9888 6468 0 net109
rlabel metal2 5424 36624 5424 36624 0 net11
rlabel metal2 10848 10248 10848 10248 0 net110
rlabel metal2 10320 13356 10320 13356 0 net111
rlabel metal2 8784 13188 8784 13188 0 net112
rlabel metal4 10320 18564 10320 18564 0 net113
rlabel metal4 6048 18480 6048 18480 0 net114
rlabel metal2 9600 35364 9600 35364 0 net115
rlabel metal2 6360 34188 6360 34188 0 net116
rlabel metal2 1560 40992 1560 40992 0 net117
rlabel metal2 8352 35448 8352 35448 0 net118
rlabel metal3 2112 4788 2112 4788 0 net119
rlabel metal3 3552 30828 3552 30828 0 net12
rlabel metal4 9504 18732 9504 18732 0 net120
rlabel metal2 10152 39480 10152 39480 0 net121
rlabel metal2 9192 37296 9192 37296 0 net122
rlabel metal2 10392 30828 10392 30828 0 net123
rlabel metal2 8904 13776 8904 13776 0 net124
rlabel metal2 10704 14700 10704 14700 0 net125
rlabel metal2 9576 14028 9576 14028 0 net126
rlabel metal2 10512 41244 10512 41244 0 net127
rlabel metal2 3336 7392 3336 7392 0 net128
rlabel metal4 8256 18816 8256 18816 0 net129
rlabel metal4 4608 19236 4608 19236 0 net13
rlabel metal4 10272 42756 10272 42756 0 net130
rlabel metal3 2112 22722 2112 22722 0 net131
rlabel metal2 9120 41874 9120 41874 0 net132
rlabel metal4 9888 42756 9888 42756 0 net133
rlabel metal2 6552 40656 6552 40656 0 net134
rlabel metal2 4056 43428 4056 43428 0 net135
rlabel metal2 6504 14196 6504 14196 0 net136
rlabel metal2 3504 33390 3504 33390 0 net137
rlabel metal2 5064 33684 5064 33684 0 net138
rlabel metal2 6312 14112 6312 14112 0 net139
rlabel metal2 4368 25452 4368 25452 0 net14
rlabel metal2 2016 18942 2016 18942 0 net140
rlabel metal2 7944 18732 7944 18732 0 net141
rlabel metal2 1752 4788 1752 4788 0 net142
rlabel metal2 1896 4284 1896 4284 0 net143
rlabel metal2 10896 22260 10896 22260 0 net144
rlabel metal2 3432 11676 3432 11676 0 net145
rlabel metal2 1848 35364 1848 35364 0 net146
rlabel metal2 6552 44436 6552 44436 0 net147
rlabel metal2 7800 44436 7800 44436 0 net148
rlabel metal2 7368 44436 7368 44436 0 net149
rlabel metal3 2832 21588 2832 21588 0 net15
rlabel metal2 5544 42924 5544 42924 0 net150
rlabel metal2 3624 43680 3624 43680 0 net151
rlabel metal2 5208 42168 5208 42168 0 net152
rlabel metal2 4392 44016 4392 44016 0 net153
rlabel metal2 9072 44940 9072 44940 0 net154
rlabel metal2 9432 44436 9432 44436 0 net155
rlabel metal2 9816 44352 9816 44352 0 net156
rlabel metal2 9192 42168 9192 42168 0 net157
rlabel metal2 7992 42168 7992 42168 0 net158
rlabel metal2 4296 42756 4296 42756 0 net159
rlabel metal2 2496 5544 2496 5544 0 net16
rlabel metal2 6936 44436 6936 44436 0 net160
rlabel metal2 6168 44436 6168 44436 0 net161
rlabel metal3 4992 44520 4992 44520 0 net162
rlabel metal2 4248 44436 4248 44436 0 net163
rlabel metal2 3144 43344 3144 43344 0 net164
rlabel metal2 5208 44352 5208 44352 0 net165
rlabel metal2 7848 11928 7848 11928 0 net166
rlabel metal2 3360 2562 3360 2562 0 net167
rlabel metal2 4656 2100 4656 2100 0 net168
rlabel metal2 3744 2688 3744 2688 0 net169
rlabel metal2 2352 19992 2352 19992 0 net17
rlabel metal2 3984 2016 3984 2016 0 net170
rlabel metal4 4992 4284 4992 4284 0 net171
rlabel metal5 2592 15624 2592 15624 0 net172
rlabel metal4 4224 1932 4224 1932 0 net173
rlabel metal2 5232 2856 5232 2856 0 net174
rlabel metal2 9480 15288 9480 15288 0 net175
rlabel metal2 10752 17304 10752 17304 0 net176
rlabel metal2 2208 1890 2208 1890 0 net177
rlabel metal2 2736 3444 2736 3444 0 net178
rlabel metal4 4896 2772 4896 2772 0 net179
rlabel metal2 2544 21420 2544 21420 0 net18
rlabel metal2 1488 2604 1488 2604 0 net180
rlabel metal4 3888 2856 3888 2856 0 net181
rlabel metal2 3648 2772 3648 2772 0 net182
rlabel metal2 10872 22848 10872 22848 0 net183
rlabel metal2 8472 17556 8472 17556 0 net184
rlabel metal2 6264 5544 6264 5544 0 net185
rlabel metal2 3984 2184 3984 2184 0 net186
rlabel metal4 10560 21756 10560 21756 0 net187
rlabel metal2 3600 16212 3600 16212 0 net188
rlabel metal2 1824 14658 1824 14658 0 net189
rlabel metal2 2208 20874 2208 20874 0 net19
rlabel metal4 8112 15708 8112 15708 0 net190
rlabel metal4 6288 15624 6288 15624 0 net191
rlabel metal4 4800 15540 4800 15540 0 net192
rlabel metal2 2208 13902 2208 13902 0 net193
rlabel metal2 3600 15540 3600 15540 0 net194
rlabel metal2 2208 14112 2208 14112 0 net195
rlabel metal3 1440 13776 1440 13776 0 net196
rlabel metal4 4608 15792 4608 15792 0 net197
rlabel metal2 2256 14700 2256 14700 0 net198
rlabel metal5 1632 16590 1632 16590 0 net199
rlabel metal2 8832 17766 8832 17766 0 net2
rlabel metal2 2304 20958 2304 20958 0 net20
rlabel metal3 4704 13188 4704 13188 0 net200
rlabel metal4 10368 38892 10368 38892 0 net201
rlabel metal3 1824 10836 1824 10836 0 net202
rlabel metal3 1440 10710 1440 10710 0 net203
rlabel metal3 2784 16380 2784 16380 0 net204
rlabel metal2 1440 11046 1440 11046 0 net205
rlabel metal2 3552 2856 3552 2856 0 net206
rlabel metal4 6912 7140 6912 7140 0 net207
rlabel metal4 11376 17976 11376 17976 0 net208
rlabel metal2 6072 16884 6072 16884 0 net209
rlabel metal2 1416 19320 1416 19320 0 net21
rlabel metal4 3984 21504 3984 21504 0 net210
rlabel metal3 4800 13272 4800 13272 0 net211
rlabel metal2 4488 13776 4488 13776 0 net212
rlabel metal2 9480 36456 9480 36456 0 net213
rlabel metal2 10728 33432 10728 33432 0 net214
rlabel metal3 8928 12138 8928 12138 0 net215
rlabel metal3 9312 10542 9312 10542 0 net216
rlabel metal2 3936 29022 3936 29022 0 net22
rlabel metal4 6864 17976 6864 17976 0 net23
rlabel metal3 8736 38766 8736 38766 0 net24
rlabel metal2 8352 34524 8352 34524 0 net25
rlabel metal3 4176 13104 4176 13104 0 net26
rlabel metal2 1728 34230 1728 34230 0 net27
rlabel metal2 8880 16296 8880 16296 0 net28
rlabel metal3 7104 25746 7104 25746 0 net29
rlabel metal2 2208 14490 2208 14490 0 net3
rlabel metal2 4320 32802 4320 32802 0 net30
rlabel metal2 4176 36624 4176 36624 0 net31
rlabel metal2 6576 29820 6576 29820 0 net32
rlabel metal2 1464 33264 1464 33264 0 net33
rlabel metal4 7056 4872 7056 4872 0 net34
rlabel metal2 1728 26712 1728 26712 0 net35
rlabel metal4 7296 19236 7296 19236 0 net36
rlabel metal2 8400 25368 8400 25368 0 net37
rlabel metal2 5184 35910 5184 35910 0 net38
rlabel metal2 4032 31290 4032 31290 0 net39
rlabel metal4 4944 7896 4944 7896 0 net4
rlabel metal2 3840 36624 3840 36624 0 net40
rlabel metal3 6624 30534 6624 30534 0 net41
rlabel metal3 1488 19824 1488 19824 0 net42
rlabel metal2 7536 19320 7536 19320 0 net43
rlabel metal2 2160 28854 2160 28854 0 net44
rlabel metal3 5664 36246 5664 36246 0 net45
rlabel metal2 3936 31374 3936 31374 0 net46
rlabel metal4 2592 34944 2592 34944 0 net47
rlabel metal2 4896 28392 4896 28392 0 net48
rlabel metal4 2544 11928 2544 11928 0 net49
rlabel metal2 4152 18564 4152 18564 0 net5
rlabel metal4 672 24360 672 24360 0 net50
rlabel metal2 2448 38136 2448 38136 0 net51
rlabel metal2 2016 34482 2016 34482 0 net52
rlabel metal2 5568 34440 5568 34440 0 net53
rlabel metal2 816 41160 816 41160 0 net54
rlabel metal2 6480 35112 6480 35112 0 net55
rlabel metal3 1104 33684 1104 33684 0 net56
rlabel metal4 1632 32802 1632 32802 0 net57
rlabel metal3 9888 41412 9888 41412 0 net58
rlabel metal2 9504 13272 9504 13272 0 net59
rlabel metal2 7872 17850 7872 17850 0 net6
rlabel metal2 10585 9408 10585 9408 0 net60
rlabel metal3 2688 32298 2688 32298 0 net61
rlabel metal2 2736 5712 2736 5712 0 net62
rlabel metal2 8256 19992 8256 19992 0 net63
rlabel metal2 9984 16296 9984 16296 0 net64
rlabel metal2 2688 28308 2688 28308 0 net65
rlabel metal2 7392 40446 7392 40446 0 net66
rlabel metal3 2784 11676 2784 11676 0 net67
rlabel metal2 2256 15456 2256 15456 0 net68
rlabel metal2 10224 29904 10224 29904 0 net69
rlabel via3 4416 20832 4416 20832 0 net7
rlabel metal2 9888 41958 9888 41958 0 net70
rlabel metal2 7320 23016 7320 23016 0 net71
rlabel metal2 7536 11760 7536 11760 0 net72
rlabel metal2 7056 20832 7056 20832 0 net73
rlabel metal2 9384 16968 9384 16968 0 net74
rlabel metal3 2592 33318 2592 33318 0 net75
rlabel metal3 2592 38640 2592 38640 0 net76
rlabel metal2 1776 35196 1776 35196 0 net77
rlabel metal2 7008 38220 7008 38220 0 net78
rlabel metal2 10128 21504 10128 21504 0 net79
rlabel metal2 3792 6468 3792 6468 0 net8
rlabel metal2 1728 42966 1728 42966 0 net80
rlabel metal2 6144 39018 6144 39018 0 net81
rlabel metal2 2304 42462 2304 42462 0 net82
rlabel metal2 8736 20874 8736 20874 0 net83
rlabel metal2 1584 11760 1584 11760 0 net84
rlabel metal2 1728 16926 1728 16926 0 net85
rlabel metal2 1824 16380 1824 16380 0 net86
rlabel metal3 720 38136 720 38136 0 net87
rlabel metal2 2496 27510 2496 27510 0 net88
rlabel metal2 2544 26880 2544 26880 0 net89
rlabel metal2 4368 20748 4368 20748 0 net9
rlabel metal2 1824 41160 1824 41160 0 net90
rlabel metal2 1440 39186 1440 39186 0 net91
rlabel metal2 2232 37464 2232 37464 0 net92
rlabel metal2 1344 32088 1344 32088 0 net93
rlabel metal2 2232 45108 2232 45108 0 net94
rlabel metal2 2712 37464 2712 37464 0 net95
rlabel metal2 3264 37506 3264 37506 0 net96
rlabel metal3 7104 17808 7104 17808 0 net97
rlabel metal2 1584 7896 1584 7896 0 net98
rlabel metal2 1296 7224 1296 7224 0 net99
<< properties >>
string FIXED_BBOX 0 0 11840 47360
<< end >>
