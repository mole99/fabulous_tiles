module W_IO (A_I_top,
    A_O_top,
    A_T_top,
    A_config_C_bit0,
    A_config_C_bit1,
    A_config_C_bit2,
    A_config_C_bit3,
    B_I_top,
    B_O_top,
    B_T_top,
    B_config_C_bit0,
    B_config_C_bit1,
    B_config_C_bit2,
    B_config_C_bit3,
    UserCLK,
    UserCLKo,
    E1BEG,
    E2BEG,
    E2BEGb,
    E6BEG,
    EE4BEG,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    W1END,
    W2END,
    W2MID,
    W6END,
    WW4END);
 output A_I_top;
 input A_O_top;
 output A_T_top;
 output A_config_C_bit0;
 output A_config_C_bit1;
 output A_config_C_bit2;
 output A_config_C_bit3;
 output B_I_top;
 input B_O_top;
 output B_T_top;
 output B_config_C_bit0;
 output B_config_C_bit1;
 output B_config_C_bit2;
 output B_config_C_bit3;
 input UserCLK;
 output UserCLKo;
 output [3:0] E1BEG;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 output [11:0] E6BEG;
 output [15:0] EE4BEG;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] W1END;
 input [7:0] W2END;
 input [7:0] W2MID;
 input [11:0] W6END;
 input [15:0] WW4END;

 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire \Inst_A_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_B_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_W_IO_switch_matrix.E1BEG0 ;
 wire \Inst_W_IO_switch_matrix.E1BEG1 ;
 wire \Inst_W_IO_switch_matrix.E1BEG2 ;
 wire \Inst_W_IO_switch_matrix.E1BEG3 ;
 wire \Inst_W_IO_switch_matrix.E2BEG0 ;
 wire \Inst_W_IO_switch_matrix.E2BEG1 ;
 wire \Inst_W_IO_switch_matrix.E2BEG2 ;
 wire \Inst_W_IO_switch_matrix.E2BEG3 ;
 wire \Inst_W_IO_switch_matrix.E2BEG4 ;
 wire \Inst_W_IO_switch_matrix.E2BEG5 ;
 wire \Inst_W_IO_switch_matrix.E2BEG6 ;
 wire \Inst_W_IO_switch_matrix.E2BEG7 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb0 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb1 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb2 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb3 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb4 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb5 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb6 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb7 ;
 wire \Inst_W_IO_switch_matrix.E6BEG0 ;
 wire \Inst_W_IO_switch_matrix.E6BEG1 ;
 wire \Inst_W_IO_switch_matrix.E6BEG10 ;
 wire \Inst_W_IO_switch_matrix.E6BEG11 ;
 wire \Inst_W_IO_switch_matrix.E6BEG2 ;
 wire \Inst_W_IO_switch_matrix.E6BEG3 ;
 wire \Inst_W_IO_switch_matrix.E6BEG4 ;
 wire \Inst_W_IO_switch_matrix.E6BEG5 ;
 wire \Inst_W_IO_switch_matrix.E6BEG6 ;
 wire \Inst_W_IO_switch_matrix.E6BEG7 ;
 wire \Inst_W_IO_switch_matrix.E6BEG8 ;
 wire \Inst_W_IO_switch_matrix.E6BEG9 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG0 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG1 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG10 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG11 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG12 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG13 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG14 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG15 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG2 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG3 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG4 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG5 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG6 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG7 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG8 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG9 ;
 wire net211;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire UserCLK_regs;
 wire clknet_0_UserCLK;
 wire clknet_1_0__leaf_UserCLK;
 wire clknet_0_UserCLK_regs;
 wire clknet_1_0__leaf_UserCLK_regs;
 wire clknet_1_1__leaf_UserCLK_regs;

 sky130_fd_sc_hd__inv_1 _032_ (.A(\Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _033_ (.A(\Inst_W_IO_ConfigMem.Inst_frame0_bit28.Q ),
    .Y(_001_));
 sky130_fd_sc_hd__inv_1 _034_ (.A(\Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _035_ (.A(\Inst_W_IO_ConfigMem.Inst_frame0_bit21.Q ),
    .Y(_003_));
 sky130_fd_sc_hd__inv_1 _036_ (.A(\Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .Y(_004_));
 sky130_fd_sc_hd__inv_1 _037_ (.A(\Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_005_));
 sky130_fd_sc_hd__mux4_1 _038_ (.A0(net40),
    .A1(net41),
    .A2(net42),
    .A3(net43),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_006_));
 sky130_fd_sc_hd__or2_1 _039_ (.A(\Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .B(_006_),
    .X(_007_));
 sky130_fd_sc_hd__mux4_1 _040_ (.A0(net59),
    .A1(net60),
    .A2(net61),
    .A3(net62),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_008_));
 sky130_fd_sc_hd__o21a_1 _041_ (.A1(_000_),
    .A2(_008_),
    .B1(\Inst_W_IO_ConfigMem.Inst_frame0_bit28.Q ),
    .X(_009_));
 sky130_fd_sc_hd__mux4_1 _042_ (.A0(net63),
    .A1(net64),
    .A2(net65),
    .A3(net66),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_010_));
 sky130_fd_sc_hd__mux4_1 _043_ (.A0(net67),
    .A1(net68),
    .A2(net69),
    .A3(net70),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _044_ (.A0(_010_),
    .A1(_011_),
    .S(\Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_012_));
 sky130_fd_sc_hd__a22o_1 _045_ (.A1(_007_),
    .A2(_009_),
    .B1(_012_),
    .B2(_001_),
    .X(net105));
 sky130_fd_sc_hd__mux4_1 _046_ (.A0(net40),
    .A1(net41),
    .A2(net42),
    .A3(net43),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_013_));
 sky130_fd_sc_hd__or2_1 _047_ (.A(\Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .B(_013_),
    .X(_014_));
 sky130_fd_sc_hd__mux4_1 _048_ (.A0(net59),
    .A1(net60),
    .A2(net61),
    .A3(net62),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_015_));
 sky130_fd_sc_hd__o21a_1 _049_ (.A1(_002_),
    .A2(_015_),
    .B1(\Inst_W_IO_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_016_));
 sky130_fd_sc_hd__mux4_1 _050_ (.A0(net63),
    .A1(net64),
    .A2(net65),
    .A3(net66),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_017_));
 sky130_fd_sc_hd__mux4_1 _051_ (.A0(net67),
    .A1(net68),
    .A2(net69),
    .A3(net70),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_018_));
 sky130_fd_sc_hd__mux2_1 _052_ (.A0(_017_),
    .A1(_018_),
    .S(\Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .X(_019_));
 sky130_fd_sc_hd__a22o_1 _053_ (.A1(_014_),
    .A2(_016_),
    .B1(_019_),
    .B2(_003_),
    .X(net99));
 sky130_fd_sc_hd__mux4_1 _054_ (.A0(net36),
    .A1(net83),
    .A2(net71),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit16.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit17.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG11 ));
 sky130_fd_sc_hd__mux4_1 _055_ (.A0(net37),
    .A1(net90),
    .A2(net74),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit14.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit15.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG10 ));
 sky130_fd_sc_hd__mux4_1 _056_ (.A0(net93),
    .A1(net86),
    .A2(net77),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit12.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit13.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG9 ));
 sky130_fd_sc_hd__mux4_1 _057_ (.A0(net94),
    .A1(net87),
    .A2(net78),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit10.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit11.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG8 ));
 sky130_fd_sc_hd__mux4_1 _058_ (.A0(net36),
    .A1(net97),
    .A2(net81),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit8.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit9.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG7 ));
 sky130_fd_sc_hd__mux4_1 _059_ (.A0(net37),
    .A1(net98),
    .A2(net82),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit6.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit7.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG6 ));
 sky130_fd_sc_hd__mux4_1 _060_ (.A0(net39),
    .A1(net91),
    .A2(net75),
    .A3(net2),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit4.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit5.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG5 ));
 sky130_fd_sc_hd__mux4_1 _061_ (.A0(net38),
    .A1(net92),
    .A2(net76),
    .A3(net1),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit2.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit3.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG4 ));
 sky130_fd_sc_hd__mux4_1 _062_ (.A0(net95),
    .A1(net88),
    .A2(net79),
    .A3(net2),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit0.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit1.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG3 ));
 sky130_fd_sc_hd__mux4_1 _063_ (.A0(net96),
    .A1(net89),
    .A2(net80),
    .A3(net1),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit30.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit31.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG2 ));
 sky130_fd_sc_hd__mux4_1 _064_ (.A0(net39),
    .A1(net84),
    .A2(net72),
    .A3(net2),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit29.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG1 ));
 sky130_fd_sc_hd__mux4_1 _065_ (.A0(net38),
    .A1(net85),
    .A2(net73),
    .A3(net1),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit26.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG0 ));
 sky130_fd_sc_hd__mux4_1 _066_ (.A0(net64),
    .A1(net68),
    .A2(net66),
    .A3(net70),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit25.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit24.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG15 ));
 sky130_fd_sc_hd__mux4_1 _067_ (.A0(net63),
    .A1(net67),
    .A2(net65),
    .A3(net69),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit23.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit22.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG14 ));
 sky130_fd_sc_hd__mux4_1 _068_ (.A0(net80),
    .A1(net73),
    .A2(net82),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit21.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit20.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG13 ));
 sky130_fd_sc_hd__mux4_1 _069_ (.A0(net74),
    .A1(net78),
    .A2(net76),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit19.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit18.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG12 ));
 sky130_fd_sc_hd__mux4_1 _070_ (.A0(net79),
    .A1(net72),
    .A2(net81),
    .A3(net2),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit17.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit16.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG11 ));
 sky130_fd_sc_hd__mux4_1 _071_ (.A0(net71),
    .A1(net77),
    .A2(net75),
    .A3(net1),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit15.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit14.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG10 ));
 sky130_fd_sc_hd__mux4_1 _072_ (.A0(net74),
    .A1(net78),
    .A2(net76),
    .A3(net80),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit13.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit12.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG9 ));
 sky130_fd_sc_hd__mux4_1 _073_ (.A0(net77),
    .A1(net81),
    .A2(net79),
    .A3(net72),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit11.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit10.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG8 ));
 sky130_fd_sc_hd__mux4_1 _074_ (.A0(net64),
    .A1(net68),
    .A2(net66),
    .A3(net70),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit9.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit8.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG7 ));
 sky130_fd_sc_hd__mux4_1 _075_ (.A0(net63),
    .A1(net67),
    .A2(net65),
    .A3(net69),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit7.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit6.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG6 ));
 sky130_fd_sc_hd__mux4_1 _076_ (.A0(net41),
    .A1(net43),
    .A2(net60),
    .A3(net62),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit5.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG5 ));
 sky130_fd_sc_hd__mux4_1 _077_ (.A0(net40),
    .A1(net42),
    .A2(net59),
    .A3(net61),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit2.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit3.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG4 ));
 sky130_fd_sc_hd__mux4_1 _078_ (.A0(net80),
    .A1(net73),
    .A2(net82),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit1.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit0.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _079_ (.A0(net74),
    .A1(net78),
    .A2(net76),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit31.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit30.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _080_ (.A0(net79),
    .A1(net72),
    .A2(net81),
    .A3(net2),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit29.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit28.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _081_ (.A0(net71),
    .A1(net77),
    .A2(net75),
    .A3(net1),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit27.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit26.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _082_ (.A0(net40),
    .A1(net83),
    .A2(net97),
    .A3(net71),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit25.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb7 ));
 sky130_fd_sc_hd__mux4_1 _083_ (.A0(net41),
    .A1(net90),
    .A2(net98),
    .A3(net74),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit22.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit23.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb6 ));
 sky130_fd_sc_hd__mux4_1 _084_ (.A0(net42),
    .A1(net91),
    .A2(net84),
    .A3(net75),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit21.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb5 ));
 sky130_fd_sc_hd__mux4_1 _085_ (.A0(net43),
    .A1(net92),
    .A2(net85),
    .A3(net76),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit18.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit19.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb4 ));
 sky130_fd_sc_hd__mux4_1 _086_ (.A0(net59),
    .A1(net93),
    .A2(net86),
    .A3(net77),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit17.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb3 ));
 sky130_fd_sc_hd__mux4_1 _087_ (.A0(net60),
    .A1(net94),
    .A2(net87),
    .A3(net78),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit15.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb2 ));
 sky130_fd_sc_hd__mux4_1 _088_ (.A0(net61),
    .A1(net95),
    .A2(net88),
    .A3(net79),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit13.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb1 ));
 sky130_fd_sc_hd__mux4_1 _089_ (.A0(net62),
    .A1(net96),
    .A2(net89),
    .A3(net80),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit11.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb0 ));
 sky130_fd_sc_hd__mux4_1 _090_ (.A0(net63),
    .A1(net83),
    .A2(net97),
    .A3(net71),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit9.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEG7 ));
 sky130_fd_sc_hd__mux4_1 _091_ (.A0(net64),
    .A1(net90),
    .A2(net98),
    .A3(net74),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit7.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEG6 ));
 sky130_fd_sc_hd__mux4_1 _092_ (.A0(net65),
    .A1(net91),
    .A2(net84),
    .A3(net75),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit5.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEG5 ));
 sky130_fd_sc_hd__mux4_1 _093_ (.A0(net66),
    .A1(net92),
    .A2(net85),
    .A3(net76),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit2.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit3.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEG4 ));
 sky130_fd_sc_hd__mux4_1 _094_ (.A0(net67),
    .A1(net93),
    .A2(net86),
    .A3(net77),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit1.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEG3 ));
 sky130_fd_sc_hd__mux4_1 _095_ (.A0(net68),
    .A1(net94),
    .A2(net87),
    .A3(net78),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame3_bit30.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame3_bit31.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _096_ (.A0(net69),
    .A1(net95),
    .A2(net88),
    .A3(net79),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame3_bit29.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _097_ (.A0(net70),
    .A1(net96),
    .A2(net89),
    .A3(net80),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame3_bit26.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame3_bit27.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEG0 ));
 sky130_fd_sc_hd__mux2_1 _098_ (.A0(net36),
    .A1(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S(\Inst_W_IO_ConfigMem.Inst_frame3_bit25.Q ),
    .X(\Inst_W_IO_switch_matrix.E1BEG3 ));
 sky130_fd_sc_hd__mux2_1 _099_ (.A0(net37),
    .A1(net2),
    .S(\Inst_W_IO_ConfigMem.Inst_frame3_bit24.Q ),
    .X(\Inst_W_IO_switch_matrix.E1BEG2 ));
 sky130_fd_sc_hd__mux2_1 _100_ (.A0(net38),
    .A1(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S(\Inst_W_IO_ConfigMem.Inst_frame3_bit23.Q ),
    .X(\Inst_W_IO_switch_matrix.E1BEG1 ));
 sky130_fd_sc_hd__mux2_1 _101_ (.A0(net39),
    .A1(net1),
    .S(\Inst_W_IO_ConfigMem.Inst_frame3_bit22.Q ),
    .X(\Inst_W_IO_switch_matrix.E1BEG0 ));
 sky130_fd_sc_hd__mux2_1 _102_ (.A0(net70),
    .A1(net41),
    .S(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .X(_020_));
 sky130_fd_sc_hd__and3b_1 _103_ (.A_N(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .B(\Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .C(net43),
    .X(_021_));
 sky130_fd_sc_hd__a211oi_1 _104_ (.A1(_004_),
    .A2(_020_),
    .B1(_021_),
    .C1(\Inst_W_IO_ConfigMem.Inst_frame0_bit22.Q ),
    .Y(_022_));
 sky130_fd_sc_hd__or3b_1 _105_ (.A(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .B(\Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .C_N(net40),
    .X(_023_));
 sky130_fd_sc_hd__o21ai_1 _106_ (.A1(net59),
    .A2(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .B1(\Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .Y(_024_));
 sky130_fd_sc_hd__nand2_1 _107_ (.A(net42),
    .B(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .Y(_025_));
 sky130_fd_sc_hd__a41o_1 _108_ (.A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit22.Q ),
    .A2(_023_),
    .A3(_024_),
    .A4(_025_),
    .B1(_022_),
    .X(net100));
 sky130_fd_sc_hd__mux2_1 _109_ (.A0(net69),
    .A1(net40),
    .S(\Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_026_));
 sky130_fd_sc_hd__and3b_1 _110_ (.A_N(\Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .B(\Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .C(net60),
    .X(_027_));
 sky130_fd_sc_hd__a211oi_1 _111_ (.A1(_005_),
    .A2(_026_),
    .B1(_027_),
    .C1(\Inst_W_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_028_));
 sky130_fd_sc_hd__or3b_1 _112_ (.A(\Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .B(\Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .C_N(net70),
    .X(_029_));
 sky130_fd_sc_hd__o21ai_1 _113_ (.A1(net61),
    .A2(\Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .B1(\Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_030_));
 sky130_fd_sc_hd__nand2_1 _114_ (.A(net59),
    .B(\Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .Y(_031_));
 sky130_fd_sc_hd__a41o_1 _115_ (.A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_029_),
    .A3(_030_),
    .A4(_031_),
    .B1(_028_),
    .X(net106));
 sky130_fd_sc_hd__dlxtp_1 _116_ (.D(net8),
    .GATE(net44),
    .Q(net101));
 sky130_fd_sc_hd__dlxtp_1 _117_ (.D(net9),
    .GATE(net44),
    .Q(net102));
 sky130_fd_sc_hd__dlxtp_1 _118_ (.D(net10),
    .GATE(net44),
    .Q(net103));
 sky130_fd_sc_hd__dlxtp_1 _119_ (.D(net11),
    .GATE(net44),
    .Q(net104));
 sky130_fd_sc_hd__dlxtp_1 _120_ (.D(net12),
    .GATE(net44),
    .Q(net107));
 sky130_fd_sc_hd__dlxtp_1 _121_ (.D(net13),
    .GATE(net44),
    .Q(net108));
 sky130_fd_sc_hd__dlxtp_1 _122_ (.D(net15),
    .GATE(net44),
    .Q(net109));
 sky130_fd_sc_hd__dlxtp_1 _123_ (.D(net16),
    .GATE(net45),
    .Q(net110));
 sky130_fd_sc_hd__dlxtp_1 _124_ (.D(net17),
    .GATE(net44),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _125_ (.D(net18),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _126_ (.D(net19),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _127_ (.D(net20),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _128_ (.D(net21),
    .GATE(net45),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _129_ (.D(net22),
    .GATE(net45),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _130_ (.D(net23),
    .GATE(net45),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _131_ (.D(net24),
    .GATE(net45),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _132_ (.D(net26),
    .GATE(net44),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _133_ (.D(net27),
    .GATE(net44),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _134_ (.D(net3),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _135_ (.D(net14),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _136_ (.D(net25),
    .GATE(net49),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _137_ (.D(net28),
    .GATE(net49),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _138_ (.D(net29),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _139_ (.D(net30),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _140_ (.D(net31),
    .GATE(net49),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _141_ (.D(net32),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _142_ (.D(net33),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _143_ (.D(net34),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _144_ (.D(net4),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _145_ (.D(net5),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _146_ (.D(net6),
    .GATE(net50),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _147_ (.D(net7),
    .GATE(net50),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _148_ (.D(net8),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _149_ (.D(net9),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _150_ (.D(net10),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _151_ (.D(net11),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _152_ (.D(net12),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _153_ (.D(net13),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _154_ (.D(net15),
    .GATE(net49),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _155_ (.D(net16),
    .GATE(net49),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _156_ (.D(net17),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _157_ (.D(net18),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _158_ (.D(net19),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _159_ (.D(net20),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _160_ (.D(net21),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _161_ (.D(net22),
    .GATE(net50),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _162_ (.D(net23),
    .GATE(net50),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _163_ (.D(net24),
    .GATE(net50),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _164_ (.D(net26),
    .GATE(net50),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _165_ (.D(net27),
    .GATE(net50),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _166_ (.D(net3),
    .GATE(net52),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _167_ (.D(net14),
    .GATE(net52),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _168_ (.D(net25),
    .GATE(net51),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _169_ (.D(net28),
    .GATE(net51),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _170_ (.D(net29),
    .GATE(net51),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _171_ (.D(net30),
    .GATE(net51),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _172_ (.D(net31),
    .GATE(net51),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _173_ (.D(net32),
    .GATE(net51),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _174_ (.D(net33),
    .GATE(net51),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _175_ (.D(net34),
    .GATE(net53),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _176_ (.D(net4),
    .GATE(net52),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _177_ (.D(net5),
    .GATE(net52),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _178_ (.D(net6),
    .GATE(net54),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _179_ (.D(net7),
    .GATE(net54),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _180_ (.D(net8),
    .GATE(net53),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _181_ (.D(net9),
    .GATE(net53),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _182_ (.D(net10),
    .GATE(net52),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _183_ (.D(net11),
    .GATE(net54),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _184_ (.D(net12),
    .GATE(net52),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _185_ (.D(net13),
    .GATE(net52),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _186_ (.D(net15),
    .GATE(net52),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _187_ (.D(net16),
    .GATE(net52),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _188_ (.D(net17),
    .GATE(net51),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _189_ (.D(net18),
    .GATE(net51),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _190_ (.D(net19),
    .GATE(net51),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _191_ (.D(net20),
    .GATE(net54),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _192_ (.D(net21),
    .GATE(net53),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _193_ (.D(net22),
    .GATE(net53),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _194_ (.D(net23),
    .GATE(net53),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _195_ (.D(net24),
    .GATE(net53),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _196_ (.D(net26),
    .GATE(net53),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _197_ (.D(net27),
    .GATE(net53),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _198_ (.D(net3),
    .GATE(net58),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _199_ (.D(net14),
    .GATE(net58),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _200_ (.D(net25),
    .GATE(net58),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _201_ (.D(net28),
    .GATE(net58),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _202_ (.D(net29),
    .GATE(net57),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _203_ (.D(net30),
    .GATE(net57),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _204_ (.D(net31),
    .GATE(net57),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _205_ (.D(net32),
    .GATE(net57),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _206_ (.D(net33),
    .GATE(net57),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _207_ (.D(net34),
    .GATE(net57),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _208_ (.D(net4),
    .GATE(net58),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _209_ (.D(net5),
    .GATE(net58),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _210_ (.D(net6),
    .GATE(net57),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _211_ (.D(net7),
    .GATE(net57),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _212_ (.D(net8),
    .GATE(net58),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _213_ (.D(net9),
    .GATE(net58),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _214_ (.D(net10),
    .GATE(net57),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _215_ (.D(net11),
    .GATE(net57),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _216_ (.D(net12),
    .GATE(net56),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _217_ (.D(net13),
    .GATE(net55),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _218_ (.D(net15),
    .GATE(net55),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _219_ (.D(net16),
    .GATE(net55),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _220_ (.D(net17),
    .GATE(net55),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _221_ (.D(net18),
    .GATE(net55),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _222_ (.D(net19),
    .GATE(net55),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _223_ (.D(net20),
    .GATE(net55),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _224_ (.D(net21),
    .GATE(net55),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _225_ (.D(net22),
    .GATE(net55),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _226_ (.D(net23),
    .GATE(net55),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _227_ (.D(net24),
    .GATE(net56),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _228_ (.D(net26),
    .GATE(net56),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _229_ (.D(net27),
    .GATE(net56),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q ));
 sky130_fd_sc_hd__dfxtp_1 _230_ (.CLK(clknet_1_0__leaf_UserCLK_regs),
    .D(net1),
    .Q(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ));
 sky130_fd_sc_hd__dfxtp_1 _231_ (.CLK(clknet_1_1__leaf_UserCLK_regs),
    .D(net2),
    .Q(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ));
 sky130_fd_sc_hd__buf_1 _232_ (.A(\Inst_W_IO_switch_matrix.E6BEG5 ),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 _233_ (.A(\Inst_W_IO_switch_matrix.E6BEG6 ),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 _234_ (.A(\Inst_W_IO_switch_matrix.E6BEG7 ),
    .X(net140));
 sky130_fd_sc_hd__buf_1 _235_ (.A(\Inst_W_IO_switch_matrix.E6BEG8 ),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 _236_ (.A(\Inst_W_IO_switch_matrix.E6BEG9 ),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 _237_ (.A(\Inst_W_IO_switch_matrix.E6BEG10 ),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 _238_ (.A(\Inst_W_IO_switch_matrix.E6BEG11 ),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 _239_ (.A(\Inst_W_IO_switch_matrix.EE4BEG0 ),
    .X(net143));
 sky130_fd_sc_hd__buf_1 _240_ (.A(\Inst_W_IO_switch_matrix.EE4BEG1 ),
    .X(net150));
 sky130_fd_sc_hd__buf_1 _241_ (.A(\Inst_W_IO_switch_matrix.EE4BEG2 ),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 _242_ (.A(\Inst_W_IO_switch_matrix.EE4BEG3 ),
    .X(net152));
 sky130_fd_sc_hd__buf_1 _243_ (.A(\Inst_W_IO_switch_matrix.EE4BEG4 ),
    .X(net153));
 sky130_fd_sc_hd__buf_1 _244_ (.A(\Inst_W_IO_switch_matrix.EE4BEG5 ),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 _245_ (.A(\Inst_W_IO_switch_matrix.EE4BEG6 ),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 _246_ (.A(\Inst_W_IO_switch_matrix.EE4BEG7 ),
    .X(net156));
 sky130_fd_sc_hd__buf_1 _247_ (.A(\Inst_W_IO_switch_matrix.EE4BEG8 ),
    .X(net157));
 sky130_fd_sc_hd__buf_1 _248_ (.A(\Inst_W_IO_switch_matrix.EE4BEG9 ),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 _249_ (.A(\Inst_W_IO_switch_matrix.EE4BEG10 ),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 _250_ (.A(\Inst_W_IO_switch_matrix.EE4BEG11 ),
    .X(net145));
 sky130_fd_sc_hd__buf_1 _251_ (.A(\Inst_W_IO_switch_matrix.EE4BEG12 ),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 _252_ (.A(\Inst_W_IO_switch_matrix.EE4BEG13 ),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 _253_ (.A(\Inst_W_IO_switch_matrix.EE4BEG14 ),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 _254_ (.A(\Inst_W_IO_switch_matrix.EE4BEG15 ),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 _255_ (.A(net3),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 _256_ (.A(net14),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 _257_ (.A(net25),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_2 _258_ (.A(net28),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 _259_ (.A(net29),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_2 _260_ (.A(net30),
    .X(net186));
 sky130_fd_sc_hd__buf_1 _261_ (.A(net31),
    .X(net187));
 sky130_fd_sc_hd__buf_1 _262_ (.A(net32),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 _263_ (.A(net33),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 _264_ (.A(net34),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 _265_ (.A(net4),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 _266_ (.A(net5),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 _267_ (.A(net6),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 _268_ (.A(net7),
    .X(net163));
 sky130_fd_sc_hd__buf_1 _269_ (.A(net8),
    .X(net164));
 sky130_fd_sc_hd__buf_1 _270_ (.A(net9),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 _271_ (.A(net10),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 _272_ (.A(net11),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 _273_ (.A(net12),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 _274_ (.A(net13),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 _275_ (.A(net15),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 _276_ (.A(net16),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_2 _277_ (.A(net17),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 _278_ (.A(net18),
    .X(net174));
 sky130_fd_sc_hd__buf_1 _279_ (.A(net19),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 _280_ (.A(net20),
    .X(net176));
 sky130_fd_sc_hd__buf_1 _281_ (.A(net21),
    .X(net177));
 sky130_fd_sc_hd__buf_1 _282_ (.A(net22),
    .X(net178));
 sky130_fd_sc_hd__buf_1 _283_ (.A(net23),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 _284_ (.A(net24),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 _285_ (.A(net26),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 _286_ (.A(net27),
    .X(net183));
 sky130_fd_sc_hd__buf_1 _287_ (.A(net58),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 _288_ (.A(net52),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 _289_ (.A(net50),
    .X(net203));
 sky130_fd_sc_hd__buf_1 _290_ (.A(net46),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 _291_ (.A(FrameStrobe[4]),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 _292_ (.A(FrameStrobe[5]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_1 _293_ (.A(FrameStrobe[6]),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 _294_ (.A(FrameStrobe[7]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 _295_ (.A(FrameStrobe[8]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_1 _296_ (.A(FrameStrobe[9]),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_1 _297_ (.A(FrameStrobe[10]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 _298_ (.A(FrameStrobe[11]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 _299_ (.A(FrameStrobe[12]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 _300_ (.A(FrameStrobe[13]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 _301_ (.A(FrameStrobe[14]),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 _302_ (.A(FrameStrobe[15]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_1 _303_ (.A(FrameStrobe[16]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 _304_ (.A(FrameStrobe[17]),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_1 _305_ (.A(FrameStrobe[18]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 _306_ (.A(FrameStrobe[19]),
    .X(net201));
 sky130_fd_sc_hd__buf_2 _307_ (.A(clknet_1_0__leaf_UserCLK),
    .X(net211));
 sky130_fd_sc_hd__buf_1 _308_ (.A(\Inst_W_IO_switch_matrix.E1BEG0 ),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 _309_ (.A(\Inst_W_IO_switch_matrix.E1BEG1 ),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 _310_ (.A(\Inst_W_IO_switch_matrix.E1BEG2 ),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 _311_ (.A(\Inst_W_IO_switch_matrix.E1BEG3 ),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 _312_ (.A(\Inst_W_IO_switch_matrix.E2BEG0 ),
    .X(net115));
 sky130_fd_sc_hd__buf_1 _313_ (.A(\Inst_W_IO_switch_matrix.E2BEG1 ),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 _314_ (.A(\Inst_W_IO_switch_matrix.E2BEG2 ),
    .X(net117));
 sky130_fd_sc_hd__buf_1 _315_ (.A(\Inst_W_IO_switch_matrix.E2BEG3 ),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 _316_ (.A(\Inst_W_IO_switch_matrix.E2BEG4 ),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 _317_ (.A(\Inst_W_IO_switch_matrix.E2BEG5 ),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 _318_ (.A(\Inst_W_IO_switch_matrix.E2BEG6 ),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 _319_ (.A(\Inst_W_IO_switch_matrix.E2BEG7 ),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 _320_ (.A(\Inst_W_IO_switch_matrix.E2BEGb0 ),
    .X(net123));
 sky130_fd_sc_hd__buf_1 _321_ (.A(\Inst_W_IO_switch_matrix.E2BEGb1 ),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 _322_ (.A(\Inst_W_IO_switch_matrix.E2BEGb2 ),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 _323_ (.A(\Inst_W_IO_switch_matrix.E2BEGb3 ),
    .X(net126));
 sky130_fd_sc_hd__buf_1 _324_ (.A(\Inst_W_IO_switch_matrix.E2BEGb4 ),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 _325_ (.A(\Inst_W_IO_switch_matrix.E2BEGb5 ),
    .X(net128));
 sky130_fd_sc_hd__buf_1 _326_ (.A(\Inst_W_IO_switch_matrix.E2BEGb6 ),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 _327_ (.A(\Inst_W_IO_switch_matrix.E2BEGb7 ),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 _328_ (.A(\Inst_W_IO_switch_matrix.E6BEG0 ),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 _329_ (.A(\Inst_W_IO_switch_matrix.E6BEG1 ),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 _330_ (.A(\Inst_W_IO_switch_matrix.E6BEG2 ),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 _331_ (.A(\Inst_W_IO_switch_matrix.E6BEG3 ),
    .X(net136));
 sky130_fd_sc_hd__buf_1 _332_ (.A(\Inst_W_IO_switch_matrix.E6BEG4 ),
    .X(net137));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_261 ();
 sky130_fd_sc_hd__buf_2 fanout44 (.A(net46),
    .X(net44));
 sky130_fd_sc_hd__buf_1 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 fanout46 (.A(FrameStrobe[3]),
    .X(net46));
 sky130_fd_sc_hd__buf_2 fanout47 (.A(net48),
    .X(net47));
 sky130_fd_sc_hd__buf_2 fanout48 (.A(net50),
    .X(net48));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout49 (.A(net50),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 fanout50 (.A(net35),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 fanout51 (.A(net54),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 fanout52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 fanout53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 fanout54 (.A(FrameStrobe[1]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__buf_1 fanout56 (.A(FrameStrobe[0]),
    .X(net56));
 sky130_fd_sc_hd__buf_2 fanout57 (.A(net58),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 fanout58 (.A(FrameStrobe[0]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(A_O_top),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(B_O_top),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(FrameData[0]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(FrameData[10]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(FrameData[11]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(FrameData[12]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(FrameData[13]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(FrameData[14]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(FrameData[15]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(FrameData[16]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(FrameData[17]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(FrameData[18]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(FrameData[19]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(FrameData[1]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(FrameData[20]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(FrameData[21]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(FrameData[22]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(FrameData[23]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(FrameData[24]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(FrameData[25]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(FrameData[26]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(FrameData[27]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(FrameData[28]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(FrameData[29]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(FrameData[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(FrameData[30]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(FrameData[31]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(FrameData[3]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(FrameData[4]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(FrameData[5]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(FrameData[6]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(FrameData[7]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(FrameData[8]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(FrameData[9]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(FrameStrobe[2]),
    .X(net35));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(W1END[0]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(W1END[1]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(W1END[2]),
    .X(net38));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(W1END[3]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(W2END[0]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(W2END[1]),
    .X(net41));
 sky130_fd_sc_hd__dlymetal6s2s_1 input42 (.A(W2END[2]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(W2END[3]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(W2END[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input45 (.A(W2END[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(W2END[6]),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 input47 (.A(W2END[7]),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 input48 (.A(W2MID[0]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input49 (.A(W2MID[1]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input50 (.A(W2MID[2]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input51 (.A(W2MID[3]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(W2MID[4]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input53 (.A(W2MID[5]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(W2MID[6]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(W2MID[7]),
    .X(net70));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(W6END[0]),
    .X(net71));
 sky130_fd_sc_hd__dlymetal6s2s_1 input57 (.A(W6END[10]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input58 (.A(W6END[11]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(W6END[1]),
    .X(net74));
 sky130_fd_sc_hd__dlymetal6s2s_1 input60 (.A(W6END[2]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(W6END[3]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(W6END[4]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(W6END[5]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(W6END[6]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(W6END[7]),
    .X(net80));
 sky130_fd_sc_hd__dlymetal6s2s_1 input66 (.A(W6END[8]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 input67 (.A(W6END[9]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input68 (.A(WW4END[0]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 input69 (.A(WW4END[10]),
    .X(net84));
 sky130_fd_sc_hd__buf_1 input70 (.A(WW4END[11]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input71 (.A(WW4END[12]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 input72 (.A(WW4END[13]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 input73 (.A(WW4END[14]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 input74 (.A(WW4END[15]),
    .X(net89));
 sky130_fd_sc_hd__buf_1 input75 (.A(WW4END[1]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input76 (.A(WW4END[2]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input77 (.A(WW4END[3]),
    .X(net92));
 sky130_fd_sc_hd__dlymetal6s2s_1 input78 (.A(WW4END[4]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 input79 (.A(WW4END[5]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 input80 (.A(WW4END[6]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(WW4END[7]),
    .X(net96));
 sky130_fd_sc_hd__buf_1 input82 (.A(WW4END[8]),
    .X(net97));
 sky130_fd_sc_hd__buf_1 input83 (.A(WW4END[9]),
    .X(net98));
 sky130_fd_sc_hd__buf_2 output84 (.A(net99),
    .X(A_I_top));
 sky130_fd_sc_hd__buf_2 output85 (.A(net100),
    .X(A_T_top));
 sky130_fd_sc_hd__buf_2 output86 (.A(net101),
    .X(A_config_C_bit0));
 sky130_fd_sc_hd__buf_2 output87 (.A(net102),
    .X(A_config_C_bit1));
 sky130_fd_sc_hd__buf_2 output88 (.A(net103),
    .X(A_config_C_bit2));
 sky130_fd_sc_hd__buf_2 output89 (.A(net104),
    .X(A_config_C_bit3));
 sky130_fd_sc_hd__buf_2 output90 (.A(net105),
    .X(B_I_top));
 sky130_fd_sc_hd__buf_2 output91 (.A(net106),
    .X(B_T_top));
 sky130_fd_sc_hd__buf_2 output92 (.A(net107),
    .X(B_config_C_bit0));
 sky130_fd_sc_hd__buf_2 output93 (.A(net108),
    .X(B_config_C_bit1));
 sky130_fd_sc_hd__buf_2 output94 (.A(net109),
    .X(B_config_C_bit2));
 sky130_fd_sc_hd__buf_2 output95 (.A(net110),
    .X(B_config_C_bit3));
 sky130_fd_sc_hd__buf_2 output96 (.A(net111),
    .X(E1BEG[0]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net112),
    .X(E1BEG[1]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net113),
    .X(E1BEG[2]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net114),
    .X(E1BEG[3]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net115),
    .X(E2BEG[0]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net116),
    .X(E2BEG[1]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net117),
    .X(E2BEG[2]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net118),
    .X(E2BEG[3]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net119),
    .X(E2BEG[4]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net120),
    .X(E2BEG[5]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net121),
    .X(E2BEG[6]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net122),
    .X(E2BEG[7]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net123),
    .X(E2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net124),
    .X(E2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net125),
    .X(E2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net126),
    .X(E2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net127),
    .X(E2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net128),
    .X(E2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net129),
    .X(E2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net130),
    .X(E2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net131),
    .X(E6BEG[0]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net132),
    .X(E6BEG[10]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net133),
    .X(E6BEG[11]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net134),
    .X(E6BEG[1]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net135),
    .X(E6BEG[2]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net136),
    .X(E6BEG[3]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net137),
    .X(E6BEG[4]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net138),
    .X(E6BEG[5]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net139),
    .X(E6BEG[6]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net140),
    .X(E6BEG[7]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net141),
    .X(E6BEG[8]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net142),
    .X(E6BEG[9]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net143),
    .X(EE4BEG[0]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net144),
    .X(EE4BEG[10]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net145),
    .X(EE4BEG[11]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net146),
    .X(EE4BEG[12]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net147),
    .X(EE4BEG[13]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net148),
    .X(EE4BEG[14]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net149),
    .X(EE4BEG[15]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net150),
    .X(EE4BEG[1]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net151),
    .X(EE4BEG[2]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net152),
    .X(EE4BEG[3]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net153),
    .X(EE4BEG[4]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net154),
    .X(EE4BEG[5]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net155),
    .X(EE4BEG[6]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net156),
    .X(EE4BEG[7]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net157),
    .X(EE4BEG[8]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net158),
    .X(EE4BEG[9]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net159),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net160),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net161),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net162),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net163),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net164),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net165),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net166),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net167),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net168),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net169),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net170),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net171),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net172),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net173),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net174),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net175),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output161 (.A(net176),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net177),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net178),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net179),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net180),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net181),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net182),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net183),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net184),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net185),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net186),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net187),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net188),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net189),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net190),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output176 (.A(net191),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output177 (.A(net192),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output178 (.A(net193),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output179 (.A(net194),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net195),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output181 (.A(net196),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output182 (.A(net197),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net198),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output184 (.A(net199),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net200),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output186 (.A(net201),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output187 (.A(net202),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output188 (.A(net203),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net204),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output190 (.A(net205),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output191 (.A(net206),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output192 (.A(net207),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output193 (.A(net208),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output194 (.A(net209),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output195 (.A(net210),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_1 output196 (.A(net211),
    .X(UserCLKo));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_regs_0_UserCLK (.A(UserCLK),
    .X(UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_UserCLK (.A(UserCLK),
    .X(clknet_0_UserCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_UserCLK (.A(clknet_0_UserCLK),
    .X(clknet_1_0__leaf_UserCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_UserCLK_regs (.A(UserCLK_regs),
    .X(clknet_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_1_0__leaf_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_1_1__leaf_UserCLK_regs));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(FrameStrobe[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(FrameStrobe[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(FrameStrobe[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(FrameStrobe[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(FrameStrobe[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(FrameStrobe[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(FrameStrobe[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(FrameStrobe[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(FrameStrobe[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(FrameStrobe[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(FrameStrobe[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(FrameStrobe[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(FrameStrobe[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(FrameStrobe[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(FrameStrobe[5]));
 sky130_fd_sc_hd__decap_8 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_5 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_5 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_93 ();
endmodule
